module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 ;
  assign n129 = ( x1 & ~x63 ) | ( x1 & x120 ) | ( ~x63 & x120 ) ;
  assign n130 = x66 ^ x13 ^ 1'b0 ;
  assign n131 = x97 & n130 ;
  assign n132 = ( x50 & x54 ) | ( x50 & ~x122 ) | ( x54 & ~x122 ) ;
  assign n133 = x62 & n132 ;
  assign n134 = ~x9 & n133 ;
  assign n135 = x104 ^ x55 ^ 1'b0 ;
  assign n136 = x45 & n135 ;
  assign n137 = ( ~x33 & x81 ) | ( ~x33 & x108 ) | ( x81 & x108 ) ;
  assign n138 = x16 & x36 ;
  assign n139 = n138 ^ x85 ^ 1'b0 ;
  assign n140 = x87 & ~n139 ;
  assign n141 = ~x39 & n140 ;
  assign n142 = x106 ^ x5 ^ 1'b0 ;
  assign n143 = x93 & n142 ;
  assign n144 = x84 ^ x43 ^ x16 ;
  assign n145 = n144 ^ x6 ^ 1'b0 ;
  assign n146 = x106 & ~n145 ;
  assign n147 = ( x21 & ~x51 ) | ( x21 & x93 ) | ( ~x51 & x93 ) ;
  assign n148 = x87 & n147 ;
  assign n149 = ~x26 & n148 ;
  assign n150 = n149 ^ x43 ^ 1'b0 ;
  assign n151 = x93 & ~n150 ;
  assign n153 = x114 ^ x78 ^ x27 ;
  assign n154 = n153 ^ x108 ^ x50 ;
  assign n152 = x45 & x51 ;
  assign n155 = n154 ^ n152 ^ 1'b0 ;
  assign n156 = ( ~x65 & n151 ) | ( ~x65 & n155 ) | ( n151 & n155 ) ;
  assign n158 = x115 ^ x36 ^ x29 ;
  assign n159 = n158 ^ x40 ^ x3 ;
  assign n157 = ( x25 & x26 ) | ( x25 & ~x112 ) | ( x26 & ~x112 ) ;
  assign n160 = n159 ^ n157 ^ x16 ;
  assign n161 = ( x41 & x74 ) | ( x41 & ~x116 ) | ( x74 & ~x116 ) ;
  assign n162 = n161 ^ n146 ^ x17 ;
  assign n163 = x70 & x74 ;
  assign n164 = n163 ^ x41 ^ 1'b0 ;
  assign n165 = ( x49 & ~x83 ) | ( x49 & n158 ) | ( ~x83 & n158 ) ;
  assign n166 = x77 ^ x23 ^ 1'b0 ;
  assign n167 = ~n165 & n166 ;
  assign n168 = ( x14 & ~x56 ) | ( x14 & x86 ) | ( ~x56 & x86 ) ;
  assign n169 = ( ~x50 & x76 ) | ( ~x50 & x92 ) | ( x76 & x92 ) ;
  assign n170 = x88 & n169 ;
  assign n171 = x72 ^ x16 ^ 1'b0 ;
  assign n172 = n157 ^ x122 ^ 1'b0 ;
  assign n173 = x107 & n172 ;
  assign n174 = ( ~x50 & x77 ) | ( ~x50 & x79 ) | ( x77 & x79 ) ;
  assign n175 = n134 ^ x44 ^ 1'b0 ;
  assign n176 = x120 & ~n175 ;
  assign n177 = x110 ^ x34 ^ 1'b0 ;
  assign n178 = n176 & n177 ;
  assign n179 = x73 ^ x45 ^ 1'b0 ;
  assign n180 = n147 & n179 ;
  assign n181 = x76 ^ x56 ^ 1'b0 ;
  assign n182 = x72 & n181 ;
  assign n183 = x118 & n182 ;
  assign n184 = ~x64 & n183 ;
  assign n185 = x19 & x30 ;
  assign n186 = n185 ^ x103 ^ 1'b0 ;
  assign n187 = ( x58 & x111 ) | ( x58 & n186 ) | ( x111 & n186 ) ;
  assign n188 = ( x62 & ~x95 ) | ( x62 & x111 ) | ( ~x95 & x111 ) ;
  assign n189 = x56 & n188 ;
  assign n190 = n189 ^ x36 ^ 1'b0 ;
  assign n191 = n190 ^ x126 ^ x117 ;
  assign n192 = ( x116 & n171 ) | ( x116 & ~n191 ) | ( n171 & ~n191 ) ;
  assign n193 = x44 & ~n164 ;
  assign n194 = n193 ^ n180 ^ 1'b0 ;
  assign n195 = x34 & x84 ;
  assign n196 = n195 ^ x101 ^ 1'b0 ;
  assign n197 = x76 ^ x49 ^ x41 ;
  assign n198 = x94 ^ x56 ^ x0 ;
  assign n199 = ( x34 & ~n197 ) | ( x34 & n198 ) | ( ~n197 & n198 ) ;
  assign n200 = x103 ^ x31 ^ 1'b0 ;
  assign n201 = n200 ^ n178 ^ 1'b0 ;
  assign n202 = n143 & ~n201 ;
  assign n203 = x19 & ~x23 ;
  assign n204 = ( ~x59 & x113 ) | ( ~x59 & n203 ) | ( x113 & n203 ) ;
  assign n205 = n204 ^ x79 ^ x18 ;
  assign n212 = x126 ^ x60 ^ 1'b0 ;
  assign n213 = x117 & n212 ;
  assign n207 = n129 ^ x86 ^ x2 ;
  assign n206 = x86 ^ x46 ^ x11 ;
  assign n208 = n207 ^ n206 ^ x96 ;
  assign n209 = n151 | n208 ;
  assign n210 = ( x99 & n156 ) | ( x99 & ~n209 ) | ( n156 & ~n209 ) ;
  assign n211 = n210 ^ n176 ^ n171 ;
  assign n214 = n213 ^ n211 ^ x72 ;
  assign n215 = x82 ^ x7 ^ 1'b0 ;
  assign n216 = x78 & n215 ;
  assign n217 = x49 & n216 ;
  assign n218 = ~n214 & n217 ;
  assign n219 = x89 ^ x33 ^ 1'b0 ;
  assign n220 = n219 ^ x24 ^ 1'b0 ;
  assign n221 = ~n218 & n220 ;
  assign n222 = ( ~x10 & x34 ) | ( ~x10 & x121 ) | ( x34 & x121 ) ;
  assign n223 = n159 & n222 ;
  assign n224 = ~x70 & n223 ;
  assign n225 = n169 ^ x114 ^ 1'b0 ;
  assign n226 = ~n224 & n225 ;
  assign n227 = n226 ^ x24 ^ 1'b0 ;
  assign n228 = n178 ^ x60 ^ x40 ;
  assign n229 = x102 & ~n190 ;
  assign n230 = ~x70 & n229 ;
  assign n231 = x104 & x119 ;
  assign n232 = n231 ^ x107 ^ 1'b0 ;
  assign n233 = ( x52 & n230 ) | ( x52 & n232 ) | ( n230 & n232 ) ;
  assign n234 = ( ~x47 & x94 ) | ( ~x47 & n233 ) | ( x94 & n233 ) ;
  assign n241 = ( x78 & ~n151 ) | ( x78 & n190 ) | ( ~n151 & n190 ) ;
  assign n235 = x126 ^ x39 ^ 1'b0 ;
  assign n236 = x66 & n235 ;
  assign n237 = n136 ^ x53 ^ x24 ;
  assign n238 = ( ~x115 & n137 ) | ( ~x115 & n237 ) | ( n137 & n237 ) ;
  assign n239 = n236 | n238 ;
  assign n240 = ~n158 & n239 ;
  assign n242 = n241 ^ n240 ^ 1'b0 ;
  assign n244 = x88 & n137 ;
  assign n245 = n244 ^ x58 ^ 1'b0 ;
  assign n243 = ~x6 & x56 ;
  assign n246 = n245 ^ n243 ^ 1'b0 ;
  assign n247 = ~n136 & n187 ;
  assign n248 = n159 ^ x77 ^ x4 ;
  assign n249 = x21 & x36 ;
  assign n250 = n248 & n249 ;
  assign n251 = ~x26 & x81 ;
  assign n252 = n251 ^ x15 ^ 1'b0 ;
  assign n253 = n184 | n252 ;
  assign n255 = ( ~x0 & x125 ) | ( ~x0 & n236 ) | ( x125 & n236 ) ;
  assign n254 = x19 & n222 ;
  assign n256 = n255 ^ n254 ^ 1'b0 ;
  assign n257 = n151 ^ x62 ^ x4 ;
  assign n258 = x79 & ~n257 ;
  assign n259 = n256 & n258 ;
  assign n260 = n230 ^ x77 ^ x60 ;
  assign n263 = x71 & n191 ;
  assign n264 = n263 ^ x93 ^ 1'b0 ;
  assign n261 = x63 & x82 ;
  assign n262 = ~n216 & n261 ;
  assign n265 = n264 ^ n262 ^ n191 ;
  assign n266 = n265 ^ n167 ^ x93 ;
  assign n267 = n198 ^ x99 ^ 1'b0 ;
  assign n268 = x125 ^ x56 ^ 1'b0 ;
  assign n269 = x108 & n268 ;
  assign n270 = ( n154 & n247 ) | ( n154 & n269 ) | ( n247 & n269 ) ;
  assign n271 = x3 & x11 ;
  assign n272 = ~n219 & n271 ;
  assign n273 = x96 & ~n171 ;
  assign n274 = n273 ^ x24 ^ 1'b0 ;
  assign n275 = n274 ^ x17 ^ 1'b0 ;
  assign n276 = n275 ^ x73 ^ 1'b0 ;
  assign n277 = n243 | n276 ;
  assign n278 = x14 & x71 ;
  assign n279 = n206 & n278 ;
  assign n280 = n279 ^ x90 ^ 1'b0 ;
  assign n281 = n280 ^ x75 ^ x10 ;
  assign n282 = x8 & n180 ;
  assign n283 = ~x113 & n282 ;
  assign n284 = n277 | n283 ;
  assign n285 = n209 | n284 ;
  assign n286 = x60 ^ x6 ^ 1'b0 ;
  assign n287 = x58 & n286 ;
  assign n288 = n188 & n287 ;
  assign n289 = ~x111 & n288 ;
  assign n290 = ( x96 & x108 ) | ( x96 & n289 ) | ( x108 & n289 ) ;
  assign n291 = ~x44 & n290 ;
  assign n292 = n219 ^ n188 ^ 1'b0 ;
  assign n293 = ( ~n178 & n291 ) | ( ~n178 & n292 ) | ( n291 & n292 ) ;
  assign n294 = x127 ^ x25 ^ x4 ;
  assign n295 = ( n129 & n224 ) | ( n129 & n294 ) | ( n224 & n294 ) ;
  assign n302 = ( ~x5 & x7 ) | ( ~x5 & x79 ) | ( x7 & x79 ) ;
  assign n303 = n302 ^ x24 ^ 1'b0 ;
  assign n304 = ~n153 & n303 ;
  assign n296 = x118 | n149 ;
  assign n299 = n155 ^ x54 ^ x52 ;
  assign n297 = n255 ^ n234 ^ 1'b0 ;
  assign n298 = x46 & ~n297 ;
  assign n300 = n299 ^ n298 ^ 1'b0 ;
  assign n301 = ~n296 & n300 ;
  assign n305 = n304 ^ n301 ^ 1'b0 ;
  assign n306 = ( x15 & x109 ) | ( x15 & n232 ) | ( x109 & n232 ) ;
  assign n307 = n134 | n306 ;
  assign n308 = n307 ^ x127 ^ x58 ;
  assign n309 = x69 ^ x46 ^ 1'b0 ;
  assign n310 = n298 & n309 ;
  assign n311 = x98 & ~n162 ;
  assign n312 = n311 ^ x53 ^ 1'b0 ;
  assign n313 = x44 & x124 ;
  assign n314 = n313 ^ x7 ^ 1'b0 ;
  assign n315 = n169 ^ x66 ^ x29 ;
  assign n316 = n159 ^ x19 ^ 1'b0 ;
  assign n317 = ~n315 & n316 ;
  assign n318 = n314 & n317 ;
  assign n319 = ( x48 & ~x94 ) | ( x48 & n241 ) | ( ~x94 & n241 ) ;
  assign n320 = ~n171 & n319 ;
  assign n321 = n320 ^ n238 ^ 1'b0 ;
  assign n322 = ( n312 & n318 ) | ( n312 & n321 ) | ( n318 & n321 ) ;
  assign n324 = x6 & x48 ;
  assign n325 = ~n191 & n324 ;
  assign n326 = x98 & ~n325 ;
  assign n327 = ~x105 & n326 ;
  assign n323 = x55 ^ x28 ^ 1'b0 ;
  assign n328 = n327 ^ n323 ^ n279 ;
  assign n336 = x47 ^ x43 ^ 1'b0 ;
  assign n337 = x85 & n336 ;
  assign n333 = ( x86 & x89 ) | ( x86 & n160 ) | ( x89 & n160 ) ;
  assign n334 = n333 ^ n134 ^ x74 ;
  assign n335 = ( x18 & x65 ) | ( x18 & ~n334 ) | ( x65 & ~n334 ) ;
  assign n330 = x41 & x93 ;
  assign n331 = ~x115 & n330 ;
  assign n329 = ( x73 & ~x101 ) | ( x73 & n204 ) | ( ~x101 & n204 ) ;
  assign n332 = n331 ^ n329 ^ x105 ;
  assign n338 = n337 ^ n335 ^ n332 ;
  assign n339 = x20 | n248 ;
  assign n340 = x44 ^ x27 ^ 1'b0 ;
  assign n341 = n339 & n340 ;
  assign n342 = n209 & n341 ;
  assign n343 = ~n337 & n342 ;
  assign n344 = x67 | n343 ;
  assign n345 = x30 & ~n149 ;
  assign n346 = n345 ^ x4 ^ 1'b0 ;
  assign n347 = ( x10 & n141 ) | ( x10 & n149 ) | ( n141 & n149 ) ;
  assign n348 = ( x49 & ~n346 ) | ( x49 & n347 ) | ( ~n346 & n347 ) ;
  assign n349 = n221 ^ n202 ^ x117 ;
  assign n350 = x55 & n136 ;
  assign n351 = x53 & n350 ;
  assign n352 = ~n239 & n351 ;
  assign n359 = n151 ^ x26 ^ 1'b0 ;
  assign n360 = ~n158 & n359 ;
  assign n357 = n186 ^ n159 ^ 1'b0 ;
  assign n353 = x53 & x83 ;
  assign n354 = n353 ^ n346 ^ 1'b0 ;
  assign n355 = ~n319 & n354 ;
  assign n356 = n355 ^ n158 ^ 1'b0 ;
  assign n358 = n357 ^ n356 ^ n302 ;
  assign n361 = n360 ^ n358 ^ n232 ;
  assign n364 = x14 & n159 ;
  assign n362 = x84 & ~n162 ;
  assign n363 = ~x81 & n362 ;
  assign n365 = n364 ^ n363 ^ x121 ;
  assign n366 = ~n361 & n365 ;
  assign n367 = n227 & n315 ;
  assign n368 = n367 ^ n180 ^ x47 ;
  assign n369 = ~x15 & x37 ;
  assign n370 = n369 ^ n184 ^ 1'b0 ;
  assign n371 = n233 ^ x82 ^ x68 ;
  assign n372 = ( x72 & x82 ) | ( x72 & n241 ) | ( x82 & n241 ) ;
  assign n373 = ( x5 & ~x88 ) | ( x5 & n237 ) | ( ~x88 & n237 ) ;
  assign n374 = n373 ^ n202 ^ x96 ;
  assign n375 = ( n371 & ~n372 ) | ( n371 & n374 ) | ( ~n372 & n374 ) ;
  assign n376 = n375 ^ x82 ^ x13 ;
  assign n377 = n141 | n376 ;
  assign n378 = n191 | n377 ;
  assign n379 = ( ~x72 & n164 ) | ( ~x72 & n378 ) | ( n164 & n378 ) ;
  assign n380 = n208 ^ x66 ^ x41 ;
  assign n381 = ~x76 & n380 ;
  assign n382 = x118 & n151 ;
  assign n383 = n382 ^ x111 ^ 1'b0 ;
  assign n384 = n151 & n241 ;
  assign n385 = n256 | n384 ;
  assign n386 = n385 ^ n213 ^ 1'b0 ;
  assign n390 = n139 | n333 ;
  assign n391 = n390 ^ n364 ^ 1'b0 ;
  assign n392 = ~n369 & n391 ;
  assign n387 = x6 & ~n158 ;
  assign n388 = n315 & n387 ;
  assign n389 = n224 | n388 ;
  assign n393 = n392 ^ n389 ^ 1'b0 ;
  assign n394 = ~n139 & n393 ;
  assign n395 = x46 & x102 ;
  assign n396 = n395 ^ x14 ^ 1'b0 ;
  assign n397 = n188 ^ x75 ^ 1'b0 ;
  assign n398 = ~n396 & n397 ;
  assign n399 = n398 ^ x2 ^ 1'b0 ;
  assign n400 = x0 & x52 ;
  assign n401 = ~n136 & n400 ;
  assign n402 = x4 & n401 ;
  assign n403 = n402 ^ x71 ^ 1'b0 ;
  assign n405 = x85 ^ x62 ^ x49 ;
  assign n404 = n153 ^ x108 ^ x25 ;
  assign n406 = n405 ^ n404 ^ n169 ;
  assign n419 = ( ~x32 & x80 ) | ( ~x32 & n199 ) | ( x80 & n199 ) ;
  assign n417 = x67 & x87 ;
  assign n418 = n417 ^ x64 ^ 1'b0 ;
  assign n407 = n213 ^ n207 ^ 1'b0 ;
  assign n408 = n333 & ~n407 ;
  assign n409 = n280 ^ n221 ^ x25 ;
  assign n410 = x42 & n409 ;
  assign n411 = n410 ^ n214 ^ 1'b0 ;
  assign n412 = n144 | n266 ;
  assign n413 = ( n228 & ~n357 ) | ( n228 & n412 ) | ( ~n357 & n412 ) ;
  assign n414 = n411 | n413 ;
  assign n415 = n408 | n414 ;
  assign n416 = n415 ^ x112 ^ 1'b0 ;
  assign n420 = n419 ^ n418 ^ n416 ;
  assign n421 = n218 ^ n180 ^ 1'b0 ;
  assign n442 = n143 & n314 ;
  assign n427 = n245 ^ x35 ^ 1'b0 ;
  assign n428 = x60 & ~n427 ;
  assign n429 = n211 & n428 ;
  assign n430 = n265 ^ x8 ^ 1'b0 ;
  assign n431 = n171 | n430 ;
  assign n436 = x123 | n431 ;
  assign n435 = ~x18 & n337 ;
  assign n437 = n436 ^ n435 ^ 1'b0 ;
  assign n438 = x0 & x91 ;
  assign n439 = n437 & n438 ;
  assign n432 = ( x7 & ~x18 ) | ( x7 & n431 ) | ( ~x18 & n431 ) ;
  assign n433 = x36 & ~n432 ;
  assign n434 = n401 & n433 ;
  assign n440 = n439 ^ n434 ^ 1'b0 ;
  assign n441 = ~n429 & n440 ;
  assign n443 = n442 ^ n441 ^ x59 ;
  assign n425 = n226 ^ x50 ^ x23 ;
  assign n423 = x69 ^ x47 ^ 1'b0 ;
  assign n424 = x43 & n423 ;
  assign n422 = n346 ^ x100 ^ 1'b0 ;
  assign n426 = n425 ^ n424 ^ n422 ;
  assign n444 = n443 ^ n426 ^ 1'b0 ;
  assign n445 = x8 & ~n444 ;
  assign n446 = x78 & ~n207 ;
  assign n447 = ~x125 & n446 ;
  assign n448 = n447 ^ x74 ^ 1'b0 ;
  assign n449 = ( n161 & ~n384 ) | ( n161 & n442 ) | ( ~n384 & n442 ) ;
  assign n450 = ~n165 & n236 ;
  assign n451 = n450 ^ n325 ^ 1'b0 ;
  assign n452 = ~n170 & n451 ;
  assign n453 = n388 | n452 ;
  assign n454 = n453 ^ n245 ^ 1'b0 ;
  assign n455 = n454 ^ x48 ^ x37 ;
  assign n456 = ~n144 & n184 ;
  assign n457 = n401 ^ n380 ^ 1'b0 ;
  assign n458 = n457 ^ n202 ^ 1'b0 ;
  assign n460 = x43 ^ x42 ^ x36 ;
  assign n459 = x64 & n167 ;
  assign n461 = n460 ^ n459 ^ 1'b0 ;
  assign n462 = n162 | n461 ;
  assign n463 = n364 ^ x37 ^ 1'b0 ;
  assign n464 = x97 & n463 ;
  assign n465 = x78 ^ x69 ^ x44 ;
  assign n466 = n465 ^ n149 ^ x96 ;
  assign n467 = n466 ^ n192 ^ x51 ;
  assign n468 = n358 & ~n467 ;
  assign n469 = n405 ^ n224 ^ n186 ;
  assign n470 = ( n143 & n468 ) | ( n143 & n469 ) | ( n468 & n469 ) ;
  assign n471 = ~x71 & n364 ;
  assign n473 = n173 ^ x79 ^ x10 ;
  assign n472 = ( x103 & ~n129 ) | ( x103 & n176 ) | ( ~n129 & n176 ) ;
  assign n474 = n473 ^ n472 ^ 1'b0 ;
  assign n475 = ~n471 & n474 ;
  assign n476 = ~n167 & n475 ;
  assign n477 = n224 ^ n137 ^ x87 ;
  assign n478 = n477 ^ n227 ^ x36 ;
  assign n479 = n422 ^ n413 ^ n375 ;
  assign n480 = x106 ^ x92 ^ 1'b0 ;
  assign n481 = x111 & n480 ;
  assign n482 = n481 ^ n350 ^ 1'b0 ;
  assign n483 = ( ~n197 & n224 ) | ( ~n197 & n293 ) | ( n224 & n293 ) ;
  assign n484 = n134 ^ x66 ^ 1'b0 ;
  assign n485 = n483 | n484 ;
  assign n488 = ( x99 & n129 ) | ( x99 & ~n236 ) | ( n129 & ~n236 ) ;
  assign n489 = n404 ^ n245 ^ 1'b0 ;
  assign n490 = n488 & ~n489 ;
  assign n486 = ( x15 & ~x36 ) | ( x15 & x105 ) | ( ~x36 & x105 ) ;
  assign n487 = ~n149 & n486 ;
  assign n491 = n490 ^ n487 ^ n349 ;
  assign n492 = ( n467 & ~n485 ) | ( n467 & n491 ) | ( ~n485 & n491 ) ;
  assign n493 = n325 ^ x47 ^ 1'b0 ;
  assign n494 = n270 & ~n493 ;
  assign n495 = n494 ^ n383 ^ 1'b0 ;
  assign n496 = n332 & n495 ;
  assign n497 = n496 ^ n357 ^ 1'b0 ;
  assign n498 = n497 ^ n257 ^ x43 ;
  assign n499 = n498 ^ x101 ^ 1'b0 ;
  assign n500 = x34 & ~n499 ;
  assign n501 = n315 ^ x88 ^ x66 ;
  assign n502 = n501 ^ n137 ^ x120 ;
  assign n503 = x112 ^ x92 ^ 1'b0 ;
  assign n504 = x94 & n503 ;
  assign n505 = ( n192 & ~n325 ) | ( n192 & n504 ) | ( ~n325 & n504 ) ;
  assign n506 = n339 ^ n236 ^ x97 ;
  assign n507 = x58 & n304 ;
  assign n508 = n507 ^ n371 ^ 1'b0 ;
  assign n509 = ( ~n245 & n365 ) | ( ~n245 & n508 ) | ( n365 & n508 ) ;
  assign n510 = ~n327 & n374 ;
  assign n511 = ~n219 & n510 ;
  assign n512 = x118 | n511 ;
  assign n519 = ( ~x13 & n236 ) | ( ~x13 & n367 ) | ( n236 & n367 ) ;
  assign n515 = x44 & x87 ;
  assign n516 = ~x118 & n515 ;
  assign n513 = x78 & ~n194 ;
  assign n514 = ~x73 & n513 ;
  assign n517 = n516 ^ n514 ^ n321 ;
  assign n518 = x114 & ~n517 ;
  assign n520 = n519 ^ n518 ^ 1'b0 ;
  assign n521 = x35 & n147 ;
  assign n522 = ~x62 & n521 ;
  assign n523 = n290 ^ x102 ^ x45 ;
  assign n524 = n522 | n523 ;
  assign n525 = n524 ^ x59 ^ 1'b0 ;
  assign n526 = n525 ^ n442 ^ 1'b0 ;
  assign n527 = ( ~x104 & n137 ) | ( ~x104 & n226 ) | ( n137 & n226 ) ;
  assign n528 = n357 & n527 ;
  assign n529 = n137 ^ x64 ^ x63 ;
  assign n530 = x15 & ~n156 ;
  assign n531 = ~x94 & n530 ;
  assign n532 = x28 & ~n531 ;
  assign n533 = ~x122 & n532 ;
  assign n534 = n529 | n533 ;
  assign n535 = n534 ^ n267 ^ 1'b0 ;
  assign n536 = n157 & n535 ;
  assign n537 = n536 ^ n434 ^ 1'b0 ;
  assign n538 = ( x17 & ~x25 ) | ( x17 & x127 ) | ( ~x25 & x127 ) ;
  assign n539 = n538 ^ x107 ^ x29 ;
  assign n540 = ( ~x42 & n149 ) | ( ~x42 & n457 ) | ( n149 & n457 ) ;
  assign n541 = n328 & ~n540 ;
  assign n542 = x41 & ~n218 ;
  assign n543 = ~n541 & n542 ;
  assign n544 = x120 ^ x66 ^ x21 ;
  assign n545 = ( x56 & x107 ) | ( x56 & n544 ) | ( x107 & n544 ) ;
  assign n546 = n167 & ~n425 ;
  assign n547 = ~x43 & n546 ;
  assign n548 = ( ~x3 & x126 ) | ( ~x3 & n547 ) | ( x126 & n547 ) ;
  assign n549 = n548 ^ n404 ^ n151 ;
  assign n550 = x34 & ~n188 ;
  assign n551 = n550 ^ x80 ^ 1'b0 ;
  assign n552 = n272 ^ x84 ^ 1'b0 ;
  assign n553 = n232 | n533 ;
  assign n554 = n162 & ~n553 ;
  assign n555 = ( x99 & n552 ) | ( x99 & ~n554 ) | ( n552 & ~n554 ) ;
  assign n556 = n283 & n555 ;
  assign n557 = n516 ^ n363 ^ x53 ;
  assign n558 = n287 & n526 ;
  assign n559 = ( ~x96 & n557 ) | ( ~x96 & n558 ) | ( n557 & n558 ) ;
  assign n564 = x17 & ~n437 ;
  assign n565 = ~n335 & n564 ;
  assign n560 = x115 & n294 ;
  assign n561 = x106 & ~n560 ;
  assign n562 = n493 & n561 ;
  assign n563 = ~n196 & n562 ;
  assign n566 = n565 ^ n563 ^ x92 ;
  assign n567 = x6 | n210 ;
  assign n568 = n224 | n567 ;
  assign n569 = n568 ^ n432 ^ 1'b0 ;
  assign n570 = n498 ^ n447 ^ x51 ;
  assign n574 = x50 | n208 ;
  assign n571 = x108 ^ x13 ^ 1'b0 ;
  assign n572 = ( x53 & n170 ) | ( x53 & ~n571 ) | ( n170 & ~n571 ) ;
  assign n573 = x22 & ~n572 ;
  assign n575 = n574 ^ n573 ^ x29 ;
  assign n576 = x30 & ~x125 ;
  assign n577 = ( x16 & n224 ) | ( x16 & n251 ) | ( n224 & n251 ) ;
  assign n578 = n576 | n577 ;
  assign n579 = n552 & ~n578 ;
  assign n580 = x49 & n257 ;
  assign n581 = n580 ^ x36 ^ 1'b0 ;
  assign n582 = ~n563 & n581 ;
  assign n583 = n582 ^ x51 ^ 1'b0 ;
  assign n584 = ( n575 & n579 ) | ( n575 & ~n583 ) | ( n579 & ~n583 ) ;
  assign n585 = x35 & x74 ;
  assign n586 = ~x31 & n585 ;
  assign n587 = n157 & ~n586 ;
  assign n588 = n587 ^ n460 ^ 1'b0 ;
  assign n589 = n361 ^ x122 ^ x48 ;
  assign n590 = ( n236 & n514 ) | ( n236 & n589 ) | ( n514 & n589 ) ;
  assign n591 = x91 & n590 ;
  assign n592 = n228 & n591 ;
  assign n593 = n455 & ~n592 ;
  assign n594 = n593 ^ n358 ^ 1'b0 ;
  assign n595 = x37 & ~x54 ;
  assign n596 = ~n293 & n595 ;
  assign n597 = n565 ^ n424 ^ n269 ;
  assign n598 = n436 & n597 ;
  assign n599 = n596 & n598 ;
  assign n603 = n307 & ~n495 ;
  assign n600 = ~n432 & n488 ;
  assign n601 = n318 & n600 ;
  assign n602 = x22 & ~n601 ;
  assign n604 = n603 ^ n602 ^ 1'b0 ;
  assign n605 = n294 ^ n173 ^ x81 ;
  assign n606 = n550 ^ n299 ^ 1'b0 ;
  assign n607 = n267 & ~n606 ;
  assign n608 = ( x49 & ~n605 ) | ( x49 & n607 ) | ( ~n605 & n607 ) ;
  assign n609 = x125 & ~n156 ;
  assign n610 = ~n608 & n609 ;
  assign n611 = n199 ^ x23 ^ 1'b0 ;
  assign n612 = ( n218 & n374 ) | ( n218 & n425 ) | ( n374 & n425 ) ;
  assign n613 = n612 ^ n575 ^ n522 ;
  assign n614 = n327 | n613 ;
  assign n615 = n614 ^ n200 ^ 1'b0 ;
  assign n616 = n615 ^ n584 ^ 1'b0 ;
  assign n617 = n611 & n616 ;
  assign n622 = x46 & x88 ;
  assign n623 = n622 ^ x25 ^ 1'b0 ;
  assign n624 = n623 ^ n571 ^ n409 ;
  assign n625 = n452 | n624 ;
  assign n618 = n412 ^ n294 ^ 1'b0 ;
  assign n619 = ( n352 & n406 ) | ( n352 & n618 ) | ( n406 & n618 ) ;
  assign n620 = n525 & ~n527 ;
  assign n621 = n619 & n620 ;
  assign n626 = n625 ^ n621 ^ 1'b0 ;
  assign n627 = ~n516 & n522 ;
  assign n628 = n437 ^ n224 ^ x28 ;
  assign n629 = ( x53 & n540 ) | ( x53 & ~n628 ) | ( n540 & ~n628 ) ;
  assign n630 = ~n627 & n629 ;
  assign n631 = ~n337 & n630 ;
  assign n636 = ( x14 & ~x101 ) | ( x14 & n136 ) | ( ~x101 & n136 ) ;
  assign n632 = ( x10 & ~x61 ) | ( x10 & n170 ) | ( ~x61 & n170 ) ;
  assign n633 = n632 ^ n574 ^ n296 ;
  assign n634 = n633 ^ x37 ^ 1'b0 ;
  assign n635 = x0 & n634 ;
  assign n637 = n636 ^ n635 ^ 1'b0 ;
  assign n638 = n209 & ~n241 ;
  assign n639 = n638 ^ x37 ^ 1'b0 ;
  assign n640 = x87 & n222 ;
  assign n641 = ~n242 & n640 ;
  assign n642 = x83 & ~n641 ;
  assign n643 = n642 ^ n505 ^ 1'b0 ;
  assign n644 = n643 ^ n613 ^ 1'b0 ;
  assign n645 = n160 ^ x37 ^ 1'b0 ;
  assign n646 = x78 & ~n645 ;
  assign n647 = n646 ^ n206 ^ 1'b0 ;
  assign n648 = n136 & n647 ;
  assign n649 = n648 ^ n481 ^ 1'b0 ;
  assign n650 = x122 | n649 ;
  assign n652 = n576 ^ n396 ^ n283 ;
  assign n653 = ~n241 & n652 ;
  assign n654 = n653 ^ n178 ^ 1'b0 ;
  assign n651 = n146 & n226 ;
  assign n655 = n654 ^ n651 ^ 1'b0 ;
  assign n656 = x81 & n655 ;
  assign n657 = n560 ^ n301 ^ 1'b0 ;
  assign n658 = n657 ^ n192 ^ x90 ;
  assign n659 = n429 ^ x127 ^ 1'b0 ;
  assign n660 = n170 ^ x102 ^ 1'b0 ;
  assign n661 = ~n269 & n660 ;
  assign n662 = n431 ^ n290 ^ 1'b0 ;
  assign n663 = ( n659 & n661 ) | ( n659 & n662 ) | ( n661 & n662 ) ;
  assign n664 = n658 | n663 ;
  assign n665 = n396 ^ x91 ^ 1'b0 ;
  assign n666 = n464 & ~n665 ;
  assign n667 = x77 & ~n168 ;
  assign n675 = ( x40 & ~n237 ) | ( x40 & n514 ) | ( ~n237 & n514 ) ;
  assign n668 = n611 ^ x111 ^ x110 ;
  assign n669 = n233 ^ n192 ^ x113 ;
  assign n670 = n669 ^ n360 ^ x62 ;
  assign n671 = n670 ^ x122 ^ 1'b0 ;
  assign n672 = n302 & n671 ;
  assign n673 = ( n432 & n668 ) | ( n432 & n672 ) | ( n668 & n672 ) ;
  assign n674 = n633 & ~n673 ;
  assign n676 = n675 ^ n674 ^ 1'b0 ;
  assign n677 = x43 & ~n274 ;
  assign n678 = n522 & n677 ;
  assign n679 = ( x80 & ~n466 ) | ( x80 & n678 ) | ( ~n466 & n678 ) ;
  assign n680 = ( n256 & n401 ) | ( n256 & n679 ) | ( n401 & n679 ) ;
  assign n681 = ( ~n370 & n415 ) | ( ~n370 & n473 ) | ( n415 & n473 ) ;
  assign n682 = x81 & ~n681 ;
  assign n683 = ~x88 & n682 ;
  assign n684 = n526 ^ x95 ^ 1'b0 ;
  assign n685 = n683 | n684 ;
  assign n686 = n331 ^ n214 ^ 1'b0 ;
  assign n687 = x64 & ~n686 ;
  assign n688 = n159 ^ x71 ^ 1'b0 ;
  assign n689 = x59 & n688 ;
  assign n690 = n689 ^ n222 ^ 1'b0 ;
  assign n691 = n687 & n690 ;
  assign n692 = ( ~x69 & x73 ) | ( ~x69 & n457 ) | ( x73 & n457 ) ;
  assign n693 = n437 ^ n320 ^ n224 ;
  assign n694 = ( x13 & n373 ) | ( x13 & n693 ) | ( n373 & n693 ) ;
  assign n695 = n692 | n694 ;
  assign n696 = ( ~x108 & x110 ) | ( ~x108 & n237 ) | ( x110 & n237 ) ;
  assign n697 = x59 & ~n696 ;
  assign n698 = n447 ^ n304 ^ 1'b0 ;
  assign n699 = n697 & ~n698 ;
  assign n700 = n245 | n422 ;
  assign n701 = n700 ^ n380 ^ 1'b0 ;
  assign n702 = x127 & n390 ;
  assign n703 = n702 ^ n298 ^ 1'b0 ;
  assign n704 = n703 ^ n421 ^ x67 ;
  assign n705 = n361 ^ n248 ^ 1'b0 ;
  assign n706 = x72 & n705 ;
  assign n707 = n706 ^ n514 ^ 1'b0 ;
  assign n708 = ~n173 & n707 ;
  assign n711 = n222 ^ n206 ^ 1'b0 ;
  assign n712 = n134 | n711 ;
  assign n709 = ~n376 & n378 ;
  assign n710 = n253 & n709 ;
  assign n713 = n712 ^ n710 ^ 1'b0 ;
  assign n714 = n544 ^ n134 ^ 1'b0 ;
  assign n715 = n714 ^ n434 ^ n357 ;
  assign n716 = n654 ^ n233 ^ 1'b0 ;
  assign n717 = ~n200 & n716 ;
  assign n718 = n612 ^ n428 ^ 1'b0 ;
  assign n719 = n131 & ~n718 ;
  assign n720 = n717 & n719 ;
  assign n721 = n720 ^ n299 ^ 1'b0 ;
  assign n722 = ( x8 & x30 ) | ( x8 & ~n672 ) | ( x30 & ~n672 ) ;
  assign n725 = n218 ^ x62 ^ x16 ;
  assign n726 = n488 & n725 ;
  assign n727 = ~x51 & n726 ;
  assign n723 = x31 | n346 ;
  assign n724 = n723 ^ n603 ^ x77 ;
  assign n728 = n727 ^ n724 ^ n379 ;
  assign n729 = n131 & ~n248 ;
  assign n730 = n729 ^ x103 ^ 1'b0 ;
  assign n731 = x96 & ~n224 ;
  assign n732 = ~x6 & n731 ;
  assign n733 = n730 | n732 ;
  assign n734 = ( x115 & n623 ) | ( x115 & ~n733 ) | ( n623 & ~n733 ) ;
  assign n735 = x124 & n694 ;
  assign n736 = ~n734 & n735 ;
  assign n737 = n663 ^ n368 ^ n250 ;
  assign n741 = x59 & ~n264 ;
  assign n742 = ~n191 & n741 ;
  assign n743 = n742 ^ n230 ^ x99 ;
  assign n738 = n446 ^ x41 ^ 1'b0 ;
  assign n739 = n738 ^ n241 ^ n191 ;
  assign n740 = n739 ^ n328 ^ 1'b0 ;
  assign n744 = n743 ^ n740 ^ x46 ;
  assign n745 = n486 ^ n165 ^ 1'b0 ;
  assign n746 = n550 | n745 ;
  assign n747 = ~x16 & x25 ;
  assign n748 = x14 & ~n747 ;
  assign n749 = ~x21 & n748 ;
  assign n750 = n746 | n749 ;
  assign n751 = n744 | n750 ;
  assign n752 = ( x96 & n307 ) | ( x96 & n696 ) | ( n307 & n696 ) ;
  assign n753 = n325 ^ x111 ^ x31 ;
  assign n754 = n207 ^ x37 ^ 1'b0 ;
  assign n755 = ( ~n752 & n753 ) | ( ~n752 & n754 ) | ( n753 & n754 ) ;
  assign n756 = n493 ^ x70 ^ 1'b0 ;
  assign n757 = n756 ^ x11 ^ 1'b0 ;
  assign n758 = ~n550 & n757 ;
  assign n759 = n758 ^ n198 ^ 1'b0 ;
  assign n760 = n722 ^ x70 ^ 1'b0 ;
  assign n761 = ( x32 & x49 ) | ( x32 & n344 ) | ( x49 & n344 ) ;
  assign n764 = n238 ^ x43 ^ 1'b0 ;
  assign n768 = ( ~x29 & x31 ) | ( ~x29 & x50 ) | ( x31 & x50 ) ;
  assign n765 = n164 | n576 ;
  assign n766 = n380 | n765 ;
  assign n767 = x115 & ~n766 ;
  assign n769 = n768 ^ n767 ^ 1'b0 ;
  assign n770 = n764 | n769 ;
  assign n762 = n668 ^ n466 ^ 1'b0 ;
  assign n763 = ~n328 & n762 ;
  assign n771 = n770 ^ n763 ^ x16 ;
  assign n772 = n693 & ~n703 ;
  assign n773 = n772 ^ n425 ^ 1'b0 ;
  assign n774 = n537 ^ x91 ^ 1'b0 ;
  assign n775 = ( x77 & n742 ) | ( x77 & n774 ) | ( n742 & n774 ) ;
  assign n776 = n516 ^ n315 ^ n269 ;
  assign n777 = n776 ^ x24 ^ x9 ;
  assign n778 = n500 ^ n366 ^ 1'b0 ;
  assign n779 = n777 & ~n778 ;
  assign n799 = n383 | n471 ;
  assign n800 = n264 & ~n799 ;
  assign n801 = n335 & ~n800 ;
  assign n802 = ~x14 & n801 ;
  assign n798 = n365 & n371 ;
  assign n794 = n227 & n277 ;
  assign n795 = n204 & ~n529 ;
  assign n796 = ~n794 & n795 ;
  assign n788 = n383 ^ x29 ^ 1'b0 ;
  assign n789 = x26 & ~n788 ;
  assign n790 = x96 & n789 ;
  assign n791 = n790 ^ x108 ^ 1'b0 ;
  assign n780 = n158 | n373 ;
  assign n781 = n780 ^ n537 ^ 1'b0 ;
  assign n782 = n304 & n633 ;
  assign n783 = n782 ^ n408 ^ 1'b0 ;
  assign n784 = n783 ^ n367 ^ 1'b0 ;
  assign n785 = n784 ^ n732 ^ 1'b0 ;
  assign n786 = n781 & ~n785 ;
  assign n787 = n786 ^ n214 ^ 1'b0 ;
  assign n792 = n791 ^ n787 ^ 1'b0 ;
  assign n793 = n357 & ~n792 ;
  assign n797 = n796 ^ n793 ^ n544 ;
  assign n803 = n802 ^ n798 ^ n797 ;
  assign n804 = n328 | n724 ;
  assign n805 = ~n208 & n298 ;
  assign n806 = n805 ^ n449 ^ 1'b0 ;
  assign n807 = ( x68 & ~n550 ) | ( x68 & n806 ) | ( ~n550 & n806 ) ;
  assign n808 = n208 | n415 ;
  assign n809 = x56 & n608 ;
  assign n810 = n637 ^ n559 ^ 1'b0 ;
  assign n811 = n576 ^ n242 ^ 1'b0 ;
  assign n812 = n810 | n811 ;
  assign n813 = n204 | n256 ;
  assign n814 = x23 & n143 ;
  assign n815 = n814 ^ n224 ^ 1'b0 ;
  assign n816 = x53 & n492 ;
  assign n817 = n548 & n816 ;
  assign n818 = n817 ^ x20 ^ 1'b0 ;
  assign n819 = n380 & ~n818 ;
  assign n820 = ( n813 & ~n815 ) | ( n813 & n819 ) | ( ~n815 & n819 ) ;
  assign n821 = ( n555 & n756 ) | ( n555 & ~n820 ) | ( n756 & ~n820 ) ;
  assign n822 = n221 ^ x88 ^ 1'b0 ;
  assign n823 = x124 & n822 ;
  assign n824 = n823 ^ n159 ^ 1'b0 ;
  assign n825 = x87 & ~n824 ;
  assign n826 = ~n149 & n825 ;
  assign n829 = n369 ^ n149 ^ x107 ;
  assign n830 = ( n253 & ~n327 ) | ( n253 & n829 ) | ( ~n327 & n829 ) ;
  assign n827 = n147 ^ x74 ^ 1'b0 ;
  assign n828 = n401 | n827 ;
  assign n831 = n830 ^ n828 ^ 1'b0 ;
  assign n832 = n680 | n831 ;
  assign n833 = n832 ^ x19 ^ 1'b0 ;
  assign n846 = n147 ^ x8 ^ 1'b0 ;
  assign n845 = ( ~x66 & n269 ) | ( ~x66 & n368 ) | ( n269 & n368 ) ;
  assign n834 = n611 ^ n256 ^ x61 ;
  assign n837 = ( x12 & ~n339 ) | ( x12 & n439 ) | ( ~n339 & n439 ) ;
  assign n835 = n687 ^ n266 ^ x69 ;
  assign n836 = x91 & ~n835 ;
  assign n838 = n837 ^ n836 ^ 1'b0 ;
  assign n839 = x55 & n632 ;
  assign n840 = n839 ^ x4 ^ 1'b0 ;
  assign n841 = n756 ^ x104 ^ x41 ;
  assign n842 = n840 & ~n841 ;
  assign n843 = n838 & n842 ;
  assign n844 = ~n834 & n843 ;
  assign n847 = n846 ^ n845 ^ n844 ;
  assign n848 = ( n170 & n283 ) | ( n170 & ~n354 ) | ( n283 & ~n354 ) ;
  assign n849 = n848 ^ n586 ^ 1'b0 ;
  assign n850 = n422 | n849 ;
  assign n851 = ( x71 & ~n165 ) | ( x71 & n224 ) | ( ~n165 & n224 ) ;
  assign n852 = n851 ^ n562 ^ n531 ;
  assign n853 = n383 | n743 ;
  assign n854 = n853 ^ n426 ^ 1'b0 ;
  assign n855 = n852 & ~n854 ;
  assign n856 = x92 | n855 ;
  assign n860 = n306 & n378 ;
  assign n861 = n860 ^ n339 ^ 1'b0 ;
  assign n862 = ( x22 & n415 ) | ( x22 & n861 ) | ( n415 & n861 ) ;
  assign n867 = n451 ^ n129 ^ x53 ;
  assign n868 = n538 ^ n173 ^ 1'b0 ;
  assign n869 = ~n867 & n868 ;
  assign n863 = n791 ^ n257 ^ 1'b0 ;
  assign n864 = x98 & x107 ;
  assign n865 = n864 ^ n260 ^ 1'b0 ;
  assign n866 = ( ~n236 & n863 ) | ( ~n236 & n865 ) | ( n863 & n865 ) ;
  assign n870 = n869 ^ n866 ^ n143 ;
  assign n871 = ( n763 & n862 ) | ( n763 & n870 ) | ( n862 & n870 ) ;
  assign n858 = ( x12 & x15 ) | ( x12 & ~x89 ) | ( x15 & ~x89 ) ;
  assign n859 = n858 ^ n692 ^ x72 ;
  assign n857 = ( ~x123 & n332 ) | ( ~x123 & n411 ) | ( n332 & n411 ) ;
  assign n872 = n871 ^ n859 ^ n857 ;
  assign n873 = ~n171 & n392 ;
  assign n874 = n416 ^ x88 ^ x32 ;
  assign n875 = ( x39 & n555 ) | ( x39 & n874 ) | ( n555 & n874 ) ;
  assign n876 = n525 & ~n612 ;
  assign n877 = n876 ^ n344 ^ 1'b0 ;
  assign n878 = n200 ^ x109 ^ 1'b0 ;
  assign n882 = x34 & x118 ;
  assign n883 = n882 ^ n259 ^ 1'b0 ;
  assign n879 = n159 & ~n198 ;
  assign n880 = ~n813 & n879 ;
  assign n881 = ( n301 & ~n522 ) | ( n301 & n880 ) | ( ~n522 & n880 ) ;
  assign n884 = n883 ^ n881 ^ n241 ;
  assign n885 = n479 & n527 ;
  assign n886 = n571 ^ x74 ^ 1'b0 ;
  assign n887 = x60 & n886 ;
  assign n888 = n887 ^ n176 ^ 1'b0 ;
  assign n889 = ( n884 & n885 ) | ( n884 & ~n888 ) | ( n885 & ~n888 ) ;
  assign n890 = n479 ^ n467 ^ 1'b0 ;
  assign n891 = ( ~n487 & n798 ) | ( ~n487 & n890 ) | ( n798 & n890 ) ;
  assign n892 = n327 | n431 ;
  assign n893 = n892 ^ n766 ^ 1'b0 ;
  assign n894 = ( ~n318 & n458 ) | ( ~n318 & n893 ) | ( n458 & n893 ) ;
  assign n895 = n442 ^ n321 ^ 1'b0 ;
  assign n896 = n280 | n383 ;
  assign n897 = n896 ^ x92 ^ 1'b0 ;
  assign n898 = n538 & ~n897 ;
  assign n899 = n487 ^ x38 ^ x24 ;
  assign n900 = x77 & ~n899 ;
  assign n901 = n160 & n900 ;
  assign n902 = x115 | n901 ;
  assign n903 = n902 ^ n845 ^ 1'b0 ;
  assign n904 = n786 ^ n327 ^ 1'b0 ;
  assign n905 = n375 & ~n904 ;
  assign n906 = n635 & ~n833 ;
  assign n910 = x16 & ~n171 ;
  assign n911 = n910 ^ x54 ^ 1'b0 ;
  assign n907 = x52 & ~n516 ;
  assign n908 = n907 ^ n158 ^ 1'b0 ;
  assign n909 = n571 & n908 ;
  assign n912 = n911 ^ n909 ^ 1'b0 ;
  assign n914 = n245 ^ x38 ^ 1'b0 ;
  assign n913 = ~n186 & n763 ;
  assign n915 = n914 ^ n913 ^ 1'b0 ;
  assign n916 = n393 ^ n318 ^ 1'b0 ;
  assign n917 = n211 ^ x93 ^ 1'b0 ;
  assign n918 = n371 ^ x102 ^ 1'b0 ;
  assign n919 = x5 & n918 ;
  assign n920 = n919 ^ n164 ^ x32 ;
  assign n921 = n920 ^ n338 ^ 1'b0 ;
  assign n922 = n422 ^ x48 ^ 1'b0 ;
  assign n923 = x92 & ~n922 ;
  assign n924 = ( x59 & n250 ) | ( x59 & ~n325 ) | ( n250 & ~n325 ) ;
  assign n925 = n924 ^ n319 ^ 1'b0 ;
  assign n926 = ( ~n921 & n923 ) | ( ~n921 & n925 ) | ( n923 & n925 ) ;
  assign n927 = n906 ^ n781 ^ n338 ;
  assign n928 = ( x44 & x97 ) | ( x44 & ~x125 ) | ( x97 & ~x125 ) ;
  assign n929 = n928 ^ x5 ^ 1'b0 ;
  assign n930 = x100 & n929 ;
  assign n931 = n930 ^ n209 ^ 1'b0 ;
  assign n932 = x15 & n931 ;
  assign n933 = n467 ^ x0 ^ 1'b0 ;
  assign n934 = n933 ^ x84 ^ 1'b0 ;
  assign n935 = n378 | n934 ;
  assign n936 = n675 ^ n281 ^ 1'b0 ;
  assign n937 = n464 & n936 ;
  assign n938 = n298 & ~n672 ;
  assign n939 = ~n560 & n938 ;
  assign n940 = n830 & n939 ;
  assign n941 = x64 & n408 ;
  assign n942 = n234 & n941 ;
  assign n943 = ( x26 & x30 ) | ( x26 & ~n625 ) | ( x30 & ~n625 ) ;
  assign n944 = x16 & ~n237 ;
  assign n945 = n944 ^ n158 ^ 1'b0 ;
  assign n946 = ( ~x17 & n401 ) | ( ~x17 & n945 ) | ( n401 & n945 ) ;
  assign n947 = n820 & ~n946 ;
  assign n948 = n289 & ~n764 ;
  assign n949 = ( x84 & x86 ) | ( x84 & n280 ) | ( x86 & n280 ) ;
  assign n950 = x110 & n949 ;
  assign n951 = ~n390 & n950 ;
  assign n952 = ( ~n325 & n383 ) | ( ~n325 & n451 ) | ( n383 & n451 ) ;
  assign n953 = n428 ^ n357 ^ 1'b0 ;
  assign n954 = n952 & n953 ;
  assign n955 = ( ~n352 & n951 ) | ( ~n352 & n954 ) | ( n951 & n954 ) ;
  assign n956 = ( n245 & n392 ) | ( n245 & n575 ) | ( n392 & n575 ) ;
  assign n957 = n481 & n956 ;
  assign n958 = n957 ^ x95 ^ 1'b0 ;
  assign n962 = n216 & n298 ;
  assign n963 = n194 & n962 ;
  assign n964 = ( n204 & n422 ) | ( n204 & n963 ) | ( n422 & n963 ) ;
  assign n959 = n243 | n601 ;
  assign n960 = n328 & ~n959 ;
  assign n961 = ~n162 & n960 ;
  assign n965 = n964 ^ n961 ^ n538 ;
  assign n966 = x126 & ~n791 ;
  assign n967 = n966 ^ n583 ^ 1'b0 ;
  assign n971 = n919 ^ n598 ^ 1'b0 ;
  assign n972 = n625 | n971 ;
  assign n968 = ( ~x55 & n161 ) | ( ~x55 & n743 ) | ( n161 & n743 ) ;
  assign n969 = ( ~x117 & n624 ) | ( ~x117 & n968 ) | ( n624 & n968 ) ;
  assign n970 = ( ~n529 & n727 ) | ( ~n529 & n969 ) | ( n727 & n969 ) ;
  assign n973 = n972 ^ n970 ^ x18 ;
  assign n974 = ~n620 & n646 ;
  assign n975 = ~n296 & n768 ;
  assign n976 = ~x3 & n975 ;
  assign n977 = n976 ^ n659 ^ 1'b0 ;
  assign n978 = n659 ^ n363 ^ 1'b0 ;
  assign n979 = n199 & n978 ;
  assign n980 = n730 ^ n366 ^ 1'b0 ;
  assign n981 = n979 & n980 ;
  assign n982 = n905 ^ n293 ^ x80 ;
  assign n983 = n982 ^ n808 ^ 1'b0 ;
  assign n984 = n473 ^ n224 ^ n182 ;
  assign n985 = n869 & n984 ;
  assign n986 = n985 ^ n980 ^ n283 ;
  assign n987 = ~n658 & n842 ;
  assign n988 = n605 ^ x31 ^ 1'b0 ;
  assign n989 = x6 & n988 ;
  assign n990 = ( ~x35 & x109 ) | ( ~x35 & n989 ) | ( x109 & n989 ) ;
  assign n991 = n584 ^ n413 ^ n348 ;
  assign n992 = n970 ^ n954 ^ n871 ;
  assign n993 = n615 ^ n472 ^ 1'b0 ;
  assign n994 = x99 & n274 ;
  assign n995 = n821 & ~n994 ;
  assign n996 = n346 & n995 ;
  assign n997 = ( n366 & ~n588 ) | ( n366 & n996 ) | ( ~n588 & n996 ) ;
  assign n998 = n784 & ~n997 ;
  assign n999 = ( n164 & ~n724 ) | ( n164 & n768 ) | ( ~n724 & n768 ) ;
  assign n1000 = ( ~n191 & n664 ) | ( ~n191 & n973 ) | ( n664 & n973 ) ;
  assign n1001 = n893 ^ n405 ^ n169 ;
  assign n1002 = n672 & n1001 ;
  assign n1003 = ( ~x115 & n139 ) | ( ~x115 & n368 ) | ( n139 & n368 ) ;
  assign n1004 = ( x92 & n327 ) | ( x92 & n350 ) | ( n327 & n350 ) ;
  assign n1005 = n923 & n1004 ;
  assign n1006 = n1005 ^ n691 ^ 1'b0 ;
  assign n1007 = n1003 | n1006 ;
  assign n1008 = ~n347 & n768 ;
  assign n1009 = n1008 ^ n703 ^ 1'b0 ;
  assign n1010 = n191 & n1009 ;
  assign n1011 = ~x42 & n1010 ;
  assign n1012 = n1011 ^ n908 ^ 1'b0 ;
  assign n1013 = n1007 | n1012 ;
  assign n1014 = ~n186 & n752 ;
  assign n1015 = n1014 ^ x66 ^ 1'b0 ;
  assign n1016 = n1015 ^ n1001 ^ 1'b0 ;
  assign n1017 = ( ~n171 & n173 ) | ( ~n171 & n257 ) | ( n173 & n257 ) ;
  assign n1018 = x59 & n1017 ;
  assign n1019 = ( x57 & ~x99 ) | ( x57 & n213 ) | ( ~x99 & n213 ) ;
  assign n1020 = x11 & ~n1019 ;
  assign n1021 = x3 & ~n739 ;
  assign n1022 = n1021 ^ n867 ^ 1'b0 ;
  assign n1023 = ( n171 & n985 ) | ( n171 & ~n1022 ) | ( n985 & ~n1022 ) ;
  assign n1024 = ( n945 & n1020 ) | ( n945 & n1023 ) | ( n1020 & n1023 ) ;
  assign n1025 = n1024 ^ n372 ^ n367 ;
  assign n1026 = ~n747 & n1025 ;
  assign n1027 = ~x28 & n1026 ;
  assign n1028 = n1027 ^ n610 ^ n422 ;
  assign n1029 = n509 & n679 ;
  assign n1030 = ~n1028 & n1029 ;
  assign n1031 = n921 ^ n647 ^ 1'b0 ;
  assign n1032 = x102 & ~n1031 ;
  assign n1033 = ( n250 & n869 ) | ( n250 & ~n1032 ) | ( n869 & ~n1032 ) ;
  assign n1034 = n846 ^ n730 ^ n182 ;
  assign n1035 = ~n994 & n1034 ;
  assign n1036 = n783 ^ n540 ^ x27 ;
  assign n1037 = n1036 ^ n830 ^ x11 ;
  assign n1038 = ( ~n250 & n482 ) | ( ~n250 & n1037 ) | ( n482 & n1037 ) ;
  assign n1039 = n316 ^ n269 ^ 1'b0 ;
  assign n1040 = x64 & ~n1039 ;
  assign n1041 = n1040 ^ n747 ^ x114 ;
  assign n1042 = n1041 ^ x19 ^ 1'b0 ;
  assign n1043 = ~n643 & n1042 ;
  assign n1044 = n821 ^ n491 ^ x56 ;
  assign n1045 = x81 & ~n1044 ;
  assign n1046 = n1045 ^ n625 ^ 1'b0 ;
  assign n1047 = x42 & n771 ;
  assign n1048 = ~n766 & n1047 ;
  assign n1049 = n357 & ~n1048 ;
  assign n1050 = n1049 ^ n464 ^ 1'b0 ;
  assign n1051 = n1050 ^ n744 ^ 1'b0 ;
  assign n1052 = ~x49 & n1051 ;
  assign n1053 = n752 ^ n221 ^ 1'b0 ;
  assign n1054 = n791 & n1053 ;
  assign n1055 = n1054 ^ n858 ^ n739 ;
  assign n1056 = n412 ^ n371 ^ 1'b0 ;
  assign n1057 = n1056 ^ n781 ^ n678 ;
  assign n1058 = n348 & ~n1057 ;
  assign n1059 = x55 & ~n490 ;
  assign n1060 = ( x10 & x37 ) | ( x10 & ~x38 ) | ( x37 & ~x38 ) ;
  assign n1061 = n1060 ^ n633 ^ x8 ;
  assign n1062 = n481 | n1061 ;
  assign n1063 = n1062 ^ n241 ^ 1'b0 ;
  assign n1064 = n893 ^ x81 ^ 1'b0 ;
  assign n1065 = x113 & n1064 ;
  assign n1066 = ( x36 & ~n607 ) | ( x36 & n863 ) | ( ~n607 & n863 ) ;
  assign n1067 = n316 ^ n265 ^ x31 ;
  assign n1068 = n1067 ^ n859 ^ 1'b0 ;
  assign n1069 = n1066 & n1068 ;
  assign n1070 = ( n331 & n350 ) | ( n331 & n863 ) | ( n350 & n863 ) ;
  assign n1071 = n1070 ^ n307 ^ x31 ;
  assign n1072 = n392 & ~n1071 ;
  assign n1073 = ( n590 & ~n617 ) | ( n590 & n899 ) | ( ~n617 & n899 ) ;
  assign n1074 = n1073 ^ n149 ^ 1'b0 ;
  assign n1075 = ~x93 & n1074 ;
  assign n1076 = n911 ^ n253 ^ n187 ;
  assign n1077 = n287 ^ n285 ^ n200 ;
  assign n1078 = n646 ^ x83 ^ 1'b0 ;
  assign n1079 = n1078 ^ n618 ^ n486 ;
  assign n1080 = ( n734 & ~n1077 ) | ( n734 & n1079 ) | ( ~n1077 & n1079 ) ;
  assign n1081 = n383 | n468 ;
  assign n1082 = x38 | n1081 ;
  assign n1083 = n165 | n1082 ;
  assign n1084 = x95 & ~n663 ;
  assign n1085 = x8 & n408 ;
  assign n1086 = n1085 ^ x20 ^ 1'b0 ;
  assign n1087 = n1086 ^ n210 ^ 1'b0 ;
  assign n1088 = n672 ^ n668 ^ n238 ;
  assign n1089 = n921 ^ n168 ^ x54 ;
  assign n1090 = ( n932 & n1088 ) | ( n932 & ~n1089 ) | ( n1088 & ~n1089 ) ;
  assign n1091 = x9 & x108 ;
  assign n1092 = ~x36 & n1091 ;
  assign n1093 = n1092 ^ n643 ^ 1'b0 ;
  assign n1094 = ~n1090 & n1093 ;
  assign n1095 = n1059 ^ n859 ^ n856 ;
  assign n1096 = ( ~x49 & n681 ) | ( ~x49 & n877 ) | ( n681 & n877 ) ;
  assign n1097 = n1096 ^ n717 ^ 1'b0 ;
  assign n1098 = ~n281 & n986 ;
  assign n1099 = x1 & n920 ;
  assign n1100 = n1099 ^ x70 ^ 1'b0 ;
  assign n1101 = n1100 ^ n753 ^ n598 ;
  assign n1102 = n919 ^ x47 ^ 1'b0 ;
  assign n1103 = n170 & n1102 ;
  assign n1104 = n766 ^ n230 ^ x59 ;
  assign n1105 = n1104 ^ n348 ^ 1'b0 ;
  assign n1106 = n1103 & n1105 ;
  assign n1107 = n1101 & n1106 ;
  assign n1108 = ( n404 & ~n448 ) | ( n404 & n1107 ) | ( ~n448 & n1107 ) ;
  assign n1109 = n354 & ~n437 ;
  assign n1110 = n873 & n1109 ;
  assign n1111 = ( n549 & n976 ) | ( n549 & n1048 ) | ( n976 & n1048 ) ;
  assign n1112 = n1110 | n1111 ;
  assign n1113 = n1108 & ~n1112 ;
  assign n1114 = ~x50 & n786 ;
  assign n1115 = n679 ^ n267 ^ 1'b0 ;
  assign n1116 = ~n984 & n1115 ;
  assign n1119 = x100 ^ x27 ^ 1'b0 ;
  assign n1120 = x72 & n1119 ;
  assign n1118 = x127 & ~n657 ;
  assign n1121 = n1120 ^ n1118 ^ 1'b0 ;
  assign n1122 = n256 | n1121 ;
  assign n1123 = n706 | n1122 ;
  assign n1124 = n1123 ^ n416 ^ n153 ;
  assign n1117 = n262 ^ n209 ^ 1'b0 ;
  assign n1125 = n1124 ^ n1117 ^ 1'b0 ;
  assign n1126 = ~n442 & n1125 ;
  assign n1127 = n632 & n1074 ;
  assign n1128 = ~n310 & n1127 ;
  assign n1129 = ( n230 & ~n544 ) | ( n230 & n815 ) | ( ~n544 & n815 ) ;
  assign n1130 = n1129 ^ n517 ^ 1'b0 ;
  assign n1131 = n149 | n1130 ;
  assign n1132 = n246 ^ n132 ^ x59 ;
  assign n1133 = n504 & ~n1132 ;
  assign n1134 = n1131 & n1133 ;
  assign n1135 = n1134 ^ n301 ^ 1'b0 ;
  assign n1136 = x44 & ~n1135 ;
  assign n1137 = ~x71 & n1136 ;
  assign n1138 = n618 & n1137 ;
  assign n1139 = ( x100 & n250 ) | ( x100 & n481 ) | ( n250 & n481 ) ;
  assign n1140 = x5 & ~n447 ;
  assign n1141 = n1140 ^ n259 ^ 1'b0 ;
  assign n1142 = n161 & n1141 ;
  assign n1143 = ~n1139 & n1142 ;
  assign n1144 = n1056 | n1143 ;
  assign n1145 = n1144 ^ n710 ^ 1'b0 ;
  assign n1146 = x62 & n854 ;
  assign n1147 = ( ~x9 & n305 ) | ( ~x9 & n577 ) | ( n305 & n577 ) ;
  assign n1148 = n692 ^ n216 ^ 1'b0 ;
  assign n1149 = n1147 | n1148 ;
  assign n1150 = n1149 ^ n899 ^ n791 ;
  assign n1151 = n917 & n1150 ;
  assign n1152 = ~n270 & n1151 ;
  assign n1153 = n781 ^ n502 ^ 1'b0 ;
  assign n1154 = n162 | n604 ;
  assign n1157 = x0 & ~n383 ;
  assign n1158 = ~n454 & n538 ;
  assign n1159 = ~x36 & n1158 ;
  assign n1160 = n1159 ^ n710 ^ 1'b0 ;
  assign n1161 = n449 & n1160 ;
  assign n1162 = n1161 ^ n1015 ^ 1'b0 ;
  assign n1163 = n1162 ^ x33 ^ 1'b0 ;
  assign n1164 = n1157 & n1163 ;
  assign n1165 = x36 & n266 ;
  assign n1166 = ~n346 & n1165 ;
  assign n1167 = ~n1164 & n1166 ;
  assign n1155 = n789 ^ n471 ^ 1'b0 ;
  assign n1156 = n202 & ~n1155 ;
  assign n1168 = n1167 ^ n1156 ^ 1'b0 ;
  assign n1169 = n1168 ^ x23 ^ 1'b0 ;
  assign n1170 = n1154 | n1169 ;
  assign n1171 = n370 ^ x44 ^ 1'b0 ;
  assign n1172 = n1171 ^ n141 ^ 1'b0 ;
  assign n1173 = n1017 ^ n245 ^ 1'b0 ;
  assign n1174 = n159 ^ x72 ^ 1'b0 ;
  assign n1175 = ~n567 & n1174 ;
  assign n1176 = ( ~n312 & n315 ) | ( ~n312 & n707 ) | ( n315 & n707 ) ;
  assign n1177 = n1175 & n1176 ;
  assign n1178 = n1177 ^ n806 ^ 1'b0 ;
  assign n1179 = n1173 & n1178 ;
  assign n1180 = n566 & n1179 ;
  assign n1181 = n352 | n363 ;
  assign n1182 = n259 & ~n1181 ;
  assign n1183 = n182 & n374 ;
  assign n1184 = n1183 ^ x54 ^ 1'b0 ;
  assign n1185 = n1184 ^ n527 ^ 1'b0 ;
  assign n1186 = n1060 ^ n1041 ^ 1'b0 ;
  assign n1187 = x62 & n1186 ;
  assign n1188 = ( ~n485 & n1185 ) | ( ~n485 & n1187 ) | ( n1185 & n1187 ) ;
  assign n1189 = n1182 | n1188 ;
  assign n1190 = ( x27 & n328 ) | ( x27 & ~n819 ) | ( n328 & ~n819 ) ;
  assign n1191 = x39 & ~n425 ;
  assign n1192 = n192 & n1191 ;
  assign n1193 = n1192 ^ n190 ^ n157 ;
  assign n1194 = n1193 ^ x47 ^ 1'b0 ;
  assign n1195 = x75 & n1067 ;
  assign n1196 = n1195 ^ n465 ^ 1'b0 ;
  assign n1197 = n1196 ^ n555 ^ 1'b0 ;
  assign n1198 = n393 & n1197 ;
  assign n1199 = n1198 ^ n437 ^ 1'b0 ;
  assign n1200 = n1199 ^ x74 ^ 1'b0 ;
  assign n1201 = ( ~n333 & n1194 ) | ( ~n333 & n1200 ) | ( n1194 & n1200 ) ;
  assign n1202 = n719 ^ n275 ^ 1'b0 ;
  assign n1203 = n386 ^ n277 ^ 1'b0 ;
  assign n1204 = n1175 & n1203 ;
  assign n1205 = n476 | n963 ;
  assign n1206 = ( x69 & n190 ) | ( x69 & n245 ) | ( n190 & n245 ) ;
  assign n1207 = n1206 ^ n1084 ^ n956 ;
  assign n1208 = ( ~x75 & n265 ) | ( ~x75 & n646 ) | ( n265 & n646 ) ;
  assign n1209 = ( x6 & ~x13 ) | ( x6 & n460 ) | ( ~x13 & n460 ) ;
  assign n1210 = n945 ^ x57 ^ 1'b0 ;
  assign n1211 = ~n1209 & n1210 ;
  assign n1212 = n533 ^ n233 ^ x8 ;
  assign n1213 = n1211 & ~n1212 ;
  assign n1214 = n1213 ^ n736 ^ 1'b0 ;
  assign n1215 = n1208 | n1214 ;
  assign n1216 = ~n529 & n537 ;
  assign n1217 = ~n1103 & n1216 ;
  assign n1218 = n707 & n1217 ;
  assign n1219 = n1017 ^ n646 ^ n573 ;
  assign n1220 = ( x75 & ~n550 ) | ( x75 & n1219 ) | ( ~n550 & n1219 ) ;
  assign n1221 = n1220 ^ n321 ^ 1'b0 ;
  assign n1222 = x108 & x112 ;
  assign n1223 = n1222 ^ n415 ^ 1'b0 ;
  assign n1224 = n1223 ^ n1097 ^ 1'b0 ;
  assign n1225 = n325 | n1224 ;
  assign n1226 = n1160 ^ n980 ^ 1'b0 ;
  assign n1227 = ( ~n856 & n1006 ) | ( ~n856 & n1226 ) | ( n1006 & n1226 ) ;
  assign n1233 = n383 | n1149 ;
  assign n1234 = n760 & ~n1233 ;
  assign n1230 = n1067 ^ x60 ^ x39 ;
  assign n1229 = ( x78 & ~n493 ) | ( x78 & n776 ) | ( ~n493 & n776 ) ;
  assign n1231 = n1230 ^ n1229 ^ 1'b0 ;
  assign n1232 = n167 & ~n1231 ;
  assign n1235 = n1234 ^ n1232 ^ n946 ;
  assign n1228 = x28 & n380 ;
  assign n1236 = n1235 ^ n1228 ^ 1'b0 ;
  assign n1237 = n214 & ~n248 ;
  assign n1238 = n1237 ^ n689 ^ 1'b0 ;
  assign n1239 = ~n554 & n923 ;
  assign n1240 = n1239 ^ n266 ^ 1'b0 ;
  assign n1241 = n197 | n1240 ;
  assign n1242 = n1241 ^ n262 ^ 1'b0 ;
  assign n1243 = n1238 | n1242 ;
  assign n1244 = n1243 ^ n1072 ^ n332 ;
  assign n1249 = n266 & n486 ;
  assign n1250 = ~n424 & n1249 ;
  assign n1245 = x34 & x91 ;
  assign n1246 = n1245 ^ x112 ^ 1'b0 ;
  assign n1247 = n605 & n744 ;
  assign n1248 = ~n1246 & n1247 ;
  assign n1251 = n1250 ^ n1248 ^ 1'b0 ;
  assign n1252 = n1251 ^ x108 ^ x30 ;
  assign n1253 = n636 ^ n477 ^ n281 ;
  assign n1254 = n1253 ^ n393 ^ n248 ;
  assign n1255 = n1035 & ~n1254 ;
  assign n1256 = n1252 & n1255 ;
  assign n1259 = n930 & n938 ;
  assign n1260 = n1259 ^ n624 ^ 1'b0 ;
  assign n1257 = n1079 ^ n607 ^ 1'b0 ;
  assign n1258 = n733 | n1257 ;
  assign n1261 = n1260 ^ n1258 ^ n569 ;
  assign n1262 = ( ~n356 & n408 ) | ( ~n356 & n732 ) | ( n408 & n732 ) ;
  assign n1263 = ( x55 & ~n472 ) | ( x55 & n525 ) | ( ~n472 & n525 ) ;
  assign n1264 = n857 & n1263 ;
  assign n1265 = ~n198 & n928 ;
  assign n1266 = n1265 ^ n708 ^ 1'b0 ;
  assign n1267 = ~n246 & n1266 ;
  assign n1268 = n1212 ^ n945 ^ 1'b0 ;
  assign n1269 = n1268 ^ n373 ^ 1'b0 ;
  assign n1270 = n1051 & n1269 ;
  assign n1271 = ~n586 & n1270 ;
  assign n1272 = n383 & ~n664 ;
  assign n1273 = ( n657 & n919 ) | ( n657 & n1104 ) | ( n919 & n1104 ) ;
  assign n1274 = n1273 ^ n349 ^ 1'b0 ;
  assign n1275 = n1251 ^ n835 ^ 1'b0 ;
  assign n1283 = n292 & n742 ;
  assign n1276 = ( n216 & ~n487 ) | ( n216 & n583 ) | ( ~n487 & n583 ) ;
  assign n1277 = ( x125 & ~n242 ) | ( x125 & n357 ) | ( ~n242 & n357 ) ;
  assign n1278 = n1277 ^ n442 ^ n287 ;
  assign n1279 = ( n633 & ~n723 ) | ( n633 & n1278 ) | ( ~n723 & n1278 ) ;
  assign n1280 = ( x60 & n198 ) | ( x60 & ~n1279 ) | ( n198 & ~n1279 ) ;
  assign n1281 = n1276 & ~n1280 ;
  assign n1282 = n296 & n1281 ;
  assign n1284 = n1283 ^ n1282 ^ 1'b0 ;
  assign n1285 = n1275 & n1284 ;
  assign n1286 = n1270 ^ n557 ^ 1'b0 ;
  assign n1287 = x22 & ~n314 ;
  assign n1288 = n1287 ^ n1100 ^ n262 ;
  assign n1289 = ( n134 & ~n210 ) | ( n134 & n753 ) | ( ~n210 & n753 ) ;
  assign n1290 = n1289 ^ n274 ^ 1'b0 ;
  assign n1291 = ( ~n1003 & n1061 ) | ( ~n1003 & n1079 ) | ( n1061 & n1079 ) ;
  assign n1292 = n146 ^ x28 ^ 1'b0 ;
  assign n1293 = n136 & n302 ;
  assign n1294 = ~n202 & n1293 ;
  assign n1295 = n1294 ^ x80 ^ x77 ;
  assign n1296 = n1295 ^ n545 ^ x38 ;
  assign n1297 = n1206 | n1296 ;
  assign n1298 = n1297 ^ n296 ^ 1'b0 ;
  assign n1299 = n1292 & ~n1298 ;
  assign n1309 = n224 & ~n800 ;
  assign n1305 = ~n749 & n952 ;
  assign n1306 = n1305 ^ x48 ^ 1'b0 ;
  assign n1300 = ~n260 & n472 ;
  assign n1301 = n1238 & n1300 ;
  assign n1302 = n375 | n1301 ;
  assign n1303 = n488 & ~n1302 ;
  assign n1304 = n1303 ^ n491 ^ 1'b0 ;
  assign n1307 = n1306 ^ n1304 ^ 1'b0 ;
  assign n1308 = ~n844 & n1307 ;
  assign n1310 = n1309 ^ n1308 ^ n703 ;
  assign n1319 = ( ~x21 & n350 ) | ( ~x21 & n656 ) | ( n350 & n656 ) ;
  assign n1311 = x113 ^ x111 ^ x15 ;
  assign n1312 = n1311 ^ n624 ^ n597 ;
  assign n1313 = n768 & ~n1312 ;
  assign n1314 = ~x52 & n1313 ;
  assign n1315 = x21 & ~n1314 ;
  assign n1316 = ~x120 & n1315 ;
  assign n1317 = n361 ^ n154 ^ 1'b0 ;
  assign n1318 = ( n318 & n1316 ) | ( n318 & ~n1317 ) | ( n1316 & ~n1317 ) ;
  assign n1320 = n1319 ^ n1318 ^ 1'b0 ;
  assign n1321 = ( n474 & n514 ) | ( n474 & n612 ) | ( n514 & n612 ) ;
  assign n1322 = n409 ^ n279 ^ 1'b0 ;
  assign n1323 = n746 | n1322 ;
  assign n1324 = n851 ^ x28 ^ 1'b0 ;
  assign n1325 = n176 & ~n295 ;
  assign n1326 = n1324 & n1325 ;
  assign n1327 = ~n915 & n1326 ;
  assign n1328 = ( x18 & ~n1260 ) | ( x18 & n1327 ) | ( ~n1260 & n1327 ) ;
  assign n1332 = n540 ^ n457 ^ n413 ;
  assign n1333 = n1332 ^ n893 ^ n316 ;
  assign n1329 = x52 & n165 ;
  assign n1330 = n1004 ^ n650 ^ 1'b0 ;
  assign n1331 = ~n1329 & n1330 ;
  assign n1334 = n1333 ^ n1331 ^ 1'b0 ;
  assign n1338 = ( x102 & n287 ) | ( x102 & ~n366 ) | ( n287 & ~n366 ) ;
  assign n1335 = n597 | n925 ;
  assign n1336 = n1335 ^ n615 ^ 1'b0 ;
  assign n1337 = n1336 ^ n1212 ^ n421 ;
  assign n1339 = n1338 ^ n1337 ^ n851 ;
  assign n1340 = n1339 ^ n945 ^ n202 ;
  assign n1341 = n734 ^ n537 ^ n149 ;
  assign n1342 = ( ~x89 & n787 ) | ( ~x89 & n1341 ) | ( n787 & n1341 ) ;
  assign n1343 = n476 ^ n439 ^ 1'b0 ;
  assign n1344 = ~n627 & n863 ;
  assign n1345 = ~n398 & n1344 ;
  assign n1346 = ( n404 & n739 ) | ( n404 & n1139 ) | ( n739 & n1139 ) ;
  assign n1347 = n789 & n1346 ;
  assign n1348 = n1347 ^ n206 ^ 1'b0 ;
  assign n1349 = ( n924 & n1345 ) | ( n924 & ~n1348 ) | ( n1345 & ~n1348 ) ;
  assign n1350 = n935 | n1349 ;
  assign n1354 = n537 ^ n320 ^ 1'b0 ;
  assign n1351 = n1302 ^ n205 ^ 1'b0 ;
  assign n1352 = n1282 | n1351 ;
  assign n1353 = n1090 | n1352 ;
  assign n1355 = n1354 ^ n1353 ^ 1'b0 ;
  assign n1356 = n572 & ~n681 ;
  assign n1357 = n1356 ^ n1015 ^ 1'b0 ;
  assign n1358 = n1219 ^ n157 ^ 1'b0 ;
  assign n1359 = n514 | n1358 ;
  assign n1360 = n1359 ^ n1092 ^ 1'b0 ;
  assign n1361 = n399 | n835 ;
  assign n1362 = ~n970 & n1361 ;
  assign n1363 = n1362 ^ n290 ^ 1'b0 ;
  assign n1364 = ( ~n262 & n1360 ) | ( ~n262 & n1363 ) | ( n1360 & n1363 ) ;
  assign n1365 = n356 & ~n366 ;
  assign n1366 = n1365 ^ n208 ^ x23 ;
  assign n1367 = n1217 | n1366 ;
  assign n1368 = n584 & ~n1367 ;
  assign n1369 = n1368 ^ n537 ^ 1'b0 ;
  assign n1370 = n143 & ~n543 ;
  assign n1371 = ( n164 & ~n1345 ) | ( n164 & n1370 ) | ( ~n1345 & n1370 ) ;
  assign n1372 = ( ~x31 & n200 ) | ( ~x31 & n421 ) | ( n200 & n421 ) ;
  assign n1373 = n1073 | n1372 ;
  assign n1374 = n447 & ~n1373 ;
  assign n1375 = x120 & ~n1374 ;
  assign n1376 = ~n1371 & n1375 ;
  assign n1377 = ( n1060 & ~n1063 ) | ( n1060 & n1376 ) | ( ~n1063 & n1376 ) ;
  assign n1378 = n1036 ^ n649 ^ 1'b0 ;
  assign n1381 = n1086 ^ n374 ^ n186 ;
  assign n1382 = n1381 ^ x53 ^ x17 ;
  assign n1383 = ( ~x102 & n151 ) | ( ~x102 & n1382 ) | ( n151 & n1382 ) ;
  assign n1384 = n1383 ^ n946 ^ n942 ;
  assign n1379 = n1324 ^ n1082 ^ n316 ;
  assign n1380 = n571 & n1379 ;
  assign n1385 = n1384 ^ n1380 ^ 1'b0 ;
  assign n1386 = ~n328 & n1385 ;
  assign n1387 = n1386 ^ n1199 ^ 1'b0 ;
  assign n1388 = n1387 ^ n789 ^ n597 ;
  assign n1389 = ( n492 & n734 ) | ( n492 & ~n1019 ) | ( n734 & ~n1019 ) ;
  assign n1390 = n319 | n1113 ;
  assign n1391 = n851 ^ n742 ^ n714 ;
  assign n1392 = n1391 ^ n472 ^ x16 ;
  assign n1393 = n367 ^ x55 ^ 1'b0 ;
  assign n1394 = n1392 & ~n1393 ;
  assign n1395 = n675 & n1394 ;
  assign n1396 = n1395 ^ n866 ^ 1'b0 ;
  assign n1397 = n204 | n692 ;
  assign n1398 = n1145 | n1359 ;
  assign n1399 = n1397 & ~n1398 ;
  assign n1400 = n563 ^ x42 ^ 1'b0 ;
  assign n1401 = n598 | n1400 ;
  assign n1402 = n1401 ^ n1240 ^ 1'b0 ;
  assign n1403 = n210 | n1402 ;
  assign n1404 = n725 | n1403 ;
  assign n1405 = ~n275 & n897 ;
  assign n1406 = ( ~n238 & n296 ) | ( ~n238 & n1405 ) | ( n296 & n1405 ) ;
  assign n1407 = n1406 ^ n655 ^ 1'b0 ;
  assign n1408 = n325 ^ n308 ^ 1'b0 ;
  assign n1409 = ~n269 & n1408 ;
  assign n1410 = x111 & n1409 ;
  assign n1411 = n1410 ^ n1312 ^ 1'b0 ;
  assign n1412 = n639 & n1247 ;
  assign n1413 = ( n221 & n262 ) | ( n221 & ~n332 ) | ( n262 & ~n332 ) ;
  assign n1414 = n1413 ^ n804 ^ 1'b0 ;
  assign n1415 = n1412 & n1414 ;
  assign n1416 = n1162 ^ n771 ^ 1'b0 ;
  assign n1417 = ( ~n1411 & n1415 ) | ( ~n1411 & n1416 ) | ( n1415 & n1416 ) ;
  assign n1418 = ( n194 & ~n969 ) | ( n194 & n1242 ) | ( ~n969 & n1242 ) ;
  assign n1419 = n301 & n1418 ;
  assign n1431 = n358 & ~n379 ;
  assign n1429 = n994 | n1002 ;
  assign n1427 = n663 ^ n208 ^ x104 ;
  assign n1426 = ~x86 & n131 ;
  assign n1428 = n1427 ^ n1426 ^ n131 ;
  assign n1430 = n1429 ^ n1428 ^ n689 ;
  assign n1420 = ( n188 & n219 ) | ( n188 & n560 ) | ( n219 & n560 ) ;
  assign n1422 = n699 ^ n431 ^ x116 ;
  assign n1421 = n618 & ~n1037 ;
  assign n1423 = n1422 ^ n1421 ^ 1'b0 ;
  assign n1424 = n1420 & ~n1423 ;
  assign n1425 = ~n582 & n1424 ;
  assign n1432 = n1431 ^ n1430 ^ n1425 ;
  assign n1433 = n675 & ~n987 ;
  assign n1434 = n1433 ^ n343 ^ 1'b0 ;
  assign n1435 = n694 & n806 ;
  assign n1437 = n1361 ^ n815 ^ 1'b0 ;
  assign n1436 = n169 & ~n940 ;
  assign n1438 = n1437 ^ n1436 ^ 1'b0 ;
  assign n1439 = ( n1079 & n1435 ) | ( n1079 & ~n1438 ) | ( n1435 & ~n1438 ) ;
  assign n1441 = n226 ^ x104 ^ x102 ;
  assign n1440 = n238 | n873 ;
  assign n1442 = n1441 ^ n1440 ^ 1'b0 ;
  assign n1443 = ( x34 & n1337 ) | ( x34 & n1442 ) | ( n1337 & n1442 ) ;
  assign n1444 = n672 & n1443 ;
  assign n1446 = n437 ^ n164 ^ 1'b0 ;
  assign n1445 = ( n981 & n1084 ) | ( n981 & ~n1392 ) | ( n1084 & ~n1392 ) ;
  assign n1447 = n1446 ^ n1445 ^ 1'b0 ;
  assign n1448 = n277 ^ x36 ^ 1'b0 ;
  assign n1449 = x2 & ~n1448 ;
  assign n1450 = n1020 ^ n872 ^ n151 ;
  assign n1451 = n547 & n1450 ;
  assign n1452 = n1003 ^ n582 ^ 1'b0 ;
  assign n1453 = n1451 | n1452 ;
  assign n1454 = n655 ^ n370 ^ 1'b0 ;
  assign n1455 = n1162 ^ n775 ^ n669 ;
  assign n1456 = ( ~n611 & n1454 ) | ( ~n611 & n1455 ) | ( n1454 & n1455 ) ;
  assign n1457 = n979 & n1456 ;
  assign n1458 = n628 & n1457 ;
  assign n1459 = ~n322 & n512 ;
  assign n1460 = ~n924 & n1459 ;
  assign n1461 = n567 ^ x21 ^ 1'b0 ;
  assign n1462 = n266 & ~n1461 ;
  assign n1463 = n1462 ^ n1422 ^ n164 ;
  assign n1464 = n584 & n1348 ;
  assign n1465 = x58 & ~n1055 ;
  assign n1466 = n1465 ^ n933 ^ 1'b0 ;
  assign n1467 = n1292 ^ n200 ^ 1'b0 ;
  assign n1468 = n1466 | n1467 ;
  assign n1472 = n154 & n1406 ;
  assign n1469 = n845 ^ n329 ^ 1'b0 ;
  assign n1470 = n689 & n1469 ;
  assign n1471 = n422 & n1470 ;
  assign n1473 = n1472 ^ n1471 ^ n786 ;
  assign n1474 = n1473 ^ n779 ^ 1'b0 ;
  assign n1475 = n1468 & n1474 ;
  assign n1476 = n732 ^ n669 ^ 1'b0 ;
  assign n1477 = n982 & n1476 ;
  assign n1478 = n1192 & n1477 ;
  assign n1479 = x19 & x98 ;
  assign n1480 = ~x111 & n1479 ;
  assign n1481 = n1480 ^ x35 ^ 1'b0 ;
  assign n1482 = n1466 & ~n1481 ;
  assign n1483 = ~n1101 & n1482 ;
  assign n1484 = n1478 & n1483 ;
  assign n1485 = x2 & n667 ;
  assign n1486 = n485 | n1138 ;
  assign n1487 = n1486 ^ n455 ^ 1'b0 ;
  assign n1488 = ( ~n901 & n1485 ) | ( ~n901 & n1487 ) | ( n1485 & n1487 ) ;
  assign n1490 = ( n132 & n224 ) | ( n132 & n1157 ) | ( n224 & n1157 ) ;
  assign n1491 = n970 ^ x127 ^ 1'b0 ;
  assign n1492 = n1490 & ~n1491 ;
  assign n1489 = ~n1044 & n1475 ;
  assign n1493 = n1492 ^ n1489 ^ 1'b0 ;
  assign n1494 = n571 ^ n511 ^ 1'b0 ;
  assign n1495 = n1494 ^ x101 ^ 1'b0 ;
  assign n1496 = n817 | n1495 ;
  assign n1497 = n154 & ~n770 ;
  assign n1498 = n1496 & n1497 ;
  assign n1499 = ( x21 & n165 ) | ( x21 & n574 ) | ( n165 & n574 ) ;
  assign n1500 = n1499 ^ n932 ^ 1'b0 ;
  assign n1501 = x88 & n1500 ;
  assign n1503 = n374 | n439 ;
  assign n1502 = x12 & n375 ;
  assign n1504 = n1503 ^ n1502 ^ 1'b0 ;
  assign n1505 = n940 ^ n352 ^ n294 ;
  assign n1506 = n1505 ^ n555 ^ 1'b0 ;
  assign n1507 = n199 & n1506 ;
  assign n1508 = n196 | n517 ;
  assign n1509 = ~n1007 & n1508 ;
  assign n1510 = n1056 ^ n596 ^ 1'b0 ;
  assign n1511 = n1510 ^ n1234 ^ x62 ;
  assign n1512 = n774 & ~n1511 ;
  assign n1513 = n803 & n1512 ;
  assign n1514 = ( n218 & ~n738 ) | ( n218 & n885 ) | ( ~n738 & n885 ) ;
  assign n1515 = n180 | n1514 ;
  assign n1516 = n1515 ^ n449 ^ n210 ;
  assign n1517 = n1366 ^ x58 ^ 1'b0 ;
  assign n1518 = ( n383 & n1446 ) | ( n383 & n1517 ) | ( n1446 & n1517 ) ;
  assign n1519 = ( n147 & n485 ) | ( n147 & n1518 ) | ( n485 & n1518 ) ;
  assign n1520 = n277 & ~n817 ;
  assign n1521 = n531 ^ x76 ^ 1'b0 ;
  assign n1522 = n717 & ~n1521 ;
  assign n1523 = ~n635 & n1522 ;
  assign n1524 = n473 | n1523 ;
  assign n1525 = n1524 ^ n304 ^ 1'b0 ;
  assign n1526 = ( x77 & ~n1019 ) | ( x77 & n1024 ) | ( ~n1019 & n1024 ) ;
  assign n1527 = n1526 ^ n603 ^ 1'b0 ;
  assign n1530 = n298 ^ n176 ^ x81 ;
  assign n1531 = n154 & ~n1530 ;
  assign n1532 = n512 & n1531 ;
  assign n1533 = ~n699 & n1532 ;
  assign n1534 = ( n777 & ~n791 ) | ( n777 & n1533 ) | ( ~n791 & n1533 ) ;
  assign n1528 = x73 & n842 ;
  assign n1529 = n1528 ^ n737 ^ 1'b0 ;
  assign n1535 = n1534 ^ n1529 ^ n911 ;
  assign n1536 = n1527 & ~n1535 ;
  assign n1537 = ~x89 & n1536 ;
  assign n1540 = n501 ^ n178 ^ 1'b0 ;
  assign n1538 = n316 & n631 ;
  assign n1539 = ~n567 & n1538 ;
  assign n1541 = n1540 ^ n1539 ^ 1'b0 ;
  assign n1552 = n512 & ~n1494 ;
  assign n1553 = ~x2 & n1552 ;
  assign n1554 = n1553 ^ n1517 ^ 1'b0 ;
  assign n1551 = x104 & ~n819 ;
  assign n1546 = ( ~n461 & n533 ) | ( ~n461 & n632 ) | ( n533 & n632 ) ;
  assign n1543 = n469 ^ n157 ^ x54 ;
  assign n1544 = x67 & ~n1543 ;
  assign n1545 = n1230 & n1544 ;
  assign n1547 = n1546 ^ n1545 ^ x84 ;
  assign n1542 = ( n452 & n517 ) | ( n452 & n1004 ) | ( n517 & n1004 ) ;
  assign n1548 = n1547 ^ n1542 ^ n194 ;
  assign n1549 = n408 & n1548 ;
  assign n1550 = n1549 ^ n543 ^ 1'b0 ;
  assign n1555 = n1554 ^ n1551 ^ n1550 ;
  assign n1556 = ( n621 & n637 ) | ( n621 & ~n695 ) | ( n637 & ~n695 ) ;
  assign n1557 = n891 & n1556 ;
  assign n1558 = ~n1445 & n1557 ;
  assign n1559 = ( n281 & n548 ) | ( n281 & n1309 ) | ( n548 & n1309 ) ;
  assign n1560 = x124 ^ x119 ^ 1'b0 ;
  assign n1561 = n269 & n1560 ;
  assign n1562 = n343 ^ n335 ^ n146 ;
  assign n1563 = n1561 & n1562 ;
  assign n1564 = n1563 ^ n840 ^ 1'b0 ;
  assign n1565 = n512 & n1564 ;
  assign n1566 = ~n1559 & n1565 ;
  assign n1567 = n366 | n1566 ;
  assign n1568 = n1567 ^ n627 ^ 1'b0 ;
  assign n1569 = n180 & n1568 ;
  assign n1570 = ( n921 & ~n1051 ) | ( n921 & n1412 ) | ( ~n1051 & n1412 ) ;
  assign n1572 = n1187 ^ n658 ^ 1'b0 ;
  assign n1573 = n472 & n1572 ;
  assign n1571 = ( n208 & n986 ) | ( n208 & ~n1182 ) | ( n986 & ~n1182 ) ;
  assign n1574 = n1573 ^ n1571 ^ n588 ;
  assign n1575 = n277 ^ x11 ^ 1'b0 ;
  assign n1576 = n132 & n1575 ;
  assign n1579 = ( x66 & n357 ) | ( x66 & ~n679 ) | ( n357 & ~n679 ) ;
  assign n1577 = n545 & n706 ;
  assign n1578 = n1577 ^ n551 ^ 1'b0 ;
  assign n1580 = n1579 ^ n1578 ^ 1'b0 ;
  assign n1585 = n441 ^ n171 ^ 1'b0 ;
  assign n1584 = n187 & ~n250 ;
  assign n1586 = n1585 ^ n1584 ^ 1'b0 ;
  assign n1582 = n539 ^ n270 ^ 1'b0 ;
  assign n1583 = n211 | n1582 ;
  assign n1581 = n1566 ^ n841 ^ n476 ;
  assign n1587 = n1586 ^ n1583 ^ n1581 ;
  assign n1588 = n1587 ^ n871 ^ 1'b0 ;
  assign n1589 = n798 ^ x69 ^ 1'b0 ;
  assign n1590 = ~n1246 & n1589 ;
  assign n1591 = n1590 ^ n965 ^ n506 ;
  assign n1592 = n1048 ^ x75 ^ 1'b0 ;
  assign n1593 = ~n971 & n1592 ;
  assign n1594 = ~n1058 & n1593 ;
  assign n1595 = n426 ^ n335 ^ 1'b0 ;
  assign n1596 = n1135 | n1595 ;
  assign n1597 = n1596 ^ n873 ^ 1'b0 ;
  assign n1598 = ( x68 & ~n264 ) | ( x68 & n1597 ) | ( ~n264 & n1597 ) ;
  assign n1599 = ~n238 & n590 ;
  assign n1600 = n1599 ^ n1554 ^ n1295 ;
  assign n1601 = ( n817 & ~n855 ) | ( n817 & n1600 ) | ( ~n855 & n1600 ) ;
  assign n1602 = n977 ^ n661 ^ n224 ;
  assign n1603 = n1602 ^ n986 ^ 1'b0 ;
  assign n1604 = x123 & n421 ;
  assign n1605 = ~n1165 & n1604 ;
  assign n1606 = n1330 & ~n1605 ;
  assign n1607 = ~n1178 & n1606 ;
  assign n1608 = ( n155 & n971 ) | ( n155 & n1338 ) | ( n971 & n1338 ) ;
  assign n1609 = n1608 ^ n398 ^ x90 ;
  assign n1610 = n1345 ^ n833 ^ 1'b0 ;
  assign n1611 = n756 & ~n1610 ;
  assign n1612 = n1611 ^ n883 ^ n848 ;
  assign n1615 = n952 ^ n829 ^ n203 ;
  assign n1613 = n946 ^ n687 ^ 1'b0 ;
  assign n1614 = n789 & ~n1613 ;
  assign n1616 = n1615 ^ n1614 ^ 1'b0 ;
  assign n1617 = n1566 ^ n253 ^ n170 ;
  assign n1618 = n1053 & ~n1617 ;
  assign n1619 = n1618 ^ n733 ^ 1'b0 ;
  assign n1620 = n1304 ^ x44 ^ 1'b0 ;
  assign n1621 = n238 | n1620 ;
  assign n1622 = n1621 ^ n1553 ^ n269 ;
  assign n1623 = n144 ^ x115 ^ x52 ;
  assign n1624 = n1623 ^ n562 ^ n331 ;
  assign n1626 = x87 ^ x14 ^ 1'b0 ;
  assign n1625 = n386 ^ x0 ^ 1'b0 ;
  assign n1627 = n1626 ^ n1625 ^ n1250 ;
  assign n1628 = ( ~n1113 & n1624 ) | ( ~n1113 & n1627 ) | ( n1624 & n1627 ) ;
  assign n1629 = n1628 ^ n1608 ^ n1176 ;
  assign n1638 = ~x18 & n1446 ;
  assign n1635 = ~n887 & n1279 ;
  assign n1636 = ( ~x25 & x63 ) | ( ~x25 & n1635 ) | ( x63 & n1635 ) ;
  assign n1637 = n1145 & ~n1636 ;
  assign n1630 = ~n448 & n1379 ;
  assign n1631 = n149 & n1630 ;
  assign n1632 = n1631 ^ n1009 ^ 1'b0 ;
  assign n1633 = n314 | n1632 ;
  assign n1634 = n1337 & ~n1633 ;
  assign n1639 = n1638 ^ n1637 ^ n1634 ;
  assign n1640 = n1288 ^ n466 ^ 1'b0 ;
  assign n1641 = n251 | n306 ;
  assign n1642 = ( x64 & ~x84 ) | ( x64 & n1641 ) | ( ~x84 & n1641 ) ;
  assign n1643 = n481 | n531 ;
  assign n1644 = n789 ^ n522 ^ n486 ;
  assign n1645 = ~n940 & n1415 ;
  assign n1646 = ( n605 & n1644 ) | ( n605 & ~n1645 ) | ( n1644 & ~n1645 ) ;
  assign n1647 = n1077 ^ n586 ^ n390 ;
  assign n1648 = x19 | n615 ;
  assign n1649 = n270 | n1648 ;
  assign n1650 = n1649 ^ n1003 ^ n301 ;
  assign n1651 = n687 & n1650 ;
  assign n1652 = ~n1647 & n1651 ;
  assign n1653 = n1652 ^ n1291 ^ 1'b0 ;
  assign n1654 = n535 & ~n822 ;
  assign n1655 = ~n552 & n881 ;
  assign n1656 = n848 & n1655 ;
  assign n1657 = n925 ^ n519 ^ 1'b0 ;
  assign n1658 = ~n970 & n1657 ;
  assign n1659 = n441 & n1658 ;
  assign n1660 = n1659 ^ n523 ^ 1'b0 ;
  assign n1661 = n226 & ~n1189 ;
  assign n1662 = x30 & n227 ;
  assign n1663 = n1662 ^ x120 ^ 1'b0 ;
  assign n1664 = n1663 ^ n1521 ^ 1'b0 ;
  assign n1669 = n544 | n659 ;
  assign n1670 = ~n473 & n770 ;
  assign n1671 = ~n1669 & n1670 ;
  assign n1672 = n1671 ^ n787 ^ 1'b0 ;
  assign n1673 = ~n984 & n1672 ;
  assign n1665 = x37 & ~n274 ;
  assign n1666 = n1665 ^ n465 ^ 1'b0 ;
  assign n1667 = ~n659 & n1630 ;
  assign n1668 = ~n1666 & n1667 ;
  assign n1674 = n1673 ^ n1668 ^ n1015 ;
  assign n1675 = n1243 | n1674 ;
  assign n1676 = n1675 ^ n1302 ^ 1'b0 ;
  assign n1677 = ~n165 & n1139 ;
  assign n1678 = n1677 ^ n639 ^ 1'b0 ;
  assign n1679 = n1678 ^ n1185 ^ 1'b0 ;
  assign n1680 = n815 & ~n942 ;
  assign n1681 = n439 & n1680 ;
  assign n1682 = n1681 ^ n1641 ^ n668 ;
  assign n1683 = ( ~n605 & n820 ) | ( ~n605 & n1028 ) | ( n820 & n1028 ) ;
  assign n1684 = n872 & n1683 ;
  assign n1685 = n1684 ^ n1152 ^ 1'b0 ;
  assign n1690 = n344 & n1157 ;
  assign n1686 = n627 ^ n535 ^ x59 ;
  assign n1687 = n1277 ^ n1024 ^ n318 ;
  assign n1688 = n1687 ^ n1448 ^ 1'b0 ;
  assign n1689 = ( n1627 & ~n1686 ) | ( n1627 & n1688 ) | ( ~n1686 & n1688 ) ;
  assign n1691 = n1690 ^ n1689 ^ n1382 ;
  assign n1692 = n488 ^ n344 ^ 1'b0 ;
  assign n1693 = n1218 ^ n394 ^ 1'b0 ;
  assign n1695 = ~n641 & n1687 ;
  assign n1696 = ( n1242 & n1693 ) | ( n1242 & ~n1695 ) | ( n1693 & ~n1695 ) ;
  assign n1694 = n492 & ~n1217 ;
  assign n1697 = n1696 ^ n1694 ^ 1'b0 ;
  assign n1698 = ( n1309 & ~n1693 ) | ( n1309 & n1697 ) | ( ~n1693 & n1697 ) ;
  assign n1699 = ~n1333 & n1647 ;
  assign n1700 = n1699 ^ n1003 ^ n956 ;
  assign n1701 = ( n659 & n1103 ) | ( n659 & n1515 ) | ( n1103 & n1515 ) ;
  assign n1702 = n997 ^ n812 ^ n767 ;
  assign n1703 = ~n1071 & n1702 ;
  assign n1704 = n1703 ^ n670 ^ 1'b0 ;
  assign n1705 = n1632 | n1704 ;
  assign n1706 = n786 ^ n667 ^ 1'b0 ;
  assign n1707 = n942 | n1706 ;
  assign n1708 = n891 & ~n1100 ;
  assign n1709 = n1707 & n1708 ;
  assign n1710 = ( n771 & n970 ) | ( n771 & ~n1024 ) | ( n970 & ~n1024 ) ;
  assign n1711 = ( n443 & n1709 ) | ( n443 & ~n1710 ) | ( n1709 & ~n1710 ) ;
  assign n1712 = ~n863 & n891 ;
  assign n1713 = ( n635 & ~n856 ) | ( n635 & n1712 ) | ( ~n856 & n1712 ) ;
  assign n1714 = ( n783 & ~n917 ) | ( n783 & n1407 ) | ( ~n917 & n1407 ) ;
  assign n1715 = ( ~x38 & n477 ) | ( ~x38 & n880 ) | ( n477 & n880 ) ;
  assign n1716 = n1715 ^ n441 ^ 1'b0 ;
  assign n1717 = n1716 ^ n945 ^ n703 ;
  assign n1718 = n168 & n1258 ;
  assign n1720 = ( n384 & n572 ) | ( n384 & ~n781 ) | ( n572 & ~n781 ) ;
  assign n1721 = n1253 ^ n398 ^ 1'b0 ;
  assign n1722 = n1720 | n1721 ;
  assign n1723 = n1722 ^ n533 ^ 1'b0 ;
  assign n1719 = ~n678 & n920 ;
  assign n1724 = n1723 ^ n1719 ^ 1'b0 ;
  assign n1725 = n1724 ^ n519 ^ n256 ;
  assign n1726 = n1715 ^ n759 ^ n458 ;
  assign n1727 = n174 & n1726 ;
  assign n1728 = n1725 & n1727 ;
  assign n1730 = ( n928 & n963 ) | ( n928 & n1134 ) | ( n963 & n1134 ) ;
  assign n1729 = ~n296 & n635 ;
  assign n1731 = n1730 ^ n1729 ^ 1'b0 ;
  assign n1732 = n1251 ^ n566 ^ 1'b0 ;
  assign n1733 = n914 ^ n251 ^ 1'b0 ;
  assign n1734 = n302 & ~n1733 ;
  assign n1735 = n1734 ^ x80 ^ 1'b0 ;
  assign n1736 = n202 & ~n346 ;
  assign n1737 = ~n817 & n1736 ;
  assign n1738 = ~n1411 & n1737 ;
  assign n1740 = n550 ^ x38 ^ 1'b0 ;
  assign n1739 = ( n158 & n1082 ) | ( n158 & ~n1543 ) | ( n1082 & ~n1543 ) ;
  assign n1741 = n1740 ^ n1739 ^ n1720 ;
  assign n1742 = n299 & ~n1107 ;
  assign n1743 = n1742 ^ n1545 ^ 1'b0 ;
  assign n1744 = n1743 ^ n1525 ^ n1425 ;
  assign n1745 = n1105 ^ n441 ^ n419 ;
  assign n1746 = x0 & n154 ;
  assign n1747 = n1745 & n1746 ;
  assign n1748 = n1074 & ~n1747 ;
  assign n1749 = ~n441 & n1748 ;
  assign n1750 = x87 & n822 ;
  assign n1751 = ~x68 & n1750 ;
  assign n1752 = ~n403 & n482 ;
  assign n1753 = n1751 & n1752 ;
  assign n1754 = n605 ^ n372 ^ x119 ;
  assign n1755 = n1753 | n1754 ;
  assign n1756 = n1167 & ~n1755 ;
  assign n1757 = ~n1656 & n1756 ;
  assign n1758 = n460 ^ x119 ^ 1'b0 ;
  assign n1759 = ( n501 & n1480 ) | ( n501 & ~n1758 ) | ( n1480 & ~n1758 ) ;
  assign n1760 = n1759 ^ x74 ^ 1'b0 ;
  assign n1761 = ( n165 & n1261 ) | ( n165 & n1420 ) | ( n1261 & n1420 ) ;
  assign n1764 = ~n184 & n260 ;
  assign n1762 = n1759 ^ x83 ^ 1'b0 ;
  assign n1763 = x20 & n1762 ;
  assign n1765 = n1764 ^ n1763 ^ n1134 ;
  assign n1766 = n831 ^ n206 ^ 1'b0 ;
  assign n1767 = ~n599 & n1766 ;
  assign n1768 = ~n810 & n1686 ;
  assign n1769 = ~n1060 & n1768 ;
  assign n1770 = ( n869 & n1141 ) | ( n869 & n1769 ) | ( n1141 & n1769 ) ;
  assign n1771 = ~n1311 & n1770 ;
  assign n1772 = ( x60 & n548 ) | ( x60 & ~n1485 ) | ( n548 & ~n1485 ) ;
  assign n1773 = n1342 ^ n1043 ^ n849 ;
  assign n1774 = ( ~n628 & n732 ) | ( ~n628 & n1341 ) | ( n732 & n1341 ) ;
  assign n1775 = n318 & ~n770 ;
  assign n1776 = ~n1123 & n1775 ;
  assign n1777 = ~x51 & x58 ;
  assign n1778 = ~n1776 & n1777 ;
  assign n1779 = n1774 & n1778 ;
  assign n1780 = n1779 ^ n206 ^ 1'b0 ;
  assign n1781 = ( ~n241 & n1685 ) | ( ~n241 & n1780 ) | ( n1685 & n1780 ) ;
  assign n1788 = n192 | n1044 ;
  assign n1789 = n1481 & ~n1788 ;
  assign n1790 = n976 | n1789 ;
  assign n1791 = n1790 ^ n590 ^ 1'b0 ;
  assign n1782 = n1061 | n1336 ;
  assign n1783 = n434 & ~n1782 ;
  assign n1784 = n1302 ^ n567 ^ 1'b0 ;
  assign n1785 = n1784 ^ n458 ^ 1'b0 ;
  assign n1786 = ( ~n1182 & n1783 ) | ( ~n1182 & n1785 ) | ( n1783 & n1785 ) ;
  assign n1787 = n973 & ~n1786 ;
  assign n1792 = n1791 ^ n1787 ^ 1'b0 ;
  assign n1793 = n1792 ^ n1084 ^ n375 ;
  assign n1794 = x46 & n1793 ;
  assign n1796 = n672 ^ n379 ^ x65 ;
  assign n1795 = ~n739 & n789 ;
  assign n1797 = n1796 ^ n1795 ^ 1'b0 ;
  assign n1798 = n1797 ^ n1055 ^ 1'b0 ;
  assign n1799 = n714 | n1442 ;
  assign n1800 = n1799 ^ n1568 ^ 1'b0 ;
  assign n1801 = x90 & n815 ;
  assign n1802 = ( n302 & n1566 ) | ( n302 & n1801 ) | ( n1566 & n1801 ) ;
  assign n1803 = n1802 ^ n425 ^ 1'b0 ;
  assign n1804 = n196 ^ x7 ^ 1'b0 ;
  assign n1805 = n1804 ^ n956 ^ x46 ;
  assign n1806 = n1516 & n1805 ;
  assign n1807 = n1282 ^ n1247 ^ n361 ;
  assign n1808 = x82 & n1058 ;
  assign n1809 = ( n685 & ~n1095 ) | ( n685 & n1743 ) | ( ~n1095 & n1743 ) ;
  assign n1810 = ( n211 & n673 ) | ( n211 & ~n1167 ) | ( n673 & ~n1167 ) ;
  assign n1811 = ( n1033 & n1551 ) | ( n1033 & ~n1810 ) | ( n1551 & ~n1810 ) ;
  assign n1812 = x96 & n1811 ;
  assign n1813 = n1809 & n1812 ;
  assign n1814 = n1384 ^ n565 ^ 1'b0 ;
  assign n1815 = n621 & n1814 ;
  assign n1816 = n1815 ^ n1203 ^ 1'b0 ;
  assign n1819 = n1184 ^ n728 ^ n241 ;
  assign n1820 = ( ~n399 & n424 ) | ( ~n399 & n1819 ) | ( n424 & n1819 ) ;
  assign n1817 = n574 ^ n136 ^ 1'b0 ;
  assign n1818 = x68 & n1817 ;
  assign n1821 = n1820 ^ n1818 ^ 1'b0 ;
  assign n1822 = ( n265 & ~n685 ) | ( n265 & n1821 ) | ( ~n685 & n1821 ) ;
  assign n1823 = n216 & n266 ;
  assign n1824 = ~n819 & n1823 ;
  assign n1826 = n1251 ^ n1032 ^ 1'b0 ;
  assign n1827 = ~n1171 & n1826 ;
  assign n1825 = x118 & n1394 ;
  assign n1828 = n1827 ^ n1825 ^ 1'b0 ;
  assign n1829 = n589 ^ n549 ^ 1'b0 ;
  assign n1830 = n1829 ^ n588 ^ x54 ;
  assign n1831 = n1647 ^ x1 ^ 1'b0 ;
  assign n1832 = ~n403 & n1831 ;
  assign n1834 = n891 ^ n369 ^ n333 ;
  assign n1833 = ( n501 & ~n856 ) | ( n501 & n1167 ) | ( ~n856 & n1167 ) ;
  assign n1835 = n1834 ^ n1833 ^ n333 ;
  assign n1838 = n899 ^ n526 ^ x48 ;
  assign n1839 = ( n992 & n1736 ) | ( n992 & n1838 ) | ( n1736 & n1838 ) ;
  assign n1837 = n1496 ^ n767 ^ n502 ;
  assign n1836 = n1409 ^ n401 ^ 1'b0 ;
  assign n1840 = n1839 ^ n1837 ^ n1836 ;
  assign n1841 = n277 ^ n194 ^ 1'b0 ;
  assign n1842 = n862 & n1841 ;
  assign n1843 = ( n669 & ~n1037 ) | ( n669 & n1842 ) | ( ~n1037 & n1842 ) ;
  assign n1844 = ~n736 & n878 ;
  assign n1845 = ~n1843 & n1844 ;
  assign n1846 = n930 ^ n752 ^ n692 ;
  assign n1847 = ~n1238 & n1846 ;
  assign n1848 = ~n626 & n1847 ;
  assign n1849 = n537 ^ n277 ^ 1'b0 ;
  assign n1850 = n393 | n1849 ;
  assign n1851 = n540 & n751 ;
  assign n1852 = n1851 ^ n569 ^ 1'b0 ;
  assign n1853 = ( ~x56 & x90 ) | ( ~x56 & n1246 ) | ( x90 & n1246 ) ;
  assign n1854 = n1853 ^ n393 ^ 1'b0 ;
  assign n1855 = n1853 | n1854 ;
  assign n1856 = ( n221 & n595 ) | ( n221 & ~n858 ) | ( n595 & ~n858 ) ;
  assign n1857 = n295 | n519 ;
  assign n1858 = n1857 ^ n469 ^ 1'b0 ;
  assign n1859 = n1858 ^ n579 ^ x23 ;
  assign n1860 = n1859 ^ n392 ^ x124 ;
  assign n1861 = n1860 ^ n1505 ^ 1'b0 ;
  assign n1862 = ( n343 & ~n1856 ) | ( n343 & n1861 ) | ( ~n1856 & n1861 ) ;
  assign n1863 = n1862 ^ n375 ^ 1'b0 ;
  assign n1864 = n1046 ^ n610 ^ 1'b0 ;
  assign n1865 = n1864 ^ n129 ^ 1'b0 ;
  assign n1866 = n1863 | n1865 ;
  assign n1867 = n1060 & n1538 ;
  assign n1870 = n647 ^ n242 ^ x51 ;
  assign n1868 = n1149 ^ n540 ^ 1'b0 ;
  assign n1869 = n1103 & n1868 ;
  assign n1871 = n1870 ^ n1869 ^ 1'b0 ;
  assign n1872 = n348 | n1871 ;
  assign n1873 = n1872 ^ n1223 ^ 1'b0 ;
  assign n1874 = n1867 & ~n1873 ;
  assign n1875 = n448 & ~n531 ;
  assign n1876 = n1875 ^ n947 ^ 1'b0 ;
  assign n1877 = x88 & ~x118 ;
  assign n1878 = n1839 & ~n1877 ;
  assign n1879 = n1878 ^ n1128 ^ 1'b0 ;
  assign n1880 = x9 & ~n314 ;
  assign n1881 = n1880 ^ n1818 ^ 1'b0 ;
  assign n1882 = n1879 & n1881 ;
  assign n1883 = n743 ^ n305 ^ 1'b0 ;
  assign n1884 = n1178 & n1883 ;
  assign n1885 = n1884 ^ n505 ^ 1'b0 ;
  assign n1886 = n441 & n1885 ;
  assign n1887 = n1131 ^ n905 ^ 1'b0 ;
  assign n1888 = n372 & n1887 ;
  assign n1889 = ~n1886 & n1888 ;
  assign n1890 = n380 ^ n275 ^ 1'b0 ;
  assign n1891 = n487 & n715 ;
  assign n1892 = n1891 ^ n1816 ^ 1'b0 ;
  assign n1893 = n1890 & n1892 ;
  assign n1894 = n794 & n1279 ;
  assign n1895 = ~n460 & n1894 ;
  assign n1896 = n1895 ^ n1538 ^ 1'b0 ;
  assign n1897 = n1896 ^ n1527 ^ n1193 ;
  assign n1898 = n1671 | n1897 ;
  assign n1899 = ( n635 & n1020 ) | ( n635 & n1229 ) | ( n1020 & n1229 ) ;
  assign n1900 = x80 & ~n1428 ;
  assign n1901 = n1899 & n1900 ;
  assign n1902 = n659 & n1901 ;
  assign n1903 = n1902 ^ n1838 ^ n354 ;
  assign n1909 = n1769 ^ n531 ^ 1'b0 ;
  assign n1904 = n239 & ~n401 ;
  assign n1905 = n714 & n1904 ;
  assign n1906 = n251 | n1905 ;
  assign n1907 = n1906 ^ n1568 ^ 1'b0 ;
  assign n1908 = x95 & ~n1907 ;
  assign n1910 = n1909 ^ n1908 ^ 1'b0 ;
  assign n1911 = n1910 ^ n1642 ^ 1'b0 ;
  assign n1912 = n1277 ^ n451 ^ 1'b0 ;
  assign n1913 = n1912 ^ n1636 ^ n915 ;
  assign n1914 = n1011 & n1220 ;
  assign n1915 = ( x66 & n738 ) | ( x66 & n916 ) | ( n738 & n916 ) ;
  assign n1916 = n1914 & ~n1915 ;
  assign n1917 = ~n160 & n357 ;
  assign n1918 = ~n815 & n1917 ;
  assign n1919 = n469 & n985 ;
  assign n1920 = n1918 & n1919 ;
  assign n1921 = n1920 ^ n1508 ^ n938 ;
  assign n1922 = ( n186 & n545 ) | ( n186 & n1644 ) | ( n545 & n1644 ) ;
  assign n1923 = ~n207 & n502 ;
  assign n1924 = n771 & ~n1923 ;
  assign n1925 = ( n820 & n1771 ) | ( n820 & n1876 ) | ( n1771 & n1876 ) ;
  assign n1926 = n1258 ^ x93 ^ 1'b0 ;
  assign n1927 = n844 | n1926 ;
  assign n1928 = n1927 ^ n730 ^ x92 ;
  assign n1929 = n1599 ^ n1212 ^ x84 ;
  assign n1930 = ( ~n237 & n953 ) | ( ~n237 & n958 ) | ( n953 & n958 ) ;
  assign n1931 = n1929 & ~n1930 ;
  assign n1932 = n1006 & n1931 ;
  assign n1936 = n216 & ~n1581 ;
  assign n1934 = x2 & ~n1673 ;
  assign n1933 = ~n533 & n1726 ;
  assign n1935 = n1934 ^ n1933 ^ 1'b0 ;
  assign n1937 = n1936 ^ n1935 ^ 1'b0 ;
  assign n1938 = n1068 | n1937 ;
  assign n1939 = n1504 ^ n346 ^ n199 ;
  assign n1940 = ( ~n285 & n1660 ) | ( ~n285 & n1939 ) | ( n1660 & n1939 ) ;
  assign n1943 = n867 ^ n454 ^ n204 ;
  assign n1944 = ( n940 & n1253 ) | ( n940 & ~n1943 ) | ( n1253 & ~n1943 ) ;
  assign n1941 = n916 | n1877 ;
  assign n1942 = n1941 ^ n965 ^ 1'b0 ;
  assign n1945 = n1944 ^ n1942 ^ 1'b0 ;
  assign n1946 = n182 | n1945 ;
  assign n1947 = n804 & n974 ;
  assign n1948 = x108 & ~n1947 ;
  assign n1949 = n1948 ^ n1538 ^ 1'b0 ;
  assign n1950 = n1949 ^ n761 ^ 1'b0 ;
  assign n1951 = n1946 | n1950 ;
  assign n1954 = ( n565 & n926 ) | ( n565 & n1822 ) | ( n926 & n1822 ) ;
  assign n1952 = n1311 ^ n1001 ^ n582 ;
  assign n1953 = ~n1754 & n1952 ;
  assign n1955 = n1954 ^ n1953 ^ 1'b0 ;
  assign n1956 = n1176 & n1348 ;
  assign n1957 = n1956 ^ n1846 ^ 1'b0 ;
  assign n1958 = n1957 ^ x97 ^ 1'b0 ;
  assign n1959 = n366 & ~n1958 ;
  assign n1960 = n149 & n1959 ;
  assign n1961 = n1960 ^ n1930 ^ 1'b0 ;
  assign n1965 = x26 & n949 ;
  assign n1966 = ~n398 & n1965 ;
  assign n1962 = n376 & ~n1663 ;
  assign n1963 = ~n804 & n1962 ;
  assign n1964 = n1963 ^ n1279 ^ 1'b0 ;
  assign n1967 = n1966 ^ n1964 ^ 1'b0 ;
  assign n1968 = n266 & ~n1967 ;
  assign n1969 = n1527 ^ n531 ^ 1'b0 ;
  assign n1973 = n598 ^ n535 ^ 1'b0 ;
  assign n1972 = x30 & ~x37 ;
  assign n1970 = n1226 ^ n316 ^ 1'b0 ;
  assign n1971 = ( x83 & ~n625 ) | ( x83 & n1970 ) | ( ~n625 & n1970 ) ;
  assign n1974 = n1973 ^ n1972 ^ n1971 ;
  assign n1976 = ( ~n199 & n830 ) | ( ~n199 & n1411 ) | ( n830 & n1411 ) ;
  assign n1977 = n661 & n1976 ;
  assign n1975 = n1001 ^ n798 ^ x118 ;
  assign n1978 = n1977 ^ n1975 ^ x87 ;
  assign n1979 = n996 & ~n1523 ;
  assign n1980 = n1707 ^ n1187 ^ n149 ;
  assign n1984 = n827 ^ n403 ^ x83 ;
  assign n1985 = n1203 | n1984 ;
  assign n1986 = n699 | n1985 ;
  assign n1981 = n1476 ^ n1220 ^ 1'b0 ;
  assign n1982 = n920 & n1981 ;
  assign n1983 = ~n232 & n1982 ;
  assign n1987 = n1986 ^ n1983 ^ 1'b0 ;
  assign n1988 = n460 | n1542 ;
  assign n1989 = n1987 & ~n1988 ;
  assign n1990 = ( n320 & n1980 ) | ( n320 & ~n1989 ) | ( n1980 & ~n1989 ) ;
  assign n1991 = n938 & n1829 ;
  assign n1992 = n1991 ^ n455 ^ 1'b0 ;
  assign n1993 = ( x59 & ~x93 ) | ( x59 & n363 ) | ( ~x93 & n363 ) ;
  assign n1994 = ( n432 & n445 ) | ( n432 & n1993 ) | ( n445 & n1993 ) ;
  assign n1995 = n1994 ^ n806 ^ 1'b0 ;
  assign n1996 = x60 & n1995 ;
  assign n1997 = n1289 & n1996 ;
  assign n1998 = ~n1912 & n1997 ;
  assign n1999 = n1998 ^ n1016 ^ n487 ;
  assign n2000 = n1999 ^ n1833 ^ n1829 ;
  assign n2001 = n829 & n1164 ;
  assign n2002 = n2001 ^ n1779 ^ 1'b0 ;
  assign n2003 = ~n1203 & n2002 ;
  assign n2004 = ( ~n1490 & n1508 ) | ( ~n1490 & n2003 ) | ( n1508 & n2003 ) ;
  assign n2005 = n209 & n1125 ;
  assign n2006 = n1620 & n2005 ;
  assign n2007 = n2006 ^ n826 ^ 1'b0 ;
  assign n2008 = n1625 ^ n294 ^ 1'b0 ;
  assign n2009 = n1110 | n2008 ;
  assign n2010 = n147 & ~n401 ;
  assign n2011 = ( n348 & n2009 ) | ( n348 & n2010 ) | ( n2009 & n2010 ) ;
  assign n2012 = ~n432 & n2011 ;
  assign n2013 = n2012 ^ n607 ^ 1'b0 ;
  assign n2014 = n1469 ^ n798 ^ n434 ;
  assign n2015 = n1278 & ~n1870 ;
  assign n2016 = n2014 & n2015 ;
  assign n2017 = n2016 ^ x3 ^ 1'b0 ;
  assign n2018 = n707 & ~n2017 ;
  assign n2019 = n349 & n1697 ;
  assign n2020 = n2019 ^ n1668 ^ n1309 ;
  assign n2021 = n1581 ^ n1168 ^ 1'b0 ;
  assign n2022 = n1499 & ~n2021 ;
  assign n2023 = n771 ^ n207 ^ 1'b0 ;
  assign n2024 = ~n153 & n2015 ;
  assign n2025 = n1205 & n2024 ;
  assign n2026 = n479 ^ n465 ^ 1'b0 ;
  assign n2027 = ~n776 & n2026 ;
  assign n2028 = n1283 ^ n668 ^ 1'b0 ;
  assign n2029 = n2027 & n2028 ;
  assign n2030 = n783 | n2029 ;
  assign n2031 = n2030 ^ n1959 ^ 1'b0 ;
  assign n2032 = n848 | n1296 ;
  assign n2033 = n2032 ^ n1346 ^ 1'b0 ;
  assign n2034 = n888 & n2033 ;
  assign n2035 = n2034 ^ n887 ^ 1'b0 ;
  assign n2036 = ( x93 & n824 ) | ( x93 & n1834 ) | ( n824 & n1834 ) ;
  assign n2041 = ( ~n895 & n1203 ) | ( ~n895 & n1490 ) | ( n1203 & n1490 ) ;
  assign n2037 = x40 ^ x0 ^ 1'b0 ;
  assign n2038 = n656 & n2037 ;
  assign n2039 = n1805 ^ n952 ^ n396 ;
  assign n2040 = n2038 & n2039 ;
  assign n2042 = n2041 ^ n2040 ^ 1'b0 ;
  assign n2043 = n1600 ^ n935 ^ 1'b0 ;
  assign n2044 = ( x94 & n1411 ) | ( x94 & ~n2043 ) | ( n1411 & ~n2043 ) ;
  assign n2045 = n1579 & n1976 ;
  assign n2046 = n2045 ^ n221 ^ 1'b0 ;
  assign n2047 = ( ~n293 & n383 ) | ( ~n293 & n1002 ) | ( n383 & n1002 ) ;
  assign n2048 = n2047 ^ n724 ^ 1'b0 ;
  assign n2049 = n171 & n1837 ;
  assign n2050 = n2049 ^ n274 ^ 1'b0 ;
  assign n2051 = n2050 ^ n1032 ^ n550 ;
  assign n2052 = n334 & ~n522 ;
  assign n2053 = n1753 & n2052 ;
  assign n2054 = n237 ^ n155 ^ 1'b0 ;
  assign n2055 = ~n971 & n2054 ;
  assign n2056 = x0 | n190 ;
  assign n2057 = ( n157 & n746 ) | ( n157 & n2056 ) | ( n746 & n2056 ) ;
  assign n2058 = n2057 ^ n1769 ^ x1 ;
  assign n2059 = ( n1280 & n2055 ) | ( n1280 & ~n2058 ) | ( n2055 & ~n2058 ) ;
  assign n2060 = n1107 ^ n713 ^ 1'b0 ;
  assign n2061 = n295 & n723 ;
  assign n2062 = n2061 ^ x24 ^ 1'b0 ;
  assign n2063 = n452 ^ n242 ^ 1'b0 ;
  assign n2064 = ~n2062 & n2063 ;
  assign n2065 = n2060 & n2064 ;
  assign n2066 = ~n230 & n365 ;
  assign n2067 = n848 & n2066 ;
  assign n2068 = n2067 ^ n2060 ^ 1'b0 ;
  assign n2069 = ~n2065 & n2068 ;
  assign n2070 = n1003 & ~n1910 ;
  assign n2071 = ( ~n390 & n1918 ) | ( ~n390 & n2070 ) | ( n1918 & n2070 ) ;
  assign n2072 = n1253 ^ x2 ^ 1'b0 ;
  assign n2073 = x37 & n2072 ;
  assign n2074 = n2073 ^ n1520 ^ 1'b0 ;
  assign n2075 = n2061 ^ n1108 ^ 1'b0 ;
  assign n2076 = x69 & n2075 ;
  assign n2084 = n178 & n979 ;
  assign n2085 = ~n1805 & n2084 ;
  assign n2086 = ( x25 & ~n1579 ) | ( x25 & n2085 ) | ( ~n1579 & n2085 ) ;
  assign n2087 = n1054 | n2086 ;
  assign n2081 = n1411 ^ n194 ^ 1'b0 ;
  assign n2077 = ( x54 & n257 ) | ( x54 & ~n260 ) | ( n257 & ~n260 ) ;
  assign n2078 = n2077 ^ n555 ^ 1'b0 ;
  assign n2079 = n1311 | n2078 ;
  assign n2080 = n1022 & ~n2079 ;
  assign n2082 = n2081 ^ n2080 ^ 1'b0 ;
  assign n2083 = n2082 ^ n1075 ^ n415 ;
  assign n2088 = n2087 ^ n2083 ^ 1'b0 ;
  assign n2094 = x124 ^ x72 ^ 1'b0 ;
  assign n2095 = ~n198 & n2094 ;
  assign n2090 = n599 ^ n434 ^ n366 ;
  assign n2091 = n1306 & n2090 ;
  assign n2092 = n497 & n2091 ;
  assign n2089 = x71 & ~n1235 ;
  assign n2093 = n2092 ^ n2089 ^ 1'b0 ;
  assign n2096 = n2095 ^ n2093 ^ n471 ;
  assign n2097 = n168 | n615 ;
  assign n2098 = n1025 ^ n202 ^ n171 ;
  assign n2099 = x10 & n2098 ;
  assign n2100 = ~n590 & n2099 ;
  assign n2101 = n2100 ^ n936 ^ n419 ;
  assign n2102 = n2101 ^ n752 ^ 1'b0 ;
  assign n2103 = ~x94 & n1415 ;
  assign n2104 = ~n2102 & n2103 ;
  assign n2105 = n2104 ^ n1365 ^ 1'b0 ;
  assign n2106 = n2097 & n2105 ;
  assign n2107 = n2096 | n2106 ;
  assign n2108 = n1586 ^ n1504 ^ n958 ;
  assign n2109 = ~n165 & n182 ;
  assign n2110 = ~n908 & n2109 ;
  assign n2111 = ( x78 & ~n462 ) | ( x78 & n2110 ) | ( ~n462 & n2110 ) ;
  assign n2112 = ( n654 & ~n1352 ) | ( n654 & n2111 ) | ( ~n1352 & n2111 ) ;
  assign n2113 = n2112 ^ n851 ^ x29 ;
  assign n2114 = x18 & ~n824 ;
  assign n2115 = ( n1219 & ~n1458 ) | ( n1219 & n2114 ) | ( ~n1458 & n2114 ) ;
  assign n2116 = ( ~n958 & n1286 ) | ( ~n958 & n2079 ) | ( n1286 & n2079 ) ;
  assign n2117 = n1697 | n2116 ;
  assign n2118 = n1097 | n2117 ;
  assign n2119 = n856 ^ n620 ^ 1'b0 ;
  assign n2123 = n1686 ^ n1592 ^ 1'b0 ;
  assign n2124 = ~n1184 & n2123 ;
  assign n2125 = n2124 ^ n841 ^ n421 ;
  assign n2120 = n412 & ~n899 ;
  assign n2121 = ~n298 & n2120 ;
  assign n2122 = ( ~x62 & n701 ) | ( ~x62 & n2121 ) | ( n701 & n2121 ) ;
  assign n2126 = n2125 ^ n2122 ^ 1'b0 ;
  assign n2127 = n2119 | n2126 ;
  assign n2128 = x95 & n227 ;
  assign n2129 = n2128 ^ x69 ^ 1'b0 ;
  assign n2130 = n129 & ~n388 ;
  assign n2131 = ( n557 & n936 ) | ( n557 & ~n2130 ) | ( n936 & ~n2130 ) ;
  assign n2132 = n2129 | n2131 ;
  assign n2135 = n420 & n989 ;
  assign n2136 = ~n834 & n2135 ;
  assign n2133 = n500 & ~n1533 ;
  assign n2134 = n2133 ^ n1296 ^ 1'b0 ;
  assign n2137 = n2136 ^ n2134 ^ 1'b0 ;
  assign n2138 = n1576 & ~n2137 ;
  assign n2139 = n1184 ^ n584 ^ n319 ;
  assign n2140 = n2139 ^ n2059 ^ n1643 ;
  assign n2141 = ~n1548 & n1561 ;
  assign n2142 = n1579 & n1914 ;
  assign n2143 = ( n219 & ~n310 ) | ( n219 & n357 ) | ( ~n310 & n357 ) ;
  assign n2144 = x64 & ~n2143 ;
  assign n2145 = n2144 ^ n319 ^ 1'b0 ;
  assign n2146 = ( n1879 & ~n2090 ) | ( n1879 & n2145 ) | ( ~n2090 & n2145 ) ;
  assign n2147 = n2125 ^ n942 ^ 1'b0 ;
  assign n2148 = n850 ^ x124 ^ 1'b0 ;
  assign n2149 = n213 & ~n2148 ;
  assign n2150 = n2149 ^ n415 ^ 1'b0 ;
  assign n2151 = n1585 ^ n681 ^ x126 ;
  assign n2152 = ( n851 & n1730 ) | ( n851 & n2151 ) | ( n1730 & n2151 ) ;
  assign n2153 = ( n1076 & n2150 ) | ( n1076 & ~n2152 ) | ( n2150 & ~n2152 ) ;
  assign n2164 = n1157 & ~n1230 ;
  assign n2165 = n2164 ^ n160 ^ 1'b0 ;
  assign n2166 = n2165 ^ n245 ^ x74 ;
  assign n2159 = n269 ^ x83 ^ 1'b0 ;
  assign n2160 = n305 & n2159 ;
  assign n2161 = ( n442 & n1733 ) | ( n442 & n2160 ) | ( n1733 & n2160 ) ;
  assign n2154 = n460 ^ n403 ^ 1'b0 ;
  assign n2155 = x93 & n1673 ;
  assign n2156 = ~n2154 & n2155 ;
  assign n2157 = n2156 ^ n198 ^ x118 ;
  assign n2158 = n1993 | n2157 ;
  assign n2162 = n2161 ^ n2158 ^ 1'b0 ;
  assign n2163 = ( n550 & ~n1896 ) | ( n550 & n2162 ) | ( ~n1896 & n2162 ) ;
  assign n2167 = n2166 ^ n2163 ^ n1379 ;
  assign n2168 = n491 ^ x80 ^ 1'b0 ;
  assign n2169 = ~n1240 & n2168 ;
  assign n2170 = n2169 ^ n838 ^ 1'b0 ;
  assign n2171 = n2038 ^ n180 ^ 1'b0 ;
  assign n2172 = ~n517 & n2171 ;
  assign n2173 = ( n826 & n2092 ) | ( n826 & n2172 ) | ( n2092 & n2172 ) ;
  assign n2174 = ( n1055 & n2170 ) | ( n1055 & n2173 ) | ( n2170 & n2173 ) ;
  assign n2175 = n1365 ^ n1227 ^ n279 ;
  assign n2176 = n940 ^ x2 ^ 1'b0 ;
  assign n2177 = n2175 & ~n2176 ;
  assign n2178 = n628 ^ n390 ^ n216 ;
  assign n2179 = ~n322 & n2178 ;
  assign n2180 = n1566 & n2179 ;
  assign n2181 = n1526 ^ n996 ^ n740 ;
  assign n2182 = n838 ^ n174 ^ 1'b0 ;
  assign n2183 = ~n218 & n1986 ;
  assign n2184 = n2183 ^ n2121 ^ 1'b0 ;
  assign n2185 = n914 ^ n198 ^ 1'b0 ;
  assign n2186 = n1534 & n2185 ;
  assign n2187 = ~x46 & n1389 ;
  assign n2188 = ~n1076 & n2187 ;
  assign n2189 = ~n227 & n420 ;
  assign n2190 = n2189 ^ n1382 ^ n1007 ;
  assign n2191 = n2190 ^ n1697 ^ x57 ;
  assign n2192 = n1152 ^ x90 ^ 1'b0 ;
  assign n2193 = x94 & n983 ;
  assign n2194 = n2193 ^ n281 ^ 1'b0 ;
  assign n2195 = ( n1053 & ~n2179 ) | ( n1053 & n2194 ) | ( ~n2179 & n2194 ) ;
  assign n2198 = ~n266 & n375 ;
  assign n2199 = ( n379 & n1517 ) | ( n379 & ~n2198 ) | ( n1517 & ~n2198 ) ;
  assign n2196 = n1673 & n1801 ;
  assign n2197 = n1006 & n2196 ;
  assign n2200 = n2199 ^ n2197 ^ 1'b0 ;
  assign n2201 = n699 ^ n190 ^ 1'b0 ;
  assign n2202 = n314 | n2201 ;
  assign n2203 = n2202 ^ n1527 ^ 1'b0 ;
  assign n2204 = n206 | n2203 ;
  assign n2205 = n2204 ^ n2175 ^ x86 ;
  assign n2206 = n1182 ^ n631 ^ 1'b0 ;
  assign n2207 = ~n572 & n2206 ;
  assign n2208 = n1896 ^ n1246 ^ 1'b0 ;
  assign n2209 = n603 & n2208 ;
  assign n2210 = ~n2131 & n2209 ;
  assign n2211 = n2207 & n2210 ;
  assign n2212 = n205 | n867 ;
  assign n2213 = n2212 ^ n442 ^ n205 ;
  assign n2215 = n1208 ^ n849 ^ 1'b0 ;
  assign n2214 = n367 & n1104 ;
  assign n2216 = n2215 ^ n2214 ^ 1'b0 ;
  assign n2217 = n1687 | n2216 ;
  assign n2218 = n2217 ^ n1175 ^ 1'b0 ;
  assign n2219 = n2006 | n2218 ;
  assign n2220 = ( x63 & ~n862 ) | ( x63 & n2219 ) | ( ~n862 & n2219 ) ;
  assign n2221 = x19 & ~n1294 ;
  assign n2222 = n2221 ^ n2170 ^ 1'b0 ;
  assign n2223 = n1147 ^ n706 ^ x51 ;
  assign n2224 = ( ~x115 & n758 ) | ( ~x115 & n1446 ) | ( n758 & n1446 ) ;
  assign n2225 = ( n575 & n826 ) | ( n575 & n2224 ) | ( n826 & n2224 ) ;
  assign n2227 = ( x119 & n1381 ) | ( x119 & ~n1769 ) | ( n1381 & ~n1769 ) ;
  assign n2228 = ( n1972 & ~n1996 ) | ( n1972 & n2227 ) | ( ~n1996 & n2227 ) ;
  assign n2226 = n210 | n1986 ;
  assign n2229 = n2228 ^ n2226 ^ 1'b0 ;
  assign n2230 = n1402 ^ n1024 ^ 1'b0 ;
  assign n2231 = n1596 | n2230 ;
  assign n2232 = n1441 | n1649 ;
  assign n2233 = n850 & n2232 ;
  assign n2234 = n1697 ^ n1096 ^ 1'b0 ;
  assign n2235 = ~n1885 & n2234 ;
  assign n2239 = ( n373 & ~n531 ) | ( n373 & n549 ) | ( ~n531 & n549 ) ;
  assign n2240 = n318 & n2239 ;
  assign n2241 = ~n1725 & n2240 ;
  assign n2242 = ~n1377 & n2241 ;
  assign n2236 = n2092 ^ n608 ^ 1'b0 ;
  assign n2237 = x85 & ~n2236 ;
  assign n2238 = n2172 & n2237 ;
  assign n2243 = n2242 ^ n2238 ^ 1'b0 ;
  assign n2244 = n771 & ~n1801 ;
  assign n2245 = n888 & ~n1400 ;
  assign n2246 = n2245 ^ n996 ^ 1'b0 ;
  assign n2247 = n2246 ^ n1171 ^ n219 ;
  assign n2250 = n457 ^ x15 ^ 1'b0 ;
  assign n2251 = n549 & ~n2250 ;
  assign n2252 = n2251 ^ n378 ^ n320 ;
  assign n2253 = n2252 ^ n149 ^ x52 ;
  assign n2248 = n485 ^ x58 ^ 1'b0 ;
  assign n2249 = n961 & ~n2248 ;
  assign n2254 = n2253 ^ n2249 ^ 1'b0 ;
  assign n2256 = n143 & ~n529 ;
  assign n2257 = ~n213 & n2256 ;
  assign n2258 = n406 & ~n1243 ;
  assign n2259 = ~n998 & n2258 ;
  assign n2260 = n2259 ^ n167 ^ 1'b0 ;
  assign n2261 = n2257 | n2260 ;
  assign n2255 = n813 & ~n1776 ;
  assign n2262 = n2261 ^ n2255 ^ n1753 ;
  assign n2263 = n1232 ^ n550 ^ 1'b0 ;
  assign n2264 = n2263 ^ n1689 ^ n625 ;
  assign n2265 = ( n595 & n977 ) | ( n595 & ~n1590 ) | ( n977 & ~n1590 ) ;
  assign n2266 = n577 ^ n167 ^ 1'b0 ;
  assign n2267 = n471 | n2266 ;
  assign n2268 = n767 | n2267 ;
  assign n2269 = n1611 | n2268 ;
  assign n2270 = n2269 ^ n693 ^ 1'b0 ;
  assign n2271 = n2265 & n2270 ;
  assign n2272 = ( n2262 & n2264 ) | ( n2262 & n2271 ) | ( n2264 & n2271 ) ;
  assign n2273 = x116 ^ x100 ^ 1'b0 ;
  assign n2274 = ( n683 & n1996 ) | ( n683 & n2273 ) | ( n1996 & n2273 ) ;
  assign n2275 = n2274 ^ n1040 ^ 1'b0 ;
  assign n2276 = n2275 ^ n468 ^ 1'b0 ;
  assign n2277 = n456 | n2276 ;
  assign n2278 = n2277 ^ n779 ^ 1'b0 ;
  assign n2279 = n2278 ^ n218 ^ x8 ;
  assign n2280 = n222 ^ x24 ^ 1'b0 ;
  assign n2281 = n2280 ^ n948 ^ 1'b0 ;
  assign n2282 = n2281 ^ n550 ^ 1'b0 ;
  assign n2283 = n214 ^ n206 ^ n171 ;
  assign n2284 = ( n550 & n989 ) | ( n550 & ~n1796 ) | ( n989 & ~n1796 ) ;
  assign n2285 = n2284 ^ n1354 ^ 1'b0 ;
  assign n2286 = ( x125 & ~n2283 ) | ( x125 & n2285 ) | ( ~n2283 & n2285 ) ;
  assign n2287 = n464 & n1538 ;
  assign n2288 = ~n2232 & n2287 ;
  assign n2289 = ( x100 & n1399 ) | ( x100 & ~n2288 ) | ( n1399 & ~n2288 ) ;
  assign n2295 = n952 ^ n611 ^ x15 ;
  assign n2296 = ( n190 & ~n401 ) | ( n190 & n2295 ) | ( ~n401 & n2295 ) ;
  assign n2297 = ( ~n429 & n715 ) | ( ~n429 & n2296 ) | ( n715 & n2296 ) ;
  assign n2298 = n2297 ^ n914 ^ x108 ;
  assign n2293 = ( n169 & ~n451 ) | ( n169 & n483 ) | ( ~n451 & n483 ) ;
  assign n2291 = n2206 ^ n1202 ^ 1'b0 ;
  assign n2292 = n866 & ~n2291 ;
  assign n2294 = n2293 ^ n2292 ^ x81 ;
  assign n2290 = n447 | n1858 ;
  assign n2299 = n2298 ^ n2294 ^ n2290 ;
  assign n2300 = n885 | n1974 ;
  assign n2301 = n1196 & n1285 ;
  assign n2302 = ( ~x77 & n238 ) | ( ~x77 & n1019 ) | ( n238 & n1019 ) ;
  assign n2303 = n971 | n2198 ;
  assign n2304 = ( x26 & n845 ) | ( x26 & n2303 ) | ( n845 & n2303 ) ;
  assign n2305 = ~n754 & n1894 ;
  assign n2306 = n1726 & ~n2305 ;
  assign n2307 = n2304 & n2306 ;
  assign n2308 = ( n608 & n1418 ) | ( n608 & ~n2307 ) | ( n1418 & ~n2307 ) ;
  assign n2309 = n2308 ^ n802 ^ n798 ;
  assign n2310 = n260 | n2309 ;
  assign n2311 = ( n945 & n2302 ) | ( n945 & ~n2310 ) | ( n2302 & ~n2310 ) ;
  assign n2312 = n1156 ^ n425 ^ 1'b0 ;
  assign n2313 = n1175 & ~n2312 ;
  assign n2314 = n2313 ^ n134 ^ 1'b0 ;
  assign n2315 = n837 | n2314 ;
  assign n2316 = n2315 ^ n1314 ^ n197 ;
  assign n2317 = n332 ^ n198 ^ 1'b0 ;
  assign n2318 = n1079 | n2317 ;
  assign n2319 = n844 & ~n2318 ;
  assign n2320 = n443 | n1020 ;
  assign n2321 = n2320 ^ n436 ^ 1'b0 ;
  assign n2322 = n1198 & n2321 ;
  assign n2323 = x23 | n1020 ;
  assign n2324 = n1462 | n2323 ;
  assign n2325 = ~n1715 & n2324 ;
  assign n2326 = ~n871 & n2246 ;
  assign n2327 = n2325 & ~n2326 ;
  assign n2328 = ~n2322 & n2327 ;
  assign n2329 = n2319 & ~n2328 ;
  assign n2330 = n381 | n1989 ;
  assign n2331 = n2330 ^ n2178 ^ 1'b0 ;
  assign n2332 = ~n164 & n1226 ;
  assign n2333 = n2332 ^ x46 ^ 1'b0 ;
  assign n2334 = x50 & n2333 ;
  assign n2335 = ~n2331 & n2334 ;
  assign n2336 = ( n775 & n889 ) | ( n775 & n967 ) | ( n889 & n967 ) ;
  assign n2337 = ( x60 & n1504 ) | ( x60 & n2336 ) | ( n1504 & n2336 ) ;
  assign n2338 = n1206 | n1280 ;
  assign n2339 = n2338 ^ n1079 ^ n522 ;
  assign n2340 = n1624 ^ n972 ^ 1'b0 ;
  assign n2341 = n291 | n1976 ;
  assign n2342 = n2340 | n2341 ;
  assign n2343 = n2342 ^ x32 ^ 1'b0 ;
  assign n2344 = ~n1349 & n2343 ;
  assign n2345 = ( n597 & n646 ) | ( n597 & ~n2257 ) | ( n646 & ~n2257 ) ;
  assign n2346 = n2179 ^ n714 ^ 1'b0 ;
  assign n2347 = n2346 ^ n1017 ^ n265 ;
  assign n2348 = ( x90 & n2345 ) | ( x90 & ~n2347 ) | ( n2345 & ~n2347 ) ;
  assign n2349 = n1135 ^ n522 ^ 1'b0 ;
  assign n2350 = ~n1451 & n2349 ;
  assign n2351 = n2350 ^ n1827 ^ 1'b0 ;
  assign n2352 = n506 | n2351 ;
  assign n2353 = ~n1105 & n1671 ;
  assign n2354 = n1314 | n2154 ;
  assign n2355 = ~n1037 & n2354 ;
  assign n2356 = n2355 ^ n171 ^ 1'b0 ;
  assign n2358 = n595 & ~n1214 ;
  assign n2359 = n2358 ^ n1776 ^ 1'b0 ;
  assign n2357 = ~n1853 & n2165 ;
  assign n2360 = n2359 ^ n2357 ^ 1'b0 ;
  assign n2361 = ( n505 & ~n2299 ) | ( n505 & n2360 ) | ( ~n2299 & n2360 ) ;
  assign n2362 = n1168 ^ n134 ^ 1'b0 ;
  assign n2363 = n632 & n2362 ;
  assign n2364 = n434 | n2363 ;
  assign n2365 = ~n964 & n2154 ;
  assign n2366 = n633 & ~n2365 ;
  assign n2367 = n841 | n2366 ;
  assign n2368 = n2367 ^ n958 ^ 1'b0 ;
  assign n2369 = n982 ^ x95 ^ 1'b0 ;
  assign n2370 = n1797 ^ n1740 ^ 1'b0 ;
  assign n2371 = n383 & ~n402 ;
  assign n2372 = n791 | n2371 ;
  assign n2373 = ( n989 & n1639 ) | ( n989 & n2372 ) | ( n1639 & n2372 ) ;
  assign n2374 = n1314 ^ n418 ^ 1'b0 ;
  assign n2375 = ~n241 & n2374 ;
  assign n2376 = n2172 ^ n1574 ^ 1'b0 ;
  assign n2377 = ( x37 & n554 ) | ( x37 & n1057 ) | ( n554 & n1057 ) ;
  assign n2378 = ( ~n178 & n2376 ) | ( ~n178 & n2377 ) | ( n2376 & n2377 ) ;
  assign n2379 = x84 & n881 ;
  assign n2380 = n2378 & n2379 ;
  assign n2381 = ( x59 & ~x123 ) | ( x59 & n291 ) | ( ~x123 & n291 ) ;
  assign n2382 = n2381 ^ n380 ^ 1'b0 ;
  assign n2383 = n1251 & ~n2382 ;
  assign n2384 = x53 & n398 ;
  assign n2385 = ~n2383 & n2384 ;
  assign n2386 = n2027 ^ n738 ^ n556 ;
  assign n2387 = n2386 ^ n1611 ^ n1383 ;
  assign n2388 = n949 & ~n1056 ;
  assign n2389 = n1060 & n2388 ;
  assign n2390 = ( n2385 & n2387 ) | ( n2385 & ~n2389 ) | ( n2387 & ~n2389 ) ;
  assign n2391 = n2390 ^ n197 ^ 1'b0 ;
  assign n2393 = n476 ^ x125 ^ 1'b0 ;
  assign n2394 = x108 & ~n2393 ;
  assign n2395 = n339 & ~n1100 ;
  assign n2396 = ~n773 & n2395 ;
  assign n2397 = n685 ^ n519 ^ 1'b0 ;
  assign n2398 = ~n2396 & n2397 ;
  assign n2399 = ( n1089 & ~n2394 ) | ( n1089 & n2398 ) | ( ~n2394 & n2398 ) ;
  assign n2392 = n2082 | n2147 ;
  assign n2400 = n2399 ^ n2392 ^ 1'b0 ;
  assign n2401 = n2139 ^ n262 ^ 1'b0 ;
  assign n2402 = ( n424 & n1280 ) | ( n424 & ~n1314 ) | ( n1280 & ~n1314 ) ;
  assign n2403 = ~n1272 & n2402 ;
  assign n2404 = n1073 & n2403 ;
  assign n2405 = n2404 ^ n490 ^ 1'b0 ;
  assign n2406 = n131 & ~n2405 ;
  assign n2407 = x93 | n1624 ;
  assign n2408 = n2407 ^ n1277 ^ 1'b0 ;
  assign n2409 = ( n488 & n1654 ) | ( n488 & n2317 ) | ( n1654 & n2317 ) ;
  assign n2410 = ~n559 & n1634 ;
  assign n2411 = n2410 ^ n592 ^ 1'b0 ;
  assign n2412 = n228 | n1976 ;
  assign n2413 = n874 & ~n2412 ;
  assign n2414 = n2413 ^ x123 ^ 1'b0 ;
  assign n2415 = n2411 & ~n2414 ;
  assign n2420 = n1813 ^ n577 ^ 1'b0 ;
  assign n2416 = n1617 | n2386 ;
  assign n2417 = n2416 ^ n1396 ^ 1'b0 ;
  assign n2418 = n373 ^ x89 ^ x39 ;
  assign n2419 = ( x115 & n2417 ) | ( x115 & n2418 ) | ( n2417 & n2418 ) ;
  assign n2421 = n2420 ^ n2419 ^ n1223 ;
  assign n2422 = n2421 ^ n1927 ^ n160 ;
  assign n2423 = n2309 ^ x2 ^ 1'b0 ;
  assign n2424 = x1 & ~n1023 ;
  assign n2425 = n1670 & n2424 ;
  assign n2426 = n2423 & ~n2425 ;
  assign n2427 = n1063 | n1240 ;
  assign n2428 = n2427 ^ n1818 ^ 1'b0 ;
  assign n2429 = n1859 & ~n2428 ;
  assign n2430 = n2429 ^ n1449 ^ n776 ;
  assign n2431 = n1754 ^ x94 ^ 1'b0 ;
  assign n2432 = n1088 | n2431 ;
  assign n2433 = n2432 ^ n375 ^ 1'b0 ;
  assign n2434 = ( n838 & n848 ) | ( n838 & ~n1076 ) | ( n848 & ~n1076 ) ;
  assign n2435 = ~n165 & n2342 ;
  assign n2436 = n1020 & n2435 ;
  assign n2437 = n1160 & ~n2436 ;
  assign n2438 = ~n2434 & n2437 ;
  assign n2439 = n1018 ^ x16 ^ 1'b0 ;
  assign n2440 = n366 | n2439 ;
  assign n2441 = n1639 & ~n2440 ;
  assign n2442 = n891 ^ n442 ^ 1'b0 ;
  assign n2443 = n2442 ^ n831 ^ 1'b0 ;
  assign n2444 = n696 | n2443 ;
  assign n2445 = n1458 | n1517 ;
  assign n2446 = n538 ^ x105 ^ 1'b0 ;
  assign n2447 = n952 & n2446 ;
  assign n2448 = n583 & n2447 ;
  assign n2449 = n2448 ^ n1523 ^ 1'b0 ;
  assign n2450 = ( ~n987 & n1720 ) | ( ~n987 & n2274 ) | ( n1720 & n2274 ) ;
  assign n2451 = n2450 ^ n2413 ^ n1190 ;
  assign n2453 = ( x61 & ~n227 ) | ( x61 & n1276 ) | ( ~n227 & n1276 ) ;
  assign n2452 = n807 & ~n1108 ;
  assign n2454 = n2453 ^ n2452 ^ n474 ;
  assign n2455 = x56 & n1450 ;
  assign n2456 = n2455 ^ n1827 ^ 1'b0 ;
  assign n2457 = n285 & ~n2456 ;
  assign n2458 = ( n617 & n903 ) | ( n617 & ~n1443 ) | ( n903 & ~n1443 ) ;
  assign n2459 = ( n487 & ~n1125 ) | ( n487 & n2045 ) | ( ~n1125 & n2045 ) ;
  assign n2460 = n808 & n893 ;
  assign n2461 = n2460 ^ n2232 ^ 1'b0 ;
  assign n2462 = n848 | n2461 ;
  assign n2463 = ~n2459 & n2462 ;
  assign n2464 = n961 & ~n1090 ;
  assign n2465 = n649 & n2464 ;
  assign n2466 = ( n487 & n1411 ) | ( n487 & n2465 ) | ( n1411 & n2465 ) ;
  assign n2467 = n1299 & n2466 ;
  assign n2468 = n1562 ^ n390 ^ x55 ;
  assign n2469 = n2295 ^ n1621 ^ 1'b0 ;
  assign n2470 = ( ~n323 & n2468 ) | ( ~n323 & n2469 ) | ( n2468 & n2469 ) ;
  assign n2471 = n1437 & n1966 ;
  assign n2472 = n2471 ^ n1556 ^ 1'b0 ;
  assign n2473 = n2472 ^ n1912 ^ x7 ;
  assign n2474 = n1476 & n2473 ;
  assign n2475 = n2474 ^ n1433 ^ 1'b0 ;
  assign n2476 = n1218 ^ n529 ^ n151 ;
  assign n2485 = n841 ^ n264 ^ x11 ;
  assign n2477 = x85 & ~n1656 ;
  assign n2478 = ~n761 & n2477 ;
  assign n2479 = n1009 & n1319 ;
  assign n2480 = n2479 ^ n829 ^ 1'b0 ;
  assign n2481 = n2480 ^ n2129 ^ 1'b0 ;
  assign n2482 = n2481 ^ n171 ^ 1'b0 ;
  assign n2483 = ~n2478 & n2482 ;
  assign n2484 = n2274 & n2483 ;
  assign n2486 = n2485 ^ n2484 ^ 1'b0 ;
  assign n2487 = n1187 & ~n2119 ;
  assign n2489 = n575 & n1765 ;
  assign n2488 = ~n1149 & n2369 ;
  assign n2490 = n2489 ^ n2488 ^ 1'b0 ;
  assign n2491 = n777 ^ n742 ^ x31 ;
  assign n2492 = n301 & n2491 ;
  assign n2493 = ~n1472 & n2492 ;
  assign n2494 = ( x115 & n1278 ) | ( x115 & n2493 ) | ( n1278 & n2493 ) ;
  assign n2495 = ( n779 & n1673 ) | ( n779 & n2494 ) | ( n1673 & n2494 ) ;
  assign n2496 = ~n2177 & n2495 ;
  assign n2497 = ( x112 & n432 ) | ( x112 & ~n681 ) | ( n432 & ~n681 ) ;
  assign n2498 = n2497 ^ n1602 ^ n895 ;
  assign n2505 = ~n618 & n694 ;
  assign n2506 = x68 & n1641 ;
  assign n2507 = n2506 ^ n393 ^ 1'b0 ;
  assign n2508 = ( n204 & n2505 ) | ( n204 & n2507 ) | ( n2505 & n2507 ) ;
  assign n2504 = n269 & n1686 ;
  assign n2499 = ( n462 & n691 ) | ( n462 & n1587 ) | ( n691 & n1587 ) ;
  assign n2500 = n1526 & ~n2499 ;
  assign n2501 = n2500 ^ n199 ^ 1'b0 ;
  assign n2502 = n2501 ^ n1954 ^ 1'b0 ;
  assign n2503 = ( n206 & n1570 ) | ( n206 & ~n2502 ) | ( n1570 & ~n2502 ) ;
  assign n2509 = n2508 ^ n2504 ^ n2503 ;
  assign n2510 = n1139 & n2394 ;
  assign n2511 = n903 & n2510 ;
  assign n2515 = n2038 ^ n1869 ^ n1060 ;
  assign n2512 = n2280 ^ n1052 ^ 1'b0 ;
  assign n2513 = n1818 & n2512 ;
  assign n2514 = ( x85 & n1416 ) | ( x85 & n2513 ) | ( n1416 & n2513 ) ;
  assign n2516 = n2515 ^ n2514 ^ 1'b0 ;
  assign n2517 = n2516 ^ n2100 ^ 1'b0 ;
  assign n2518 = n2511 | n2517 ;
  assign n2519 = ~n1267 & n1505 ;
  assign n2520 = n2518 & n2519 ;
  assign n2521 = n669 ^ n188 ^ 1'b0 ;
  assign n2522 = ( ~x127 & n1157 ) | ( ~x127 & n1381 ) | ( n1157 & n1381 ) ;
  assign n2523 = ( n692 & n2521 ) | ( n692 & n2522 ) | ( n2521 & n2522 ) ;
  assign n2524 = n1123 ^ n247 ^ 1'b0 ;
  assign n2525 = n2524 ^ n2342 ^ 1'b0 ;
  assign n2526 = n734 & ~n2525 ;
  assign n2527 = n2526 ^ x12 ^ 1'b0 ;
  assign n2536 = ( x108 & n1620 ) | ( x108 & n2283 ) | ( n1620 & n2283 ) ;
  assign n2537 = n1295 ^ x10 ^ 1'b0 ;
  assign n2538 = n2537 ^ n746 ^ 1'b0 ;
  assign n2539 = n2536 & ~n2538 ;
  assign n2533 = n1858 ^ n500 ^ 1'b0 ;
  assign n2534 = n301 & n2533 ;
  assign n2528 = ( ~n242 & n422 ) | ( ~n242 & n424 ) | ( n422 & n424 ) ;
  assign n2529 = n1723 | n2528 ;
  assign n2530 = n2529 ^ x52 ^ 1'b0 ;
  assign n2531 = n1394 ^ n214 ^ 1'b0 ;
  assign n2532 = n2530 & n2531 ;
  assign n2535 = n2534 ^ n2532 ^ n753 ;
  assign n2540 = n2539 ^ n2535 ^ 1'b0 ;
  assign n2541 = n2081 & ~n2540 ;
  assign n2542 = ( x122 & n703 ) | ( x122 & ~n952 ) | ( n703 & ~n952 ) ;
  assign n2543 = n998 | n2542 ;
  assign n2544 = n319 & ~n1100 ;
  assign n2545 = ( n2541 & n2543 ) | ( n2541 & n2544 ) | ( n2543 & n2544 ) ;
  assign n2546 = ~n162 & n442 ;
  assign n2547 = n2546 ^ n522 ^ 1'b0 ;
  assign n2548 = n2547 ^ x62 ^ 1'b0 ;
  assign n2549 = n2190 & n2548 ;
  assign n2550 = n2077 | n2549 ;
  assign n2551 = n998 & ~n1687 ;
  assign n2552 = n2551 ^ n2071 ^ 1'b0 ;
  assign n2553 = ~n835 & n1907 ;
  assign n2556 = n194 | n837 ;
  assign n2557 = n2027 | n2556 ;
  assign n2555 = n2305 ^ n1455 ^ x50 ;
  assign n2558 = n2557 ^ n2555 ^ 1'b0 ;
  assign n2559 = n2558 ^ n800 ^ n599 ;
  assign n2554 = n1441 | n1853 ;
  assign n2560 = n2559 ^ n2554 ^ 1'b0 ;
  assign n2561 = n2560 ^ n756 ^ 1'b0 ;
  assign n2562 = n1441 ^ n1101 ^ n281 ;
  assign n2563 = n2111 ^ n723 ^ n461 ;
  assign n2564 = ( n683 & ~n2562 ) | ( n683 & n2563 ) | ( ~n2562 & n2563 ) ;
  assign n2565 = n442 | n2564 ;
  assign n2566 = n1330 & ~n2085 ;
  assign n2567 = n2566 ^ n822 ^ 1'b0 ;
  assign n2568 = n1969 & ~n2567 ;
  assign n2572 = ( ~n464 & n563 ) | ( ~n464 & n1856 ) | ( n563 & n1856 ) ;
  assign n2569 = n1089 & n1198 ;
  assign n2570 = n1629 ^ x68 ^ 1'b0 ;
  assign n2571 = n2569 & n2570 ;
  assign n2573 = n2572 ^ n2571 ^ n2465 ;
  assign n2575 = n2265 ^ n1381 ^ 1'b0 ;
  assign n2576 = x47 & ~n2575 ;
  assign n2577 = x107 & n2576 ;
  assign n2578 = n2577 ^ n708 ^ 1'b0 ;
  assign n2574 = ~n1464 & n2263 ;
  assign n2579 = n2578 ^ n2574 ^ 1'b0 ;
  assign n2585 = n1554 ^ n447 ^ n393 ;
  assign n2582 = n2190 ^ n1196 ^ 1'b0 ;
  assign n2583 = n1443 | n2582 ;
  assign n2584 = n1056 & ~n2583 ;
  assign n2580 = ~n1774 & n2383 ;
  assign n2581 = n914 & n2580 ;
  assign n2586 = n2585 ^ n2584 ^ n2581 ;
  assign n2587 = n1939 ^ n291 ^ 1'b0 ;
  assign n2588 = n476 | n2229 ;
  assign n2589 = n2587 | n2588 ;
  assign n2590 = n2426 ^ n2007 ^ n1366 ;
  assign n2596 = n260 ^ x94 ^ 1'b0 ;
  assign n2597 = n2571 & ~n2596 ;
  assign n2594 = x39 & n863 ;
  assign n2595 = n2594 ^ n1244 ^ 1'b0 ;
  assign n2591 = n1494 ^ n486 ^ 1'b0 ;
  assign n2592 = n2091 & ~n2591 ;
  assign n2593 = ( x7 & n1439 ) | ( x7 & n2592 ) | ( n1439 & n2592 ) ;
  assign n2598 = n2597 ^ n2595 ^ n2593 ;
  assign n2599 = n1843 ^ n1819 ^ 1'b0 ;
  assign n2600 = ( n408 & ~n986 ) | ( n408 & n2534 ) | ( ~n986 & n2534 ) ;
  assign n2601 = n979 & n2600 ;
  assign n2602 = ~n2599 & n2601 ;
  assign n2603 = ( ~n627 & n659 ) | ( ~n627 & n715 ) | ( n659 & n715 ) ;
  assign n2606 = n588 ^ n457 ^ x8 ;
  assign n2607 = n2606 ^ n787 ^ 1'b0 ;
  assign n2608 = n1308 & n1585 ;
  assign n2609 = ( n361 & n2607 ) | ( n361 & n2608 ) | ( n2607 & n2608 ) ;
  assign n2604 = n678 ^ x62 ^ 1'b0 ;
  assign n2605 = n1199 | n2604 ;
  assign n2610 = n2609 ^ n2605 ^ n1660 ;
  assign n2611 = ~n2603 & n2610 ;
  assign n2612 = ~n905 & n2611 ;
  assign n2613 = n157 & ~n699 ;
  assign n2614 = ~n409 & n1165 ;
  assign n2615 = n1076 | n2614 ;
  assign n2616 = n728 & n1077 ;
  assign n2621 = n968 ^ x110 ^ 1'b0 ;
  assign n2622 = n2151 & ~n2410 ;
  assign n2623 = ~n2621 & n2622 ;
  assign n2617 = ~n559 & n650 ;
  assign n2618 = n2617 ^ n1986 ^ 1'b0 ;
  assign n2619 = ( n1400 & ~n1979 ) | ( n1400 & n2618 ) | ( ~n1979 & n2618 ) ;
  assign n2620 = ~n1862 & n2619 ;
  assign n2624 = n2623 ^ n2620 ^ 1'b0 ;
  assign n2625 = n445 & n972 ;
  assign n2626 = n2462 ^ x22 ^ 1'b0 ;
  assign n2627 = ( x24 & ~n1117 ) | ( x24 & n1918 ) | ( ~n1117 & n1918 ) ;
  assign n2628 = n2627 ^ n1793 ^ 1'b0 ;
  assign n2629 = ~n2626 & n2628 ;
  assign n2630 = x122 & ~n2511 ;
  assign n2631 = n1425 & n2630 ;
  assign n2632 = ~n837 & n2631 ;
  assign n2633 = n296 ^ n199 ^ 1'b0 ;
  assign n2634 = x97 & ~n2633 ;
  assign n2635 = n448 & n2634 ;
  assign n2636 = ~n2178 & n2635 ;
  assign n2637 = ( ~n810 & n1856 ) | ( ~n810 & n2636 ) | ( n1856 & n2636 ) ;
  assign n2638 = n2637 ^ n2046 ^ n332 ;
  assign n2639 = n689 & n1032 ;
  assign n2640 = x63 | n1572 ;
  assign n2641 = n2391 & n2640 ;
  assign n2642 = ( n928 & n1516 ) | ( n928 & n1966 ) | ( n1516 & n1966 ) ;
  assign n2643 = n1587 ^ n1555 ^ 1'b0 ;
  assign n2644 = n2642 | n2643 ;
  assign n2645 = n2644 ^ n1687 ^ n404 ;
  assign n2646 = n1890 & n2173 ;
  assign n2647 = ( n933 & ~n2645 ) | ( n933 & n2646 ) | ( ~n2645 & n2646 ) ;
  assign n2650 = n1912 & n2124 ;
  assign n2648 = n987 ^ n734 ^ n310 ;
  assign n2649 = n2648 ^ n476 ^ n156 ;
  assign n2651 = n2650 ^ n2649 ^ 1'b0 ;
  assign n2652 = n1001 & n2651 ;
  assign n2653 = n2652 ^ n548 ^ 1'b0 ;
  assign n2654 = ( x56 & ~n1311 ) | ( x56 & n2116 ) | ( ~n1311 & n2116 ) ;
  assign n2655 = n394 ^ n335 ^ 1'b0 ;
  assign n2656 = n779 & n1757 ;
  assign n2657 = ~n589 & n2656 ;
  assign n2658 = ( n428 & n429 ) | ( n428 & ~n1084 ) | ( n429 & ~n1084 ) ;
  assign n2659 = n557 | n579 ;
  assign n2660 = n420 & n1117 ;
  assign n2661 = n1275 & n2660 ;
  assign n2662 = ~n2532 & n2661 ;
  assign n2663 = ( n399 & ~n627 ) | ( n399 & n2662 ) | ( ~n627 & n2662 ) ;
  assign n2664 = n2663 ^ n1922 ^ 1'b0 ;
  assign n2665 = ~n2659 & n2664 ;
  assign n2666 = n1527 ^ n296 ^ n255 ;
  assign n2667 = ( ~n812 & n1108 ) | ( ~n812 & n2162 ) | ( n1108 & n2162 ) ;
  assign n2668 = n318 ^ n199 ^ 1'b0 ;
  assign n2669 = n956 & ~n2668 ;
  assign n2670 = ~n1450 & n2669 ;
  assign n2671 = n187 & ~n1033 ;
  assign n2672 = x6 & ~n1897 ;
  assign n2673 = ~x115 & n2672 ;
  assign n2674 = n188 & n1842 ;
  assign n2675 = ( n1820 & ~n2006 ) | ( n1820 & n2674 ) | ( ~n2006 & n2674 ) ;
  assign n2676 = ( ~n1092 & n2673 ) | ( ~n1092 & n2675 ) | ( n2673 & n2675 ) ;
  assign n2679 = n1880 ^ n1238 ^ 1'b0 ;
  assign n2677 = n386 & ~n1013 ;
  assign n2678 = n1190 & n2677 ;
  assign n2680 = n2679 ^ n2678 ^ 1'b0 ;
  assign n2681 = ~n1807 & n2680 ;
  assign n2682 = n256 ^ n156 ^ x96 ;
  assign n2683 = n2178 & ~n2682 ;
  assign n2684 = ~n277 & n1178 ;
  assign n2685 = n2684 ^ n664 ^ 1'b0 ;
  assign n2686 = n2683 & ~n2685 ;
  assign n2687 = n603 ^ n182 ^ 1'b0 ;
  assign n2688 = n2687 ^ n1132 ^ x107 ;
  assign n2689 = ( n891 & ~n1786 ) | ( n891 & n2679 ) | ( ~n1786 & n2679 ) ;
  assign n2696 = n1189 & n1763 ;
  assign n2697 = ~n1426 & n2696 ;
  assign n2693 = n1869 ^ n1258 ^ n180 ;
  assign n2690 = ~n1617 & n2029 ;
  assign n2691 = n2690 ^ n1229 ^ 1'b0 ;
  assign n2692 = n2296 & ~n2691 ;
  assign n2694 = n2693 ^ n2692 ^ n1860 ;
  assign n2695 = n472 & n2694 ;
  assign n2698 = n2697 ^ n2695 ^ 1'b0 ;
  assign n2699 = n1314 | n2698 ;
  assign n2700 = n768 & n1846 ;
  assign n2701 = n1003 & n2700 ;
  assign n2702 = ( n833 & ~n1763 ) | ( n833 & n2701 ) | ( ~n1763 & n2701 ) ;
  assign n2703 = n2702 ^ n2115 ^ n1268 ;
  assign n2707 = ( n170 & n1668 ) | ( n170 & n2160 ) | ( n1668 & n2160 ) ;
  assign n2704 = x117 & ~n2252 ;
  assign n2705 = n2704 ^ n1645 ^ x6 ;
  assign n2706 = n2705 ^ n2555 ^ n157 ;
  assign n2708 = n2707 ^ n2706 ^ 1'b0 ;
  assign n2709 = n2336 | n2708 ;
  assign n2710 = n419 & ~n673 ;
  assign n2711 = ~n329 & n2710 ;
  assign n2712 = n2711 ^ n2565 ^ n1801 ;
  assign n2713 = n2665 & n2712 ;
  assign n2717 = n1213 & n1422 ;
  assign n2714 = ~n1184 & n2534 ;
  assign n2715 = n2714 ^ n928 ^ 1'b0 ;
  assign n2716 = n143 & ~n2715 ;
  assign n2718 = n2717 ^ n2716 ^ 1'b0 ;
  assign n2719 = ~n234 & n2280 ;
  assign n2720 = n1776 & n2719 ;
  assign n2721 = n2036 & ~n2720 ;
  assign n2722 = n2718 & n2721 ;
  assign n2723 = n2722 ^ n2693 ^ n1666 ;
  assign n2728 = n2090 ^ n467 ^ x123 ;
  assign n2726 = n1396 & ~n1518 ;
  assign n2724 = n539 | n887 ;
  assign n2725 = n786 & n2724 ;
  assign n2727 = n2726 ^ n2725 ^ 1'b0 ;
  assign n2729 = n2728 ^ n2727 ^ n1175 ;
  assign n2732 = ~n241 & n610 ;
  assign n2730 = n358 | n1397 ;
  assign n2731 = n352 | n2730 ;
  assign n2733 = n2732 ^ n2731 ^ 1'b0 ;
  assign n2737 = n2562 ^ n594 ^ n289 ;
  assign n2735 = n1123 & ~n2092 ;
  assign n2736 = n1132 & ~n2735 ;
  assign n2734 = n511 & n2394 ;
  assign n2738 = n2737 ^ n2736 ^ n2734 ;
  assign n2739 = n1505 & n1617 ;
  assign n2740 = n2215 & n2739 ;
  assign n2741 = x3 & ~n971 ;
  assign n2742 = n767 & n2741 ;
  assign n2743 = n153 & ~n2409 ;
  assign n2744 = n2100 ^ n537 ^ n416 ;
  assign n2745 = ( ~n1165 & n2310 ) | ( ~n1165 & n2744 ) | ( n2310 & n2744 ) ;
  assign n2746 = n1561 ^ n850 ^ n216 ;
  assign n2747 = x35 & n2746 ;
  assign n2748 = ~n936 & n2747 ;
  assign n2749 = n2748 ^ n1156 ^ n448 ;
  assign n2750 = n2749 ^ n1061 ^ 1'b0 ;
  assign n2751 = x13 & ~n2750 ;
  assign n2752 = ( n2097 & n2550 ) | ( n2097 & ~n2751 ) | ( n2550 & ~n2751 ) ;
  assign n2753 = n162 | n1340 ;
  assign n2754 = n1503 | n2753 ;
  assign n2755 = n713 & ~n1712 ;
  assign n2756 = n2755 ^ n1274 ^ 1'b0 ;
  assign n2757 = n2756 ^ n877 ^ x82 ;
  assign n2759 = n1198 ^ n255 ^ 1'b0 ;
  assign n2760 = n1187 & n2759 ;
  assign n2758 = n502 & ~n1508 ;
  assign n2761 = n2760 ^ n2758 ^ n580 ;
  assign n2762 = n1645 ^ n1405 ^ 1'b0 ;
  assign n2763 = n2394 ^ n1615 ^ 1'b0 ;
  assign n2764 = n2763 ^ n2642 ^ n1542 ;
  assign n2766 = ( ~x93 & n320 ) | ( ~x93 & n1379 ) | ( n320 & n1379 ) ;
  assign n2767 = n2766 ^ n815 ^ n531 ;
  assign n2768 = n2767 ^ n1444 ^ 1'b0 ;
  assign n2765 = n545 & n2549 ;
  assign n2769 = n2768 ^ n2765 ^ 1'b0 ;
  assign n2770 = n1597 ^ n1494 ^ n265 ;
  assign n2772 = n1428 ^ n1056 ^ n786 ;
  assign n2773 = n2257 ^ n1405 ^ 1'b0 ;
  assign n2774 = n1615 ^ n733 ^ n646 ;
  assign n2775 = n2774 ^ n1198 ^ 1'b0 ;
  assign n2776 = ~n1419 & n2775 ;
  assign n2777 = n1232 & n2776 ;
  assign n2778 = ~n2773 & n2777 ;
  assign n2779 = ( ~n533 & n2772 ) | ( ~n533 & n2778 ) | ( n2772 & n2778 ) ;
  assign n2771 = x19 & n1741 ;
  assign n2780 = n2779 ^ n2771 ^ 1'b0 ;
  assign n2781 = n557 ^ n237 ^ n164 ;
  assign n2782 = n253 & n2781 ;
  assign n2783 = ( ~n2770 & n2780 ) | ( ~n2770 & n2782 ) | ( n2780 & n2782 ) ;
  assign n2784 = n1543 ^ n1473 ^ n506 ;
  assign n2785 = n947 | n1732 ;
  assign n2786 = n1978 ^ n1417 ^ n887 ;
  assign n2787 = n2786 ^ n1357 ^ n379 ;
  assign n2788 = n972 & ~n2787 ;
  assign n2789 = ( ~x116 & n1035 ) | ( ~x116 & n2059 ) | ( n1035 & n2059 ) ;
  assign n2790 = n1020 & ~n2789 ;
  assign n2800 = x9 & n983 ;
  assign n2801 = n2800 ^ n226 ^ 1'b0 ;
  assign n2792 = n612 ^ x43 ^ x11 ;
  assign n2793 = n2792 ^ n821 ^ n787 ;
  assign n2791 = ~n547 & n666 ;
  assign n2794 = n2793 ^ n2791 ^ 1'b0 ;
  assign n2795 = ~n2065 & n2794 ;
  assign n2796 = ~n1581 & n2795 ;
  assign n2797 = n1032 ^ n971 ^ 1'b0 ;
  assign n2798 = n2797 ^ n2199 ^ n1976 ;
  assign n2799 = ( x44 & n2796 ) | ( x44 & ~n2798 ) | ( n2796 & ~n2798 ) ;
  assign n2802 = n2801 ^ n2799 ^ 1'b0 ;
  assign n2803 = n605 & ~n708 ;
  assign n2804 = n1920 & n2803 ;
  assign n2805 = n1909 ^ n1077 ^ n717 ;
  assign n2806 = n2161 ^ n1799 ^ 1'b0 ;
  assign n2807 = n2805 | n2806 ;
  assign n2808 = ( n290 & ~n1467 ) | ( n290 & n2807 ) | ( ~n1467 & n2807 ) ;
  assign n2809 = n218 | n696 ;
  assign n2810 = n248 & ~n2809 ;
  assign n2811 = ( n990 & n2618 ) | ( n990 & n2810 ) | ( n2618 & n2810 ) ;
  assign n2812 = n490 & n2811 ;
  assign n2813 = n454 & n2812 ;
  assign n2814 = x119 & ~n2813 ;
  assign n2815 = n2814 ^ n535 ^ 1'b0 ;
  assign n2816 = ( n2804 & n2808 ) | ( n2804 & ~n2815 ) | ( n2808 & ~n2815 ) ;
  assign n2817 = ~n154 & n1095 ;
  assign n2819 = n1294 ^ n721 ^ n485 ;
  assign n2818 = n1048 ^ n967 ^ n663 ;
  assign n2820 = n2819 ^ n2818 ^ 1'b0 ;
  assign n2821 = n2820 ^ n1726 ^ 1'b0 ;
  assign n2822 = n548 & ~n1707 ;
  assign n2823 = n2792 & ~n2822 ;
  assign n2824 = n375 & ~n862 ;
  assign n2825 = ~n452 & n2537 ;
  assign n2826 = n2824 & n2825 ;
  assign n2827 = n2826 ^ n1304 ^ 1'b0 ;
  assign n2830 = n1342 ^ n1132 ^ n635 ;
  assign n2828 = n447 ^ x113 ^ 1'b0 ;
  assign n2829 = ~n1583 & n2828 ;
  assign n2831 = n2830 ^ n2829 ^ 1'b0 ;
  assign n2832 = n1916 & n2160 ;
  assign n2833 = n2832 ^ n230 ^ 1'b0 ;
  assign n2834 = ( n298 & n366 ) | ( n298 & ~n1784 ) | ( n366 & ~n1784 ) ;
  assign n2835 = ~n1296 & n2834 ;
  assign n2836 = ~x103 & n2835 ;
  assign n2840 = n2110 ^ n1455 ^ n558 ;
  assign n2837 = n2129 ^ n1510 ^ 1'b0 ;
  assign n2838 = n1899 & n2837 ;
  assign n2839 = n2838 ^ n1072 ^ 1'b0 ;
  assign n2841 = n2840 ^ n2839 ^ 1'b0 ;
  assign n2842 = n2836 & n2841 ;
  assign n2843 = n1328 & n1616 ;
  assign n2844 = n800 & ~n2352 ;
  assign n2845 = n924 & n932 ;
  assign n2846 = n365 | n743 ;
  assign n2847 = n2845 & n2846 ;
  assign n2848 = n1013 ^ n618 ^ n158 ;
  assign n2849 = ( ~n454 & n2847 ) | ( ~n454 & n2848 ) | ( n2847 & n2848 ) ;
  assign n2850 = ~n485 & n2842 ;
  assign n2851 = n802 & n2850 ;
  assign n2852 = n661 & ~n1254 ;
  assign n2853 = n2852 ^ n2197 ^ 1'b0 ;
  assign n2856 = ( ~n969 & n1278 ) | ( ~n969 & n1905 ) | ( n1278 & n1905 ) ;
  assign n2854 = ( x70 & ~n605 ) | ( x70 & n699 ) | ( ~n605 & n699 ) ;
  assign n2855 = x90 & n2854 ;
  assign n2857 = n2856 ^ n2855 ^ n154 ;
  assign n2858 = n2857 ^ n786 ^ 1'b0 ;
  assign n2859 = x104 ^ x88 ^ x57 ;
  assign n2860 = ( x112 & n346 ) | ( x112 & ~n654 ) | ( n346 & ~n654 ) ;
  assign n2861 = n2860 ^ n208 ^ 1'b0 ;
  assign n2862 = n2443 & ~n2861 ;
  assign n2863 = ( n681 & n2859 ) | ( n681 & n2862 ) | ( n2859 & n2862 ) ;
  assign n2867 = n1846 ^ x116 ^ x100 ;
  assign n2864 = n1501 & n2274 ;
  assign n2865 = ~x35 & n2864 ;
  assign n2866 = n170 & ~n2865 ;
  assign n2868 = n2867 ^ n2866 ^ 1'b0 ;
  assign n2869 = n294 & n1827 ;
  assign n2870 = n2869 ^ n2418 ^ 1'b0 ;
  assign n2871 = ( x5 & n2868 ) | ( x5 & n2870 ) | ( n2868 & n2870 ) ;
  assign n2873 = x21 & ~n970 ;
  assign n2874 = ~n989 & n2873 ;
  assign n2872 = n413 ^ n144 ^ 1'b0 ;
  assign n2875 = n2874 ^ n2872 ^ n1934 ;
  assign n2876 = n2130 ^ n1886 ^ x40 ;
  assign n2877 = n2876 ^ n2659 ^ 1'b0 ;
  assign n2878 = n2361 & ~n2877 ;
  assign n2879 = n649 | n1505 ;
  assign n2880 = n2879 ^ n245 ^ 1'b0 ;
  assign n2881 = n388 | n2880 ;
  assign n2884 = n924 ^ n815 ^ 1'b0 ;
  assign n2885 = ( n356 & n940 ) | ( n356 & n2884 ) | ( n940 & n2884 ) ;
  assign n2882 = ( n348 & ~n924 ) | ( n348 & n1346 ) | ( ~n924 & n1346 ) ;
  assign n2883 = n2882 ^ n1448 ^ n973 ;
  assign n2886 = n2885 ^ n2883 ^ n366 ;
  assign n2887 = n2511 ^ n899 ^ 1'b0 ;
  assign n2888 = n1298 ^ n597 ^ 1'b0 ;
  assign n2889 = ~n831 & n2888 ;
  assign n2890 = n2889 ^ n2299 ^ 1'b0 ;
  assign n2891 = n1735 | n2890 ;
  assign n2892 = n1830 | n2626 ;
  assign n2893 = n2892 ^ n1274 ^ 1'b0 ;
  assign n2894 = n1288 & ~n2893 ;
  assign n2895 = ~n1243 & n1252 ;
  assign n2896 = n2411 & ~n2895 ;
  assign n2897 = n2757 ^ n2116 ^ n1687 ;
  assign n2898 = n1801 ^ n715 ^ n487 ;
  assign n2899 = n2898 ^ n1603 ^ 1'b0 ;
  assign n2900 = ( x2 & n290 ) | ( x2 & ~n2453 ) | ( n290 & ~n2453 ) ;
  assign n2901 = n647 ^ x57 ^ 1'b0 ;
  assign n2902 = n2901 ^ n1961 ^ 1'b0 ;
  assign n2903 = n2900 & n2902 ;
  assign n2904 = n691 & n1162 ;
  assign n2905 = n724 & n2904 ;
  assign n2906 = n1516 | n2905 ;
  assign n2907 = n2906 ^ n2309 ^ 1'b0 ;
  assign n2908 = n1443 | n2907 ;
  assign n2909 = n1913 | n2597 ;
  assign n2910 = n2909 ^ n1149 ^ 1'b0 ;
  assign n2911 = n2811 ^ n1935 ^ n1280 ;
  assign n2912 = ( n1277 & n1810 ) | ( n1277 & n2911 ) | ( n1810 & n2911 ) ;
  assign n2915 = ( n329 & n2085 ) | ( n329 & n2323 ) | ( n2085 & n2323 ) ;
  assign n2916 = n2915 ^ n255 ^ 1'b0 ;
  assign n2917 = n2085 | n2916 ;
  assign n2918 = ( ~n1282 & n2079 ) | ( ~n1282 & n2917 ) | ( n2079 & n2917 ) ;
  assign n2913 = n2810 ^ n1422 ^ n893 ;
  assign n2914 = n2913 ^ n522 ^ 1'b0 ;
  assign n2919 = n2918 ^ n2914 ^ n383 ;
  assign n2920 = ~n1819 & n1890 ;
  assign n2921 = ~n1898 & n2920 ;
  assign n2922 = ( ~n199 & n2862 ) | ( ~n199 & n2921 ) | ( n2862 & n2921 ) ;
  assign n2923 = ( ~x84 & n1345 ) | ( ~x84 & n2160 ) | ( n1345 & n2160 ) ;
  assign n2924 = n2923 ^ n2308 ^ 1'b0 ;
  assign n2925 = n2922 | n2924 ;
  assign n2926 = n2807 ^ n2573 ^ n550 ;
  assign n2927 = ( n1494 & ~n1846 ) | ( n1494 & n1858 ) | ( ~n1846 & n1858 ) ;
  assign n2928 = n447 | n2927 ;
  assign n2929 = n999 | n2928 ;
  assign n2930 = n837 | n2310 ;
  assign n2931 = n2062 & ~n2930 ;
  assign n2932 = n367 | n541 ;
  assign n2933 = ~n681 & n919 ;
  assign n2934 = n2933 ^ n527 ^ 1'b0 ;
  assign n2935 = n1957 | n2934 ;
  assign n2936 = n2338 & ~n2935 ;
  assign n2937 = ( x45 & n1688 ) | ( x45 & ~n2600 ) | ( n1688 & ~n2600 ) ;
  assign n2938 = ( x33 & n1448 ) | ( x33 & ~n2937 ) | ( n1448 & ~n2937 ) ;
  assign n2939 = n2938 ^ n1730 ^ n589 ;
  assign n2940 = n260 & ~n2939 ;
  assign n2941 = n2936 & n2940 ;
  assign n2945 = n456 & ~n1427 ;
  assign n2946 = n522 | n2945 ;
  assign n2947 = n302 | n2946 ;
  assign n2948 = n2947 ^ n1185 ^ n608 ;
  assign n2942 = n2381 ^ n378 ^ 1'b0 ;
  assign n2943 = n1905 | n2942 ;
  assign n2944 = ( ~n668 & n885 ) | ( ~n668 & n2943 ) | ( n885 & n2943 ) ;
  assign n2949 = n2948 ^ n2944 ^ n2929 ;
  assign n2950 = n2045 ^ n1864 ^ 1'b0 ;
  assign n2951 = ~n866 & n1123 ;
  assign n2952 = n1092 | n2951 ;
  assign n2953 = n1811 | n2952 ;
  assign n2954 = x35 & n2953 ;
  assign n2955 = n160 & n2954 ;
  assign n2957 = n161 & n1176 ;
  assign n2958 = n2957 ^ n764 ^ 1'b0 ;
  assign n2959 = ( ~n636 & n2796 ) | ( ~n636 & n2958 ) | ( n2796 & n2958 ) ;
  assign n2960 = n2728 ^ n1982 ^ 1'b0 ;
  assign n2961 = ~n2959 & n2960 ;
  assign n2962 = n2961 ^ n1274 ^ 1'b0 ;
  assign n2963 = n2962 ^ n701 ^ 1'b0 ;
  assign n2956 = n2381 ^ n1279 ^ n468 ;
  assign n2964 = n2963 ^ n2956 ^ 1'b0 ;
  assign n2965 = n2792 ^ n2659 ^ n248 ;
  assign n2966 = n310 & n603 ;
  assign n2967 = n2965 & n2966 ;
  assign n2968 = n2967 ^ n2845 ^ n2101 ;
  assign n2973 = n2683 ^ n2006 ^ 1'b0 ;
  assign n2974 = n1951 | n2973 ;
  assign n2969 = ( ~n1139 & n1272 ) | ( ~n1139 & n2081 ) | ( n1272 & n2081 ) ;
  assign n2970 = n2969 ^ n2283 ^ n751 ;
  assign n2971 = n2970 ^ n1449 ^ 1'b0 ;
  assign n2972 = n1337 & n2971 ;
  assign n2975 = n2974 ^ n2972 ^ n1689 ;
  assign n2976 = n379 | n2086 ;
  assign n2977 = n2976 ^ n1561 ^ 1'b0 ;
  assign n2978 = n1378 ^ n661 ^ n408 ;
  assign n2979 = n2978 ^ n2899 ^ 1'b0 ;
  assign n2980 = ~n631 & n2979 ;
  assign n2981 = n539 | n1060 ;
  assign n2982 = ( n508 & n1334 ) | ( n508 & n2981 ) | ( n1334 & n2981 ) ;
  assign n2983 = n1848 ^ x17 ^ 1'b0 ;
  assign n2984 = n498 | n2983 ;
  assign n2985 = n2097 | n2984 ;
  assign n2986 = n692 ^ n230 ^ 1'b0 ;
  assign n2987 = ~n559 & n2986 ;
  assign n2988 = n1334 ^ n715 ^ 1'b0 ;
  assign n2989 = ( ~x123 & n2987 ) | ( ~x123 & n2988 ) | ( n2987 & n2988 ) ;
  assign n2990 = n2522 ^ n1913 ^ 1'b0 ;
  assign n2991 = x40 & ~n247 ;
  assign n2992 = n2991 ^ n1157 ^ 1'b0 ;
  assign n2993 = ( n865 & n1779 ) | ( n865 & ~n2992 ) | ( n1779 & ~n2992 ) ;
  assign n2994 = ( n972 & ~n1283 ) | ( n972 & n1636 ) | ( ~n1283 & n1636 ) ;
  assign n2995 = n1437 & n2994 ;
  assign n2996 = n1075 & n2995 ;
  assign n2998 = n689 ^ x102 ^ 1'b0 ;
  assign n2997 = ~n1044 & n1501 ;
  assign n2999 = n2998 ^ n2997 ^ 1'b0 ;
  assign n3000 = n2048 | n2999 ;
  assign n3001 = n3000 ^ x103 ^ 1'b0 ;
  assign n3002 = n191 & ~n1392 ;
  assign n3003 = ( x70 & n1619 ) | ( x70 & n1679 ) | ( n1619 & n1679 ) ;
  assign n3004 = ( n2673 & n3002 ) | ( n2673 & ~n3003 ) | ( n3002 & ~n3003 ) ;
  assign n3005 = x92 | n971 ;
  assign n3006 = n1084 | n1417 ;
  assign n3007 = x36 | n3006 ;
  assign n3008 = ~n984 & n3007 ;
  assign n3009 = n3005 & n3008 ;
  assign n3010 = n1714 & n3009 ;
  assign n3024 = n903 ^ n629 ^ 1'b0 ;
  assign n3018 = n2959 ^ n1897 ^ n1084 ;
  assign n3020 = n838 & ~n1156 ;
  assign n3019 = ( n323 & n1943 ) | ( n323 & ~n2160 ) | ( n1943 & ~n2160 ) ;
  assign n3021 = n3020 ^ n3019 ^ 1'b0 ;
  assign n3022 = ~n2401 & n3021 ;
  assign n3023 = ~n3018 & n3022 ;
  assign n3025 = n3024 ^ n3023 ^ 1'b0 ;
  assign n3011 = n488 & ~n603 ;
  assign n3012 = ~n467 & n2434 ;
  assign n3013 = n3011 & n3012 ;
  assign n3014 = n3013 ^ n1311 ^ 1'b0 ;
  assign n3015 = n930 & n3014 ;
  assign n3016 = x101 & ~n756 ;
  assign n3017 = n3015 & ~n3016 ;
  assign n3026 = n3025 ^ n3017 ^ 1'b0 ;
  assign n3027 = ( x117 & ~n479 ) | ( x117 & n2945 ) | ( ~n479 & n2945 ) ;
  assign n3028 = n3027 ^ n256 ^ 1'b0 ;
  assign n3029 = ( n178 & ~n1364 ) | ( n178 & n2307 ) | ( ~n1364 & n2307 ) ;
  assign n3030 = n3029 ^ n661 ^ 1'b0 ;
  assign n3031 = x117 & n2634 ;
  assign n3032 = n3031 ^ n1294 ^ n187 ;
  assign n3033 = ( n1095 & ~n2569 ) | ( n1095 & n3032 ) | ( ~n2569 & n3032 ) ;
  assign n3034 = n2162 & n3033 ;
  assign n3035 = n3030 & n3034 ;
  assign n3036 = n3035 ^ n1725 ^ 1'b0 ;
  assign n3037 = n625 & ~n2653 ;
  assign n3039 = n623 | n3016 ;
  assign n3040 = x14 | n3039 ;
  assign n3041 = n3040 ^ n872 ^ 1'b0 ;
  assign n3042 = x0 & n3041 ;
  assign n3043 = ~n2359 & n3042 ;
  assign n3044 = n1987 & n3043 ;
  assign n3038 = n167 & ~n1481 ;
  assign n3045 = n3044 ^ n3038 ^ 1'b0 ;
  assign n3046 = ~n209 & n2834 ;
  assign n3047 = n3046 ^ n2819 ^ 1'b0 ;
  assign n3051 = n531 | n1139 ;
  assign n3050 = n1232 ^ n1229 ^ 1'b0 ;
  assign n3048 = n2772 ^ n829 ^ 1'b0 ;
  assign n3049 = ~n2156 & n3048 ;
  assign n3052 = n3051 ^ n3050 ^ n3049 ;
  assign n3053 = n3052 ^ n866 ^ 1'b0 ;
  assign n3054 = x60 & n3053 ;
  assign n3055 = n205 & ~n952 ;
  assign n3056 = n3055 ^ n1602 ^ x50 ;
  assign n3058 = n364 & ~n1433 ;
  assign n3059 = n3058 ^ n1363 ^ 1'b0 ;
  assign n3060 = n3059 ^ n679 ^ n560 ;
  assign n3061 = n3046 ^ n809 ^ 1'b0 ;
  assign n3062 = n3060 & ~n3061 ;
  assign n3057 = ~x57 & n2601 ;
  assign n3063 = n3062 ^ n3057 ^ 1'b0 ;
  assign n3064 = n869 & ~n1152 ;
  assign n3065 = n3064 ^ x3 ^ 1'b0 ;
  assign n3066 = n1879 & ~n3065 ;
  assign n3067 = ~n141 & n3066 ;
  assign n3068 = ( ~n431 & n1374 ) | ( ~n431 & n3067 ) | ( n1374 & n3067 ) ;
  assign n3069 = n322 ^ n234 ^ x119 ;
  assign n3070 = n3069 ^ n1101 ^ x42 ;
  assign n3071 = n2925 ^ n2869 ^ n321 ;
  assign n3072 = ~x94 & n672 ;
  assign n3073 = n2058 | n3072 ;
  assign n3074 = n1381 | n3073 ;
  assign n3075 = n1880 ^ n764 ^ 1'b0 ;
  assign n3076 = ( ~n1214 & n2878 ) | ( ~n1214 & n3075 ) | ( n2878 & n3075 ) ;
  assign n3077 = n1428 & n1966 ;
  assign n3079 = ~n405 & n416 ;
  assign n3080 = n3079 ^ n672 ^ 1'b0 ;
  assign n3078 = n357 & n2895 ;
  assign n3081 = n3080 ^ n3078 ^ 1'b0 ;
  assign n3082 = n147 & ~n437 ;
  assign n3083 = n3082 ^ x75 ^ 1'b0 ;
  assign n3084 = ( n1087 & ~n1810 ) | ( n1087 & n3083 ) | ( ~n1810 & n3083 ) ;
  assign n3085 = n2421 & n3084 ;
  assign n3086 = n3085 ^ n1587 ^ 1'b0 ;
  assign n3087 = ( n167 & ~n298 ) | ( n167 & n1410 ) | ( ~n298 & n1410 ) ;
  assign n3088 = n2505 & n3087 ;
  assign n3089 = n3088 ^ x3 ^ 1'b0 ;
  assign n3090 = n550 | n3089 ;
  assign n3091 = n3090 ^ n1279 ^ 1'b0 ;
  assign n3092 = x127 & n986 ;
  assign n3093 = ~x48 & n3092 ;
  assign n3094 = n3093 ^ n149 ^ 1'b0 ;
  assign n3095 = ~n3091 & n3094 ;
  assign n3096 = n1229 ^ n334 ^ 1'b0 ;
  assign n3097 = ( ~n283 & n2057 ) | ( ~n283 & n2295 ) | ( n2057 & n2295 ) ;
  assign n3098 = ~n267 & n3097 ;
  assign n3099 = ( n1804 & n3096 ) | ( n1804 & ~n3098 ) | ( n3096 & ~n3098 ) ;
  assign n3100 = n1387 ^ n1116 ^ n299 ;
  assign n3101 = n973 & n3100 ;
  assign n3102 = ( n147 & ~n392 ) | ( n147 & n2033 ) | ( ~n392 & n2033 ) ;
  assign n3103 = n3102 ^ n2272 ^ n454 ;
  assign n3104 = n1566 ^ n586 ^ 1'b0 ;
  assign n3105 = ( n728 & n2676 ) | ( n728 & n3104 ) | ( n2676 & n3104 ) ;
  assign n3109 = n1132 ^ n227 ^ 1'b0 ;
  assign n3106 = n1104 ^ n465 ^ 1'b0 ;
  assign n3107 = n517 | n3106 ;
  assign n3108 = n3107 ^ n2121 ^ 1'b0 ;
  assign n3110 = n3109 ^ n3108 ^ n1028 ;
  assign n3111 = n2657 ^ n1590 ^ n595 ;
  assign n3112 = n2797 ^ n1236 ^ n699 ;
  assign n3113 = n3112 ^ n456 ^ 1'b0 ;
  assign n3114 = n2342 & ~n3113 ;
  assign n3115 = n3114 ^ n320 ^ 1'b0 ;
  assign n3116 = n1084 & ~n3115 ;
  assign n3117 = n947 ^ n447 ^ 1'b0 ;
  assign n3118 = n2729 & ~n3117 ;
  assign n3119 = ~n528 & n1348 ;
  assign n3120 = n1910 & n3119 ;
  assign n3121 = n1942 ^ n1423 ^ 1'b0 ;
  assign n3122 = ~n1478 & n1686 ;
  assign n3123 = ~n2152 & n3122 ;
  assign n3124 = n485 ^ x17 ^ 1'b0 ;
  assign n3125 = n3124 ^ n260 ^ 1'b0 ;
  assign n3126 = n1139 & n3125 ;
  assign n3127 = n408 & ~n953 ;
  assign n3128 = ~n3126 & n3127 ;
  assign n3129 = x47 & ~n327 ;
  assign n3130 = n425 & n3129 ;
  assign n3131 = ( ~n222 & n1019 ) | ( ~n222 & n3130 ) | ( n1019 & n3130 ) ;
  assign n3132 = n3131 ^ n1334 ^ 1'b0 ;
  assign n3133 = ( n1139 & n1989 ) | ( n1139 & ~n3132 ) | ( n1989 & ~n3132 ) ;
  assign n3134 = x126 & ~n266 ;
  assign n3135 = ( n766 & ~n2715 ) | ( n766 & n3134 ) | ( ~n2715 & n3134 ) ;
  assign n3136 = ( n538 & n1443 ) | ( n538 & n1464 ) | ( n1443 & n1464 ) ;
  assign n3137 = n161 & n3136 ;
  assign n3138 = n474 & n1781 ;
  assign n3139 = n3138 ^ n2129 ^ 1'b0 ;
  assign n3140 = n3139 ^ n1777 ^ 1'b0 ;
  assign n3141 = n3137 | n3140 ;
  assign n3142 = n2320 | n3141 ;
  assign n3144 = n2143 ^ n1796 ^ n739 ;
  assign n3143 = n1165 & ~n2965 ;
  assign n3145 = n3144 ^ n3143 ^ 1'b0 ;
  assign n3146 = n1733 ^ n1080 ^ n1059 ;
  assign n3147 = n3146 ^ n1172 ^ 1'b0 ;
  assign n3148 = n1638 & n3147 ;
  assign n3149 = ( n134 & ~n361 ) | ( n134 & n1405 ) | ( ~n361 & n1405 ) ;
  assign n3150 = n3149 ^ n1338 ^ 1'b0 ;
  assign n3151 = n3148 & n3150 ;
  assign n3152 = n2059 | n2189 ;
  assign n3153 = n2559 ^ n1041 ^ n856 ;
  assign n3154 = n2671 ^ x71 ^ 1'b0 ;
  assign n3155 = ~n344 & n558 ;
  assign n3156 = n1427 & n3155 ;
  assign n3157 = n1369 ^ n187 ^ 1'b0 ;
  assign n3158 = n3156 | n3157 ;
  assign n3159 = n1699 & n1767 ;
  assign n3160 = n3159 ^ n1086 ^ 1'b0 ;
  assign n3162 = ( n301 & n664 ) | ( n301 & ~n938 ) | ( n664 & ~n938 ) ;
  assign n3161 = n2383 ^ n325 ^ n315 ;
  assign n3163 = n3162 ^ n3161 ^ n1909 ;
  assign n3164 = ( n3158 & n3160 ) | ( n3158 & ~n3163 ) | ( n3160 & ~n3163 ) ;
  assign n3165 = n2782 ^ n1162 ^ 1'b0 ;
  assign n3166 = n3165 ^ n2911 ^ n1885 ;
  assign n3167 = n3166 ^ n2627 ^ n2292 ;
  assign n3169 = n500 ^ x65 ^ 1'b0 ;
  assign n3170 = n2569 ^ n1786 ^ 1'b0 ;
  assign n3171 = n1143 | n3170 ;
  assign n3172 = n488 & n670 ;
  assign n3173 = n1225 & n3172 ;
  assign n3174 = ( n567 & n1842 ) | ( n567 & ~n3173 ) | ( n1842 & ~n3173 ) ;
  assign n3175 = ~n893 & n3174 ;
  assign n3176 = ( n3169 & ~n3171 ) | ( n3169 & n3175 ) | ( ~n3171 & n3175 ) ;
  assign n3168 = n3146 ^ n2726 ^ n1171 ;
  assign n3177 = n3176 ^ n3168 ^ 1'b0 ;
  assign n3178 = n1707 ^ n742 ^ x111 ;
  assign n3179 = n2416 | n3178 ;
  assign n3180 = n2668 | n3179 ;
  assign n3181 = n3180 ^ n607 ^ 1'b0 ;
  assign n3182 = n1638 & n3181 ;
  assign n3183 = n3182 ^ n1663 ^ 1'b0 ;
  assign n3186 = n1188 ^ n852 ^ n627 ;
  assign n3187 = n357 & ~n1603 ;
  assign n3188 = n3186 & n3187 ;
  assign n3184 = n582 & n1801 ;
  assign n3185 = ~n2532 & n3184 ;
  assign n3189 = n3188 ^ n3185 ^ n1511 ;
  assign n3190 = n1466 | n3189 ;
  assign n3191 = ~x72 & n143 ;
  assign n3192 = ( n1625 & ~n1881 ) | ( n1625 & n3191 ) | ( ~n1881 & n3191 ) ;
  assign n3193 = n1062 & n3192 ;
  assign n3194 = ~n2634 & n3193 ;
  assign n3195 = ( n2113 & ~n2921 ) | ( n2113 & n3194 ) | ( ~n2921 & n3194 ) ;
  assign n3196 = n3049 ^ x115 ^ 1'b0 ;
  assign n3197 = n1397 | n3196 ;
  assign n3198 = ( n1928 & n2417 ) | ( n1928 & ~n2847 ) | ( n2417 & ~n2847 ) ;
  assign n3199 = ~n2579 & n3198 ;
  assign n3200 = n3197 & n3199 ;
  assign n3201 = n555 & ~n1250 ;
  assign n3202 = n3201 ^ n1902 ^ 1'b0 ;
  assign n3203 = n1319 & n2674 ;
  assign n3204 = n3203 ^ n1627 ^ 1'b0 ;
  assign n3205 = n3204 ^ n1553 ^ 1'b0 ;
  assign n3206 = ( n221 & ~n2988 ) | ( n221 & n3205 ) | ( ~n2988 & n3205 ) ;
  assign n3207 = ( n3200 & ~n3202 ) | ( n3200 & n3206 ) | ( ~n3202 & n3206 ) ;
  assign n3208 = ~n1807 & n2802 ;
  assign n3209 = n3208 ^ n3104 ^ 1'b0 ;
  assign n3210 = ~n471 & n984 ;
  assign n3211 = ( n161 & n1223 ) | ( n161 & n2607 ) | ( n1223 & n2607 ) ;
  assign n3212 = n3211 ^ n1588 ^ n247 ;
  assign n3213 = n3212 ^ n2141 ^ 1'b0 ;
  assign n3221 = ( n160 & n668 ) | ( n160 & n1162 ) | ( n668 & n1162 ) ;
  assign n3214 = ~n506 & n783 ;
  assign n3215 = n264 | n3214 ;
  assign n3216 = n728 & ~n3215 ;
  assign n3217 = ~n2792 & n3216 ;
  assign n3218 = ( x89 & n1685 ) | ( x89 & n3217 ) | ( n1685 & n3217 ) ;
  assign n3219 = n3218 ^ n1922 ^ 1'b0 ;
  assign n3220 = ~n451 & n3219 ;
  assign n3222 = n3221 ^ n3220 ^ n691 ;
  assign n3223 = ( n219 & ~n2011 ) | ( n219 & n2679 ) | ( ~n2011 & n2679 ) ;
  assign n3224 = ( ~n1764 & n2768 ) | ( ~n1764 & n3223 ) | ( n2768 & n3223 ) ;
  assign n3225 = n997 | n2018 ;
  assign n3226 = n763 & ~n1037 ;
  assign n3227 = n1860 & n3226 ;
  assign n3228 = n1785 | n3227 ;
  assign n3229 = n3228 ^ n1449 ^ n1096 ;
  assign n3230 = ~x86 & n3229 ;
  assign n3231 = n611 ^ n421 ^ 1'b0 ;
  assign n3232 = ~n1533 & n3231 ;
  assign n3233 = n3232 ^ n2211 ^ 1'b0 ;
  assign n3234 = n253 | n3233 ;
  assign n3235 = n1226 ^ n269 ^ x71 ;
  assign n3236 = ~n1481 & n3235 ;
  assign n3237 = n3236 ^ n845 ^ 1'b0 ;
  assign n3238 = ( ~n2355 & n2371 ) | ( ~n2355 & n3237 ) | ( n2371 & n3237 ) ;
  assign n3240 = n1838 ^ n658 ^ 1'b0 ;
  assign n3239 = ( n1230 & n2138 ) | ( n1230 & n2971 ) | ( n2138 & n2971 ) ;
  assign n3241 = n3240 ^ n3239 ^ 1'b0 ;
  assign n3242 = n1236 & ~n3241 ;
  assign n3247 = ( n916 & n934 ) | ( n916 & ~n2939 ) | ( n934 & ~n2939 ) ;
  assign n3248 = n1898 & n2509 ;
  assign n3249 = n3247 & n3248 ;
  assign n3243 = n184 ^ n171 ^ 1'b0 ;
  assign n3244 = n2418 & ~n3243 ;
  assign n3245 = ~n1992 & n3244 ;
  assign n3246 = n156 & n3245 ;
  assign n3250 = n3249 ^ n3246 ^ 1'b0 ;
  assign n3251 = ~n683 & n3250 ;
  assign n3252 = ~n683 & n1348 ;
  assign n3253 = n555 & ~n1427 ;
  assign n3254 = n490 & n3253 ;
  assign n3255 = n3254 ^ n312 ^ 1'b0 ;
  assign n3256 = ( x7 & ~n329 ) | ( x7 & n3255 ) | ( ~n329 & n3255 ) ;
  assign n3257 = x11 | n817 ;
  assign n3258 = n1496 ^ n1185 ^ n815 ;
  assign n3259 = n3258 ^ n1472 ^ n1320 ;
  assign n3260 = ( n132 & n3257 ) | ( n132 & ~n3259 ) | ( n3257 & ~n3259 ) ;
  assign n3261 = n3260 ^ x92 ^ 1'b0 ;
  assign n3262 = ~n3256 & n3261 ;
  assign n3263 = n187 & n2541 ;
  assign n3264 = n3263 ^ n1333 ^ 1'b0 ;
  assign n3265 = n1449 | n1955 ;
  assign n3266 = n877 & ~n1264 ;
  assign n3267 = ( n1607 & ~n2204 ) | ( n1607 & n3266 ) | ( ~n2204 & n3266 ) ;
  assign n3268 = n2711 & ~n3267 ;
  assign n3269 = n598 | n1154 ;
  assign n3270 = n3268 & ~n3269 ;
  assign n3271 = ( n710 & n1246 ) | ( n710 & n1279 ) | ( n1246 & n1279 ) ;
  assign n3272 = x85 | n3271 ;
  assign n3273 = ( ~x69 & n1121 ) | ( ~x69 & n3272 ) | ( n1121 & n3272 ) ;
  assign n3274 = ( n588 & n1444 ) | ( n588 & ~n2187 ) | ( n1444 & ~n2187 ) ;
  assign n3275 = ~n3273 & n3274 ;
  assign n3276 = n3275 ^ n707 ^ 1'b0 ;
  assign n3277 = n1365 ^ x114 ^ 1'b0 ;
  assign n3278 = n352 | n3277 ;
  assign n3279 = n724 & n3278 ;
  assign n3280 = n3013 ^ x59 ^ 1'b0 ;
  assign n3281 = n1736 & ~n3280 ;
  assign n3282 = ( n708 & ~n2453 ) | ( n708 & n3281 ) | ( ~n2453 & n3281 ) ;
  assign n3283 = n624 & ~n1040 ;
  assign n3284 = n644 | n3283 ;
  assign n3285 = n3284 ^ n987 ^ 1'b0 ;
  assign n3288 = ~n1776 & n2793 ;
  assign n3286 = ( x48 & ~x64 ) | ( x48 & n456 ) | ( ~x64 & n456 ) ;
  assign n3287 = n3286 ^ n1234 ^ 1'b0 ;
  assign n3289 = n3288 ^ n3287 ^ n1989 ;
  assign n3290 = ( n537 & n3285 ) | ( n537 & n3289 ) | ( n3285 & n3289 ) ;
  assign n3291 = n1178 ^ n756 ^ 1'b0 ;
  assign n3292 = n3291 ^ n525 ^ 1'b0 ;
  assign n3293 = n986 & n3292 ;
  assign n3294 = n420 ^ x11 ^ 1'b0 ;
  assign n3295 = ~n3214 & n3294 ;
  assign n3296 = n1043 & ~n1139 ;
  assign n3297 = ( ~n3174 & n3295 ) | ( ~n3174 & n3296 ) | ( n3295 & n3296 ) ;
  assign n3298 = ~n434 & n1211 ;
  assign n3299 = n3298 ^ n1848 ^ 1'b0 ;
  assign n3300 = n1538 ^ n1319 ^ 1'b0 ;
  assign n3301 = ~n742 & n3300 ;
  assign n3302 = n485 ^ n376 ^ 1'b0 ;
  assign n3303 = ~n1018 & n3302 ;
  assign n3304 = n3303 ^ n1129 ^ n520 ;
  assign n3305 = n3301 & ~n3304 ;
  assign n3306 = n3305 ^ n2632 ^ 1'b0 ;
  assign n3307 = ( ~x18 & n157 ) | ( ~x18 & n2297 ) | ( n157 & n2297 ) ;
  assign n3308 = n176 & n3049 ;
  assign n3309 = ~n2692 & n3308 ;
  assign n3310 = ~n3307 & n3309 ;
  assign n3311 = n1776 | n2569 ;
  assign n3312 = n262 & n846 ;
  assign n3313 = n3312 ^ n1554 ^ 1'b0 ;
  assign n3314 = ~n447 & n3313 ;
  assign n3315 = n3151 ^ n3142 ^ 1'b0 ;
  assign n3316 = n1139 ^ n540 ^ x69 ;
  assign n3317 = n3316 ^ n905 ^ 1'b0 ;
  assign n3318 = ~n2233 & n3317 ;
  assign n3319 = ( ~x17 & n323 ) | ( ~x17 & n2679 ) | ( n323 & n2679 ) ;
  assign n3320 = n3304 ^ n1646 ^ 1'b0 ;
  assign n3321 = n3319 | n3320 ;
  assign n3322 = n1807 & ~n3321 ;
  assign n3325 = ~x52 & n1196 ;
  assign n3323 = n2232 & ~n2557 ;
  assign n3324 = ( ~n1201 & n3109 ) | ( ~n1201 & n3323 ) | ( n3109 & n3323 ) ;
  assign n3326 = n3325 ^ n3324 ^ n747 ;
  assign n3327 = x32 & ~n1838 ;
  assign n3328 = n3327 ^ n472 ^ 1'b0 ;
  assign n3329 = n2875 | n3328 ;
  assign n3330 = n3326 & ~n3329 ;
  assign n3331 = n2303 ^ n623 ^ n141 ;
  assign n3332 = n3331 ^ n1707 ^ 1'b0 ;
  assign n3333 = n3332 ^ n3272 ^ 1'b0 ;
  assign n3334 = ( n990 & n3089 ) | ( n990 & ~n3333 ) | ( n3089 & ~n3333 ) ;
  assign n3335 = n1807 | n2170 ;
  assign n3336 = n608 ^ n523 ^ 1'b0 ;
  assign n3337 = n2386 | n3336 ;
  assign n3338 = n2863 | n3337 ;
  assign n3339 = n3338 ^ n2839 ^ 1'b0 ;
  assign n3340 = n3207 | n3339 ;
  assign n3341 = ( n158 & ~n529 ) | ( n158 & n1860 ) | ( ~n529 & n1860 ) ;
  assign n3342 = n2596 ^ n1448 ^ 1'b0 ;
  assign n3343 = n3341 | n3342 ;
  assign n3344 = n704 & ~n1947 ;
  assign n3345 = n2779 & n3344 ;
  assign n3346 = ( n2638 & ~n3343 ) | ( n2638 & n3345 ) | ( ~n3343 & n3345 ) ;
  assign n3347 = n898 ^ n831 ^ 1'b0 ;
  assign n3353 = n1456 ^ n473 ^ 1'b0 ;
  assign n3354 = n3042 & ~n3353 ;
  assign n3348 = x19 | n871 ;
  assign n3349 = n820 | n3348 ;
  assign n3350 = n2000 ^ x119 ^ 1'b0 ;
  assign n3351 = n1697 | n3350 ;
  assign n3352 = ( n1986 & ~n3349 ) | ( n1986 & n3351 ) | ( ~n3349 & n3351 ) ;
  assign n3355 = n3354 ^ n3352 ^ 1'b0 ;
  assign n3356 = n245 | n2945 ;
  assign n3357 = n706 | n3356 ;
  assign n3358 = n3357 ^ n401 ^ 1'b0 ;
  assign n3359 = n3358 ^ n1289 ^ x121 ;
  assign n3360 = ( ~n1038 & n1692 ) | ( ~n1038 & n3359 ) | ( n1692 & n3359 ) ;
  assign n3361 = n1411 ^ n576 ^ 1'b0 ;
  assign n3362 = n339 & ~n3361 ;
  assign n3363 = ~n2789 & n3362 ;
  assign n3364 = n942 & ~n2801 ;
  assign n3365 = n241 ^ x25 ^ 1'b0 ;
  assign n3366 = n2223 & ~n3365 ;
  assign n3367 = n1027 ^ n626 ^ x98 ;
  assign n3368 = n756 & ~n1167 ;
  assign n3369 = n3368 ^ n1686 ^ 1'b0 ;
  assign n3370 = n3367 & ~n3369 ;
  assign n3371 = n3370 ^ n1891 ^ 1'b0 ;
  assign n3372 = n454 | n810 ;
  assign n3373 = n1624 & ~n3372 ;
  assign n3374 = n3373 ^ n2934 ^ n1858 ;
  assign n3375 = n3374 ^ n3013 ^ n371 ;
  assign n3376 = n3375 ^ n817 ^ 1'b0 ;
  assign n3377 = n187 | n808 ;
  assign n3378 = n3377 ^ n2793 ^ n2199 ;
  assign n3379 = ( n1879 & n2108 ) | ( n1879 & ~n3378 ) | ( n2108 & ~n3378 ) ;
  assign n3380 = ( n3371 & n3376 ) | ( n3371 & ~n3379 ) | ( n3376 & ~n3379 ) ;
  assign n3383 = n1082 ^ n464 ^ 1'b0 ;
  assign n3381 = n492 & ~n710 ;
  assign n3382 = n1253 & n3381 ;
  assign n3384 = n3383 ^ n3382 ^ n1984 ;
  assign n3385 = ~n1316 & n3384 ;
  assign n3386 = n1032 ^ n360 ^ n160 ;
  assign n3387 = n1940 ^ x21 ^ 1'b0 ;
  assign n3388 = n3386 & ~n3387 ;
  assign n3389 = n2371 ^ n1999 ^ 1'b0 ;
  assign n3390 = n1190 & n1814 ;
  assign n3391 = n1352 | n3390 ;
  assign n3395 = n858 & n2178 ;
  assign n3396 = n3395 ^ n442 ^ 1'b0 ;
  assign n3392 = n1400 | n1695 ;
  assign n3393 = n3392 ^ n479 ^ 1'b0 ;
  assign n3394 = ( n859 & ~n2494 ) | ( n859 & n3393 ) | ( ~n2494 & n3393 ) ;
  assign n3397 = n3396 ^ n3394 ^ 1'b0 ;
  assign n3398 = n157 & ~n3397 ;
  assign n3399 = n1929 ^ n1006 ^ n977 ;
  assign n3400 = n1316 ^ n334 ^ 1'b0 ;
  assign n3401 = n265 | n3400 ;
  assign n3402 = ( ~n1555 & n3399 ) | ( ~n1555 & n3401 ) | ( n3399 & n3401 ) ;
  assign n3403 = ( n1811 & ~n3223 ) | ( n1811 & n3402 ) | ( ~n3223 & n3402 ) ;
  assign n3406 = ( ~n213 & n875 ) | ( ~n213 & n2297 ) | ( n875 & n2297 ) ;
  assign n3404 = n550 & ~n1036 ;
  assign n3405 = n3404 ^ n559 ^ 1'b0 ;
  assign n3407 = n3406 ^ n3405 ^ 1'b0 ;
  assign n3408 = n1028 ^ n458 ^ 1'b0 ;
  assign n3409 = n597 | n3408 ;
  assign n3410 = ( ~x118 & n392 ) | ( ~x118 & n1894 ) | ( n392 & n1894 ) ;
  assign n3411 = n3410 ^ n974 ^ 1'b0 ;
  assign n3412 = n3411 ^ n1653 ^ 1'b0 ;
  assign n3413 = n1060 & ~n3412 ;
  assign n3414 = n3413 ^ n2689 ^ 1'b0 ;
  assign n3415 = ~n3409 & n3414 ;
  assign n3416 = ( ~n1359 & n2713 ) | ( ~n1359 & n2922 ) | ( n2713 & n2922 ) ;
  assign n3417 = ( n920 & n1113 ) | ( n920 & n2449 ) | ( n1113 & n2449 ) ;
  assign n3418 = n2063 ^ n1309 ^ n608 ;
  assign n3419 = n3418 ^ n2242 ^ n537 ;
  assign n3424 = n468 | n2792 ;
  assign n3422 = n1579 ^ n318 ^ x55 ;
  assign n3421 = n1405 ^ n696 ^ 1'b0 ;
  assign n3420 = n2472 ^ n1404 ^ n784 ;
  assign n3423 = n3422 ^ n3421 ^ n3420 ;
  assign n3425 = n3424 ^ n3423 ^ 1'b0 ;
  assign n3426 = ~n3419 & n3425 ;
  assign n3427 = n754 & ~n2035 ;
  assign n3428 = n3427 ^ n176 ^ 1'b0 ;
  assign n3429 = n3428 ^ n826 ^ 1'b0 ;
  assign n3430 = n1132 ^ n343 ^ 1'b0 ;
  assign n3431 = n334 & n3430 ;
  assign n3432 = n3431 ^ n1226 ^ 1'b0 ;
  assign n3435 = n2092 ^ x92 ^ 1'b0 ;
  assign n3436 = ~n468 & n3435 ;
  assign n3433 = n1573 ^ n866 ^ 1'b0 ;
  assign n3434 = n1104 & ~n3433 ;
  assign n3437 = n3436 ^ n3434 ^ 1'b0 ;
  assign n3438 = ( ~n470 & n1764 ) | ( ~n470 & n2674 ) | ( n1764 & n2674 ) ;
  assign n3439 = ( n253 & ~n2965 ) | ( n253 & n3438 ) | ( ~n2965 & n3438 ) ;
  assign n3440 = ( ~n3432 & n3437 ) | ( ~n3432 & n3439 ) | ( n3437 & n3439 ) ;
  assign n3441 = n722 ^ n194 ^ x50 ;
  assign n3442 = n3441 ^ n1077 ^ 1'b0 ;
  assign n3443 = n1629 | n2632 ;
  assign n3444 = ( ~n1252 & n1578 ) | ( ~n1252 & n2596 ) | ( n1578 & n2596 ) ;
  assign n3445 = n1781 & ~n1786 ;
  assign n3446 = ~n3444 & n3445 ;
  assign n3447 = n2818 ^ n447 ^ 1'b0 ;
  assign n3448 = n1033 ^ n946 ^ 1'b0 ;
  assign n3449 = ( ~n2468 & n3396 ) | ( ~n2468 & n3448 ) | ( n3396 & n3448 ) ;
  assign n3450 = n157 | n3449 ;
  assign n3451 = ( x31 & ~n424 ) | ( x31 & n783 ) | ( ~n424 & n783 ) ;
  assign n3452 = n3451 ^ n402 ^ 1'b0 ;
  assign n3453 = ~n1460 & n3452 ;
  assign n3454 = n3453 ^ n504 ^ 1'b0 ;
  assign n3455 = n2992 ^ n1547 ^ n703 ;
  assign n3456 = n1223 ^ n363 ^ 1'b0 ;
  assign n3457 = n3455 & ~n3456 ;
  assign n3458 = n685 | n1171 ;
  assign n3459 = n615 & ~n3458 ;
  assign n3460 = n3433 ^ n1647 ^ 1'b0 ;
  assign n3461 = n1410 & ~n3460 ;
  assign n3462 = ( n202 & n3459 ) | ( n202 & ~n3461 ) | ( n3459 & ~n3461 ) ;
  assign n3463 = n3462 ^ n912 ^ n893 ;
  assign n3464 = n3457 & n3463 ;
  assign n3465 = n3464 ^ n2481 ^ 1'b0 ;
  assign n3466 = x63 & n1469 ;
  assign n3467 = ~n1525 & n3466 ;
  assign n3471 = ( ~n238 & n384 ) | ( ~n238 & n1100 ) | ( n384 & n1100 ) ;
  assign n3468 = n3130 ^ x60 ^ 1'b0 ;
  assign n3469 = n2006 | n3468 ;
  assign n3470 = n3451 & ~n3469 ;
  assign n3472 = n3471 ^ n3470 ^ 1'b0 ;
  assign n3473 = n214 & n3472 ;
  assign n3474 = n3376 ^ n531 ^ 1'b0 ;
  assign n3475 = n3473 & ~n3474 ;
  assign n3476 = ( ~n699 & n1167 ) | ( ~n699 & n2665 ) | ( n1167 & n2665 ) ;
  assign n3479 = ~n1357 & n3072 ;
  assign n3477 = n2834 ^ n544 ^ 1'b0 ;
  assign n3478 = n666 & n3477 ;
  assign n3480 = n3479 ^ n3478 ^ 1'b0 ;
  assign n3481 = n1337 | n2480 ;
  assign n3482 = ( n197 & n321 ) | ( n197 & ~n364 ) | ( n321 & ~n364 ) ;
  assign n3483 = n1519 ^ n1455 ^ n663 ;
  assign n3484 = ( n924 & n3482 ) | ( n924 & n3483 ) | ( n3482 & n3483 ) ;
  assign n3485 = n3484 ^ n1449 ^ n1150 ;
  assign n3486 = ~n3481 & n3485 ;
  assign n3487 = ~n730 & n1490 ;
  assign n3488 = ~n3059 & n3487 ;
  assign n3489 = ( n844 & ~n1730 ) | ( n844 & n3488 ) | ( ~n1730 & n3488 ) ;
  assign n3490 = n455 & n807 ;
  assign n3491 = n3490 ^ n3362 ^ 1'b0 ;
  assign n3492 = ( n1139 & n3489 ) | ( n1139 & n3491 ) | ( n3489 & n3491 ) ;
  assign n3493 = n310 & n411 ;
  assign n3494 = x103 | n997 ;
  assign n3495 = x45 & n1673 ;
  assign n3496 = ~n3494 & n3495 ;
  assign n3497 = ~n3283 & n3496 ;
  assign n3498 = n3497 ^ n2202 ^ n1206 ;
  assign n3499 = n3498 ^ n1051 ^ 1'b0 ;
  assign n3500 = ( n1534 & ~n2557 ) | ( n1534 & n2947 ) | ( ~n2557 & n2947 ) ;
  assign n3501 = ( n425 & n1051 ) | ( n425 & ~n3500 ) | ( n1051 & ~n3500 ) ;
  assign n3502 = n2500 ^ n1769 ^ x72 ;
  assign n3503 = ( ~n2836 & n3501 ) | ( ~n2836 & n3502 ) | ( n3501 & n3502 ) ;
  assign n3504 = n3437 ^ n381 ^ 1'b0 ;
  assign n3505 = n3504 ^ n1628 ^ 1'b0 ;
  assign n3506 = n846 ^ n657 ^ n376 ;
  assign n3507 = n1723 & ~n3506 ;
  assign n3508 = ~n1409 & n3507 ;
  assign n3509 = ( ~n544 & n579 ) | ( ~n544 & n1086 ) | ( n579 & n1086 ) ;
  assign n3510 = ( n2095 & n3508 ) | ( n2095 & n3509 ) | ( n3508 & n3509 ) ;
  assign n3511 = n3354 ^ n1701 ^ n497 ;
  assign n3513 = n573 & n3031 ;
  assign n3512 = n275 | n2702 ;
  assign n3514 = n3513 ^ n3512 ^ 1'b0 ;
  assign n3515 = n1566 ^ n1138 ^ 1'b0 ;
  assign n3516 = ~n1529 & n3515 ;
  assign n3517 = n1661 & n3516 ;
  assign n3518 = n1082 ^ n804 ^ 1'b0 ;
  assign n3519 = n161 & ~n3518 ;
  assign n3520 = n3519 ^ n2104 ^ 1'b0 ;
  assign n3521 = n1268 | n3520 ;
  assign n3522 = n3517 | n3521 ;
  assign n3523 = n3514 & ~n3522 ;
  assign n3524 = ( n2705 & ~n3121 ) | ( n2705 & n3523 ) | ( ~n3121 & n3523 ) ;
  assign n3525 = n2715 | n3306 ;
  assign n3526 = n998 ^ n921 ^ 1'b0 ;
  assign n3527 = n559 | n3526 ;
  assign n3528 = n706 | n1202 ;
  assign n3529 = n2774 & ~n3528 ;
  assign n3530 = n584 & ~n1234 ;
  assign n3532 = n467 | n676 ;
  assign n3531 = n1796 & n2088 ;
  assign n3533 = n3532 ^ n3531 ^ 1'b0 ;
  assign n3534 = n354 & n2692 ;
  assign n3535 = ~n2008 & n3534 ;
  assign n3536 = ~n3533 & n3535 ;
  assign n3537 = n1032 & ~n1717 ;
  assign n3538 = n3537 ^ n3050 ^ 1'b0 ;
  assign n3539 = ~n1352 & n2536 ;
  assign n3540 = n3539 ^ n2074 ^ 1'b0 ;
  assign n3541 = n3538 | n3540 ;
  assign n3542 = n3541 ^ n1740 ^ 1'b0 ;
  assign n3543 = n2112 ^ n531 ^ 1'b0 ;
  assign n3544 = n3543 ^ n3334 ^ n1084 ;
  assign n3545 = n661 & ~n3100 ;
  assign n3546 = n984 & n3545 ;
  assign n3547 = ~n2204 & n2507 ;
  assign n3548 = ( x0 & ~n1726 ) | ( x0 & n3547 ) | ( ~n1726 & n3547 ) ;
  assign n3549 = x40 & ~n2220 ;
  assign n3550 = n379 & n3549 ;
  assign n3551 = n1246 ^ n508 ^ x28 ;
  assign n3552 = n3551 ^ n2722 ^ n759 ;
  assign n3553 = ( n338 & n482 ) | ( n338 & ~n1369 ) | ( n482 & ~n1369 ) ;
  assign n3556 = n3301 ^ n1733 ^ n1490 ;
  assign n3557 = ( ~n349 & n3488 ) | ( ~n349 & n3556 ) | ( n3488 & n3556 ) ;
  assign n3555 = ~n2870 & n3217 ;
  assign n3554 = n1640 ^ n544 ^ n250 ;
  assign n3558 = n3557 ^ n3555 ^ n3554 ;
  assign n3559 = ( n3552 & ~n3553 ) | ( n3552 & n3558 ) | ( ~n3553 & n3558 ) ;
  assign n3560 = n1870 ^ n318 ^ 1'b0 ;
  assign n3569 = ( n580 & n1209 ) | ( n580 & n3424 ) | ( n1209 & n3424 ) ;
  assign n3570 = n2033 & n2971 ;
  assign n3571 = ~n3569 & n3570 ;
  assign n3572 = n3571 ^ n1501 ^ 1'b0 ;
  assign n3561 = ( n230 & n488 ) | ( n230 & n1412 ) | ( n488 & n1412 ) ;
  assign n3562 = ( n715 & n1272 ) | ( n715 & n3561 ) | ( n1272 & n3561 ) ;
  assign n3563 = n3562 ^ n636 ^ 1'b0 ;
  assign n3564 = n3563 ^ x24 ^ 1'b0 ;
  assign n3565 = n1957 ^ n611 ^ n483 ;
  assign n3566 = ( n1849 & n1909 ) | ( n1849 & n3565 ) | ( n1909 & n3565 ) ;
  assign n3567 = n3566 ^ n3481 ^ n1384 ;
  assign n3568 = n3564 & n3567 ;
  assign n3573 = n3572 ^ n3568 ^ 1'b0 ;
  assign n3574 = n314 & ~n1317 ;
  assign n3575 = ( ~n1374 & n1653 ) | ( ~n1374 & n3574 ) | ( n1653 & n3574 ) ;
  assign n3576 = ( n1162 & ~n1286 ) | ( n1162 & n1521 ) | ( ~n1286 & n1521 ) ;
  assign n3577 = ~n1905 & n2505 ;
  assign n3578 = n3577 ^ n1125 ^ 1'b0 ;
  assign n3579 = n1636 ^ n464 ^ 1'b0 ;
  assign n3580 = ( n219 & ~n274 ) | ( n219 & n3579 ) | ( ~n274 & n3579 ) ;
  assign n3581 = ( ~n644 & n3578 ) | ( ~n644 & n3580 ) | ( n3578 & n3580 ) ;
  assign n3582 = ~n3100 & n3581 ;
  assign n3583 = n3582 ^ n1946 ^ n1640 ;
  assign n3584 = n1858 ^ n479 ^ n132 ;
  assign n3585 = ( n613 & n3583 ) | ( n613 & ~n3584 ) | ( n3583 & ~n3584 ) ;
  assign n3586 = n1333 ^ x34 ^ 1'b0 ;
  assign n3587 = n2295 | n3586 ;
  assign n3588 = ( ~n293 & n1578 ) | ( ~n293 & n2179 ) | ( n1578 & n2179 ) ;
  assign n3589 = n1498 | n2352 ;
  assign n3590 = n2131 | n3589 ;
  assign n3591 = ~n1274 & n3590 ;
  assign n3592 = ~n3588 & n3591 ;
  assign n3594 = n658 ^ n363 ^ 1'b0 ;
  assign n3595 = n2294 & n3594 ;
  assign n3593 = n806 | n3555 ;
  assign n3596 = n3595 ^ n3593 ^ 1'b0 ;
  assign n3597 = ( x63 & n325 ) | ( x63 & n605 ) | ( n325 & n605 ) ;
  assign n3598 = n3597 ^ n1851 ^ 1'b0 ;
  assign n3599 = ( n1391 & n1438 ) | ( n1391 & ~n1903 ) | ( n1438 & ~n1903 ) ;
  assign n3600 = ( n2702 & n3598 ) | ( n2702 & ~n3599 ) | ( n3598 & ~n3599 ) ;
  assign n3601 = n209 ^ n139 ^ 1'b0 ;
  assign n3602 = n1171 | n3601 ;
  assign n3603 = n2139 & ~n3602 ;
  assign n3604 = n3603 ^ n1975 ^ 1'b0 ;
  assign n3605 = ( n3442 & n3600 ) | ( n3442 & n3604 ) | ( n3600 & n3604 ) ;
  assign n3606 = n2834 ^ n2340 ^ x37 ;
  assign n3607 = n194 & n3606 ;
  assign n3608 = n3607 ^ n1581 ^ n1193 ;
  assign n3609 = n3496 ^ n3281 ^ 1'b0 ;
  assign n3610 = ~n454 & n3609 ;
  assign n3611 = ( n2507 & ~n2653 ) | ( n2507 & n2808 ) | ( ~n2653 & n2808 ) ;
  assign n3612 = n1907 ^ n1828 ^ n1100 ;
  assign n3613 = ( n332 & n1785 ) | ( n332 & n2339 ) | ( n1785 & n2339 ) ;
  assign n3614 = n1731 ^ n1392 ^ n490 ;
  assign n3615 = n3614 ^ n743 ^ 1'b0 ;
  assign n3616 = ~n2416 & n3615 ;
  assign n3617 = n3616 ^ n1624 ^ n861 ;
  assign n3618 = n1930 | n3617 ;
  assign n3619 = n3613 & ~n3618 ;
  assign n3620 = ( n577 & ~n3345 ) | ( n577 & n3619 ) | ( ~n3345 & n3619 ) ;
  assign n3621 = n1490 ^ n1391 ^ 1'b0 ;
  assign n3622 = n3621 ^ n1650 ^ 1'b0 ;
  assign n3624 = n1801 | n3328 ;
  assign n3625 = n1720 & n2898 ;
  assign n3626 = ( n1434 & ~n3624 ) | ( n1434 & n3625 ) | ( ~n3624 & n3625 ) ;
  assign n3627 = ~n2354 & n3390 ;
  assign n3628 = ~n3626 & n3627 ;
  assign n3623 = ~n770 & n2420 ;
  assign n3629 = n3628 ^ n3623 ^ 1'b0 ;
  assign n3630 = n807 ^ n293 ^ 1'b0 ;
  assign n3631 = n3255 ^ n3077 ^ 1'b0 ;
  assign n3639 = n316 & ~n348 ;
  assign n3640 = n3639 ^ n442 ^ 1'b0 ;
  assign n3641 = n3640 ^ n2328 ^ n2143 ;
  assign n3642 = n2363 ^ n1982 ^ 1'b0 ;
  assign n3643 = ( n2334 & n3641 ) | ( n2334 & n3642 ) | ( n3641 & n3642 ) ;
  assign n3632 = n1027 & ~n1920 ;
  assign n3633 = ( ~n167 & n2766 ) | ( ~n167 & n3632 ) | ( n2766 & n3632 ) ;
  assign n3634 = n874 ^ x9 ^ 1'b0 ;
  assign n3635 = n3634 ^ n206 ^ 1'b0 ;
  assign n3636 = n3635 ^ n2417 ^ 1'b0 ;
  assign n3637 = n327 & ~n3636 ;
  assign n3638 = n3633 | n3637 ;
  assign n3644 = n3643 ^ n3638 ^ 1'b0 ;
  assign n3645 = n1517 ^ n1420 ^ 1'b0 ;
  assign n3646 = n3645 ^ n3383 ^ n3254 ;
  assign n3647 = ~n628 & n915 ;
  assign n3648 = ~n2724 & n3647 ;
  assign n3649 = ( ~n680 & n1268 ) | ( ~n680 & n2340 ) | ( n1268 & n2340 ) ;
  assign n3650 = ~n3358 & n3649 ;
  assign n3651 = n3212 ^ n2766 ^ 1'b0 ;
  assign n3652 = n3650 & ~n3651 ;
  assign n3653 = n3652 ^ n2027 ^ 1'b0 ;
  assign n3654 = ~n3648 & n3653 ;
  assign n3655 = n1211 & ~n1235 ;
  assign n3656 = n2522 ^ n2480 ^ x37 ;
  assign n3657 = ( n1862 & ~n2184 ) | ( n1862 & n3656 ) | ( ~n2184 & n3656 ) ;
  assign n3658 = n3657 ^ n3546 ^ 1'b0 ;
  assign n3660 = n953 ^ n402 ^ 1'b0 ;
  assign n3659 = ~n207 & n2834 ;
  assign n3661 = n3660 ^ n3659 ^ 1'b0 ;
  assign n3662 = n1198 & ~n3455 ;
  assign n3663 = n812 ^ x62 ^ 1'b0 ;
  assign n3664 = n3662 | n3663 ;
  assign n3665 = n3664 ^ n1004 ^ 1'b0 ;
  assign n3666 = n3287 & ~n3665 ;
  assign n3667 = n2344 ^ n2050 ^ 1'b0 ;
  assign n3668 = n3666 & n3667 ;
  assign n3669 = ~n3661 & n3668 ;
  assign n3670 = ~n986 & n3669 ;
  assign n3671 = n2447 ^ n1548 ^ 1'b0 ;
  assign n3672 = ~n2178 & n3671 ;
  assign n3676 = x93 & n1426 ;
  assign n3677 = n3676 ^ n652 ^ 1'b0 ;
  assign n3678 = ( ~n160 & n2014 ) | ( ~n160 & n3677 ) | ( n2014 & n3677 ) ;
  assign n3673 = n161 & ~n1341 ;
  assign n3674 = n3673 ^ n1037 ^ 1'b0 ;
  assign n3675 = ~n1037 & n3674 ;
  assign n3679 = n3678 ^ n3675 ^ 1'b0 ;
  assign n3680 = n3679 ^ n1333 ^ n643 ;
  assign n3681 = n808 ^ n370 ^ 1'b0 ;
  assign n3682 = n1883 | n3681 ;
  assign n3683 = ~n727 & n2014 ;
  assign n3684 = ~x86 & n3683 ;
  assign n3685 = ( ~n357 & n517 ) | ( ~n357 & n2376 ) | ( n517 & n2376 ) ;
  assign n3686 = ( ~n2473 & n3684 ) | ( ~n2473 & n3685 ) | ( n3684 & n3685 ) ;
  assign n3687 = n3686 ^ n2851 ^ x77 ;
  assign n3688 = ~n874 & n2383 ;
  assign n3689 = n3688 ^ n3506 ^ n1658 ;
  assign n3690 = n643 | n1329 ;
  assign n3691 = x12 | n3690 ;
  assign n3692 = n3691 ^ n1208 ^ n412 ;
  assign n3693 = n3689 & n3692 ;
  assign n3694 = ~n2634 & n3693 ;
  assign n3695 = n784 & ~n2671 ;
  assign n3696 = n1597 & n3695 ;
  assign n3697 = ~n3694 & n3696 ;
  assign n3698 = ( n1612 & ~n2493 ) | ( n1612 & n3424 ) | ( ~n2493 & n3424 ) ;
  assign n3699 = n3674 ^ n1304 ^ n529 ;
  assign n3700 = ( ~n2423 & n3572 ) | ( ~n2423 & n3699 ) | ( n3572 & n3699 ) ;
  assign n3701 = n1640 | n3700 ;
  assign n3702 = n1028 & ~n1209 ;
  assign n3703 = ~n2160 & n3702 ;
  assign n3704 = n1129 ^ n967 ^ 1'b0 ;
  assign n3705 = ~n3214 & n3704 ;
  assign n3706 = n3703 & n3705 ;
  assign n3712 = n1555 ^ n1083 ^ 1'b0 ;
  assign n3708 = x97 & ~n465 ;
  assign n3709 = n3708 ^ n2340 ^ 1'b0 ;
  assign n3710 = n470 & ~n3709 ;
  assign n3707 = ~n2303 & n3191 ;
  assign n3711 = n3710 ^ n3707 ^ 1'b0 ;
  assign n3713 = n3712 ^ n3711 ^ 1'b0 ;
  assign n3718 = n1194 & n2623 ;
  assign n3714 = n2033 & ~n3070 ;
  assign n3715 = ~n267 & n3714 ;
  assign n3716 = ~n473 & n3715 ;
  assign n3717 = n945 & ~n3716 ;
  assign n3719 = n3718 ^ n3717 ^ 1'b0 ;
  assign n3720 = ( ~n384 & n1518 ) | ( ~n384 & n1637 ) | ( n1518 & n1637 ) ;
  assign n3721 = n3720 ^ n2774 ^ n2153 ;
  assign n3722 = n1838 | n3721 ;
  assign n3723 = ( n1434 & n1679 ) | ( n1434 & ~n2173 ) | ( n1679 & ~n2173 ) ;
  assign n3724 = n454 & n3723 ;
  assign n3725 = n218 & n983 ;
  assign n3726 = n1003 | n1695 ;
  assign n3727 = n1413 & ~n3726 ;
  assign n3728 = ~n2195 & n3727 ;
  assign n3729 = ( n1558 & n3386 ) | ( n1558 & n3517 ) | ( n3386 & n3517 ) ;
  assign n3730 = n3728 & ~n3729 ;
  assign n3731 = n3725 & n3730 ;
  assign n3732 = n1426 ^ n855 ^ n270 ;
  assign n3733 = ~n331 & n3732 ;
  assign n3734 = n3731 & n3733 ;
  assign n3736 = n550 ^ n301 ^ 1'b0 ;
  assign n3735 = n1444 & ~n1587 ;
  assign n3737 = n3736 ^ n3735 ^ 1'b0 ;
  assign n3738 = ( x81 & n1217 ) | ( x81 & ~n1301 ) | ( n1217 & ~n1301 ) ;
  assign n3739 = n3738 ^ n1418 ^ x55 ;
  assign n3740 = n3739 ^ n613 ^ n227 ;
  assign n3741 = ( ~n844 & n1642 ) | ( ~n844 & n2494 ) | ( n1642 & n2494 ) ;
  assign n3742 = n783 | n1861 ;
  assign n3743 = n3741 & n3742 ;
  assign n3744 = n3740 & n3743 ;
  assign n3745 = n293 ^ n287 ^ 1'b0 ;
  assign n3746 = n1484 | n3745 ;
  assign n3747 = n3746 ^ n1986 ^ 1'b0 ;
  assign n3748 = ( n1753 & n3161 ) | ( n1753 & ~n3747 ) | ( n3161 & ~n3747 ) ;
  assign n3749 = n1852 ^ n1114 ^ n477 ;
  assign n3750 = n3749 ^ n1212 ^ n1189 ;
  assign n3751 = n1921 & ~n3750 ;
  assign n3752 = ( n171 & ~n2161 ) | ( n171 & n3751 ) | ( ~n2161 & n3751 ) ;
  assign n3753 = n2076 ^ n1225 ^ n1060 ;
  assign n3754 = ( ~n728 & n1074 ) | ( ~n728 & n3753 ) | ( n1074 & n3753 ) ;
  assign n3755 = n873 | n2865 ;
  assign n3756 = n502 & ~n3755 ;
  assign n3757 = n3756 ^ n3084 ^ n1212 ;
  assign n3762 = n861 ^ n656 ^ 1'b0 ;
  assign n3760 = x48 & n1647 ;
  assign n3761 = ~n188 & n3760 ;
  assign n3758 = n987 & n1173 ;
  assign n3759 = n3758 ^ n200 ^ 1'b0 ;
  assign n3763 = n3762 ^ n3761 ^ n3759 ;
  assign n3764 = n3763 ^ n199 ^ 1'b0 ;
  assign n3765 = n1974 ^ n1574 ^ 1'b0 ;
  assign n3766 = n2867 | n3765 ;
  assign n3767 = n1996 & ~n3766 ;
  assign n3768 = ~n1840 & n3767 ;
  assign n3769 = ( ~n1143 & n2655 ) | ( ~n1143 & n3768 ) | ( n2655 & n3768 ) ;
  assign n3773 = n2460 ^ n1802 ^ 1'b0 ;
  assign n3774 = n1003 | n3773 ;
  assign n3770 = ( n206 & n1156 ) | ( n206 & ~n2606 ) | ( n1156 & ~n2606 ) ;
  assign n3771 = n3770 ^ n717 ^ 1'b0 ;
  assign n3772 = n971 | n3771 ;
  assign n3775 = n3774 ^ n3772 ^ 1'b0 ;
  assign n3776 = n3709 ^ n3515 ^ n1743 ;
  assign n3777 = n3629 & n3776 ;
  assign n3778 = ( ~n157 & n368 ) | ( ~n157 & n1070 ) | ( n368 & n1070 ) ;
  assign n3779 = ~n703 & n3778 ;
  assign n3780 = ~n3432 & n3779 ;
  assign n3781 = n3560 ^ n983 ^ 1'b0 ;
  assign n3782 = n3583 ^ n314 ^ 1'b0 ;
  assign n3783 = n2522 | n3782 ;
  assign n3784 = n3783 ^ n2860 ^ 1'b0 ;
  assign n3785 = n3656 ^ n989 ^ 1'b0 ;
  assign n3786 = n1839 & n3785 ;
  assign n3787 = n428 ^ n380 ^ x118 ;
  assign n3788 = ( n531 & ~n747 ) | ( n531 & n3787 ) | ( ~n747 & n3787 ) ;
  assign n3789 = n2072 | n3214 ;
  assign n3790 = n3789 ^ n970 ^ 1'b0 ;
  assign n3791 = ~n927 & n3569 ;
  assign n3792 = n149 & ~n1583 ;
  assign n3793 = n3792 ^ n697 ^ 1'b0 ;
  assign n3794 = x115 | n208 ;
  assign n3795 = n3794 ^ n2596 ^ 1'b0 ;
  assign n3796 = ~n1366 & n3795 ;
  assign n3797 = n2717 ^ n457 ^ 1'b0 ;
  assign n3798 = n3406 ^ n431 ^ 1'b0 ;
  assign n3799 = n1159 & n2571 ;
  assign n3800 = n504 & n1002 ;
  assign n3801 = n3799 & n3800 ;
  assign n3802 = n2295 ^ n1094 ^ 1'b0 ;
  assign n3803 = n1270 & n1896 ;
  assign n3804 = ~n2386 & n3803 ;
  assign n3805 = ~x57 & n3804 ;
  assign n3806 = n3802 & n3805 ;
  assign n3807 = n842 ^ n149 ^ 1'b0 ;
  assign n3808 = n3807 ^ n2463 ^ 1'b0 ;
  assign n3809 = ( ~n863 & n3183 ) | ( ~n863 & n3808 ) | ( n3183 & n3808 ) ;
  assign n3810 = n618 & ~n1993 ;
  assign n3811 = n3810 ^ n402 ^ 1'b0 ;
  assign n3812 = n611 & ~n3811 ;
  assign n3813 = n2181 & ~n2939 ;
  assign n3814 = n3813 ^ n2025 ^ 1'b0 ;
  assign n3815 = n3812 | n3814 ;
  assign n3816 = n3815 ^ n1270 ^ n855 ;
  assign n3817 = ( n1020 & ~n1656 ) | ( n1020 & n2555 ) | ( ~n1656 & n2555 ) ;
  assign n3818 = ~n402 & n1343 ;
  assign n3819 = n3817 & n3818 ;
  assign n3820 = n1547 & ~n3819 ;
  assign n3821 = n3820 ^ x62 ^ 1'b0 ;
  assign n3822 = n1370 & n3821 ;
  assign n3823 = ( ~n174 & n1590 ) | ( ~n174 & n2799 ) | ( n1590 & n2799 ) ;
  assign n3828 = n3694 ^ n2251 ^ n1481 ;
  assign n3827 = n2631 ^ n2564 ^ 1'b0 ;
  assign n3825 = n2424 | n2776 ;
  assign n3824 = ( n1223 & ~n2006 ) | ( n1223 & n2697 ) | ( ~n2006 & n2697 ) ;
  assign n3826 = n3825 ^ n3824 ^ n755 ;
  assign n3829 = n3828 ^ n3827 ^ n3826 ;
  assign n3830 = n167 | n3100 ;
  assign n3832 = ( n678 & ~n1004 ) | ( n678 & n1818 ) | ( ~n1004 & n1818 ) ;
  assign n3831 = n2901 & ~n3811 ;
  assign n3833 = n3832 ^ n3831 ^ n203 ;
  assign n3834 = n3833 ^ n449 ^ 1'b0 ;
  assign n3835 = n3450 & ~n3834 ;
  assign n3836 = n2882 & ~n3835 ;
  assign n3837 = n495 & ~n3632 ;
  assign n3838 = n3496 | n3837 ;
  assign n3849 = n232 | n1182 ;
  assign n3850 = n3849 ^ n672 ^ 1'b0 ;
  assign n3841 = n132 | n294 ;
  assign n3839 = n1686 & n2516 ;
  assign n3840 = ~n694 & n3839 ;
  assign n3842 = n3841 ^ n3840 ^ n3341 ;
  assign n3843 = n169 & n2960 ;
  assign n3844 = n3843 ^ n479 ^ 1'b0 ;
  assign n3845 = ~n1419 & n3844 ;
  assign n3846 = n3845 ^ n262 ^ 1'b0 ;
  assign n3847 = n3842 | n3846 ;
  assign n3848 = n3847 ^ n555 ^ x18 ;
  assign n3851 = n3850 ^ n3848 ^ n2541 ;
  assign n3852 = x92 & ~n1007 ;
  assign n3853 = n3852 ^ n1496 ^ 1'b0 ;
  assign n3854 = ~n755 & n3853 ;
  assign n3855 = ~n2304 & n3045 ;
  assign n3856 = n1863 & n3855 ;
  assign n3862 = n3496 ^ n196 ^ 1'b0 ;
  assign n3863 = n3862 ^ n1801 ^ 1'b0 ;
  assign n3864 = ~n2083 & n3863 ;
  assign n3857 = n1617 ^ n595 ^ n455 ;
  assign n3858 = n3688 ^ n3441 ^ n227 ;
  assign n3859 = n3858 ^ n979 ^ 1'b0 ;
  assign n3860 = n3055 & ~n3859 ;
  assign n3861 = n3857 & n3860 ;
  assign n3865 = n3864 ^ n3861 ^ x57 ;
  assign n3866 = n1887 & n3443 ;
  assign n3867 = n3866 ^ n1581 ^ 1'b0 ;
  assign n3868 = n1794 | n2481 ;
  assign n3869 = n1270 | n3868 ;
  assign n3870 = n1121 ^ n238 ^ 1'b0 ;
  assign n3871 = n840 ^ n487 ^ 1'b0 ;
  assign n3872 = n204 & ~n3871 ;
  assign n3873 = n3872 ^ n3507 ^ 1'b0 ;
  assign n3874 = n2283 & n3873 ;
  assign n3875 = n3874 ^ n3869 ^ 1'b0 ;
  assign n3876 = n3870 & n3875 ;
  assign n3877 = ~n3869 & n3876 ;
  assign n3878 = n3120 | n3684 ;
  assign n3879 = n3878 ^ n2789 ^ 1'b0 ;
  assign n3880 = n3877 | n3879 ;
  assign n3881 = n3880 ^ n3580 ^ 1'b0 ;
  assign n3882 = n227 & ~n576 ;
  assign n3883 = ~n3169 & n3882 ;
  assign n3884 = n3070 | n3883 ;
  assign n3885 = n3884 ^ n1199 ^ 1'b0 ;
  assign n3886 = n1410 & ~n3885 ;
  assign n3887 = n1223 & n3886 ;
  assign n3888 = ( n662 & n1460 ) | ( n662 & n2224 ) | ( n1460 & n2224 ) ;
  assign n3889 = ( n1661 & ~n2572 ) | ( n1661 & n3888 ) | ( ~n2572 & n3888 ) ;
  assign n3890 = n3889 ^ n2070 ^ n1845 ;
  assign n3891 = n636 & n2521 ;
  assign n3892 = n3891 ^ n867 ^ 1'b0 ;
  assign n3893 = n1784 & ~n3892 ;
  assign n3894 = n1893 ^ x5 ^ 1'b0 ;
  assign n3895 = n647 ^ n260 ^ x93 ;
  assign n3896 = n574 ^ n511 ^ 1'b0 ;
  assign n3897 = ( n1378 & n3895 ) | ( n1378 & ~n3896 ) | ( n3895 & ~n3896 ) ;
  assign n3899 = x127 & n1480 ;
  assign n3898 = n1282 | n2758 ;
  assign n3900 = n3899 ^ n3898 ^ 1'b0 ;
  assign n3901 = n1585 ^ n1077 ^ 1'b0 ;
  assign n3902 = ~n3900 & n3901 ;
  assign n3903 = n1336 ^ n1141 ^ n251 ;
  assign n3904 = n1666 & n3903 ;
  assign n3905 = n3904 ^ n1686 ^ n979 ;
  assign n3906 = n2949 & n3905 ;
  assign n3907 = ~n3902 & n3906 ;
  assign n3908 = n830 | n3089 ;
  assign n3909 = n703 & ~n3908 ;
  assign n3910 = n3362 ^ n2104 ^ 1'b0 ;
  assign n3911 = n3909 | n3910 ;
  assign n3912 = n2552 ^ n269 ^ 1'b0 ;
  assign n3913 = n3911 | n3912 ;
  assign n3914 = n1764 & ~n3913 ;
  assign n3915 = n363 & n3914 ;
  assign n3916 = ~n211 & n1559 ;
  assign n3917 = ~n2057 & n3916 ;
  assign n3918 = n1272 | n3917 ;
  assign n3919 = n1548 | n3918 ;
  assign n3920 = n3919 ^ n1266 ^ 1'b0 ;
  assign n3921 = n2508 & n3920 ;
  assign n3922 = ~n275 & n316 ;
  assign n3923 = n3922 ^ n576 ^ 1'b0 ;
  assign n3924 = n3923 ^ n1348 ^ n1076 ;
  assign n3925 = n539 | n3924 ;
  assign n3926 = n1388 & ~n2340 ;
  assign n3927 = n1290 & ~n2563 ;
  assign n3931 = ~n808 & n3553 ;
  assign n3932 = ~n838 & n3931 ;
  assign n3933 = n2404 | n3932 ;
  assign n3934 = n3933 ^ n3288 ^ 1'b0 ;
  assign n3928 = n676 ^ x52 ^ 1'b0 ;
  assign n3929 = ~n1185 & n3928 ;
  assign n3930 = n3929 ^ n2606 ^ 1'b0 ;
  assign n3935 = n3934 ^ n3930 ^ n202 ;
  assign n3937 = n1134 | n1619 ;
  assign n3938 = n1743 | n3937 ;
  assign n3936 = ~n1205 & n1821 ;
  assign n3939 = n3938 ^ n3936 ^ 1'b0 ;
  assign n3940 = n2587 | n3939 ;
  assign n3941 = ~n493 & n1236 ;
  assign n3942 = n3941 ^ n2581 ^ 1'b0 ;
  assign n3943 = n1342 ^ n204 ^ 1'b0 ;
  assign n3944 = n3943 ^ n1205 ^ 1'b0 ;
  assign n3945 = ( n380 & n1785 ) | ( n380 & n2798 ) | ( n1785 & n2798 ) ;
  assign n3946 = n3945 ^ n1079 ^ x1 ;
  assign n3947 = ~n2835 & n3946 ;
  assign n3948 = ( ~n1364 & n1777 ) | ( ~n1364 & n2539 ) | ( n1777 & n2539 ) ;
  assign n3949 = ( n2200 & n3099 ) | ( n2200 & ~n3948 ) | ( n3099 & ~n3948 ) ;
  assign n3950 = n1247 ^ n264 ^ 1'b0 ;
  assign n3951 = ( n164 & ~n537 ) | ( n164 & n3950 ) | ( ~n537 & n3950 ) ;
  assign n3952 = ~n1851 & n3951 ;
  assign n3953 = n3664 ^ n1485 ^ 1'b0 ;
  assign n3954 = n2676 & n3953 ;
  assign n3955 = n3954 ^ n1898 ^ 1'b0 ;
  assign n3956 = ( n3020 & n3817 ) | ( n3020 & n3826 ) | ( n3817 & n3826 ) ;
  assign n3957 = n2528 ^ n1131 ^ 1'b0 ;
  assign n3958 = n132 & n3957 ;
  assign n3959 = n3958 ^ n569 ^ 1'b0 ;
  assign n3960 = n3959 ^ n1252 ^ 1'b0 ;
  assign n3961 = n3956 | n3960 ;
  assign n3962 = n1032 ^ n1002 ^ 1'b0 ;
  assign n3963 = n2778 ^ n1738 ^ 1'b0 ;
  assign n3964 = ~n685 & n3963 ;
  assign n3965 = n3964 ^ n2711 ^ n1074 ;
  assign n3966 = n3965 ^ n1413 ^ 1'b0 ;
  assign n3967 = n915 | n968 ;
  assign n3968 = n875 | n3967 ;
  assign n3970 = n2499 ^ n936 ^ 1'b0 ;
  assign n3969 = n1509 | n2605 ;
  assign n3971 = n3970 ^ n3969 ^ 1'b0 ;
  assign n3972 = ( n3246 & n3968 ) | ( n3246 & ~n3971 ) | ( n3968 & ~n3971 ) ;
  assign n3973 = n1894 ^ n334 ^ 1'b0 ;
  assign n3974 = n2398 ^ n1472 ^ n1410 ;
  assign n3975 = n3974 ^ n1104 ^ n796 ;
  assign n3976 = n2587 | n3975 ;
  assign n3981 = x101 & ~n1046 ;
  assign n3982 = n3981 ^ n831 ^ 1'b0 ;
  assign n3983 = n3982 ^ x63 ^ 1'b0 ;
  assign n3984 = n2160 & n3983 ;
  assign n3985 = n3984 ^ x13 ^ 1'b0 ;
  assign n3978 = n1059 | n1290 ;
  assign n3979 = n316 | n3978 ;
  assign n3977 = n2522 ^ n1591 ^ x111 ;
  assign n3980 = n3979 ^ n3977 ^ 1'b0 ;
  assign n3986 = n3985 ^ n3980 ^ 1'b0 ;
  assign n3989 = x70 & n943 ;
  assign n3990 = n3989 ^ n1689 ^ 1'b0 ;
  assign n3987 = n2401 | n2518 ;
  assign n3988 = n3987 ^ n2305 ^ 1'b0 ;
  assign n3991 = n3990 ^ n3988 ^ 1'b0 ;
  assign n3992 = ~n2683 & n2895 ;
  assign n3993 = n1117 & n2224 ;
  assign n3994 = n3993 ^ n1312 ^ 1'b0 ;
  assign n3995 = n167 & ~n1061 ;
  assign n3996 = n3995 ^ n1647 ^ 1'b0 ;
  assign n3997 = n3536 ^ n3378 ^ 1'b0 ;
  assign n3998 = ~n3996 & n3997 ;
  assign n3999 = ~n3016 & n3998 ;
  assign n4000 = ( n774 & n3994 ) | ( n774 & ~n3999 ) | ( n3994 & ~n3999 ) ;
  assign n4001 = n474 & n789 ;
  assign n4002 = ~n1801 & n4001 ;
  assign n4003 = n1503 ^ n396 ^ 1'b0 ;
  assign n4004 = n1915 | n4003 ;
  assign n4005 = n3761 ^ n3459 ^ n3015 ;
  assign n4006 = ( n844 & ~n4004 ) | ( n844 & n4005 ) | ( ~n4004 & n4005 ) ;
  assign n4007 = n2460 & n2860 ;
  assign n4008 = n4007 ^ n3416 ^ n1454 ;
  assign n4009 = n2313 & n2473 ;
  assign n4010 = n4009 ^ n1838 ^ 1'b0 ;
  assign n4011 = ~n867 & n2179 ;
  assign n4012 = n4011 ^ n1162 ^ 1'b0 ;
  assign n4013 = ( n205 & ~n3124 ) | ( n205 & n4012 ) | ( ~n3124 & n4012 ) ;
  assign n4014 = n4013 ^ n287 ^ 1'b0 ;
  assign n4015 = n4014 ^ n2262 ^ n2153 ;
  assign n4016 = n299 & n4015 ;
  assign n4017 = ~n4010 & n4016 ;
  assign n4020 = ~n134 & n2900 ;
  assign n4021 = n3621 & n4020 ;
  assign n4018 = ~n1072 & n2692 ;
  assign n4019 = n4018 ^ n3536 ^ 1'b0 ;
  assign n4022 = n4021 ^ n4019 ^ n3844 ;
  assign n4023 = n4022 ^ n2376 ^ n689 ;
  assign n4024 = n691 & ~n1535 ;
  assign n4025 = n4024 ^ n943 ^ 1'b0 ;
  assign n4026 = n3285 | n4025 ;
  assign n4030 = n632 ^ n528 ^ 1'b0 ;
  assign n4027 = n878 & n1319 ;
  assign n4028 = n759 & n4027 ;
  assign n4029 = n4028 ^ n1669 ^ n838 ;
  assign n4031 = n4030 ^ n4029 ^ 1'b0 ;
  assign n4032 = n1936 | n4031 ;
  assign n4033 = n1469 ^ n813 ^ 1'b0 ;
  assign n4034 = n4033 ^ n2654 ^ n2090 ;
  assign n4037 = ~n1697 & n2251 ;
  assign n4038 = n4037 ^ n2824 ^ 1'b0 ;
  assign n4035 = n3903 ^ n883 ^ 1'b0 ;
  assign n4036 = n1430 & ~n4035 ;
  assign n4039 = n4038 ^ n4036 ^ n2553 ;
  assign n4042 = n655 & ~n1630 ;
  assign n4040 = ~n1718 & n2587 ;
  assign n4041 = n2468 & n4040 ;
  assign n4043 = n4042 ^ n4041 ^ n1573 ;
  assign n4044 = ( n1774 & ~n1935 ) | ( n1774 & n4043 ) | ( ~n1935 & n4043 ) ;
  assign n4045 = n889 ^ n775 ^ 1'b0 ;
  assign n4046 = n1316 | n3671 ;
  assign n4047 = n4046 ^ n2562 ^ 1'b0 ;
  assign n4048 = ~n601 & n4047 ;
  assign n4049 = ( ~n1429 & n2653 ) | ( ~n1429 & n4048 ) | ( n2653 & n4048 ) ;
  assign n4050 = n4045 & ~n4049 ;
  assign n4051 = n3087 ^ n1629 ^ n1406 ;
  assign n4052 = ( x22 & n760 ) | ( x22 & ~n2881 ) | ( n760 & ~n2881 ) ;
  assign n4053 = ( ~n3031 & n3473 ) | ( ~n3031 & n4052 ) | ( n3473 & n4052 ) ;
  assign n4054 = n1417 ^ n984 ^ 1'b0 ;
  assign n4055 = n3152 & ~n4054 ;
  assign n4056 = ~n3384 & n4055 ;
  assign n4057 = ~n4053 & n4056 ;
  assign n4058 = n4057 ^ n4030 ^ n2390 ;
  assign n4059 = x38 & ~n985 ;
  assign n4060 = n4059 ^ n3858 ^ n1068 ;
  assign n4061 = x77 | n1399 ;
  assign n4062 = n2416 ^ n492 ^ 1'b0 ;
  assign n4063 = n2836 & n3953 ;
  assign n4064 = ( x0 & n4062 ) | ( x0 & n4063 ) | ( n4062 & n4063 ) ;
  assign n4065 = n301 & ~n831 ;
  assign n4066 = n4065 ^ n3664 ^ 1'b0 ;
  assign n4067 = n4066 ^ n3134 ^ n1154 ;
  assign n4068 = ( n732 & ~n848 ) | ( n732 & n1586 ) | ( ~n848 & n1586 ) ;
  assign n4069 = n4068 ^ n1100 ^ n813 ;
  assign n4070 = ( n208 & n4067 ) | ( n208 & ~n4069 ) | ( n4067 & ~n4069 ) ;
  assign n4071 = n141 & n4070 ;
  assign n4072 = ( n1069 & n1273 ) | ( n1069 & n2368 ) | ( n1273 & n2368 ) ;
  assign n4073 = ( n570 & ~n1221 ) | ( n570 & n1893 ) | ( ~n1221 & n1893 ) ;
  assign n4074 = n4073 ^ n3341 ^ 1'b0 ;
  assign n4075 = ~n2787 & n4074 ;
  assign n4076 = n809 & n3050 ;
  assign n4077 = n4076 ^ n915 ^ 1'b0 ;
  assign n4078 = n4077 ^ n791 ^ n563 ;
  assign n4079 = n897 & n4078 ;
  assign n4080 = n643 & n4079 ;
  assign n4081 = ( n1885 & n2061 ) | ( n1885 & ~n4080 ) | ( n2061 & ~n4080 ) ;
  assign n4082 = n378 | n2244 ;
  assign n4083 = n3606 ^ n1388 ^ n451 ;
  assign n4084 = ( n2779 & n4082 ) | ( n2779 & ~n4083 ) | ( n4082 & ~n4083 ) ;
  assign n4086 = n3075 ^ n2197 ^ n1654 ;
  assign n4085 = n266 & ~n2673 ;
  assign n4087 = n4086 ^ n4085 ^ n1165 ;
  assign n4088 = n1196 & n2165 ;
  assign n4089 = n4088 ^ n296 ^ 1'b0 ;
  assign n4090 = ( n1271 & n3455 ) | ( n1271 & ~n4089 ) | ( n3455 & ~n4089 ) ;
  assign n4091 = x57 & n2543 ;
  assign n4092 = ( n2071 & n4090 ) | ( n2071 & ~n4091 ) | ( n4090 & ~n4091 ) ;
  assign n4093 = n165 | n2965 ;
  assign n4094 = n837 | n1198 ;
  assign n4095 = n4094 ^ n2558 ^ 1'b0 ;
  assign n4096 = n994 | n4095 ;
  assign n4103 = n1221 ^ n322 ^ 1'b0 ;
  assign n4104 = n545 & ~n3579 ;
  assign n4105 = n4103 & n4104 ;
  assign n4097 = ( n248 & ~n544 ) | ( n248 & n1870 ) | ( ~n544 & n1870 ) ;
  assign n4098 = n4097 ^ n3144 ^ n696 ;
  assign n4100 = ( n739 & ~n905 ) | ( n739 & n1578 ) | ( ~n905 & n1578 ) ;
  assign n4099 = ( ~n1686 & n1913 ) | ( ~n1686 & n4020 ) | ( n1913 & n4020 ) ;
  assign n4101 = n4100 ^ n4099 ^ n1223 ;
  assign n4102 = n4098 & n4101 ;
  assign n4106 = n4105 ^ n4102 ^ 1'b0 ;
  assign n4107 = ( n2805 & ~n4096 ) | ( n2805 & n4106 ) | ( ~n4096 & n4106 ) ;
  assign n4108 = n1468 ^ n455 ^ n363 ;
  assign n4109 = n908 & ~n2008 ;
  assign n4110 = n1062 & ~n3592 ;
  assign n4111 = ( n136 & n822 ) | ( n136 & ~n1564 ) | ( n822 & ~n1564 ) ;
  assign n4112 = ~n1716 & n4111 ;
  assign n4113 = ~n421 & n4112 ;
  assign n4114 = n2419 & n4113 ;
  assign n4115 = ~n2104 & n3252 ;
  assign n4116 = n3885 ^ n2752 ^ 1'b0 ;
  assign n4117 = n2915 | n3787 ;
  assign n4118 = n191 | n4117 ;
  assign n4119 = ~n2381 & n2746 ;
  assign n4120 = ~n393 & n4119 ;
  assign n4121 = ( n2838 & n4118 ) | ( n2838 & n4120 ) | ( n4118 & n4120 ) ;
  assign n4122 = n3191 ^ n2939 ^ 1'b0 ;
  assign n4123 = n4121 & ~n4122 ;
  assign n4124 = ~n1223 & n4123 ;
  assign n4125 = n4124 ^ n2921 ^ n1298 ;
  assign n4126 = n323 & n356 ;
  assign n4127 = ~n374 & n4126 ;
  assign n4128 = n3330 | n4127 ;
  assign n4129 = n4128 ^ n2897 ^ 1'b0 ;
  assign n4130 = n861 | n1376 ;
  assign n4131 = n1984 & ~n4130 ;
  assign n4132 = ( n2104 & n3787 ) | ( n2104 & ~n4131 ) | ( n3787 & ~n4131 ) ;
  assign n4133 = n4132 ^ n592 ^ x40 ;
  assign n4134 = n4133 ^ n3297 ^ 1'b0 ;
  assign n4135 = ~n1751 & n1819 ;
  assign n4136 = n1580 ^ n1283 ^ n167 ;
  assign n4137 = n777 | n4136 ;
  assign n4138 = n4137 ^ n878 ^ n650 ;
  assign n4139 = ~n413 & n3470 ;
  assign n4140 = ( n4135 & n4138 ) | ( n4135 & ~n4139 ) | ( n4138 & ~n4139 ) ;
  assign n4141 = ( ~n2010 & n3374 ) | ( ~n2010 & n4140 ) | ( n3374 & n4140 ) ;
  assign n4142 = n2849 & ~n3719 ;
  assign n4143 = n2438 ^ n1939 ^ 1'b0 ;
  assign n4144 = n773 & n4143 ;
  assign n4145 = ~x21 & n599 ;
  assign n4146 = ~n2114 & n3174 ;
  assign n4147 = n4146 ^ n199 ^ 1'b0 ;
  assign n4148 = n4147 ^ n873 ^ 1'b0 ;
  assign n4149 = n3671 ^ n3071 ^ 1'b0 ;
  assign n4150 = n2198 | n4149 ;
  assign n4151 = n4150 ^ n743 ^ 1'b0 ;
  assign n4152 = n2547 & n4151 ;
  assign n4153 = n2067 | n2197 ;
  assign n4154 = n1910 & ~n4153 ;
  assign n4155 = x127 & ~n4154 ;
  assign n4156 = ( n1096 & n2160 ) | ( n1096 & ~n2377 ) | ( n2160 & ~n2377 ) ;
  assign n4158 = n1559 ^ n1555 ^ 1'b0 ;
  assign n4157 = n1866 & ~n3787 ;
  assign n4159 = n4158 ^ n4157 ^ 1'b0 ;
  assign n4160 = x11 & ~n4159 ;
  assign n4161 = ~n1076 & n2184 ;
  assign n4162 = n4161 ^ n196 ^ 1'b0 ;
  assign n4163 = n766 ^ n747 ^ x113 ;
  assign n4164 = n4163 ^ n3162 ^ n877 ;
  assign n4165 = n4164 ^ x63 ^ 1'b0 ;
  assign n4166 = n4165 ^ n2487 ^ n295 ;
  assign n4167 = n4166 ^ n1747 ^ n636 ;
  assign n4168 = n4162 & n4167 ;
  assign n4169 = n2625 & n4168 ;
  assign n4170 = n4160 & ~n4169 ;
  assign n4171 = n4156 & n4170 ;
  assign n4174 = ~n155 & n372 ;
  assign n4172 = n800 ^ n162 ^ x9 ;
  assign n4173 = n3835 & ~n4172 ;
  assign n4175 = n4174 ^ n4173 ^ 1'b0 ;
  assign n4189 = x89 & n1032 ;
  assign n4190 = n4189 ^ n1534 ^ 1'b0 ;
  assign n4187 = n144 & n1887 ;
  assign n4184 = n2732 ^ n1027 ^ n473 ;
  assign n4185 = x32 & n4184 ;
  assign n4186 = n884 & ~n4185 ;
  assign n4188 = n4187 ^ n4186 ^ 1'b0 ;
  assign n4191 = n4190 ^ n4188 ^ 1'b0 ;
  assign n4192 = n1077 & ~n4191 ;
  assign n4180 = ( ~n1208 & n1381 ) | ( ~n1208 & n1887 ) | ( n1381 & n1887 ) ;
  assign n4181 = n4180 ^ n1822 ^ n158 ;
  assign n4182 = ~n1278 & n4181 ;
  assign n4177 = n464 ^ n151 ^ 1'b0 ;
  assign n4178 = n1652 ^ n846 ^ 1'b0 ;
  assign n4179 = n4177 & ~n4178 ;
  assign n4183 = n4182 ^ n4179 ^ 1'b0 ;
  assign n4176 = n1204 ^ n803 ^ 1'b0 ;
  assign n4193 = n4192 ^ n4183 ^ n4176 ;
  assign n4194 = n963 | n1982 ;
  assign n4195 = n4194 ^ n3175 ^ n1253 ;
  assign n4196 = n358 | n2971 ;
  assign n4197 = n4196 ^ n265 ^ 1'b0 ;
  assign n4198 = ~n4195 & n4197 ;
  assign n4199 = n949 & ~n3507 ;
  assign n4200 = n4199 ^ n3496 ^ n916 ;
  assign n4201 = n4200 ^ n2572 ^ 1'b0 ;
  assign n4202 = n3631 & n4201 ;
  assign n4203 = n1591 ^ n251 ^ 1'b0 ;
  assign n4204 = n744 & n3062 ;
  assign n4205 = ~n4203 & n4204 ;
  assign n4206 = n1546 & n4205 ;
  assign n4207 = ~n1820 & n2901 ;
  assign n4208 = n560 ^ n323 ^ 1'b0 ;
  assign n4209 = n4067 ^ n2975 ^ 1'b0 ;
  assign n4210 = n4208 | n4209 ;
  assign n4211 = n803 | n3357 ;
  assign n4212 = n4211 ^ n2808 ^ n1065 ;
  assign n4213 = n2623 & n4212 ;
  assign n4214 = n4213 ^ n3209 ^ 1'b0 ;
  assign n4215 = n2810 | n4214 ;
  assign n4216 = n1138 | n1296 ;
  assign n4217 = n4216 ^ n2152 ^ n1381 ;
  assign n4218 = n4217 ^ n462 ^ x40 ;
  assign n4219 = ( ~n1204 & n3260 ) | ( ~n1204 & n4218 ) | ( n3260 & n4218 ) ;
  assign n4220 = n1901 ^ n431 ^ 1'b0 ;
  assign n4221 = n3134 ^ n1946 ^ n899 ;
  assign n4222 = ~n2549 & n4221 ;
  assign n4223 = n3592 ^ n2693 ^ 1'b0 ;
  assign n4224 = n4222 & ~n4223 ;
  assign n4225 = x72 & n1346 ;
  assign n4226 = n4225 ^ n447 ^ 1'b0 ;
  assign n4227 = n2178 & n4226 ;
  assign n4229 = x74 & ~n2404 ;
  assign n4230 = ~n1278 & n4229 ;
  assign n4231 = n3999 & ~n4230 ;
  assign n4228 = n1707 & n2842 ;
  assign n4232 = n4231 ^ n4228 ^ n3316 ;
  assign n4238 = ( n1429 & n2491 ) | ( n1429 & n3598 ) | ( n2491 & n3598 ) ;
  assign n4235 = n1846 & n2057 ;
  assign n4236 = n2065 & n4235 ;
  assign n4237 = n4236 ^ n318 ^ 1'b0 ;
  assign n4239 = n4238 ^ n4237 ^ 1'b0 ;
  assign n4233 = n2469 ^ n926 ^ 1'b0 ;
  assign n4234 = n4233 ^ n1295 ^ n1050 ;
  assign n4240 = n4239 ^ n4234 ^ 1'b0 ;
  assign n4241 = n2272 ^ n1167 ^ 1'b0 ;
  assign n4242 = ~n2722 & n4241 ;
  assign n4243 = n319 ^ x75 ^ 1'b0 ;
  assign n4244 = n2701 & ~n4243 ;
  assign n4245 = n522 & n4244 ;
  assign n4246 = ( n1286 & n1289 ) | ( n1286 & ~n3459 ) | ( n1289 & ~n3459 ) ;
  assign n4247 = n4246 ^ n4012 ^ n308 ;
  assign n4248 = n2199 ^ n2146 ^ x63 ;
  assign n4249 = n4247 | n4248 ;
  assign n4250 = n4249 ^ n1302 ^ 1'b0 ;
  assign n4251 = n1422 ^ n1346 ^ n1316 ;
  assign n4252 = n3112 ^ n2432 ^ 1'b0 ;
  assign n4253 = ~n4251 & n4252 ;
  assign n4254 = n4253 ^ n1534 ^ n1050 ;
  assign n4255 = n4254 ^ n1230 ^ n1018 ;
  assign n4256 = n144 | n3011 ;
  assign n4257 = ( x80 & ~n237 ) | ( x80 & n4256 ) | ( ~n237 & n4256 ) ;
  assign n4258 = n998 & ~n3748 ;
  assign n4259 = n4258 ^ n838 ^ 1'b0 ;
  assign n4260 = n4259 ^ x111 ^ 1'b0 ;
  assign n4261 = ( n1451 & n4257 ) | ( n1451 & n4260 ) | ( n4257 & n4260 ) ;
  assign n4264 = n796 ^ x11 ^ 1'b0 ;
  assign n4265 = n1816 & ~n4264 ;
  assign n4262 = n1467 ^ n416 ^ 1'b0 ;
  assign n4263 = n4262 ^ n679 ^ n422 ;
  assign n4266 = n4265 ^ n4263 ^ 1'b0 ;
  assign n4267 = n1007 ^ n708 ^ 1'b0 ;
  assign n4268 = n625 & n3253 ;
  assign n4269 = n1314 & n4268 ;
  assign n4270 = n2453 ^ n1498 ^ 1'b0 ;
  assign n4271 = ( n4267 & ~n4269 ) | ( n4267 & n4270 ) | ( ~n4269 & n4270 ) ;
  assign n4272 = n246 & ~n2091 ;
  assign n4273 = n3563 ^ n1023 ^ 1'b0 ;
  assign n4274 = x96 & n4273 ;
  assign n4275 = n1835 & n4274 ;
  assign n4276 = n3354 ^ n2344 ^ 1'b0 ;
  assign n4277 = ~n2984 & n4276 ;
  assign n4278 = ( n1598 & n2489 ) | ( n1598 & ~n4036 ) | ( n2489 & ~n4036 ) ;
  assign n4279 = n3428 ^ n2726 ^ 1'b0 ;
  assign n4280 = ~n851 & n1095 ;
  assign n4281 = n4280 ^ x42 ^ 1'b0 ;
  assign n4282 = x113 & n2768 ;
  assign n4296 = ( n1175 & ~n2065 ) | ( n1175 & n3396 ) | ( ~n2065 & n3396 ) ;
  assign n4283 = n1366 & ~n1601 ;
  assign n4284 = n4267 & ~n4283 ;
  assign n4285 = ~n1062 & n4284 ;
  assign n4286 = n2735 ^ x91 ^ 1'b0 ;
  assign n4287 = n4286 ^ n3934 ^ n2612 ;
  assign n4288 = n1079 ^ n987 ^ 1'b0 ;
  assign n4289 = n982 & ~n4288 ;
  assign n4290 = n883 & ~n4289 ;
  assign n4291 = n4290 ^ n2261 ^ 1'b0 ;
  assign n4292 = n3374 & ~n4291 ;
  assign n4293 = ~n154 & n4292 ;
  assign n4294 = ~n4287 & n4293 ;
  assign n4295 = n4285 | n4294 ;
  assign n4297 = n4296 ^ n4295 ^ 1'b0 ;
  assign n4298 = ~n1286 & n1883 ;
  assign n4299 = n812 & n4298 ;
  assign n4300 = n4299 ^ n2618 ^ 1'b0 ;
  assign n4301 = n4300 ^ n1328 ^ 1'b0 ;
  assign n4302 = n1923 & n4301 ;
  assign n4303 = n2444 ^ n866 ^ 1'b0 ;
  assign n4304 = n1071 | n4303 ;
  assign n4305 = ( n2310 & n4302 ) | ( n2310 & ~n4304 ) | ( n4302 & ~n4304 ) ;
  assign n4306 = n728 | n4216 ;
  assign n4307 = n3895 ^ n1749 ^ 1'b0 ;
  assign n4308 = n4307 ^ n390 ^ 1'b0 ;
  assign n4309 = n3450 ^ n1068 ^ 1'b0 ;
  assign n4310 = ~n4308 & n4309 ;
  assign n4311 = n3955 & n4310 ;
  assign n4312 = n2342 & n3616 ;
  assign n4313 = n4312 ^ n535 ^ 1'b0 ;
  assign n4314 = n1437 & ~n4313 ;
  assign n4315 = ~n4137 & n4314 ;
  assign n4317 = n608 ^ n269 ^ 1'b0 ;
  assign n4318 = n621 & n4317 ;
  assign n4319 = n4090 & n4318 ;
  assign n4320 = n426 & n4319 ;
  assign n4321 = ( n256 & n1310 ) | ( n256 & n4320 ) | ( n1310 & n4320 ) ;
  assign n4316 = x74 & ~n1629 ;
  assign n4322 = n4321 ^ n4316 ^ n310 ;
  assign n4323 = n4322 ^ n3640 ^ 1'b0 ;
  assign n4324 = x50 & ~n3569 ;
  assign n4325 = n4324 ^ n3278 ^ 1'b0 ;
  assign n4329 = n760 ^ n194 ^ 1'b0 ;
  assign n4326 = ~n940 & n1702 ;
  assign n4327 = ~n744 & n4326 ;
  assign n4328 = n4327 ^ n699 ^ x35 ;
  assign n4330 = n4329 ^ n4328 ^ 1'b0 ;
  assign n4331 = n3043 & n4330 ;
  assign n4332 = n4331 ^ n3323 ^ 1'b0 ;
  assign n4333 = x18 | n4332 ;
  assign n4334 = n2703 | n4333 ;
  assign n4335 = n842 | n2605 ;
  assign n4336 = n2901 ^ n2522 ^ 1'b0 ;
  assign n4340 = n3056 ^ n1531 ^ 1'b0 ;
  assign n4337 = n1837 & n2279 ;
  assign n4338 = ~n3707 & n4337 ;
  assign n4339 = ( ~x74 & n1591 ) | ( ~x74 & n4338 ) | ( n1591 & n4338 ) ;
  assign n4341 = n4340 ^ n4339 ^ n1934 ;
  assign n4342 = ~n1434 & n2348 ;
  assign n4343 = n4342 ^ n2581 ^ 1'b0 ;
  assign n4344 = ( n191 & n469 ) | ( n191 & n3212 ) | ( n469 & n3212 ) ;
  assign n4345 = n3542 ^ n1125 ^ 1'b0 ;
  assign n4346 = n4344 & n4345 ;
  assign n4347 = n4194 ^ n2889 ^ n987 ;
  assign n4348 = ( x118 & ~n2543 ) | ( x118 & n3215 ) | ( ~n2543 & n3215 ) ;
  assign n4357 = ( ~n3020 & n4007 ) | ( ~n3020 & n4086 ) | ( n4007 & n4086 ) ;
  assign n4349 = n2735 ^ n527 ^ 1'b0 ;
  assign n4350 = n2338 ^ n1886 ^ 1'b0 ;
  assign n4351 = n3031 & ~n4350 ;
  assign n4352 = ~n3766 & n4351 ;
  assign n4353 = n4349 & n4352 ;
  assign n4354 = ( ~n2453 & n2781 ) | ( ~n2453 & n4353 ) | ( n2781 & n4353 ) ;
  assign n4355 = n4354 ^ n1020 ^ 1'b0 ;
  assign n4356 = n2578 & n4355 ;
  assign n4358 = n4357 ^ n4356 ^ 1'b0 ;
  assign n4359 = n4348 & n4358 ;
  assign n4360 = n4359 ^ n928 ^ 1'b0 ;
  assign n4361 = ~n2971 & n4360 ;
  assign n4362 = ( n657 & ~n1263 ) | ( n657 & n3778 ) | ( ~n1263 & n3778 ) ;
  assign n4363 = n1590 | n4362 ;
  assign n4364 = ( n1032 & n1921 ) | ( n1032 & n2782 ) | ( n1921 & n2782 ) ;
  assign n4365 = n740 & n4364 ;
  assign n4366 = n4107 ^ n3749 ^ 1'b0 ;
  assign n4367 = n3581 & n4366 ;
  assign n4369 = n3178 | n3625 ;
  assign n4370 = n4369 ^ n283 ^ 1'b0 ;
  assign n4371 = ( n1830 & n4192 ) | ( n1830 & ~n4370 ) | ( n4192 & ~n4370 ) ;
  assign n4372 = x65 & n4371 ;
  assign n4373 = n4372 ^ n1400 ^ 1'b0 ;
  assign n4368 = n236 & ~n1193 ;
  assign n4374 = n4373 ^ n4368 ^ 1'b0 ;
  assign n4375 = n2237 ^ n134 ^ 1'b0 ;
  assign n4376 = n4374 | n4375 ;
  assign n4377 = n1372 ^ n1100 ^ n522 ;
  assign n4378 = ~n168 & n4377 ;
  assign n4379 = n3252 ^ n1736 ^ n314 ;
  assign n4380 = ( n437 & n761 ) | ( n437 & n4132 ) | ( n761 & n4132 ) ;
  assign n4381 = x87 & ~n4380 ;
  assign n4382 = n4381 ^ n1160 ^ 1'b0 ;
  assign n4383 = n798 ^ n732 ^ n322 ;
  assign n4384 = ( n1207 & n3625 ) | ( n1207 & ~n4383 ) | ( n3625 & ~n4383 ) ;
  assign n4385 = n4177 ^ n1261 ^ 1'b0 ;
  assign n4386 = n4384 & ~n4385 ;
  assign n4396 = x106 | n2006 ;
  assign n4392 = ( n1022 & n1215 ) | ( n1022 & n1864 ) | ( n1215 & n1864 ) ;
  assign n4387 = n1311 ^ n1013 ^ n305 ;
  assign n4388 = n4387 ^ n3996 ^ 1'b0 ;
  assign n4389 = n3051 | n4388 ;
  assign n4390 = ( n294 & n2498 ) | ( n294 & ~n4389 ) | ( n2498 & ~n4389 ) ;
  assign n4391 = ( n232 & ~n3254 ) | ( n232 & n4390 ) | ( ~n3254 & n4390 ) ;
  assign n4393 = n4392 ^ n4391 ^ n2950 ;
  assign n4394 = n4393 ^ n3521 ^ n3192 ;
  assign n4395 = n1287 & ~n4394 ;
  assign n4397 = n4396 ^ n4395 ^ 1'b0 ;
  assign n4398 = n2615 | n4397 ;
  assign n4399 = n4386 & ~n4398 ;
  assign n4401 = n246 & ~n323 ;
  assign n4402 = ( n570 & n1554 ) | ( n570 & n4401 ) | ( n1554 & n4401 ) ;
  assign n4400 = n691 & n1849 ;
  assign n4403 = n4402 ^ n4400 ^ 1'b0 ;
  assign n4404 = ~n2295 & n2788 ;
  assign n4405 = n3889 & n4404 ;
  assign n4406 = n4405 ^ n3505 ^ 1'b0 ;
  assign n4407 = n3200 ^ n675 ^ 1'b0 ;
  assign n4408 = n681 | n4407 ;
  assign n4409 = n2296 ^ n1622 ^ 1'b0 ;
  assign n4410 = n2187 | n4336 ;
  assign n4411 = n2090 & n3314 ;
  assign n4412 = n4410 & n4411 ;
  assign n4414 = n1966 & ~n2535 ;
  assign n4413 = n2515 ^ n2165 ^ n646 ;
  assign n4415 = n4414 ^ n4413 ^ n1360 ;
  assign n4416 = n4415 ^ n974 ^ n889 ;
  assign n4417 = n4416 ^ n692 ^ 1'b0 ;
  assign n4418 = n2447 ^ n2301 ^ 1'b0 ;
  assign n4419 = n4418 ^ n573 ^ 1'b0 ;
  assign n4420 = n3979 & ~n4419 ;
  assign n4421 = n422 & n4420 ;
  assign n4422 = ( ~n1143 & n3124 ) | ( ~n1143 & n4421 ) | ( n3124 & n4421 ) ;
  assign n4423 = n2898 & n3934 ;
  assign n4424 = n4423 ^ n3140 ^ n948 ;
  assign n4425 = n4424 ^ n3837 ^ 1'b0 ;
  assign n4426 = n1054 & n4425 ;
  assign n4427 = n3418 ^ n2657 ^ 1'b0 ;
  assign n4428 = ~n1243 & n3354 ;
  assign n4429 = n4428 ^ n436 ^ 1'b0 ;
  assign n4430 = n1783 ^ n509 ^ 1'b0 ;
  assign n4431 = n4430 ^ n4282 ^ 1'b0 ;
  assign n4432 = n4429 | n4431 ;
  assign n4433 = ~n1568 & n1774 ;
  assign n4434 = ( n612 & ~n2207 ) | ( n612 & n4433 ) | ( ~n2207 & n4433 ) ;
  assign n4440 = n1599 ^ n1221 ^ n773 ;
  assign n4435 = ~n196 & n915 ;
  assign n4436 = n4435 ^ n2692 ^ 1'b0 ;
  assign n4437 = n618 & ~n4436 ;
  assign n4438 = n4437 ^ n4018 ^ 1'b0 ;
  assign n4439 = n2154 & n4438 ;
  assign n4441 = n4440 ^ n4439 ^ 1'b0 ;
  assign n4442 = n4121 ^ n2676 ^ 1'b0 ;
  assign n4443 = n3111 & n4442 ;
  assign n4444 = n1428 | n2377 ;
  assign n4445 = n1611 | n4444 ;
  assign n4446 = n1505 ^ n426 ^ 1'b0 ;
  assign n4447 = n2645 | n4446 ;
  assign n4448 = n1343 | n4447 ;
  assign n4449 = n2704 ^ n1275 ^ n784 ;
  assign n4450 = ( ~x83 & n3845 ) | ( ~x83 & n4449 ) | ( n3845 & n4449 ) ;
  assign n4454 = n2790 | n3611 ;
  assign n4451 = n4316 ^ n3468 ^ 1'b0 ;
  assign n4452 = ( n824 & ~n1250 ) | ( n824 & n4451 ) | ( ~n1250 & n4451 ) ;
  assign n4453 = n4090 & n4452 ;
  assign n4455 = n4454 ^ n4453 ^ 1'b0 ;
  assign n4456 = n2676 ^ n1913 ^ 1'b0 ;
  assign n4457 = ~n883 & n1024 ;
  assign n4458 = n4457 ^ n3001 ^ 1'b0 ;
  assign n4459 = ( n2623 & n4401 ) | ( n2623 & ~n4458 ) | ( n4401 & ~n4458 ) ;
  assign n4460 = n2839 & ~n3635 ;
  assign n4461 = ~n920 & n4460 ;
  assign n4462 = n4461 ^ n4281 ^ x31 ;
  assign n4463 = ( n1382 & n2092 ) | ( n1382 & n3517 ) | ( n2092 & n3517 ) ;
  assign n4464 = n4463 ^ n196 ^ 1'b0 ;
  assign n4465 = n1707 & ~n4464 ;
  assign n4466 = n2294 ^ n1900 ^ 1'b0 ;
  assign n4467 = n776 ^ n466 ^ 1'b0 ;
  assign n4468 = ~n206 & n4467 ;
  assign n4469 = n4466 & ~n4468 ;
  assign n4470 = n1922 ^ n1773 ^ 1'b0 ;
  assign n4471 = n1553 & ~n4470 ;
  assign n4472 = n4469 & n4471 ;
  assign n4473 = n2390 ^ n1468 ^ 1'b0 ;
  assign n4474 = n808 | n4473 ;
  assign n4475 = n1439 & n1818 ;
  assign n4480 = n1287 ^ n482 ^ 1'b0 ;
  assign n4481 = ~n641 & n4480 ;
  assign n4482 = ( ~n1939 & n2242 ) | ( ~n1939 & n4481 ) | ( n2242 & n4481 ) ;
  assign n4476 = n897 ^ n277 ^ 1'b0 ;
  assign n4477 = ( n1590 & n4127 ) | ( n1590 & n4476 ) | ( n4127 & n4476 ) ;
  assign n4478 = n4477 ^ n710 ^ 1'b0 ;
  assign n4479 = ~n3670 & n4478 ;
  assign n4483 = n4482 ^ n4479 ^ n2687 ;
  assign n4485 = ( ~n434 & n508 ) | ( ~n434 & n2723 ) | ( n508 & n2723 ) ;
  assign n4484 = ( n1427 & ~n1658 ) | ( n1427 & n4418 ) | ( ~n1658 & n4418 ) ;
  assign n4486 = n4485 ^ n4484 ^ 1'b0 ;
  assign n4487 = ( ~n1090 & n2091 ) | ( ~n1090 & n4486 ) | ( n2091 & n4486 ) ;
  assign n4488 = n1053 & n2565 ;
  assign n4489 = ( n603 & n2046 ) | ( n603 & ~n4488 ) | ( n2046 & ~n4488 ) ;
  assign n4491 = n2143 ^ n469 ^ n371 ;
  assign n4492 = n888 & ~n4491 ;
  assign n4490 = n2778 | n3020 ;
  assign n4493 = n4492 ^ n4490 ^ 1'b0 ;
  assign n4494 = n4493 ^ n4466 ^ 1'b0 ;
  assign n4495 = ~n1258 & n2283 ;
  assign n4496 = n4495 ^ n3945 ^ 1'b0 ;
  assign n4497 = n4496 ^ n4033 ^ x63 ;
  assign n4498 = ( ~n1687 & n4100 ) | ( ~n1687 & n4497 ) | ( n4100 & n4497 ) ;
  assign n4499 = n4498 ^ n1632 ^ 1'b0 ;
  assign n4500 = n4494 & n4499 ;
  assign n4501 = ( n144 & n293 ) | ( n144 & ~n2927 ) | ( n293 & ~n2927 ) ;
  assign n4502 = ( ~n1543 & n3899 ) | ( ~n1543 & n4501 ) | ( n3899 & n4501 ) ;
  assign n4503 = n4502 ^ n4259 ^ n2223 ;
  assign n4504 = n495 & ~n2848 ;
  assign n4505 = ~n2549 & n4504 ;
  assign n4506 = n132 | n845 ;
  assign n4507 = n2434 & n4506 ;
  assign n4508 = n3016 & n4507 ;
  assign n4509 = n4508 ^ n2660 ^ n1230 ;
  assign n4510 = n4509 ^ n4385 ^ n2522 ;
  assign n4511 = ~n1361 & n4510 ;
  assign n4512 = n704 & ~n758 ;
  assign n4513 = n1287 | n4512 ;
  assign n4514 = n813 & ~n861 ;
  assign n4515 = n4514 ^ n838 ^ 1'b0 ;
  assign n4516 = ( n582 & ~n1172 ) | ( n582 & n4515 ) | ( ~n1172 & n4515 ) ;
  assign n4517 = n4516 ^ n3033 ^ 1'b0 ;
  assign n4522 = n2048 | n2600 ;
  assign n4523 = ~n874 & n4522 ;
  assign n4524 = ~n3519 & n4523 ;
  assign n4518 = ( n2114 & n2274 ) | ( n2114 & n2396 ) | ( n2274 & n2396 ) ;
  assign n4519 = n869 & n1581 ;
  assign n4520 = n1973 & n4519 ;
  assign n4521 = ( n1188 & ~n4518 ) | ( n1188 & n4520 ) | ( ~n4518 & n4520 ) ;
  assign n4525 = n4524 ^ n4521 ^ n4445 ;
  assign n4526 = n1385 ^ n1032 ^ n230 ;
  assign n4527 = n2550 & ~n3552 ;
  assign n4528 = n3656 ^ n2119 ^ n1827 ;
  assign n4529 = ~n872 & n2311 ;
  assign n4530 = ( n865 & ~n1490 ) | ( n865 & n1861 ) | ( ~n1490 & n1861 ) ;
  assign n4531 = n689 & n3477 ;
  assign n4532 = ~n4530 & n4531 ;
  assign n4533 = n1964 & n2587 ;
  assign n4534 = ~n167 & n4533 ;
  assign n4535 = n2413 ^ n1323 ^ 1'b0 ;
  assign n4536 = ( n1660 & n2231 ) | ( n1660 & ~n2507 ) | ( n2231 & ~n2507 ) ;
  assign n4537 = ~n2360 & n4536 ;
  assign n4538 = n4537 ^ n1251 ^ 1'b0 ;
  assign n4539 = ( n4534 & n4535 ) | ( n4534 & n4538 ) | ( n4535 & n4538 ) ;
  assign n4540 = n412 & ~n604 ;
  assign n4541 = n2264 & n4540 ;
  assign n4542 = n4541 ^ n241 ^ 1'b0 ;
  assign n4543 = ~n4539 & n4542 ;
  assign n4544 = n3367 ^ n947 ^ 1'b0 ;
  assign n4545 = ( n363 & n871 ) | ( n363 & ~n1023 ) | ( n871 & ~n1023 ) ;
  assign n4546 = n3885 ^ n1187 ^ 1'b0 ;
  assign n4547 = n728 ^ n318 ^ 1'b0 ;
  assign n4548 = n4546 | n4547 ;
  assign n4549 = x48 & ~n411 ;
  assign n4550 = n4549 ^ n1095 ^ 1'b0 ;
  assign n4551 = n3945 ^ n2774 ^ 1'b0 ;
  assign n4552 = ~n2424 & n4551 ;
  assign n4553 = ( n3238 & n4550 ) | ( n3238 & n4552 ) | ( n4550 & n4552 ) ;
  assign n4558 = n4184 ^ x88 ^ 1'b0 ;
  assign n4554 = ( n352 & n477 ) | ( n352 & n1277 ) | ( n477 & n1277 ) ;
  assign n4555 = n4554 ^ n1621 ^ n1329 ;
  assign n4556 = n562 | n4555 ;
  assign n4557 = n2778 & ~n4556 ;
  assign n4559 = n4558 ^ n4557 ^ 1'b0 ;
  assign n4560 = x6 & n4559 ;
  assign n4561 = n3256 & n4560 ;
  assign n4562 = x120 & ~n4561 ;
  assign n4563 = ~n4553 & n4562 ;
  assign n4564 = n1830 ^ n683 ^ 1'b0 ;
  assign n4565 = n4564 ^ n4539 ^ 1'b0 ;
  assign n4566 = n1943 | n4565 ;
  assign n4567 = n4563 | n4566 ;
  assign n4568 = n3454 ^ n419 ^ 1'b0 ;
  assign n4569 = ~n139 & n4568 ;
  assign n4571 = ( ~n806 & n1475 ) | ( ~n806 & n1876 ) | ( n1475 & n1876 ) ;
  assign n4570 = x32 & ~n1296 ;
  assign n4572 = n4571 ^ n4570 ^ 1'b0 ;
  assign n4573 = ( n2100 & n3121 ) | ( n2100 & ~n3747 ) | ( n3121 & ~n3747 ) ;
  assign n4574 = n3480 ^ n2975 ^ n325 ;
  assign n4576 = n641 & n1449 ;
  assign n4577 = ( n687 & ~n1870 ) | ( n687 & n4576 ) | ( ~n1870 & n4576 ) ;
  assign n4575 = n375 & n3277 ;
  assign n4578 = n4577 ^ n4575 ^ 1'b0 ;
  assign n4579 = ( n1753 & ~n3787 ) | ( n1753 & n4290 ) | ( ~n3787 & n4290 ) ;
  assign n4580 = ~x25 & n4579 ;
  assign n4581 = n2440 | n4580 ;
  assign n4582 = n4581 ^ n727 ^ 1'b0 ;
  assign n4583 = n4386 ^ n3556 ^ n2452 ;
  assign n4584 = n4583 ^ n3883 ^ n555 ;
  assign n4585 = ( n329 & n4582 ) | ( n329 & n4584 ) | ( n4582 & n4584 ) ;
  assign n4586 = ~n1521 & n2740 ;
  assign n4587 = n4586 ^ n514 ^ 1'b0 ;
  assign n4588 = n1311 ^ n654 ^ n149 ;
  assign n4589 = ( n842 & ~n2985 ) | ( n842 & n4588 ) | ( ~n2985 & n4588 ) ;
  assign n4590 = n3684 ^ n1411 ^ 1'b0 ;
  assign n4591 = n1006 | n4590 ;
  assign n4592 = n4591 ^ n1264 ^ 1'b0 ;
  assign n4593 = n4332 | n4592 ;
  assign n4594 = ( x45 & ~n697 ) | ( x45 & n1100 ) | ( ~n697 & n1100 ) ;
  assign n4595 = n4594 ^ n2098 ^ n1121 ;
  assign n4596 = n4595 ^ n1244 ^ 1'b0 ;
  assign n4597 = ~n4593 & n4596 ;
  assign n4599 = n2978 ^ n2315 ^ n1487 ;
  assign n4598 = n2114 | n4005 ;
  assign n4600 = n4599 ^ n4598 ^ n2200 ;
  assign n4601 = x66 & n1070 ;
  assign n4602 = n4601 ^ n687 ^ 1'b0 ;
  assign n4603 = n4602 ^ n141 ^ x7 ;
  assign n4604 = n4092 & ~n4603 ;
  assign n4605 = ~n2345 & n4604 ;
  assign n4606 = n2951 & n3008 ;
  assign n4607 = n880 | n3996 ;
  assign n4608 = n4606 | n4607 ;
  assign n4609 = n549 & n4290 ;
  assign n4610 = n2732 ^ n1135 ^ 1'b0 ;
  assign n4611 = n2835 & ~n4610 ;
  assign n4612 = ~n4509 & n4611 ;
  assign n4613 = n1312 & n4612 ;
  assign n4614 = ( n4608 & ~n4609 ) | ( n4608 & n4613 ) | ( ~n4609 & n4613 ) ;
  assign n4615 = n320 | n3290 ;
  assign n4619 = n2162 ^ n1946 ^ 1'b0 ;
  assign n4616 = n598 ^ x92 ^ 1'b0 ;
  assign n4617 = n4616 ^ n2043 ^ 1'b0 ;
  assign n4618 = n3759 & ~n4617 ;
  assign n4620 = n4619 ^ n4618 ^ 1'b0 ;
  assign n4621 = ~n1905 & n4620 ;
  assign n4622 = n2919 | n4524 ;
  assign n4623 = n134 & ~n2670 ;
  assign n4624 = ~n1422 & n4623 ;
  assign n4625 = n2718 ^ n2334 ^ n880 ;
  assign n4626 = n4625 ^ x66 ^ 1'b0 ;
  assign n4627 = n4626 ^ n4344 ^ 1'b0 ;
  assign n4628 = n4627 ^ n974 ^ 1'b0 ;
  assign n4629 = ( n2059 & n2421 ) | ( n2059 & n4628 ) | ( n2421 & n4628 ) ;
  assign n4634 = ( n259 & ~n1405 ) | ( n259 & n1590 ) | ( ~n1405 & n1590 ) ;
  assign n4630 = n3732 ^ n1756 ^ n775 ;
  assign n4631 = n2693 ^ n1514 ^ 1'b0 ;
  assign n4632 = n4630 & ~n4631 ;
  assign n4633 = n4632 ^ n452 ^ 1'b0 ;
  assign n4635 = n4634 ^ n4633 ^ 1'b0 ;
  assign n4636 = n4635 ^ n1899 ^ 1'b0 ;
  assign n4637 = ( ~n789 & n1754 ) | ( ~n789 & n3022 ) | ( n1754 & n3022 ) ;
  assign n4638 = n1332 & ~n2459 ;
  assign n4639 = n4638 ^ n4383 ^ 1'b0 ;
  assign n4640 = ( n689 & n881 ) | ( n689 & n2724 ) | ( n881 & n2724 ) ;
  assign n4641 = n1938 ^ x75 ^ x17 ;
  assign n4643 = n360 & ~n830 ;
  assign n4644 = n429 & n4643 ;
  assign n4642 = n2470 & ~n3046 ;
  assign n4645 = n4644 ^ n4642 ^ 1'b0 ;
  assign n4646 = n4645 ^ n3351 ^ 1'b0 ;
  assign n4647 = n4641 & ~n4646 ;
  assign n4648 = ~n454 & n4647 ;
  assign n4653 = ( x19 & ~n1040 ) | ( x19 & n1426 ) | ( ~n1040 & n1426 ) ;
  assign n4654 = n970 | n4653 ;
  assign n4655 = n4654 ^ n306 ^ 1'b0 ;
  assign n4649 = n880 | n1656 ;
  assign n4650 = n372 | n4649 ;
  assign n4651 = n4650 ^ n4552 ^ 1'b0 ;
  assign n4652 = n728 & n4651 ;
  assign n4656 = n4655 ^ n4652 ^ 1'b0 ;
  assign n4657 = n1666 | n3077 ;
  assign n4664 = ~n2687 & n4067 ;
  assign n4665 = ~n945 & n4664 ;
  assign n4658 = ~n822 & n1894 ;
  assign n4659 = n4658 ^ n2152 ^ 1'b0 ;
  assign n4660 = ~n2194 & n4659 ;
  assign n4661 = n1235 ^ n381 ^ 1'b0 ;
  assign n4662 = ~n4033 & n4661 ;
  assign n4663 = ~n4660 & n4662 ;
  assign n4666 = n4665 ^ n4663 ^ n3128 ;
  assign n4667 = n2614 ^ n432 ^ 1'b0 ;
  assign n4668 = n4651 & n4667 ;
  assign n4669 = ~n333 & n4668 ;
  assign n4670 = n380 & ~n4669 ;
  assign n4671 = ~n4666 & n4670 ;
  assign n4672 = n318 & n1407 ;
  assign n4673 = n4672 ^ n511 ^ 1'b0 ;
  assign n4674 = n1165 ^ n949 ^ 1'b0 ;
  assign n4675 = ~n604 & n4674 ;
  assign n4676 = n182 & n4675 ;
  assign n4677 = ~n4673 & n4676 ;
  assign n4678 = n2763 & n4677 ;
  assign n4679 = n4458 ^ n1698 ^ n1611 ;
  assign n4680 = n3725 ^ n2489 ^ 1'b0 ;
  assign n4681 = n2271 & n4470 ;
  assign n4682 = n1615 & n4681 ;
  assign n4683 = n4680 & n4682 ;
  assign n4685 = x24 & ~n1131 ;
  assign n4686 = n4685 ^ n615 ^ 1'b0 ;
  assign n4684 = n1866 ^ n1275 ^ 1'b0 ;
  assign n4687 = n4686 ^ n4684 ^ 1'b0 ;
  assign n4688 = n1889 | n4687 ;
  assign n4689 = n2663 | n4688 ;
  assign n4690 = n4689 ^ n2860 ^ n1449 ;
  assign n4691 = ( n1287 & n1596 ) | ( n1287 & ~n2015 ) | ( n1596 & ~n2015 ) ;
  assign n4692 = ( x77 & n1017 ) | ( x77 & ~n1628 ) | ( n1017 & ~n1628 ) ;
  assign n4693 = n3035 & ~n4692 ;
  assign n4694 = n3325 ^ n3272 ^ 1'b0 ;
  assign n4695 = ~n358 & n3410 ;
  assign n4696 = n4695 ^ n2174 ^ 1'b0 ;
  assign n4697 = ( n2915 & n4418 ) | ( n2915 & n4696 ) | ( n4418 & n4696 ) ;
  assign n4698 = n1533 | n2425 ;
  assign n4699 = n4698 ^ n2528 ^ 1'b0 ;
  assign n4700 = n2507 & n4699 ;
  assign n4701 = ( n914 & n2428 ) | ( n914 & n3018 ) | ( n2428 & n3018 ) ;
  assign n4702 = n2360 & ~n4701 ;
  assign n4703 = ( n316 & n569 ) | ( n316 & ~n1864 ) | ( n569 & ~n1864 ) ;
  assign n4704 = n2368 & n4703 ;
  assign n4705 = n4704 ^ n2174 ^ n719 ;
  assign n4706 = n4705 ^ n2951 ^ 1'b0 ;
  assign n4710 = n2978 ^ n908 ^ 1'b0 ;
  assign n4711 = n2836 | n4710 ;
  assign n4712 = ( n1830 & n4371 ) | ( n1830 & ~n4711 ) | ( n4371 & ~n4711 ) ;
  assign n4707 = n1280 | n2409 ;
  assign n4708 = n4707 ^ n3942 ^ 1'b0 ;
  assign n4709 = ~n2936 & n4708 ;
  assign n4713 = n4712 ^ n4709 ^ 1'b0 ;
  assign n4714 = n1547 ^ n667 ^ x89 ;
  assign n4715 = n4714 ^ n1976 ^ n1626 ;
  assign n4716 = x117 & n4715 ;
  assign n4717 = n619 & ~n1777 ;
  assign n4718 = n3132 | n4717 ;
  assign n4719 = n3542 & n4552 ;
  assign n4721 = n1645 & ~n2965 ;
  assign n4722 = n4721 ^ n821 ^ 1'b0 ;
  assign n4720 = ~n1274 & n4521 ;
  assign n4723 = n4722 ^ n4720 ^ 1'b0 ;
  assign n4724 = n2121 | n3722 ;
  assign n4725 = x106 | n4724 ;
  assign n4726 = ~n4723 & n4725 ;
  assign n4727 = n3500 ^ n1669 ^ n1277 ;
  assign n4731 = n2587 | n3598 ;
  assign n4730 = n2015 | n2485 ;
  assign n4728 = n2992 ^ n1556 ^ 1'b0 ;
  assign n4729 = n4449 & ~n4728 ;
  assign n4732 = n4731 ^ n4730 ^ n4729 ;
  assign n4733 = n2460 ^ n523 ^ 1'b0 ;
  assign n4734 = n203 & n4733 ;
  assign n4735 = n1202 & n4734 ;
  assign n4736 = ( n3290 & n4406 ) | ( n3290 & n4735 ) | ( n4406 & n4735 ) ;
  assign n4737 = n4096 ^ n925 ^ 1'b0 ;
  assign n4738 = n3181 & n4737 ;
  assign n4739 = n4738 ^ n4563 ^ 1'b0 ;
  assign n4740 = ~n2394 & n3926 ;
  assign n4741 = n1798 ^ n1472 ^ 1'b0 ;
  assign n4742 = ( n1793 & ~n3811 ) | ( n1793 & n3841 ) | ( ~n3811 & n3841 ) ;
  assign n4743 = n4742 ^ n2322 ^ 1'b0 ;
  assign n4744 = n4743 ^ n331 ^ x12 ;
  assign n4746 = n1145 ^ n919 ^ 1'b0 ;
  assign n4747 = n1338 & ~n4746 ;
  assign n4745 = n3130 ^ n1942 ^ 1'b0 ;
  assign n4748 = n4747 ^ n4745 ^ 1'b0 ;
  assign n4749 = n2684 & ~n4748 ;
  assign n4750 = n4749 ^ n3417 ^ n1478 ;
  assign n4751 = n1600 ^ n972 ^ 1'b0 ;
  assign n4752 = n3949 ^ n1468 ^ x69 ;
  assign n4753 = n307 & ~n2170 ;
  assign n4754 = ~n469 & n4753 ;
  assign n4759 = n2313 ^ x38 ^ 1'b0 ;
  assign n4760 = n2606 & n4759 ;
  assign n4761 = ( n1264 & n3089 ) | ( n1264 & n3968 ) | ( n3089 & n3968 ) ;
  assign n4762 = n4760 & n4761 ;
  assign n4755 = n2332 & ~n2560 ;
  assign n4756 = n4755 ^ n845 ^ 1'b0 ;
  assign n4757 = n1020 | n2796 ;
  assign n4758 = n4756 & n4757 ;
  assign n4763 = n4762 ^ n4758 ^ 1'b0 ;
  assign n4764 = n2898 & n4763 ;
  assign n4765 = ( ~n701 & n4754 ) | ( ~n701 & n4764 ) | ( n4754 & n4764 ) ;
  assign n4766 = n3396 ^ n1894 ^ n1069 ;
  assign n4767 = ~n348 & n2274 ;
  assign n4768 = n4767 ^ n338 ^ 1'b0 ;
  assign n4769 = ( x42 & n3019 ) | ( x42 & ~n4768 ) | ( n3019 & ~n4768 ) ;
  assign n4770 = n4769 ^ n490 ^ n456 ;
  assign n4771 = n4770 ^ n1472 ^ 1'b0 ;
  assign n4772 = n409 ^ x93 ^ 1'b0 ;
  assign n4773 = n4772 ^ n488 ^ 1'b0 ;
  assign n4774 = n3378 | n4773 ;
  assign n4775 = ~n2978 & n4774 ;
  assign n4776 = n3781 ^ n3713 ^ 1'b0 ;
  assign n4777 = n4775 | n4776 ;
  assign n4778 = n3286 ^ n1023 ^ n176 ;
  assign n4779 = ( ~x31 & n2889 ) | ( ~x31 & n4778 ) | ( n2889 & n4778 ) ;
  assign n4780 = ~n2284 & n3792 ;
  assign n4781 = n4780 ^ n654 ^ 1'b0 ;
  assign n4782 = n3491 | n4781 ;
  assign n4783 = n1493 | n4782 ;
  assign n4784 = n3189 ^ n3186 ^ 1'b0 ;
  assign n4785 = n4784 ^ n3436 ^ 1'b0 ;
  assign n4786 = x94 & ~n4785 ;
  assign n4787 = ~n1540 & n2114 ;
  assign n4788 = n2181 & n2205 ;
  assign n4789 = n4788 ^ n3328 ^ 1'b0 ;
  assign n4790 = n4789 ^ x80 ^ 1'b0 ;
  assign n4791 = ~n4787 & n4790 ;
  assign n4792 = n4791 ^ n2027 ^ n157 ;
  assign n4793 = n1903 & ~n4792 ;
  assign n4794 = n1670 & n1880 ;
  assign n4795 = n1551 & n4794 ;
  assign n4796 = n4558 | n4795 ;
  assign n4797 = n4796 ^ n1024 ^ 1'b0 ;
  assign n4798 = n2436 ^ n528 ^ 1'b0 ;
  assign n4799 = n4797 & n4798 ;
  assign n4800 = ( ~n299 & n914 ) | ( ~n299 & n1060 ) | ( n914 & n1060 ) ;
  assign n4801 = n4800 ^ n2121 ^ 1'b0 ;
  assign n4802 = n4799 & n4801 ;
  assign n4803 = n4050 ^ n831 ^ 1'b0 ;
  assign n4804 = n846 & n4803 ;
  assign n4805 = ( n3540 & ~n4432 ) | ( n3540 & n4733 ) | ( ~n4432 & n4733 ) ;
  assign n4806 = n1097 & ~n2915 ;
  assign n4807 = n4806 ^ n316 ^ 1'b0 ;
  assign n4808 = x66 & ~n4807 ;
  assign n4809 = n1656 & n4808 ;
  assign n4810 = ~n3417 & n4809 ;
  assign n4811 = ~n2030 & n2655 ;
  assign n4812 = ~n3393 & n4811 ;
  assign n4813 = n1062 & n4812 ;
  assign n4814 = n4813 ^ n1843 ^ 1'b0 ;
  assign n4817 = x65 ^ x1 ^ 1'b0 ;
  assign n4818 = n428 & n4817 ;
  assign n4815 = n646 | n2511 ;
  assign n4816 = n4492 & n4815 ;
  assign n4819 = n4818 ^ n4816 ^ n4735 ;
  assign n4820 = n3271 ^ n676 ^ n329 ;
  assign n4821 = ( ~n222 & n3903 ) | ( ~n222 & n4820 ) | ( n3903 & n4820 ) ;
  assign n4822 = ( ~n768 & n1485 ) | ( ~n768 & n3750 ) | ( n1485 & n3750 ) ;
  assign n4823 = n4821 & ~n4822 ;
  assign n4824 = ~n2217 & n4675 ;
  assign n4825 = n4824 ^ x58 ^ 1'b0 ;
  assign n4826 = n169 & ~n1745 ;
  assign n4827 = n401 & n4826 ;
  assign n4828 = n552 & ~n4827 ;
  assign n4829 = n1856 & n4828 ;
  assign n4830 = ~n4825 & n4829 ;
  assign n4831 = ( n4396 & n4823 ) | ( n4396 & ~n4830 ) | ( n4823 & ~n4830 ) ;
  assign n4836 = n3432 ^ n2440 ^ 1'b0 ;
  assign n4832 = n2116 | n2585 ;
  assign n4833 = x118 & ~n4832 ;
  assign n4834 = n4833 ^ n2198 ^ 1'b0 ;
  assign n4835 = n1445 & n4834 ;
  assign n4837 = n4836 ^ n4835 ^ 1'b0 ;
  assign n4838 = ( ~n3606 & n4097 ) | ( ~n3606 & n4837 ) | ( n4097 & n4837 ) ;
  assign n4839 = n2294 & ~n3383 ;
  assign n4840 = n2963 ^ n2732 ^ 1'b0 ;
  assign n4841 = n4067 ^ n2112 ^ n563 ;
  assign n4842 = n4840 & n4841 ;
  assign n4843 = n3214 | n3396 ;
  assign n4844 = n4843 ^ n1394 ^ 1'b0 ;
  assign n4845 = n4844 ^ n3738 ^ 1'b0 ;
  assign n4846 = ~n206 & n4845 ;
  assign n4847 = n885 & n4846 ;
  assign n4848 = n4847 ^ n2636 ^ 1'b0 ;
  assign n4850 = n3160 ^ n1278 ^ 1'b0 ;
  assign n4849 = n3740 ^ n676 ^ 1'b0 ;
  assign n4851 = n4850 ^ n4849 ^ 1'b0 ;
  assign n4852 = n985 & ~n2136 ;
  assign n4853 = ~n2265 & n4852 ;
  assign n4856 = n1441 | n3569 ;
  assign n4857 = n501 | n4856 ;
  assign n4854 = n3950 ^ n2870 ^ 1'b0 ;
  assign n4855 = n2470 | n4854 ;
  assign n4858 = n4857 ^ n4855 ^ 1'b0 ;
  assign n4859 = ( n1018 & n4853 ) | ( n1018 & n4858 ) | ( n4853 & n4858 ) ;
  assign n4860 = n4859 ^ n2938 ^ 1'b0 ;
  assign n4861 = n1160 & n4860 ;
  assign n4862 = ( ~n2855 & n3123 ) | ( ~n2855 & n4861 ) | ( n3123 & n4861 ) ;
  assign n4863 = n4183 ^ n285 ^ 1'b0 ;
  assign n4864 = n4219 & ~n4863 ;
  assign n4867 = n4756 ^ n3289 ^ n221 ;
  assign n4868 = x44 & n4867 ;
  assign n4869 = n2859 & n4868 ;
  assign n4865 = ( n927 & n1143 ) | ( n927 & ~n1306 ) | ( n1143 & ~n1306 ) ;
  assign n4866 = n3699 | n4865 ;
  assign n4870 = n4869 ^ n4866 ^ 1'b0 ;
  assign n4871 = n1581 ^ x74 ^ x45 ;
  assign n4872 = ~n3885 & n4871 ;
  assign n4873 = n2851 ^ n1308 ^ 1'b0 ;
  assign n4874 = n1345 | n1615 ;
  assign n4875 = n392 & n887 ;
  assign n4876 = n967 | n4875 ;
  assign n4877 = ( ~x30 & n420 ) | ( ~x30 & n2521 ) | ( n420 & n2521 ) ;
  assign n4878 = n492 & n3206 ;
  assign n4879 = n4063 & n4878 ;
  assign n4880 = ~n4877 & n4879 ;
  assign n4881 = n1555 & n2051 ;
  assign n4882 = ( n169 & n314 ) | ( n169 & ~n1196 ) | ( n314 & ~n1196 ) ;
  assign n4883 = ~n582 & n3822 ;
  assign n4889 = n2505 ^ n1880 ^ n1055 ;
  assign n4888 = n1291 | n1542 ;
  assign n4884 = ( n1240 & ~n1487 ) | ( n1240 & n4390 ) | ( ~n1487 & n4390 ) ;
  assign n4885 = ( n2181 & n2272 ) | ( n2181 & ~n4884 ) | ( n2272 & ~n4884 ) ;
  assign n4886 = n793 & n4885 ;
  assign n4887 = n197 & n4886 ;
  assign n4890 = n4889 ^ n4888 ^ n4887 ;
  assign n4891 = ~n1312 & n3656 ;
  assign n4892 = n4891 ^ n4344 ^ n1079 ;
  assign n4893 = n371 & n981 ;
  assign n4894 = n3709 & n4893 ;
  assign n4895 = n2480 & n4894 ;
  assign n4896 = n4402 ^ n2947 ^ 1'b0 ;
  assign n4897 = ~n544 & n1094 ;
  assign n4898 = n442 & ~n3633 ;
  assign n4899 = n4898 ^ n738 ^ 1'b0 ;
  assign n4900 = ( n3026 & n4897 ) | ( n3026 & ~n4899 ) | ( n4897 & ~n4899 ) ;
  assign n4901 = n2770 ^ n992 ^ 1'b0 ;
  assign n4902 = ~n4272 & n4901 ;
  assign n4903 = n3828 | n4046 ;
  assign n4904 = n4903 ^ n3240 ^ 1'b0 ;
  assign n4905 = ~n349 & n4904 ;
  assign n4906 = n2163 ^ n1896 ^ 1'b0 ;
  assign n4907 = n1055 | n4906 ;
  assign n4908 = n1966 & ~n4810 ;
  assign n4909 = n4233 ^ n2682 ^ 1'b0 ;
  assign n4910 = n411 | n4909 ;
  assign n4911 = n4910 ^ n3583 ^ 1'b0 ;
  assign n4912 = n1023 & ~n4911 ;
  assign n4913 = n170 & n4912 ;
  assign n4914 = n4913 ^ n1314 ^ 1'b0 ;
  assign n4915 = ( ~n1032 & n1683 ) | ( ~n1032 & n3367 ) | ( n1683 & n3367 ) ;
  assign n4916 = ~n1570 & n4915 ;
  assign n4917 = n4916 ^ n3590 ^ 1'b0 ;
  assign n4918 = n4914 | n4917 ;
  assign n4919 = ~n3854 & n3940 ;
  assign n4920 = n2339 & n4919 ;
  assign n4921 = n266 & ~n707 ;
  assign n4922 = x2 & ~n4921 ;
  assign n4923 = ~n589 & n4922 ;
  assign n4924 = n4923 ^ n894 ^ 1'b0 ;
  assign n4925 = n2417 & ~n4924 ;
  assign n4926 = n2227 & n4925 ;
  assign n4927 = n4926 ^ n2740 ^ 1'b0 ;
  assign n4928 = n4602 ^ x7 ^ 1'b0 ;
  assign n4929 = n3734 ^ n2641 ^ 1'b0 ;
  assign n4930 = n4928 | n4929 ;
  assign n4940 = n203 & ~n3694 ;
  assign n4941 = n4940 ^ x118 ^ 1'b0 ;
  assign n4942 = n4941 ^ n1058 ^ x119 ;
  assign n4943 = ( n1234 & n1666 ) | ( n1234 & ~n4942 ) | ( n1666 & ~n4942 ) ;
  assign n4939 = n2937 | n3223 ;
  assign n4931 = n3441 & n3507 ;
  assign n4932 = n4140 & n4931 ;
  assign n4933 = n1110 & n1198 ;
  assign n4934 = ~n136 & n1084 ;
  assign n4935 = n4934 ^ n332 ^ 1'b0 ;
  assign n4936 = n4933 & ~n4935 ;
  assign n4937 = n4932 & n4936 ;
  assign n4938 = ~n689 & n4937 ;
  assign n4944 = n4943 ^ n4939 ^ n4938 ;
  assign n4945 = n1733 ^ n1352 ^ 1'b0 ;
  assign n4946 = ( n171 & n1451 ) | ( n171 & n4945 ) | ( n1451 & n4945 ) ;
  assign n4947 = n1345 | n4873 ;
  assign n4948 = n4947 ^ n1384 ^ 1'b0 ;
  assign n4949 = ( n1279 & n1507 ) | ( n1279 & n2242 ) | ( n1507 & n2242 ) ;
  assign n4950 = ( n1213 & n3940 ) | ( n1213 & ~n4949 ) | ( n3940 & ~n4949 ) ;
  assign n4951 = ~n1751 & n2011 ;
  assign n4952 = ~x43 & n4951 ;
  assign n4957 = x44 | n557 ;
  assign n4958 = n4957 ^ n2065 ^ 1'b0 ;
  assign n4959 = n4912 & ~n4958 ;
  assign n4953 = ( n826 & ~n897 ) | ( n826 & n935 ) | ( ~n897 & n935 ) ;
  assign n4954 = ~n921 & n1623 ;
  assign n4955 = n1608 & n4954 ;
  assign n4956 = ( n878 & ~n4953 ) | ( n878 & n4955 ) | ( ~n4953 & n4955 ) ;
  assign n4960 = n4959 ^ n4956 ^ 1'b0 ;
  assign n4961 = n2004 ^ n157 ^ 1'b0 ;
  assign n4962 = n4865 ^ n184 ^ 1'b0 ;
  assign n4963 = n4736 & n4962 ;
  assign n4964 = n4961 & n4963 ;
  assign n4965 = n1951 ^ n194 ^ 1'b0 ;
  assign n4966 = n2735 | n4965 ;
  assign n4967 = ( n274 & n477 ) | ( n274 & n2072 ) | ( n477 & n2072 ) ;
  assign n4968 = n4967 ^ n4671 ^ 1'b0 ;
  assign n4969 = n242 & ~n4968 ;
  assign n4970 = ( n3860 & n4966 ) | ( n3860 & ~n4969 ) | ( n4966 & ~n4969 ) ;
  assign n4971 = ~n2447 & n3763 ;
  assign n4972 = n2167 ^ n1201 ^ 1'b0 ;
  assign n4973 = n4971 & n4972 ;
  assign n4974 = n2652 ^ n2522 ^ n2307 ;
  assign n4975 = n2198 | n2375 ;
  assign n4976 = n512 | n4975 ;
  assign n4977 = n3371 ^ x125 ^ 1'b0 ;
  assign n4978 = n4976 & ~n4977 ;
  assign n4979 = n4978 ^ n3238 ^ 1'b0 ;
  assign n4980 = ~n210 & n4501 ;
  assign n4981 = ~n3343 & n4418 ;
  assign n4982 = n2499 & n4981 ;
  assign n4983 = n2967 ^ n2498 ^ 1'b0 ;
  assign n4984 = n4982 | n4983 ;
  assign n4985 = n4980 | n4984 ;
  assign n4986 = n363 & ~n4985 ;
  assign n4987 = ( n4974 & n4979 ) | ( n4974 & n4986 ) | ( n4979 & n4986 ) ;
  assign n4988 = n579 | n1418 ;
  assign n4989 = n4988 ^ n2085 ^ 1'b0 ;
  assign n4990 = n3429 & n4989 ;
  assign n4991 = n1763 & n4990 ;
  assign n4992 = n4991 ^ n2532 ^ 1'b0 ;
  assign n4993 = n2284 ^ n2015 ^ x74 ;
  assign n4994 = n4993 ^ n2383 ^ 1'b0 ;
  assign n4995 = ~n3029 & n4994 ;
  assign n4996 = ( n474 & ~n2192 ) | ( n474 & n4039 ) | ( ~n2192 & n4039 ) ;
  assign n4997 = n386 & ~n2728 ;
  assign n4998 = n4997 ^ n866 ^ x108 ;
  assign n4999 = n4998 ^ n1009 ^ 1'b0 ;
  assign n5000 = n3909 ^ n2242 ^ n838 ;
  assign n5001 = n1704 ^ n1650 ^ n1043 ;
  assign n5002 = ( ~n505 & n5000 ) | ( ~n505 & n5001 ) | ( n5000 & n5001 ) ;
  assign n5003 = n5002 ^ n169 ^ 1'b0 ;
  assign n5004 = n3028 | n5003 ;
  assign n5005 = n4487 ^ n4237 ^ 1'b0 ;
  assign n5006 = n4342 ^ n1534 ^ 1'b0 ;
  assign n5007 = n1171 | n1439 ;
  assign n5008 = n5007 ^ n3946 ^ 1'b0 ;
  assign n5009 = n167 & n5008 ;
  assign n5010 = ~n3784 & n5009 ;
  assign n5011 = n4091 ^ x83 ^ 1'b0 ;
  assign n5015 = n213 & ~n2262 ;
  assign n5016 = n5015 ^ n2951 ^ 1'b0 ;
  assign n5012 = n717 | n3266 ;
  assign n5013 = n5012 ^ n1262 ^ 1'b0 ;
  assign n5014 = n5013 ^ n2136 ^ n877 ;
  assign n5017 = n5016 ^ n5014 ^ n3797 ;
  assign n5018 = ( n2489 & n2627 ) | ( n2489 & n4468 ) | ( n2627 & n4468 ) ;
  assign n5019 = n5018 ^ x55 ^ 1'b0 ;
  assign n5020 = n5017 & n5019 ;
  assign n5021 = n310 & ~n3795 ;
  assign n5022 = n2882 & n5021 ;
  assign n5023 = ( n2668 & n2758 ) | ( n2668 & ~n3812 ) | ( n2758 & ~n3812 ) ;
  assign n5024 = n2882 | n5023 ;
  assign n5025 = n3509 ^ n1263 ^ 1'b0 ;
  assign n5026 = n1740 ^ n246 ^ 1'b0 ;
  assign n5027 = n1692 | n2207 ;
  assign n5028 = n5026 | n5027 ;
  assign n5029 = ~n1838 & n5028 ;
  assign n5030 = n227 & n5029 ;
  assign n5031 = n2781 & ~n5030 ;
  assign n5032 = n5031 ^ n954 ^ 1'b0 ;
  assign n5033 = n1735 | n5032 ;
  assign n5034 = n5033 ^ n3102 ^ 1'b0 ;
  assign n5035 = ~n2200 & n5034 ;
  assign n5039 = n1324 | n3578 ;
  assign n5040 = n1639 & ~n5039 ;
  assign n5037 = n2317 ^ x51 ^ 1'b0 ;
  assign n5038 = n5037 ^ n4172 ^ n501 ;
  assign n5041 = n5040 ^ n5038 ^ n219 ;
  assign n5036 = ~n1219 & n3301 ;
  assign n5042 = n5041 ^ n5036 ^ n603 ;
  assign n5043 = n984 & n1894 ;
  assign n5044 = n5043 ^ n1449 ^ 1'b0 ;
  assign n5045 = n5044 ^ n1739 ^ n1219 ;
  assign n5046 = n5045 ^ n2076 ^ 1'b0 ;
  assign n5047 = n3013 | n5046 ;
  assign n5049 = ~n1212 & n1705 ;
  assign n5048 = x108 | n1088 ;
  assign n5050 = n5049 ^ n5048 ^ 1'b0 ;
  assign n5051 = ( x2 & n5047 ) | ( x2 & ~n5050 ) | ( n5047 & ~n5050 ) ;
  assign n5052 = ~n717 & n1531 ;
  assign n5053 = n668 ^ n658 ^ x60 ;
  assign n5054 = ( n2965 & ~n5052 ) | ( n2965 & n5053 ) | ( ~n5052 & n5053 ) ;
  assign n5055 = n1568 | n5054 ;
  assign n5056 = n3002 | n5055 ;
  assign n5057 = n3154 & n5056 ;
  assign n5058 = x126 ^ x98 ^ 1'b0 ;
  assign n5059 = ( ~x18 & n2774 ) | ( ~x18 & n4230 ) | ( n2774 & n4230 ) ;
  assign n5060 = n555 & ~n4449 ;
  assign n5061 = n5060 ^ n1349 ^ 1'b0 ;
  assign n5062 = ~n5059 & n5061 ;
  assign n5063 = n1399 & n5062 ;
  assign n5064 = n1765 ^ n1027 ^ n525 ;
  assign n5065 = ( n888 & ~n2819 ) | ( n888 & n3281 ) | ( ~n2819 & n3281 ) ;
  assign n5066 = n3095 & n5065 ;
  assign n5067 = n5066 ^ n2041 ^ 1'b0 ;
  assign n5068 = ( n2299 & n5064 ) | ( n2299 & n5067 ) | ( n5064 & n5067 ) ;
  assign n5069 = ( n1551 & n4390 ) | ( n1551 & ~n5068 ) | ( n4390 & ~n5068 ) ;
  assign n5070 = n552 | n652 ;
  assign n5071 = ( n321 & n1661 ) | ( n321 & ~n3632 ) | ( n1661 & ~n3632 ) ;
  assign n5072 = n5071 ^ n3276 ^ 1'b0 ;
  assign n5073 = n5070 & ~n5072 ;
  assign n5074 = n5073 ^ n4059 ^ 1'b0 ;
  assign n5075 = n4494 & n5074 ;
  assign n5076 = n1308 & ~n2036 ;
  assign n5077 = n5076 ^ n3318 ^ 1'b0 ;
  assign n5078 = n2798 & n3083 ;
  assign n5079 = ( n2269 & n2984 ) | ( n2269 & n3260 ) | ( n2984 & n3260 ) ;
  assign n5080 = n5079 ^ n3448 ^ 1'b0 ;
  assign n5081 = ( n4982 & ~n5078 ) | ( n4982 & n5080 ) | ( ~n5078 & n5080 ) ;
  assign n5082 = n3030 ^ n1096 ^ 1'b0 ;
  assign n5083 = n293 & n4099 ;
  assign n5084 = n2368 ^ n2111 ^ n2004 ;
  assign n5085 = n3144 | n5084 ;
  assign n5086 = n5083 & ~n5085 ;
  assign n5087 = n917 & ~n5086 ;
  assign n5088 = ~n5082 & n5087 ;
  assign n5089 = n4028 ^ n2391 ^ n522 ;
  assign n5090 = n1999 ^ n549 ^ 1'b0 ;
  assign n5091 = n676 & ~n5090 ;
  assign n5092 = n880 | n925 ;
  assign n5093 = n5092 ^ n2214 ^ 1'b0 ;
  assign n5094 = n5093 ^ n2334 ^ n1383 ;
  assign n5095 = ( n1343 & n3962 ) | ( n1343 & ~n5094 ) | ( n3962 & ~n5094 ) ;
  assign n5096 = n2585 & ~n5095 ;
  assign n5097 = n2792 ^ n1263 ^ 1'b0 ;
  assign n5098 = n5097 ^ n3463 ^ n147 ;
  assign n5099 = ( n2687 & n3386 ) | ( n2687 & ~n5098 ) | ( n3386 & ~n5098 ) ;
  assign n5100 = ~n468 & n3112 ;
  assign n5101 = ~n2342 & n5100 ;
  assign n5102 = n5101 ^ n194 ^ 1'b0 ;
  assign n5103 = n5102 ^ n2366 ^ 1'b0 ;
  assign n5104 = ( n617 & n744 ) | ( n617 & ~n787 ) | ( n744 & ~n787 ) ;
  assign n5105 = n2058 & ~n3096 ;
  assign n5106 = n1915 & n5105 ;
  assign n5107 = x59 & ~n5106 ;
  assign n5108 = ~n1420 & n5107 ;
  assign n5109 = n3219 | n5108 ;
  assign n5110 = n5109 ^ n3374 ^ n2758 ;
  assign n5111 = n5110 ^ n3325 ^ 1'b0 ;
  assign n5112 = n5104 & n5111 ;
  assign n5114 = n4387 ^ n883 ^ n617 ;
  assign n5113 = ( x118 & n1075 ) | ( x118 & ~n3169 ) | ( n1075 & ~n3169 ) ;
  assign n5115 = n5114 ^ n5113 ^ 1'b0 ;
  assign n5116 = n537 & ~n2400 ;
  assign n5117 = ~n3448 & n5116 ;
  assign n5121 = n548 ^ n390 ^ n155 ;
  assign n5122 = n5121 ^ n3055 ^ n357 ;
  assign n5118 = ( n479 & n2003 ) | ( n479 & ~n2572 ) | ( n2003 & ~n2572 ) ;
  assign n5119 = ~n639 & n5118 ;
  assign n5120 = n3424 & n5119 ;
  assign n5123 = n5122 ^ n5120 ^ n2911 ;
  assign n5124 = n2092 ^ n1443 ^ 1'b0 ;
  assign n5125 = n1317 ^ n766 ^ 1'b0 ;
  assign n5126 = n2720 | n5125 ;
  assign n5127 = ( n2921 & ~n4539 ) | ( n2921 & n5126 ) | ( ~n4539 & n5126 ) ;
  assign n5128 = n2239 & n5127 ;
  assign n5129 = n4423 ^ n2039 ^ 1'b0 ;
  assign n5132 = ( n903 & n1467 ) | ( n903 & ~n1713 ) | ( n1467 & ~n1713 ) ;
  assign n5130 = n2542 ^ n328 ^ 1'b0 ;
  assign n5131 = n2265 & n5130 ;
  assign n5133 = n5132 ^ n5131 ^ n432 ;
  assign n5134 = n3707 ^ n3596 ^ n1653 ;
  assign n5135 = n4062 | n5134 ;
  assign n5136 = n5135 ^ n2939 ^ 1'b0 ;
  assign n5137 = n4344 ^ n3221 ^ n196 ;
  assign n5138 = ~n1827 & n3564 ;
  assign n5139 = ~n1232 & n5138 ;
  assign n5140 = ( n2654 & ~n3888 ) | ( n2654 & n5139 ) | ( ~n3888 & n5139 ) ;
  assign n5141 = ~n5137 & n5140 ;
  assign n5142 = n5136 & n5141 ;
  assign n5143 = n3790 | n4616 ;
  assign n5144 = n2440 ^ n1251 ^ 1'b0 ;
  assign n5145 = n3828 ^ n2832 ^ 1'b0 ;
  assign n5146 = n1590 & n5145 ;
  assign n5147 = n5146 ^ n3183 ^ 1'b0 ;
  assign n5148 = n5147 ^ n1337 ^ n469 ;
  assign n5149 = ~n809 & n1078 ;
  assign n5150 = n4287 ^ n958 ^ 1'b0 ;
  assign n5151 = n5149 | n5150 ;
  assign n5152 = ( n1575 & n3362 ) | ( n1575 & n5151 ) | ( n3362 & n5151 ) ;
  assign n5153 = n1368 | n2478 ;
  assign n5154 = ( n844 & n3264 ) | ( n844 & ~n5153 ) | ( n3264 & ~n5153 ) ;
  assign n5155 = n2792 ^ n2450 ^ 1'b0 ;
  assign n5156 = n3258 | n5155 ;
  assign n5157 = ~n2867 & n5156 ;
  assign n5159 = n893 & n3303 ;
  assign n5158 = n541 & ~n3109 ;
  assign n5160 = n5159 ^ n5158 ^ 1'b0 ;
  assign n5161 = n5160 ^ n1690 ^ 1'b0 ;
  assign n5162 = n4481 & n5161 ;
  assign n5163 = n5157 & n5162 ;
  assign n5164 = n1776 ^ n710 ^ n318 ;
  assign n5165 = ( x56 & n3544 ) | ( x56 & n5164 ) | ( n3544 & n5164 ) ;
  assign n5166 = ( ~n296 & n2342 ) | ( ~n296 & n4593 ) | ( n2342 & n4593 ) ;
  assign n5167 = n3296 ^ n2654 ^ n221 ;
  assign n5168 = n3602 ^ n1326 ^ x77 ;
  assign n5169 = n5168 ^ n1821 ^ x70 ;
  assign n5170 = n2131 ^ n182 ^ x42 ;
  assign n5171 = ( n935 & n2394 ) | ( n935 & n5170 ) | ( n2394 & n5170 ) ;
  assign n5172 = ( n5167 & ~n5169 ) | ( n5167 & n5171 ) | ( ~n5169 & n5171 ) ;
  assign n5173 = ~n416 & n887 ;
  assign n5174 = n5173 ^ n3600 ^ n2869 ;
  assign n5175 = n2621 ^ n306 ^ 1'b0 ;
  assign n5176 = n5175 ^ n3921 ^ n2242 ;
  assign n5177 = n2947 ^ n1187 ^ 1'b0 ;
  assign n5178 = x54 & ~n4550 ;
  assign n5179 = n1390 | n3845 ;
  assign n5180 = ~n2100 & n2315 ;
  assign n5181 = ~n5179 & n5180 ;
  assign n5182 = ( n5177 & n5178 ) | ( n5177 & n5181 ) | ( n5178 & n5181 ) ;
  assign n5190 = n1187 & ~n1471 ;
  assign n5191 = n1471 & n5190 ;
  assign n5192 = n2644 | n4388 ;
  assign n5193 = n2644 & ~n5192 ;
  assign n5194 = n1961 & ~n5193 ;
  assign n5195 = n5191 & n5194 ;
  assign n5183 = ~n196 & n1754 ;
  assign n5184 = ~n3580 & n5183 ;
  assign n5185 = n316 & ~n586 ;
  assign n5186 = n5184 & n5185 ;
  assign n5187 = n4120 ^ n3465 ^ 1'b0 ;
  assign n5188 = n2840 & ~n5187 ;
  assign n5189 = ( n2082 & ~n5186 ) | ( n2082 & n5188 ) | ( ~n5186 & n5188 ) ;
  assign n5196 = n5195 ^ n5189 ^ 1'b0 ;
  assign n5197 = n1205 | n1913 ;
  assign n5198 = n5197 ^ n3363 ^ 1'b0 ;
  assign n5199 = n149 & ~n2017 ;
  assign n5200 = ~n5198 & n5199 ;
  assign n5201 = n3660 ^ n563 ^ 1'b0 ;
  assign n5202 = n2896 ^ n1616 ^ 1'b0 ;
  assign n5203 = n2560 ^ n753 ^ n563 ;
  assign n5205 = n4383 ^ n3348 ^ 1'b0 ;
  assign n5206 = ~n2104 & n5205 ;
  assign n5207 = n4135 & n5206 ;
  assign n5208 = n5207 ^ n1754 ^ 1'b0 ;
  assign n5204 = n482 & n1643 ;
  assign n5209 = n5208 ^ n5204 ^ 1'b0 ;
  assign n5210 = ( n3105 & ~n3784 ) | ( n3105 & n5209 ) | ( ~n3784 & n5209 ) ;
  assign n5211 = n767 | n4877 ;
  assign n5212 = ( ~n752 & n3940 ) | ( ~n752 & n5211 ) | ( n3940 & n5211 ) ;
  assign n5213 = ~n1513 & n2962 ;
  assign n5214 = n994 & n2681 ;
  assign n5215 = n5214 ^ n2875 ^ n1028 ;
  assign n5216 = n333 & ~n2027 ;
  assign n5217 = n2442 | n4401 ;
  assign n5218 = n1702 | n5217 ;
  assign n5219 = n5218 ^ n2111 ^ n1446 ;
  assign n5220 = n5219 ^ n2655 ^ n2147 ;
  assign n5221 = ( n2823 & n3069 ) | ( n2823 & n5220 ) | ( n3069 & n5220 ) ;
  assign n5222 = n5151 ^ n4014 ^ n3869 ;
  assign n5224 = ~n257 & n466 ;
  assign n5223 = n4787 ^ n1308 ^ 1'b0 ;
  assign n5225 = n5224 ^ n5223 ^ 1'b0 ;
  assign n5226 = n5225 ^ n3723 ^ 1'b0 ;
  assign n5227 = n5222 | n5226 ;
  assign n5228 = n2051 & n2998 ;
  assign n5229 = n812 & ~n1668 ;
  assign n5230 = n5229 ^ n1982 ^ n1650 ;
  assign n5231 = ~n569 & n5230 ;
  assign n5232 = n5231 ^ n2687 ^ 1'b0 ;
  assign n5233 = n5228 | n5232 ;
  assign n5234 = n3307 ^ n3027 ^ x40 ;
  assign n5235 = ( n821 & n2894 ) | ( n821 & n3857 ) | ( n2894 & n3857 ) ;
  assign n5236 = n5234 & n5235 ;
  assign n5237 = ~n2578 & n5236 ;
  assign n5238 = n2191 ^ n2083 ^ n851 ;
  assign n5239 = n4036 & ~n5238 ;
  assign n5240 = n5239 ^ n4361 ^ n693 ;
  assign n5241 = ~n1580 & n3581 ;
  assign n5242 = n3820 & n5241 ;
  assign n5243 = n5242 ^ n198 ^ 1'b0 ;
  assign n5244 = ~n1000 & n5243 ;
  assign n5245 = n5244 ^ n211 ^ 1'b0 ;
  assign n5248 = n1271 ^ n672 ^ 1'b0 ;
  assign n5249 = n5248 ^ n1611 ^ n230 ;
  assign n5246 = ~n3562 & n4045 ;
  assign n5247 = ( ~n1581 & n2204 ) | ( ~n1581 & n5246 ) | ( n2204 & n5246 ) ;
  assign n5250 = n5249 ^ n5247 ^ 1'b0 ;
  assign n5251 = ~n2490 & n5250 ;
  assign n5253 = n283 | n2623 ;
  assign n5254 = n3246 & ~n5253 ;
  assign n5252 = ~n953 & n4466 ;
  assign n5255 = n5254 ^ n5252 ^ 1'b0 ;
  assign n5256 = ~n366 & n3604 ;
  assign n5262 = ( n1175 & n3185 ) | ( n1175 & n3205 ) | ( n3185 & n3205 ) ;
  assign n5259 = n2354 & n2760 ;
  assign n5260 = n5259 ^ n315 ^ 1'b0 ;
  assign n5257 = n1311 ^ n991 ^ n937 ;
  assign n5258 = n2592 & n5257 ;
  assign n5261 = n5260 ^ n5258 ^ 1'b0 ;
  assign n5263 = n5262 ^ n5261 ^ n2998 ;
  assign n5265 = n1513 ^ n272 ^ 1'b0 ;
  assign n5264 = ~n1015 & n2514 ;
  assign n5266 = n5265 ^ n5264 ^ 1'b0 ;
  assign n5267 = ~n1940 & n5266 ;
  assign n5268 = ( n2322 & n3283 ) | ( n2322 & ~n5267 ) | ( n3283 & ~n5267 ) ;
  assign n5269 = ~n460 & n481 ;
  assign n5270 = ~n2835 & n5269 ;
  assign n5271 = n5270 ^ n3756 ^ n1840 ;
  assign n5273 = ( x2 & n1745 ) | ( x2 & n2971 ) | ( n1745 & n2971 ) ;
  assign n5272 = ( n650 & n1754 ) | ( n650 & n3296 ) | ( n1754 & n3296 ) ;
  assign n5274 = n5273 ^ n5272 ^ x10 ;
  assign n5275 = n5274 ^ n1510 ^ n255 ;
  assign n5276 = ( ~n1406 & n1423 ) | ( ~n1406 & n2671 ) | ( n1423 & n2671 ) ;
  assign n5277 = n4559 & n4822 ;
  assign n5278 = ( ~n129 & n1462 ) | ( ~n129 & n4123 ) | ( n1462 & n4123 ) ;
  assign n5279 = n5278 ^ n198 ^ 1'b0 ;
  assign n5280 = n5277 | n5279 ;
  assign n5281 = ~n2353 & n2832 ;
  assign n5282 = ( n2558 & ~n2785 ) | ( n2558 & n5281 ) | ( ~n2785 & n5281 ) ;
  assign n5283 = n5282 ^ n1986 ^ n961 ;
  assign n5284 = n5283 ^ n3560 ^ n3178 ;
  assign n5285 = n1529 | n2481 ;
  assign n5286 = n2744 | n5285 ;
  assign n5287 = n2965 ^ n2000 ^ n1000 ;
  assign n5288 = n809 & ~n3772 ;
  assign n5289 = n5288 ^ n657 ^ 1'b0 ;
  assign n5290 = ( n3955 & n5287 ) | ( n3955 & ~n5289 ) | ( n5287 & ~n5289 ) ;
  assign n5294 = n4302 ^ n2112 ^ 1'b0 ;
  assign n5292 = n989 & n4858 ;
  assign n5293 = n5292 ^ n390 ^ 1'b0 ;
  assign n5291 = ( n2199 & n2381 ) | ( n2199 & ~n4602 ) | ( n2381 & ~n4602 ) ;
  assign n5295 = n5294 ^ n5293 ^ n5291 ;
  assign n5296 = n3165 ^ n2257 ^ 1'b0 ;
  assign n5297 = x25 & ~n5296 ;
  assign n5298 = n1276 ^ n912 ^ 1'b0 ;
  assign n5299 = n5298 ^ n4939 ^ 1'b0 ;
  assign n5300 = n666 & n5299 ;
  assign n5301 = ( n2114 & ~n2296 ) | ( n2114 & n4222 ) | ( ~n2296 & n4222 ) ;
  assign n5302 = n5301 ^ n1418 ^ 1'b0 ;
  assign n5303 = n3067 ^ n1534 ^ n819 ;
  assign n5304 = ( ~n643 & n3134 ) | ( ~n643 & n5303 ) | ( n3134 & n5303 ) ;
  assign n5305 = n2884 ^ n384 ^ n228 ;
  assign n5306 = ~n3903 & n5305 ;
  assign n5307 = n5304 & n5306 ;
  assign n5308 = n5302 & n5307 ;
  assign n5309 = n5308 ^ n3011 ^ n236 ;
  assign n5310 = ~n3255 & n5309 ;
  assign n5311 = n5310 ^ n2671 ^ 1'b0 ;
  assign n5312 = ( n1114 & n3641 ) | ( n1114 & ~n5311 ) | ( n3641 & ~n5311 ) ;
  assign n5313 = n5153 ^ n3380 ^ 1'b0 ;
  assign n5314 = ( n1866 & n3750 ) | ( n1866 & ~n4768 ) | ( n3750 & ~n4768 ) ;
  assign n5315 = n2406 & ~n4715 ;
  assign n5316 = n5315 ^ x17 ^ 1'b0 ;
  assign n5317 = n5314 | n5316 ;
  assign n5318 = n5317 ^ n555 ^ 1'b0 ;
  assign n5319 = ( ~n1382 & n4747 ) | ( ~n1382 & n5318 ) | ( n4747 & n5318 ) ;
  assign n5320 = n5095 & ~n5319 ;
  assign n5321 = n1020 | n1492 ;
  assign n5322 = ( n2569 & n3242 ) | ( n2569 & ~n5321 ) | ( n3242 & ~n5321 ) ;
  assign n5323 = n3812 ^ n3255 ^ n1472 ;
  assign n5324 = n5323 ^ n2882 ^ 1'b0 ;
  assign n5325 = n4328 & ~n5324 ;
  assign n5326 = ~n5322 & n5325 ;
  assign n5327 = ~n547 & n1743 ;
  assign n5328 = n5327 ^ x15 ^ 1'b0 ;
  assign n5329 = ( n3346 & ~n4688 ) | ( n3346 & n5328 ) | ( ~n4688 & n5328 ) ;
  assign n5330 = n1409 ^ n888 ^ 1'b0 ;
  assign n5331 = n2056 & n5330 ;
  assign n5332 = n1976 ^ x2 ^ 1'b0 ;
  assign n5333 = n1901 & n5332 ;
  assign n5334 = n5333 ^ n2215 ^ 1'b0 ;
  assign n5335 = n2317 ^ x18 ^ 1'b0 ;
  assign n5336 = n3759 & ~n5335 ;
  assign n5337 = n5336 ^ n3072 ^ 1'b0 ;
  assign n5338 = n5334 | n5337 ;
  assign n5339 = n383 | n4998 ;
  assign n5340 = n5339 ^ n2140 ^ n2083 ;
  assign n5341 = ( n1458 & n1954 ) | ( n1458 & ~n5340 ) | ( n1954 & ~n5340 ) ;
  assign n5342 = n4253 ^ n3977 ^ n1820 ;
  assign n5343 = ( ~n4754 & n5341 ) | ( ~n4754 & n5342 ) | ( n5341 & n5342 ) ;
  assign n5344 = n753 & n4438 ;
  assign n5345 = ~n4233 & n5344 ;
  assign n5353 = ( n186 & n1067 ) | ( n186 & ~n1546 ) | ( n1067 & ~n1546 ) ;
  assign n5346 = n1617 | n2691 ;
  assign n5347 = n773 | n5346 ;
  assign n5348 = n5347 ^ n3020 ^ 1'b0 ;
  assign n5349 = n1076 | n5348 ;
  assign n5350 = n1668 | n5349 ;
  assign n5351 = ( ~n1253 & n2179 ) | ( ~n1253 & n5350 ) | ( n2179 & n5350 ) ;
  assign n5352 = ~n3840 & n5351 ;
  assign n5354 = n5353 ^ n5352 ^ 1'b0 ;
  assign n5355 = ~n3247 & n4296 ;
  assign n5356 = ( n1587 & n1641 ) | ( n1587 & ~n2468 ) | ( n1641 & ~n2468 ) ;
  assign n5357 = ~n1467 & n5356 ;
  assign n5358 = n584 & n5357 ;
  assign n5359 = n347 | n5358 ;
  assign n5360 = n5359 ^ n460 ^ 1'b0 ;
  assign n5361 = ( n1773 & ~n3599 ) | ( n1773 & n5360 ) | ( ~n3599 & n5360 ) ;
  assign n5362 = n2610 | n5361 ;
  assign n5365 = ( x63 & n935 ) | ( x63 & ~n3244 ) | ( n935 & ~n3244 ) ;
  assign n5363 = n2599 & n2987 ;
  assign n5364 = n5363 ^ n516 ^ 1'b0 ;
  assign n5366 = n5365 ^ n5364 ^ n1712 ;
  assign n5367 = n2542 ^ n1199 ^ 1'b0 ;
  assign n5368 = n5367 ^ n1914 ^ 1'b0 ;
  assign n5369 = ( n3485 & n4905 ) | ( n3485 & ~n5368 ) | ( n4905 & ~n5368 ) ;
  assign n5375 = n925 ^ n786 ^ 1'b0 ;
  assign n5370 = n375 & ~n1463 ;
  assign n5371 = n2962 | n5248 ;
  assign n5372 = ~n1551 & n5371 ;
  assign n5373 = n5372 ^ n894 ^ 1'b0 ;
  assign n5374 = ( n188 & n5370 ) | ( n188 & ~n5373 ) | ( n5370 & ~n5373 ) ;
  assign n5376 = n5375 ^ n5374 ^ 1'b0 ;
  assign n5377 = n695 ^ x119 ^ 1'b0 ;
  assign n5378 = n2929 | n5377 ;
  assign n5379 = n5378 ^ n2564 ^ 1'b0 ;
  assign n5380 = ( n2308 & ~n3288 ) | ( n2308 & n3579 ) | ( ~n3288 & n3579 ) ;
  assign n5381 = n5380 ^ n2294 ^ n2020 ;
  assign n5382 = n3253 ^ n2608 ^ 1'b0 ;
  assign n5383 = n5382 ^ n4752 ^ 1'b0 ;
  assign n5384 = n221 & ~n5383 ;
  assign n5386 = ( ~x19 & x40 ) | ( ~x19 & n1445 ) | ( x40 & n1445 ) ;
  assign n5385 = n2232 ^ x100 ^ 1'b0 ;
  assign n5387 = n5386 ^ n5385 ^ n4956 ;
  assign n5388 = n5387 ^ n996 ^ n413 ;
  assign n5390 = n1449 & n3661 ;
  assign n5391 = n5390 ^ n554 ^ x29 ;
  assign n5389 = n4443 ^ n1098 ^ 1'b0 ;
  assign n5392 = n5391 ^ n5389 ^ n2908 ;
  assign n5393 = n5392 ^ n2010 ^ 1'b0 ;
  assign n5394 = n462 | n5393 ;
  assign n5395 = ( n296 & n378 ) | ( n296 & ~n3484 ) | ( n378 & ~n3484 ) ;
  assign n5397 = n333 & n2340 ;
  assign n5396 = n2194 ^ n1970 ^ 1'b0 ;
  assign n5398 = n5397 ^ n5396 ^ 1'b0 ;
  assign n5399 = ( ~n3556 & n5395 ) | ( ~n3556 & n5398 ) | ( n5395 & n5398 ) ;
  assign n5400 = n3027 ^ n432 ^ 1'b0 ;
  assign n5401 = n1062 & ~n5400 ;
  assign n5402 = n1200 & n5401 ;
  assign n5403 = ( n2259 & n5399 ) | ( n2259 & ~n5402 ) | ( n5399 & ~n5402 ) ;
  assign n5404 = n5403 ^ n2315 ^ 1'b0 ;
  assign n5405 = n3167 & n5404 ;
  assign n5406 = ~n1108 & n1711 ;
  assign n5407 = ~n1912 & n5406 ;
  assign n5408 = ( ~n331 & n2832 ) | ( ~n331 & n5407 ) | ( n2832 & n5407 ) ;
  assign n5409 = n5408 ^ n4917 ^ 1'b0 ;
  assign n5410 = ~n4259 & n5409 ;
  assign n5411 = n5302 ^ n2325 ^ n1244 ;
  assign n5412 = n977 | n5411 ;
  assign n5413 = n3761 ^ n2192 ^ 1'b0 ;
  assign n5414 = n926 & ~n5413 ;
  assign n5415 = n5414 ^ n956 ^ 1'b0 ;
  assign n5416 = n5415 ^ n4318 ^ 1'b0 ;
  assign n5417 = n5115 ^ n1758 ^ 1'b0 ;
  assign n5418 = ( ~n232 & n3554 ) | ( ~n232 & n4251 ) | ( n3554 & n4251 ) ;
  assign n5419 = x75 & ~n1723 ;
  assign n5420 = ~n5418 & n5419 ;
  assign n5421 = n3051 ^ n1340 ^ 1'b0 ;
  assign n5422 = ~n3694 & n5421 ;
  assign n5423 = ~x110 & n5422 ;
  assign n5424 = n5420 | n5423 ;
  assign n5425 = n5424 ^ n4582 ^ 1'b0 ;
  assign n5426 = n3584 & ~n5425 ;
  assign n5427 = n5426 ^ n881 ^ 1'b0 ;
  assign n5428 = n393 ^ n234 ^ x74 ;
  assign n5429 = n5428 ^ n4904 ^ n821 ;
  assign n5431 = n2810 ^ n2179 ^ n697 ;
  assign n5430 = ~n1030 & n2436 ;
  assign n5432 = n5431 ^ n5430 ^ n3235 ;
  assign n5433 = n2636 | n5432 ;
  assign n5434 = n3864 & ~n4844 ;
  assign n5436 = n658 | n1618 ;
  assign n5435 = n4164 & ~n5273 ;
  assign n5437 = n5436 ^ n5435 ^ 1'b0 ;
  assign n5438 = n5434 & ~n5437 ;
  assign n5442 = ( n2251 & ~n3792 ) | ( n2251 & n5211 ) | ( ~n3792 & n5211 ) ;
  assign n5440 = n2522 ^ n1346 ^ n672 ;
  assign n5439 = n5260 ^ n2167 ^ 1'b0 ;
  assign n5441 = n5440 ^ n5439 ^ n3194 ;
  assign n5443 = n5442 ^ n5441 ^ 1'b0 ;
  assign n5444 = n5438 | n5443 ;
  assign n5445 = n5444 ^ n1376 ^ 1'b0 ;
  assign n5446 = n5433 & ~n5445 ;
  assign n5447 = n4822 ^ n3715 ^ 1'b0 ;
  assign n5449 = n1439 | n1756 ;
  assign n5448 = n3046 ^ n2060 ^ x86 ;
  assign n5450 = n5449 ^ n5448 ^ n1211 ;
  assign n5451 = n5450 ^ n4934 ^ n2457 ;
  assign n5452 = x119 & n4877 ;
  assign n5453 = n5452 ^ n1290 ^ 1'b0 ;
  assign n5454 = ( x61 & ~n1905 ) | ( x61 & n3091 ) | ( ~n1905 & n3091 ) ;
  assign n5455 = n1208 ^ n783 ^ 1'b0 ;
  assign n5456 = n396 | n1448 ;
  assign n5457 = n5456 ^ n3190 ^ 1'b0 ;
  assign n5458 = ( n3319 & n5455 ) | ( n3319 & ~n5457 ) | ( n5455 & ~n5457 ) ;
  assign n5459 = x41 & ~n2300 ;
  assign n5460 = n5458 & n5459 ;
  assign n5461 = ( n5453 & n5454 ) | ( n5453 & n5460 ) | ( n5454 & n5460 ) ;
  assign n5462 = n147 & ~n5160 ;
  assign n5463 = ~n1867 & n5462 ;
  assign n5464 = ~n1568 & n2315 ;
  assign n5465 = n5464 ^ n1526 ^ 1'b0 ;
  assign n5466 = n5463 & ~n5465 ;
  assign n5471 = ( ~n472 & n2129 ) | ( ~n472 & n3045 ) | ( n2129 & n3045 ) ;
  assign n5467 = n4362 ^ n3649 ^ 1'b0 ;
  assign n5468 = n3161 | n5467 ;
  assign n5469 = ( n2003 & n3470 ) | ( n2003 & n3889 ) | ( n3470 & n3889 ) ;
  assign n5470 = ( n1444 & ~n5468 ) | ( n1444 & n5469 ) | ( ~n5468 & n5469 ) ;
  assign n5472 = n5471 ^ n5470 ^ 1'b0 ;
  assign n5473 = n3235 ^ n2776 ^ 1'b0 ;
  assign n5474 = ( n1732 & ~n2134 ) | ( n1732 & n2895 ) | ( ~n2134 & n2895 ) ;
  assign n5475 = ( n2782 & n5473 ) | ( n2782 & ~n5474 ) | ( n5473 & ~n5474 ) ;
  assign n5476 = n3441 ^ n243 ^ 1'b0 ;
  assign n5477 = n1044 | n5476 ;
  assign n5478 = n1043 | n5477 ;
  assign n5479 = n4082 & n5478 ;
  assign n5480 = n2895 & n4267 ;
  assign n5481 = n199 & ~n272 ;
  assign n5482 = ~x58 & n5481 ;
  assign n5483 = n1654 | n5482 ;
  assign n5484 = n5483 ^ n942 ^ 1'b0 ;
  assign n5485 = n2223 & n5484 ;
  assign n5486 = n5480 & ~n5485 ;
  assign n5487 = n1976 ^ n1803 ^ 1'b0 ;
  assign n5488 = ~n1974 & n5487 ;
  assign n5489 = n5446 ^ n4246 ^ 1'b0 ;
  assign n5490 = n5488 & ~n5489 ;
  assign n5491 = n2817 & ~n3961 ;
  assign n5492 = n5491 ^ n2989 ^ n1814 ;
  assign n5493 = n2528 ^ n1673 ^ n335 ;
  assign n5494 = n612 | n2307 ;
  assign n5495 = n5494 ^ n1761 ^ 1'b0 ;
  assign n5496 = n5493 & ~n5495 ;
  assign n5497 = n5496 ^ n3013 ^ 1'b0 ;
  assign n5498 = n2192 & n5497 ;
  assign n5499 = n1422 | n3484 ;
  assign n5500 = n5056 | n5499 ;
  assign n5501 = ~n2087 & n5500 ;
  assign n5502 = ~n366 & n5501 ;
  assign n5503 = n5502 ^ n1366 ^ 1'b0 ;
  assign n5504 = ~n620 & n2227 ;
  assign n5505 = n5504 ^ n1966 ^ 1'b0 ;
  assign n5506 = n5505 ^ n1264 ^ 1'b0 ;
  assign n5507 = n514 & ~n976 ;
  assign n5508 = n5507 ^ n1167 ^ n210 ;
  assign n5509 = ( x118 & ~n1683 ) | ( x118 & n2098 ) | ( ~n1683 & n2098 ) ;
  assign n5510 = n5397 ^ n4396 ^ n781 ;
  assign n5511 = ~n392 & n2650 ;
  assign n5512 = n2830 ^ n2006 ^ n147 ;
  assign n5513 = n4837 | n5512 ;
  assign n5514 = n3812 ^ n1839 ^ n1108 ;
  assign n5515 = n4655 & ~n5514 ;
  assign n5516 = n1838 & n5515 ;
  assign n5518 = x112 & ~n2025 ;
  assign n5519 = ~n1691 & n5518 ;
  assign n5520 = n5519 ^ n1114 ^ 1'b0 ;
  assign n5521 = ( n601 & n1553 ) | ( n601 & ~n2659 ) | ( n1553 & ~n2659 ) ;
  assign n5522 = n5521 ^ n1758 ^ n211 ;
  assign n5523 = n2699 & n5522 ;
  assign n5524 = n4508 ^ n1784 ^ x2 ;
  assign n5525 = ( n5520 & n5523 ) | ( n5520 & ~n5524 ) | ( n5523 & ~n5524 ) ;
  assign n5517 = ~n1323 & n3403 ;
  assign n5526 = n5525 ^ n5517 ^ 1'b0 ;
  assign n5530 = ~n3211 & n4289 ;
  assign n5531 = n2432 | n5530 ;
  assign n5532 = n3644 | n5531 ;
  assign n5533 = n2160 ^ n2036 ^ 1'b0 ;
  assign n5534 = ~n2826 & n5533 ;
  assign n5535 = n5534 ^ n2269 ^ 1'b0 ;
  assign n5536 = n798 & ~n5535 ;
  assign n5537 = ~n5532 & n5536 ;
  assign n5528 = ~n318 & n620 ;
  assign n5527 = n3393 ^ n2313 ^ 1'b0 ;
  assign n5529 = n5528 ^ n5527 ^ 1'b0 ;
  assign n5538 = n5537 ^ n5529 ^ 1'b0 ;
  assign n5539 = ( ~n708 & n2153 ) | ( ~n708 & n3840 ) | ( n2153 & n3840 ) ;
  assign n5540 = n691 & ~n5539 ;
  assign n5541 = n5540 ^ n4378 ^ 1'b0 ;
  assign n5542 = n3307 ^ n1361 ^ n713 ;
  assign n5543 = ( n597 & n1426 ) | ( n597 & ~n2165 ) | ( n1426 & ~n2165 ) ;
  assign n5544 = n5543 ^ n2387 ^ 1'b0 ;
  assign n5545 = ( n3144 & n5542 ) | ( n3144 & n5544 ) | ( n5542 & n5544 ) ;
  assign n5546 = ( x3 & n2136 ) | ( x3 & n5174 ) | ( n2136 & n5174 ) ;
  assign n5547 = n3682 ^ n3441 ^ n1046 ;
  assign n5548 = n971 ^ n848 ^ 1'b0 ;
  assign n5549 = x12 & n5548 ;
  assign n5550 = ~n424 & n5549 ;
  assign n5551 = n5550 ^ n1426 ^ 1'b0 ;
  assign n5552 = n5547 | n5551 ;
  assign n5553 = n3540 | n5552 ;
  assign n5554 = n5553 ^ n424 ^ 1'b0 ;
  assign n5557 = n4367 ^ n315 ^ 1'b0 ;
  assign n5555 = n3025 ^ n1000 ^ 1'b0 ;
  assign n5556 = n2436 | n5555 ;
  assign n5558 = n5557 ^ n5556 ^ 1'b0 ;
  assign n5559 = ~n1758 & n5558 ;
  assign n5560 = n4518 ^ n292 ^ 1'b0 ;
  assign n5561 = n2377 ^ x94 ^ 1'b0 ;
  assign n5562 = ( n1733 & n2059 ) | ( n1733 & n3689 ) | ( n2059 & n3689 ) ;
  assign n5574 = n363 | n1676 ;
  assign n5575 = n1203 & ~n5574 ;
  assign n5576 = n490 & n5575 ;
  assign n5577 = n1928 | n5576 ;
  assign n5578 = n3636 & ~n5577 ;
  assign n5563 = n2389 & n4852 ;
  assign n5564 = n5563 ^ n2972 ^ n1397 ;
  assign n5565 = n1809 | n5564 ;
  assign n5566 = n5565 ^ n4769 ^ 1'b0 ;
  assign n5567 = ( n703 & ~n1608 ) | ( n703 & n3131 ) | ( ~n1608 & n3131 ) ;
  assign n5568 = n2728 & ~n5567 ;
  assign n5569 = n5568 ^ n2198 ^ 1'b0 ;
  assign n5570 = n4127 ^ n2748 ^ 1'b0 ;
  assign n5571 = ~n3579 & n5570 ;
  assign n5572 = n516 & n5571 ;
  assign n5573 = ( n5566 & n5569 ) | ( n5566 & ~n5572 ) | ( n5569 & ~n5572 ) ;
  assign n5579 = n5578 ^ n5573 ^ n5116 ;
  assign n5580 = ( n1357 & ~n1429 ) | ( n1357 & n2729 ) | ( ~n1429 & n2729 ) ;
  assign n5581 = n264 ^ x37 ^ 1'b0 ;
  assign n5582 = n1371 & ~n5581 ;
  assign n5583 = n1622 & ~n3380 ;
  assign n5584 = ~n5582 & n5583 ;
  assign n5585 = ( n3899 & n4307 ) | ( n3899 & n5584 ) | ( n4307 & n5584 ) ;
  assign n5586 = n3553 ^ n2905 ^ n1612 ;
  assign n5587 = n3973 ^ n2178 ^ n1472 ;
  assign n5590 = ( n948 & n4492 ) | ( n948 & ~n5098 ) | ( n4492 & ~n5098 ) ;
  assign n5588 = ( n597 & ~n1695 ) | ( n597 & n4655 ) | ( ~n1695 & n4655 ) ;
  assign n5589 = ~n5170 & n5588 ;
  assign n5591 = n5590 ^ n5589 ^ 1'b0 ;
  assign n5594 = n1993 ^ n1157 ^ 1'b0 ;
  assign n5595 = n199 & ~n5594 ;
  assign n5596 = n5595 ^ n3331 ^ n1704 ;
  assign n5592 = n2732 ^ n1070 ^ 1'b0 ;
  assign n5593 = ~n1170 & n5592 ;
  assign n5597 = n5596 ^ n5593 ^ 1'b0 ;
  assign n5598 = ( n1555 & n3362 ) | ( n1555 & ~n4679 ) | ( n3362 & ~n4679 ) ;
  assign n5599 = n5597 & n5598 ;
  assign n5600 = ~n5591 & n5599 ;
  assign n5601 = n2242 & ~n3946 ;
  assign n5602 = n2960 & ~n4199 ;
  assign n5603 = n5601 & n5602 ;
  assign n5604 = n5603 ^ n2987 ^ n454 ;
  assign n5605 = ( ~n262 & n3421 ) | ( ~n262 & n4255 ) | ( n3421 & n4255 ) ;
  assign n5606 = n2688 ^ n1364 ^ x56 ;
  assign n5607 = ~n1674 & n5606 ;
  assign n5608 = n5607 ^ n2851 ^ 1'b0 ;
  assign n5609 = n4101 ^ n1143 ^ n797 ;
  assign n5610 = n5231 ^ n4397 ^ 1'b0 ;
  assign n5611 = n5609 & ~n5610 ;
  assign n5612 = n5611 ^ n5349 ^ 1'b0 ;
  assign n5620 = n1267 | n3348 ;
  assign n5621 = n4387 & ~n5620 ;
  assign n5615 = x90 & n308 ;
  assign n5616 = n1840 & ~n3027 ;
  assign n5617 = n5615 | n5616 ;
  assign n5618 = n2366 & ~n5617 ;
  assign n5619 = n2931 | n5618 ;
  assign n5622 = n5621 ^ n5619 ^ 1'b0 ;
  assign n5613 = n3358 ^ n1654 ^ 1'b0 ;
  assign n5614 = ~n439 & n5613 ;
  assign n5623 = n5622 ^ n5614 ^ n2272 ;
  assign n5624 = ~n895 & n5251 ;
  assign n5625 = ~n415 & n5624 ;
  assign n5626 = n5170 | n5235 ;
  assign n5627 = n808 & n977 ;
  assign n5628 = n659 ^ n357 ^ 1'b0 ;
  assign n5629 = ~n5627 & n5628 ;
  assign n5630 = ( n695 & ~n2668 ) | ( n695 & n4704 ) | ( ~n2668 & n4704 ) ;
  assign n5631 = n3649 & ~n5630 ;
  assign n5632 = n5631 ^ n2377 ^ 1'b0 ;
  assign n5633 = ( n2406 & ~n5629 ) | ( n2406 & n5632 ) | ( ~n5629 & n5632 ) ;
  assign n5634 = n3576 ^ n1781 ^ n1270 ;
  assign n5635 = n2114 | n5634 ;
  assign n5637 = n3205 & ~n4980 ;
  assign n5638 = n5637 ^ n2671 ^ 1'b0 ;
  assign n5636 = n1767 & ~n2277 ;
  assign n5639 = n5638 ^ n5636 ^ 1'b0 ;
  assign n5640 = n5639 ^ n3362 ^ 1'b0 ;
  assign n5641 = n2267 ^ n2101 ^ n1472 ;
  assign n5642 = ~n4094 & n5641 ;
  assign n5643 = n5642 ^ n4086 ^ 1'b0 ;
  assign n5644 = ( n2535 & ~n2691 ) | ( n2535 & n5643 ) | ( ~n2691 & n5643 ) ;
  assign n5645 = ( n646 & ~n3321 ) | ( n646 & n5644 ) | ( ~n3321 & n5644 ) ;
  assign n5646 = n2653 ^ n242 ^ 1'b0 ;
  assign n5647 = ~n3069 & n5646 ;
  assign n5648 = n5647 ^ x70 ^ 1'b0 ;
  assign n5649 = n1731 & n5648 ;
  assign n5651 = ~n1132 & n5211 ;
  assign n5652 = n5651 ^ n251 ^ 1'b0 ;
  assign n5650 = n3227 ^ n920 ^ n157 ;
  assign n5653 = n5652 ^ n5650 ^ 1'b0 ;
  assign n5654 = n5649 & n5653 ;
  assign n5655 = n1635 ^ n890 ^ n672 ;
  assign n5656 = n4832 ^ n3547 ^ 1'b0 ;
  assign n5657 = n5655 & n5656 ;
  assign n5658 = n349 & n1378 ;
  assign n5659 = n5658 ^ n3588 ^ 1'b0 ;
  assign n5660 = ( n871 & n1439 ) | ( n871 & n5659 ) | ( n1439 & n5659 ) ;
  assign n5661 = ~n1783 & n4090 ;
  assign n5662 = n951 ^ x115 ^ 1'b0 ;
  assign n5663 = ( n5591 & ~n5661 ) | ( n5591 & n5662 ) | ( ~n5661 & n5662 ) ;
  assign n5664 = ~x108 & n883 ;
  assign n5665 = n5664 ^ n3581 ^ n3420 ;
  assign n5666 = ( n1131 & n2388 ) | ( n1131 & n5665 ) | ( n2388 & n5665 ) ;
  assign n5669 = n443 & ~n3212 ;
  assign n5670 = n5669 ^ n1160 ^ 1'b0 ;
  assign n5671 = n5670 ^ n1055 ^ 1'b0 ;
  assign n5672 = n4577 & n5671 ;
  assign n5673 = n5672 ^ n5218 ^ n1262 ;
  assign n5667 = ( n479 & n2839 ) | ( n479 & n3917 ) | ( n2839 & n3917 ) ;
  assign n5668 = n352 | n5667 ;
  assign n5674 = n5673 ^ n5668 ^ 1'b0 ;
  assign n5675 = ( n4008 & n5666 ) | ( n4008 & ~n5674 ) | ( n5666 & ~n5674 ) ;
  assign n5676 = ( n3728 & n4252 ) | ( n3728 & ~n4275 ) | ( n4252 & ~n4275 ) ;
  assign n5677 = n1094 & n2811 ;
  assign n5678 = n5677 ^ n1514 ^ 1'b0 ;
  assign n5679 = ( n1319 & ~n2539 ) | ( n1319 & n5678 ) | ( ~n2539 & n5678 ) ;
  assign n5680 = n5679 ^ n3035 ^ n2579 ;
  assign n5681 = n2908 | n3924 ;
  assign n5682 = ( n2300 & n5680 ) | ( n2300 & n5681 ) | ( n5680 & n5681 ) ;
  assign n5683 = n3998 & n5682 ;
  assign n5684 = n445 | n1758 ;
  assign n5685 = n5684 ^ n1184 ^ 1'b0 ;
  assign n5686 = n3513 ^ n2774 ^ n2198 ;
  assign n5687 = ~n4722 & n5686 ;
  assign n5688 = n1864 | n4004 ;
  assign n5689 = n5688 ^ n4085 ^ 1'b0 ;
  assign n5690 = n5689 ^ n1435 ^ n445 ;
  assign n5691 = n5434 & n5690 ;
  assign n5692 = n5428 ^ n4492 ^ n1819 ;
  assign n5693 = n4466 ^ n2513 ^ 1'b0 ;
  assign n5694 = n464 & n5693 ;
  assign n5700 = ( n584 & n813 ) | ( n584 & n4396 ) | ( n813 & n4396 ) ;
  assign n5695 = n2421 ^ n590 ^ n467 ;
  assign n5696 = n3567 & n5695 ;
  assign n5697 = n5696 ^ n5156 ^ 1'b0 ;
  assign n5698 = n5697 ^ n154 ^ 1'b0 ;
  assign n5699 = n5143 | n5698 ;
  assign n5701 = n5700 ^ n5699 ^ 1'b0 ;
  assign n5702 = n4760 ^ n4308 ^ n4100 ;
  assign n5703 = ~n2354 & n3583 ;
  assign n5704 = n5703 ^ n1321 ^ 1'b0 ;
  assign n5705 = ( ~n786 & n5702 ) | ( ~n786 & n5704 ) | ( n5702 & n5704 ) ;
  assign n5706 = ~n2927 & n3471 ;
  assign n5707 = n755 & n1185 ;
  assign n5708 = ( n678 & n1811 ) | ( n678 & n5707 ) | ( n1811 & n5707 ) ;
  assign n5709 = n4340 ^ n4030 ^ n270 ;
  assign n5710 = ~n2722 & n5661 ;
  assign n5711 = ~n2387 & n5710 ;
  assign n5713 = n384 & ~n4280 ;
  assign n5712 = n815 & ~n2170 ;
  assign n5714 = n5713 ^ n5712 ^ n190 ;
  assign n5715 = n5714 ^ n5579 ^ 1'b0 ;
  assign n5716 = n4691 ^ n3491 ^ 1'b0 ;
  assign n5717 = n1087 & n1609 ;
  assign n5718 = n3543 | n5717 ;
  assign n5719 = ( ~n1247 & n2344 ) | ( ~n1247 & n5718 ) | ( n2344 & n5718 ) ;
  assign n5720 = n5719 ^ n4892 ^ 1'b0 ;
  assign n5721 = ~n316 & n744 ;
  assign n5722 = n1656 & ~n1712 ;
  assign n5723 = ~n5721 & n5722 ;
  assign n5724 = ( ~n1764 & n2272 ) | ( ~n1764 & n5723 ) | ( n2272 & n5723 ) ;
  assign n5725 = n2385 ^ n1802 ^ 1'b0 ;
  assign n5726 = n559 | n5725 ;
  assign n5727 = n5726 ^ n1068 ^ 1'b0 ;
  assign n5728 = n1046 | n2608 ;
  assign n5729 = n5728 ^ n2914 ^ 1'b0 ;
  assign n5730 = n5727 & n5729 ;
  assign n5731 = ~n3100 & n3597 ;
  assign n5732 = n5731 ^ n724 ^ 1'b0 ;
  assign n5733 = n5714 ^ n2578 ^ 1'b0 ;
  assign n5734 = n1176 & ~n5733 ;
  assign n5735 = n1287 & n3498 ;
  assign n5736 = ( n358 & n3264 ) | ( n358 & n3686 ) | ( n3264 & n3686 ) ;
  assign n5737 = n3295 & ~n5736 ;
  assign n5738 = n5177 & n5737 ;
  assign n5739 = n1454 & n2296 ;
  assign n5740 = ~n3506 & n5234 ;
  assign n5741 = n5740 ^ n1839 ^ 1'b0 ;
  assign n5742 = ( ~n610 & n5739 ) | ( ~n610 & n5741 ) | ( n5739 & n5741 ) ;
  assign n5743 = ( n199 & ~n2299 ) | ( n199 & n5742 ) | ( ~n2299 & n5742 ) ;
  assign n5744 = n1899 & n1964 ;
  assign n5745 = n5744 ^ n1905 ^ 1'b0 ;
  assign n5746 = ( ~n1157 & n1718 ) | ( ~n1157 & n5745 ) | ( n1718 & n5745 ) ;
  assign n5747 = x37 & ~n1204 ;
  assign n5748 = n3488 & n5747 ;
  assign n5749 = n5748 ^ n4967 ^ 1'b0 ;
  assign n5750 = ~n3532 & n5749 ;
  assign n5751 = n4731 & n5750 ;
  assign n5759 = n3406 ^ n1876 ^ n501 ;
  assign n5760 = ( n280 & ~n2955 ) | ( n280 & n5759 ) | ( ~n2955 & n5759 ) ;
  assign n5766 = n1510 | n4252 ;
  assign n5761 = n4894 ^ n2879 ^ 1'b0 ;
  assign n5762 = n1527 & ~n5761 ;
  assign n5763 = n5762 ^ n5395 ^ n721 ;
  assign n5764 = n5763 ^ n4497 ^ n1430 ;
  assign n5765 = ( n3451 & n3797 ) | ( n3451 & n5764 ) | ( n3797 & n5764 ) ;
  assign n5767 = n5766 ^ n5765 ^ 1'b0 ;
  assign n5768 = ~n5760 & n5767 ;
  assign n5752 = n1780 ^ n1170 ^ 1'b0 ;
  assign n5753 = n522 & n5752 ;
  assign n5754 = n398 & n3643 ;
  assign n5755 = ~n5753 & n5754 ;
  assign n5756 = n2572 ^ n693 ^ x81 ;
  assign n5757 = n5756 ^ n4272 ^ n1213 ;
  assign n5758 = ~n5755 & n5757 ;
  assign n5769 = n5768 ^ n5758 ^ 1'b0 ;
  assign n5770 = x101 & ~n3653 ;
  assign n5771 = n5770 ^ n3550 ^ 1'b0 ;
  assign n5772 = ( n3346 & ~n5246 ) | ( n3346 & n5771 ) | ( ~n5246 & n5771 ) ;
  assign n5773 = ( ~n537 & n1019 ) | ( ~n537 & n2598 ) | ( n1019 & n2598 ) ;
  assign n5774 = n2767 | n5773 ;
  assign n5775 = ~n519 & n4260 ;
  assign n5776 = n5775 ^ n604 ^ 1'b0 ;
  assign n5777 = ~n5774 & n5776 ;
  assign n5778 = ~n4045 & n5777 ;
  assign n5779 = ( n357 & ~n574 ) | ( n357 & n2608 ) | ( ~n574 & n2608 ) ;
  assign n5780 = n5779 ^ n891 ^ n852 ;
  assign n5781 = ~n2891 & n3874 ;
  assign n5782 = n2300 & n5781 ;
  assign n5783 = n4800 | n5782 ;
  assign n5784 = n5783 ^ n5554 ^ 1'b0 ;
  assign n5788 = ( n1670 & n1999 ) | ( n1670 & n3633 ) | ( n1999 & n3633 ) ;
  assign n5785 = n3909 ^ n2265 ^ n1644 ;
  assign n5786 = n5785 ^ n4491 ^ 1'b0 ;
  assign n5787 = n5786 ^ n2074 ^ n1656 ;
  assign n5789 = n5788 ^ n5787 ^ 1'b0 ;
  assign n5790 = n474 & ~n1747 ;
  assign n5791 = n5790 ^ x99 ^ 1'b0 ;
  assign n5792 = n5791 ^ n2340 ^ n2246 ;
  assign n5793 = ( n452 & n786 ) | ( n452 & ~n5792 ) | ( n786 & ~n5792 ) ;
  assign n5800 = n491 ^ n458 ^ n246 ;
  assign n5801 = ~n1715 & n5800 ;
  assign n5799 = n3131 & ~n4171 ;
  assign n5794 = n3087 ^ n595 ^ 1'b0 ;
  assign n5795 = ~n2737 & n5794 ;
  assign n5796 = n5795 ^ n5766 ^ n1733 ;
  assign n5797 = n2514 & ~n3887 ;
  assign n5798 = ( n5623 & n5796 ) | ( n5623 & ~n5797 ) | ( n5796 & ~n5797 ) ;
  assign n5802 = n5801 ^ n5799 ^ n5798 ;
  assign n5803 = ( n2288 & n3844 ) | ( n2288 & n5431 ) | ( n3844 & n5431 ) ;
  assign n5804 = n3740 ^ n1583 ^ 1'b0 ;
  assign n5805 = n3139 ^ n1073 ^ n269 ;
  assign n5806 = ( n473 & n1309 ) | ( n473 & ~n5805 ) | ( n1309 & ~n5805 ) ;
  assign n5807 = n5806 ^ x80 ^ 1'b0 ;
  assign n5808 = n5661 ^ n4334 ^ n2819 ;
  assign n5809 = x13 & n500 ;
  assign n5810 = n1478 & n5809 ;
  assign n5811 = ( n347 & n504 ) | ( n347 & ~n2600 ) | ( n504 & ~n2600 ) ;
  assign n5812 = ~n5810 & n5811 ;
  assign n5813 = n366 & n1556 ;
  assign n5814 = n3440 & n5813 ;
  assign n5815 = n188 & n1739 ;
  assign n5816 = n2071 ^ n1764 ^ 1'b0 ;
  assign n5817 = n5815 & n5816 ;
  assign n5818 = n2981 & ~n4092 ;
  assign n5819 = n4103 ^ n2684 ^ n442 ;
  assign n5820 = n2343 & n2744 ;
  assign n5821 = ~n5819 & n5820 ;
  assign n5822 = n2493 ^ n1046 ^ x57 ;
  assign n5823 = n5822 ^ n541 ^ 1'b0 ;
  assign n5824 = n4485 ^ n3145 ^ 1'b0 ;
  assign n5825 = ( n817 & n5132 ) | ( n817 & n5824 ) | ( n5132 & n5824 ) ;
  assign n5826 = n5825 ^ n5041 ^ n3746 ;
  assign n5827 = n2453 ^ n2013 ^ 1'b0 ;
  assign n5828 = n3295 & n4998 ;
  assign n5829 = ~n2265 & n5828 ;
  assign n5830 = n4466 ^ n411 ^ 1'b0 ;
  assign n5831 = n1449 & ~n5830 ;
  assign n5832 = n4349 ^ n2175 ^ n447 ;
  assign n5833 = ( n203 & ~n5831 ) | ( n203 & n5832 ) | ( ~n5831 & n5832 ) ;
  assign n5835 = n4800 ^ n1406 ^ n403 ;
  assign n5836 = n5835 ^ n5377 ^ 1'b0 ;
  assign n5834 = n1361 & ~n3558 ;
  assign n5837 = n5836 ^ n5834 ^ 1'b0 ;
  assign n5838 = n4910 ^ n2264 ^ 1'b0 ;
  assign n5839 = ~n747 & n5838 ;
  assign n5840 = ~n178 & n2098 ;
  assign n5841 = n3099 | n5840 ;
  assign n5842 = n5841 ^ n2058 ^ 1'b0 ;
  assign n5843 = n3483 | n5842 ;
  assign n5844 = ~n1874 & n5843 ;
  assign n5845 = n5839 & ~n5844 ;
  assign n5846 = n5845 ^ n1897 ^ 1'b0 ;
  assign n5847 = n1771 ^ n1173 ^ 1'b0 ;
  assign n5848 = ~n2612 & n5847 ;
  assign n5849 = ~n1460 & n5026 ;
  assign n5850 = n5849 ^ x39 ^ 1'b0 ;
  assign n5851 = n5848 & n5850 ;
  assign n5852 = n1336 ^ n144 ^ 1'b0 ;
  assign n5853 = n3510 & n5852 ;
  assign n5854 = x123 & n5853 ;
  assign n5855 = ~n793 & n5854 ;
  assign n5857 = ( ~n161 & n436 ) | ( ~n161 & n1632 ) | ( n436 & n1632 ) ;
  assign n5856 = n287 & n2189 ;
  assign n5858 = n5857 ^ n5856 ^ 1'b0 ;
  assign n5859 = ~n1989 & n5858 ;
  assign n5860 = ~n867 & n5859 ;
  assign n5861 = n4046 & n5860 ;
  assign n5862 = n1145 ^ n361 ^ 1'b0 ;
  assign n5863 = n5861 & n5862 ;
  assign n5864 = x83 & n2692 ;
  assign n5865 = n1298 ^ n1199 ^ 1'b0 ;
  assign n5866 = n442 & n1108 ;
  assign n5867 = n5865 & ~n5866 ;
  assign n5868 = n3606 & n5097 ;
  assign n5869 = n2387 ^ n2299 ^ 1'b0 ;
  assign n5870 = x93 & ~n5869 ;
  assign n5871 = n5870 ^ n5450 ^ 1'b0 ;
  assign n5872 = n2625 | n5871 ;
  assign n5873 = n4163 ^ n1896 ^ n1189 ;
  assign n5874 = ~n824 & n5873 ;
  assign n5875 = n5874 ^ n4393 ^ 1'b0 ;
  assign n5876 = n5219 ^ n3840 ^ 1'b0 ;
  assign n5877 = n1542 & n5876 ;
  assign n5878 = ~n1277 & n5877 ;
  assign n5879 = n1731 & n3059 ;
  assign n5880 = n5879 ^ n1061 ^ 1'b0 ;
  assign n5881 = ( n5836 & ~n5878 ) | ( n5836 & n5880 ) | ( ~n5878 & n5880 ) ;
  assign n5882 = n4630 & n5687 ;
  assign n5883 = n5882 ^ x63 ^ 1'b0 ;
  assign n5884 = n1276 & ~n4728 ;
  assign n5885 = n5884 ^ n710 ^ 1'b0 ;
  assign n5886 = n224 & n955 ;
  assign n5887 = n5885 & n5886 ;
  assign n5888 = n5347 ^ n734 ^ n421 ;
  assign n5889 = n5888 ^ n4172 ^ n1979 ;
  assign n5892 = n664 | n2906 ;
  assign n5893 = n227 | n5892 ;
  assign n5894 = n5893 ^ n5530 ^ n5000 ;
  assign n5890 = ( ~n246 & n1104 ) | ( ~n246 & n2242 ) | ( n1104 & n2242 ) ;
  assign n5891 = x116 & ~n5890 ;
  assign n5895 = n5894 ^ n5891 ^ 1'b0 ;
  assign n5896 = ~n5889 & n5895 ;
  assign n5899 = n3319 ^ n1683 ^ 1'b0 ;
  assign n5897 = n406 ^ x44 ^ 1'b0 ;
  assign n5898 = n2082 | n5897 ;
  assign n5900 = n5899 ^ n5898 ^ n1798 ;
  assign n5901 = n5629 ^ n457 ^ 1'b0 ;
  assign n5902 = ~n361 & n5901 ;
  assign n5903 = ( ~n267 & n875 ) | ( ~n267 & n5902 ) | ( n875 & n5902 ) ;
  assign n5904 = n3357 ^ n770 ^ 1'b0 ;
  assign n5905 = n5904 ^ n5840 ^ n412 ;
  assign n5906 = n5905 ^ x22 ^ x6 ;
  assign n5907 = ( ~n2142 & n4401 ) | ( ~n2142 & n5906 ) | ( n4401 & n5906 ) ;
  assign n5908 = ~n1075 & n2960 ;
  assign n5909 = n5908 ^ n3337 ^ 1'b0 ;
  assign n5910 = ( n1473 & n5907 ) | ( n1473 & ~n5909 ) | ( n5907 & ~n5909 ) ;
  assign n5911 = ( n1762 & n5903 ) | ( n1762 & n5910 ) | ( n5903 & n5910 ) ;
  assign n5912 = n3093 ^ n1292 ^ 1'b0 ;
  assign n5913 = n4094 | n5912 ;
  assign n5914 = n2585 ^ n1253 ^ 1'b0 ;
  assign n5915 = n5914 ^ n1301 ^ 1'b0 ;
  assign n5916 = n5915 ^ n1251 ^ 1'b0 ;
  assign n5917 = n5096 & n5916 ;
  assign n5918 = x53 & ~n207 ;
  assign n5919 = n1108 & n5918 ;
  assign n5920 = n1278 & ~n3631 ;
  assign n5921 = n5634 & ~n5920 ;
  assign n5922 = n5921 ^ n4211 ^ 1'b0 ;
  assign n5923 = n1696 & n5922 ;
  assign n5924 = n5923 ^ n576 ^ 1'b0 ;
  assign n5925 = n5919 | n5924 ;
  assign n5931 = n3820 & n5353 ;
  assign n5932 = n5931 ^ n2516 ^ 1'b0 ;
  assign n5927 = n661 & ~n3374 ;
  assign n5928 = n5927 ^ n1572 ^ 1'b0 ;
  assign n5926 = n2956 & n4226 ;
  assign n5929 = n5928 ^ n5926 ^ 1'b0 ;
  assign n5930 = n2674 & ~n5929 ;
  assign n5933 = n5932 ^ n5930 ^ 1'b0 ;
  assign n5934 = n643 | n5259 ;
  assign n5935 = n5934 ^ n1057 ^ 1'b0 ;
  assign n5936 = n3551 & ~n5935 ;
  assign n5937 = n1691 ^ n599 ^ 1'b0 ;
  assign n5938 = n5278 ^ n4650 ^ n3867 ;
  assign n5939 = n840 ^ n763 ^ n541 ;
  assign n5946 = n5230 ^ n2534 ^ 1'b0 ;
  assign n5947 = n5488 & n5946 ;
  assign n5948 = n2385 & n5947 ;
  assign n5940 = n5432 ^ n993 ^ 1'b0 ;
  assign n5941 = n422 ^ n307 ^ 1'b0 ;
  assign n5942 = n3598 ^ n3497 ^ n2947 ;
  assign n5943 = n2534 & ~n5942 ;
  assign n5944 = n5941 & n5943 ;
  assign n5945 = ( n714 & ~n5940 ) | ( n714 & n5944 ) | ( ~n5940 & n5944 ) ;
  assign n5949 = n5948 ^ n5945 ^ n1769 ;
  assign n5950 = ~n1695 & n4606 ;
  assign n5951 = ~n3666 & n5950 ;
  assign n5952 = n2285 & n3282 ;
  assign n5953 = n5952 ^ n4889 ^ n2607 ;
  assign n5954 = n3575 ^ n2107 ^ n1957 ;
  assign n5955 = n821 | n1011 ;
  assign n5956 = ( x127 & n2802 ) | ( x127 & ~n3841 ) | ( n2802 & ~n3841 ) ;
  assign n5957 = n2449 & n3634 ;
  assign n5958 = n5957 ^ n3010 ^ 1'b0 ;
  assign n5959 = n5782 ^ n2869 ^ 1'b0 ;
  assign n5960 = ~n3239 & n5959 ;
  assign n5961 = ( n1006 & n1413 ) | ( n1006 & n2773 ) | ( n1413 & n2773 ) ;
  assign n5962 = n182 & ~n3091 ;
  assign n5963 = ~n5961 & n5962 ;
  assign n5965 = n154 & n3109 ;
  assign n5966 = n5965 ^ n2121 ^ n1910 ;
  assign n5967 = n5966 ^ n2356 ^ 1'b0 ;
  assign n5968 = ~n5618 & n5665 ;
  assign n5969 = ~n5967 & n5968 ;
  assign n5964 = ~n977 & n3896 ;
  assign n5970 = n5969 ^ n5964 ^ 1'b0 ;
  assign n5971 = ( ~n4230 & n5360 ) | ( ~n4230 & n5655 ) | ( n5360 & n5655 ) ;
  assign n5972 = n2426 ^ n349 ^ 1'b0 ;
  assign n5973 = ~n3613 & n5972 ;
  assign n5974 = n1083 & ~n2416 ;
  assign n5975 = n5974 ^ n5223 ^ 1'b0 ;
  assign n5976 = n5975 ^ n2027 ^ n1874 ;
  assign n5977 = n1184 & n3777 ;
  assign n5978 = n3073 ^ n141 ^ 1'b0 ;
  assign n5979 = ~n1580 & n5978 ;
  assign n5980 = n5979 ^ n1251 ^ 1'b0 ;
  assign n5981 = n2332 & n5980 ;
  assign n5982 = ~n1592 & n5981 ;
  assign n5983 = n3213 | n5982 ;
  assign n5984 = n5983 ^ n2297 ^ 1'b0 ;
  assign n5985 = n3105 | n5984 ;
  assign n5986 = n5985 ^ n3132 ^ 1'b0 ;
  assign n5987 = n403 | n4917 ;
  assign n5988 = n5986 | n5987 ;
  assign n5989 = x54 & ~n803 ;
  assign n5990 = ~n4310 & n5989 ;
  assign n5991 = n620 | n2470 ;
  assign n5992 = n5991 ^ n3503 ^ 1'b0 ;
  assign n5993 = ( n627 & n2489 ) | ( n627 & ~n3173 ) | ( n2489 & ~n3173 ) ;
  assign n5994 = n406 & ~n2316 ;
  assign n5995 = ~n298 & n5994 ;
  assign n5996 = n5993 & n5995 ;
  assign n5997 = n1236 ^ n149 ^ 1'b0 ;
  assign n5998 = n5997 ^ n1131 ^ 1'b0 ;
  assign n5999 = ~n5996 & n5998 ;
  assign n6001 = ~n2083 & n3399 ;
  assign n6002 = n6001 ^ n1591 ^ 1'b0 ;
  assign n6000 = n260 & ~n2432 ;
  assign n6003 = n6002 ^ n6000 ^ 1'b0 ;
  assign n6004 = n5865 ^ n2478 ^ 1'b0 ;
  assign n6005 = n999 & n4265 ;
  assign n6007 = ( ~x3 & n2391 ) | ( ~x3 & n3051 ) | ( n2391 & n3051 ) ;
  assign n6008 = n838 ^ n572 ^ 1'b0 ;
  assign n6009 = n6008 ^ n874 ^ 1'b0 ;
  assign n6010 = n2342 & ~n6009 ;
  assign n6011 = n5437 | n5575 ;
  assign n6012 = n6010 | n6011 ;
  assign n6013 = ( ~n3075 & n6007 ) | ( ~n3075 & n6012 ) | ( n6007 & n6012 ) ;
  assign n6006 = ~n1326 & n5289 ;
  assign n6014 = n6013 ^ n6006 ^ 1'b0 ;
  assign n6021 = ( ~n1538 & n2348 ) | ( ~n1538 & n3905 ) | ( n2348 & n3905 ) ;
  assign n6015 = n4832 ^ n2113 ^ 1'b0 ;
  assign n6016 = ~n3073 & n6015 ;
  assign n6017 = n6016 ^ n2679 ^ 1'b0 ;
  assign n6018 = n2375 & ~n6017 ;
  assign n6019 = ~n462 & n6018 ;
  assign n6020 = n3328 & n6019 ;
  assign n6022 = n6021 ^ n6020 ^ 1'b0 ;
  assign n6023 = n5521 ^ n1915 ^ 1'b0 ;
  assign n6024 = n2840 ^ n2077 ^ 1'b0 ;
  assign n6025 = x108 & ~n6024 ;
  assign n6026 = n6025 ^ n293 ^ 1'b0 ;
  assign n6027 = n508 | n5274 ;
  assign n6028 = ~n533 & n6027 ;
  assign n6029 = n6028 ^ n3442 ^ 1'b0 ;
  assign n6030 = n331 ^ n312 ^ 1'b0 ;
  assign n6031 = n3029 ^ n996 ^ 1'b0 ;
  assign n6032 = n6031 ^ n2344 ^ 1'b0 ;
  assign n6033 = n6030 & n6032 ;
  assign n6034 = n6033 ^ n1503 ^ 1'b0 ;
  assign n6035 = n6034 ^ n4214 ^ n4083 ;
  assign n6036 = n4441 & n5000 ;
  assign n6037 = n1044 ^ n241 ^ 1'b0 ;
  assign n6038 = n4808 & n6037 ;
  assign n6039 = ~n4989 & n6038 ;
  assign n6040 = n6039 ^ n5170 ^ 1'b0 ;
  assign n6041 = ( ~x69 & n1213 ) | ( ~x69 & n3633 ) | ( n1213 & n3633 ) ;
  assign n6042 = n3579 ^ n3004 ^ 1'b0 ;
  assign n6043 = ( n1354 & n6041 ) | ( n1354 & ~n6042 ) | ( n6041 & ~n6042 ) ;
  assign n6044 = n2998 ^ n1585 ^ 1'b0 ;
  assign n6045 = n3331 & n6044 ;
  assign n6046 = ( ~n1290 & n2322 ) | ( ~n1290 & n3491 ) | ( n2322 & n3491 ) ;
  assign n6048 = n1051 ^ n131 ^ 1'b0 ;
  assign n6049 = ( n923 & n2647 ) | ( n923 & n3100 ) | ( n2647 & n3100 ) ;
  assign n6050 = ~n6048 & n6049 ;
  assign n6047 = n2059 | n2213 ;
  assign n6051 = n6050 ^ n6047 ^ 1'b0 ;
  assign n6052 = n6046 & ~n6051 ;
  assign n6053 = ~n6045 & n6052 ;
  assign n6054 = ~n1682 & n2608 ;
  assign n6055 = ~n3379 & n6054 ;
  assign n6056 = n6053 | n6055 ;
  assign n6057 = n6056 ^ n5795 ^ 1'b0 ;
  assign n6058 = n2275 & ~n6057 ;
  assign n6059 = n570 | n3532 ;
  assign n6060 = ( ~n1044 & n5287 ) | ( ~n1044 & n6059 ) | ( n5287 & n6059 ) ;
  assign n6061 = ~n1932 & n6060 ;
  assign n6062 = ~n6058 & n6061 ;
  assign n6075 = ( n481 & n1635 ) | ( n481 & n2854 ) | ( n1635 & n2854 ) ;
  assign n6076 = n2285 & n6075 ;
  assign n6077 = ~n6075 & n6076 ;
  assign n6074 = n3698 ^ n3471 ^ 1'b0 ;
  assign n6064 = n2798 & ~n3527 ;
  assign n6065 = n2542 & n6064 ;
  assign n6063 = ( ~n406 & n1337 ) | ( ~n406 & n2215 ) | ( n1337 & n2215 ) ;
  assign n6066 = n6065 ^ n6063 ^ n2563 ;
  assign n6067 = n5261 ^ n2070 ^ 1'b0 ;
  assign n6068 = ( n1046 & n6066 ) | ( n1046 & ~n6067 ) | ( n6066 & ~n6067 ) ;
  assign n6070 = n134 | n2671 ;
  assign n6071 = n1849 & ~n6070 ;
  assign n6069 = n3133 & n5287 ;
  assign n6072 = n6071 ^ n6069 ^ 1'b0 ;
  assign n6073 = ( n3784 & n6068 ) | ( n3784 & ~n6072 ) | ( n6068 & ~n6072 ) ;
  assign n6078 = n6077 ^ n6074 ^ n6073 ;
  assign n6079 = x84 | n873 ;
  assign n6080 = n4373 & ~n6079 ;
  assign n6081 = n734 & ~n5432 ;
  assign n6082 = n6081 ^ n1819 ^ 1'b0 ;
  assign n6083 = n6082 ^ n4888 ^ 1'b0 ;
  assign n6084 = n4138 ^ n2992 ^ n1072 ;
  assign n6085 = ( ~n895 & n2715 ) | ( ~n895 & n3609 ) | ( n2715 & n3609 ) ;
  assign n6086 = n6084 & ~n6085 ;
  assign n6087 = n4327 | n6086 ;
  assign n6088 = n6083 & ~n6087 ;
  assign n6089 = n3903 ^ n1352 ^ n1317 ;
  assign n6090 = n6089 ^ n348 ^ 1'b0 ;
  assign n6091 = n3847 | n6090 ;
  assign n6101 = n5298 ^ n2709 ^ 1'b0 ;
  assign n6095 = n5935 ^ n3130 ^ n2913 ;
  assign n6096 = n6095 ^ n4103 ^ n3242 ;
  assign n6097 = n3235 & ~n6096 ;
  assign n6098 = n6097 ^ n1272 ^ 1'b0 ;
  assign n6092 = n559 | n1834 ;
  assign n6093 = x89 & n6092 ;
  assign n6094 = n495 & ~n6093 ;
  assign n6099 = n6098 ^ n6094 ^ 1'b0 ;
  assign n6100 = n6099 ^ n3930 ^ n1911 ;
  assign n6102 = n6101 ^ n6100 ^ 1'b0 ;
  assign n6103 = ( ~n1160 & n1548 ) | ( ~n1160 & n2001 ) | ( n1548 & n2001 ) ;
  assign n6104 = ( x99 & ~n4177 ) | ( x99 & n6103 ) | ( ~n4177 & n6103 ) ;
  assign n6105 = ( n298 & ~n392 ) | ( n298 & n1623 ) | ( ~n392 & n1623 ) ;
  assign n6106 = n490 & n6105 ;
  assign n6107 = n6104 & n6106 ;
  assign n6108 = n289 | n577 ;
  assign n6109 = n1976 & ~n6108 ;
  assign n6110 = n738 | n6109 ;
  assign n6111 = n6107 & ~n6110 ;
  assign n6112 = n6111 ^ n2947 ^ 1'b0 ;
  assign n6113 = ( ~n579 & n3703 ) | ( ~n579 & n5493 ) | ( n3703 & n5493 ) ;
  assign n6114 = ~n1687 & n4325 ;
  assign n6115 = n6113 & ~n6114 ;
  assign n6116 = n4599 & n6115 ;
  assign n6117 = n5728 ^ n3528 ^ 1'b0 ;
  assign n6118 = n182 | n6117 ;
  assign n6119 = ( n708 & n4904 ) | ( n708 & n6118 ) | ( n4904 & n6118 ) ;
  assign n6120 = n2490 ^ n2288 ^ x52 ;
  assign n6121 = n6119 & ~n6120 ;
  assign n6125 = n744 & ~n2296 ;
  assign n6122 = n4710 ^ n3700 ^ 1'b0 ;
  assign n6123 = ( n1538 & n2528 ) | ( n1538 & n6122 ) | ( n2528 & n6122 ) ;
  assign n6124 = n6123 ^ n6075 ^ n511 ;
  assign n6126 = n6125 ^ n6124 ^ n5701 ;
  assign n6127 = ( n1478 & n2780 ) | ( n1478 & n2906 ) | ( n2780 & n2906 ) ;
  assign n6128 = n4907 ^ n3544 ^ 1'b0 ;
  assign n6129 = ( x64 & n2284 ) | ( x64 & n2944 ) | ( n2284 & n2944 ) ;
  assign n6130 = n6129 ^ n232 ^ 1'b0 ;
  assign n6131 = n3998 ^ x67 ^ 1'b0 ;
  assign n6132 = n6130 | n6131 ;
  assign n6133 = n3246 & ~n6132 ;
  assign n6134 = n1780 | n6133 ;
  assign n6135 = n394 & ~n1580 ;
  assign n6136 = n3215 ^ n723 ^ 1'b0 ;
  assign n6137 = ( n1069 & ~n3264 ) | ( n1069 & n6136 ) | ( ~n3264 & n6136 ) ;
  assign n6138 = x80 | n579 ;
  assign n6139 = n2100 & n6138 ;
  assign n6140 = ( n1361 & n1419 ) | ( n1361 & n6139 ) | ( n1419 & n6139 ) ;
  assign n6141 = n1643 & ~n6140 ;
  assign n6142 = n6137 & n6141 ;
  assign n6143 = n2703 ^ n1097 ^ 1'b0 ;
  assign n6144 = n4196 ^ n3375 ^ 1'b0 ;
  assign n6145 = n6144 ^ n827 ^ 1'b0 ;
  assign n6146 = ( ~n935 & n1639 ) | ( ~n935 & n1731 ) | ( n1639 & n1731 ) ;
  assign n6147 = n6146 ^ n2042 ^ 1'b0 ;
  assign n6148 = n6147 ^ n4639 ^ n1623 ;
  assign n6149 = n4085 & n5440 ;
  assign n6150 = n2426 & n6149 ;
  assign n6151 = n6150 ^ n4524 ^ n3301 ;
  assign n6152 = n6151 ^ n5745 ^ 1'b0 ;
  assign n6153 = n2943 | n6152 ;
  assign n6154 = n1761 & ~n3133 ;
  assign n6155 = ~n2625 & n2815 ;
  assign n6156 = n5097 & n6155 ;
  assign n6157 = n4697 & ~n6156 ;
  assign n6158 = n6157 ^ n5572 ^ 1'b0 ;
  assign n6159 = ( n691 & ~n1190 ) | ( n691 & n1402 ) | ( ~n1190 & n1402 ) ;
  assign n6160 = n6159 ^ n3544 ^ 1'b0 ;
  assign n6161 = ~n3433 & n6160 ;
  assign n6162 = ( ~n307 & n405 ) | ( ~n307 & n813 ) | ( n405 & n813 ) ;
  assign n6163 = n6162 ^ n1794 ^ 1'b0 ;
  assign n6164 = n5339 ^ n2947 ^ x30 ;
  assign n6165 = ~n5616 & n6164 ;
  assign n6166 = ~n3183 & n6165 ;
  assign n6167 = ~n6163 & n6166 ;
  assign n6168 = n2453 ^ n1726 ^ 1'b0 ;
  assign n6169 = ( n1036 & n1586 ) | ( n1036 & ~n2401 ) | ( n1586 & ~n2401 ) ;
  assign n6170 = n4611 & n6169 ;
  assign n6171 = ( n1808 & n6168 ) | ( n1808 & n6170 ) | ( n6168 & n6170 ) ;
  assign n6172 = n6171 ^ n6164 ^ n2956 ;
  assign n6173 = n6172 ^ n4344 ^ n3022 ;
  assign n6174 = n1861 & ~n6173 ;
  assign n6175 = n6174 ^ n1688 ^ 1'b0 ;
  assign n6176 = ( n857 & ~n4256 ) | ( n857 & n5840 ) | ( ~n4256 & n5840 ) ;
  assign n6177 = n5243 & ~n6176 ;
  assign n6178 = n4424 & n6177 ;
  assign n6179 = n3775 & ~n6178 ;
  assign n6180 = n6179 ^ n2820 ^ 1'b0 ;
  assign n6181 = n2303 | n4214 ;
  assign n6182 = n6180 & ~n6181 ;
  assign n6183 = ( n3622 & n3633 ) | ( n3622 & ~n3940 ) | ( n3633 & ~n3940 ) ;
  assign n6184 = n418 & ~n2813 ;
  assign n6185 = n571 & n6184 ;
  assign n6186 = n890 & ~n6185 ;
  assign n6187 = ( n3696 & ~n3870 ) | ( n3696 & n6186 ) | ( ~n3870 & n6186 ) ;
  assign n6188 = n151 & ~n4401 ;
  assign n6189 = n1390 & n6188 ;
  assign n6190 = n6189 ^ n2400 ^ 1'b0 ;
  assign n6191 = n1260 ^ n383 ^ 1'b0 ;
  assign n6192 = ( n4132 & n4494 ) | ( n4132 & n6191 ) | ( n4494 & n6191 ) ;
  assign n6193 = ( n2624 & ~n4741 ) | ( n2624 & n6192 ) | ( ~n4741 & n6192 ) ;
  assign n6194 = n6190 | n6193 ;
  assign n6198 = n4405 ^ n2181 ^ x59 ;
  assign n6195 = n2539 ^ n1555 ^ 1'b0 ;
  assign n6196 = ~n1480 & n6195 ;
  assign n6197 = ( ~n809 & n1048 ) | ( ~n809 & n6196 ) | ( n1048 & n6196 ) ;
  assign n6199 = n6198 ^ n6197 ^ n3772 ;
  assign n6200 = n967 | n5479 ;
  assign n6201 = n6200 ^ n4765 ^ 1'b0 ;
  assign n6202 = n6126 ^ n4226 ^ 1'b0 ;
  assign n6203 = ( ~n1067 & n4163 ) | ( ~n1067 & n5374 ) | ( n4163 & n5374 ) ;
  assign n6204 = n4176 & n5570 ;
  assign n6205 = n2297 ^ n1242 ^ 1'b0 ;
  assign n6206 = n1067 & n6205 ;
  assign n6207 = ~n5546 & n6206 ;
  assign n6208 = n3734 ^ x49 ^ x4 ;
  assign n6209 = n1199 ^ n1057 ^ 1'b0 ;
  assign n6210 = n2095 ^ x78 ^ 1'b0 ;
  assign n6211 = n6210 ^ n176 ^ 1'b0 ;
  assign n6212 = n6211 ^ n2621 ^ 1'b0 ;
  assign n6213 = n2452 ^ n2060 ^ 1'b0 ;
  assign n6214 = n6213 ^ x52 ^ 1'b0 ;
  assign n6215 = ( n1333 & n3710 ) | ( n1333 & ~n6214 ) | ( n3710 & ~n6214 ) ;
  assign n6216 = n5270 ^ n4871 ^ n2296 ;
  assign n6217 = n6216 ^ n356 ^ n323 ;
  assign n6218 = n6065 ^ n3614 ^ n1853 ;
  assign n6219 = n2199 ^ n265 ^ 1'b0 ;
  assign n6220 = n4060 & n6219 ;
  assign n6221 = n6220 ^ n4087 ^ 1'b0 ;
  assign n6222 = n6218 & n6221 ;
  assign n6223 = n6222 ^ n3264 ^ 1'b0 ;
  assign n6224 = n2074 ^ n1390 ^ 1'b0 ;
  assign n6225 = n5686 | n6224 ;
  assign n6226 = n5160 & ~n6225 ;
  assign n6227 = n6226 ^ n408 ^ 1'b0 ;
  assign n6228 = n296 | n2217 ;
  assign n6229 = n1636 & ~n6228 ;
  assign n6230 = ~n831 & n3324 ;
  assign n6231 = n3911 ^ n3126 ^ n2151 ;
  assign n6232 = n2886 ^ n334 ^ 1'b0 ;
  assign n6233 = n4238 ^ n314 ^ 1'b0 ;
  assign n6234 = n612 | n6233 ;
  assign n6235 = n6234 ^ n493 ^ 1'b0 ;
  assign n6238 = ~n1180 & n1548 ;
  assign n6239 = n6238 ^ n1583 ^ 1'b0 ;
  assign n6236 = n2408 ^ n2072 ^ x113 ;
  assign n6237 = n1000 | n6236 ;
  assign n6240 = n6239 ^ n6237 ^ 1'b0 ;
  assign n6242 = n497 | n1721 ;
  assign n6243 = x94 & ~n6242 ;
  assign n6241 = n4820 ^ n3945 ^ 1'b0 ;
  assign n6244 = n6243 ^ n6241 ^ 1'b0 ;
  assign n6245 = n4014 ^ n681 ^ 1'b0 ;
  assign n6246 = n1080 & ~n1252 ;
  assign n6247 = n880 & ~n3909 ;
  assign n6248 = n4226 | n6247 ;
  assign n6249 = n6246 & n6248 ;
  assign n6250 = n599 & n888 ;
  assign n6251 = n5746 | n6250 ;
  assign n6252 = n6249 & ~n6251 ;
  assign n6255 = n685 | n1215 ;
  assign n6256 = n6255 ^ n1962 ^ 1'b0 ;
  assign n6253 = n1023 & n3281 ;
  assign n6254 = ~n869 & n6253 ;
  assign n6257 = n6256 ^ n6254 ^ 1'b0 ;
  assign n6258 = n1966 ^ x23 ^ 1'b0 ;
  assign n6259 = n6258 ^ n704 ^ 1'b0 ;
  assign n6260 = n6257 & n6259 ;
  assign n6262 = n4251 ^ n1324 ^ 1'b0 ;
  assign n6261 = n1017 ^ n255 ^ n178 ;
  assign n6263 = n6262 ^ n6261 ^ n1630 ;
  assign n6264 = ( n989 & ~n3661 ) | ( n989 & n6247 ) | ( ~n3661 & n6247 ) ;
  assign n6265 = ~n3955 & n6264 ;
  assign n6266 = ~n6263 & n6265 ;
  assign n6267 = ( n315 & ~n1889 ) | ( n315 & n6266 ) | ( ~n1889 & n6266 ) ;
  assign n6268 = n5438 ^ n3214 ^ n1302 ;
  assign n6273 = n3853 ^ n1203 ^ 1'b0 ;
  assign n6270 = n2739 & n5381 ;
  assign n6271 = n6270 ^ n1669 ^ 1'b0 ;
  assign n6269 = n2376 & n2717 ;
  assign n6272 = n6271 ^ n6269 ^ 1'b0 ;
  assign n6274 = n6273 ^ n6272 ^ n2119 ;
  assign n6275 = n6274 ^ n5985 ^ n810 ;
  assign n6276 = n1065 ^ n1032 ^ 1'b0 ;
  assign n6277 = ( ~n2493 & n6266 ) | ( ~n2493 & n6276 ) | ( n6266 & n6276 ) ;
  assign n6278 = n2822 ^ n972 ^ 1'b0 ;
  assign n6279 = n528 | n6278 ;
  assign n6280 = ( n171 & n5109 ) | ( n171 & n6279 ) | ( n5109 & n6279 ) ;
  assign n6281 = n3946 ^ n511 ^ 1'b0 ;
  assign n6282 = n308 | n6281 ;
  assign n6283 = n6282 ^ n1432 ^ 1'b0 ;
  assign n6284 = n2967 & n6283 ;
  assign n6285 = n171 & n898 ;
  assign n6286 = n6285 ^ n3297 ^ 1'b0 ;
  assign n6287 = n4634 ^ n3716 ^ n1089 ;
  assign n6288 = n6287 ^ n5985 ^ n4703 ;
  assign n6289 = n6288 ^ n2359 ^ 1'b0 ;
  assign n6290 = ( n1658 & ~n3612 ) | ( n1658 & n3975 ) | ( ~n3612 & n3975 ) ;
  assign n6298 = ( n486 & n707 ) | ( n486 & n1813 ) | ( n707 & n1813 ) ;
  assign n6299 = n6298 ^ n3059 ^ n493 ;
  assign n6291 = ( ~n749 & n1561 ) | ( ~n749 & n1635 ) | ( n1561 & n1635 ) ;
  assign n6294 = ( n509 & ~n1054 ) | ( n509 & n5211 ) | ( ~n1054 & n5211 ) ;
  assign n6292 = n890 ^ n219 ^ 1'b0 ;
  assign n6293 = ~n2511 & n6292 ;
  assign n6295 = n6294 ^ n6293 ^ n4658 ;
  assign n6296 = ( ~n429 & n6291 ) | ( ~n429 & n6295 ) | ( n6291 & n6295 ) ;
  assign n6297 = ~n1416 & n6296 ;
  assign n6300 = n6299 ^ n6297 ^ n5163 ;
  assign n6301 = n2962 ^ n2430 ^ n1736 ;
  assign n6302 = n6300 & n6301 ;
  assign n6303 = ~n3791 & n6302 ;
  assign n6309 = n3341 ^ n2295 ^ 1'b0 ;
  assign n6310 = n6309 ^ n1535 ^ n813 ;
  assign n6311 = n6310 ^ n1951 ^ n689 ;
  assign n6304 = ( n2215 & n3653 ) | ( n2215 & n3820 ) | ( n3653 & n3820 ) ;
  assign n6305 = n2251 & n2751 ;
  assign n6306 = n6305 ^ n2541 ^ 1'b0 ;
  assign n6307 = n6304 & ~n6306 ;
  assign n6308 = ~n2838 & n6307 ;
  assign n6312 = n6311 ^ n6308 ^ n5678 ;
  assign n6313 = n1850 & ~n5296 ;
  assign n6314 = ~n3379 & n6313 ;
  assign n6315 = ( n529 & n6312 ) | ( n529 & ~n6314 ) | ( n6312 & ~n6314 ) ;
  assign n6319 = ( n2844 & n3787 ) | ( n2844 & ~n4853 ) | ( n3787 & ~n4853 ) ;
  assign n6316 = n2704 ^ n1020 ^ n556 ;
  assign n6317 = n6316 ^ n4749 ^ n1277 ;
  assign n6318 = n277 | n6317 ;
  assign n6320 = n6319 ^ n6318 ^ 1'b0 ;
  assign n6321 = n5593 ^ x76 ^ 1'b0 ;
  assign n6322 = ( n383 & n964 ) | ( n383 & ~n5749 ) | ( n964 & ~n5749 ) ;
  assign n6323 = n1566 | n3137 ;
  assign n6324 = n4440 & ~n6323 ;
  assign n6325 = ( n2945 & n6322 ) | ( n2945 & ~n6324 ) | ( n6322 & ~n6324 ) ;
  assign n6326 = n6325 ^ n5578 ^ n1804 ;
  assign n6331 = ( ~x122 & n1520 ) | ( ~x122 & n2913 ) | ( n1520 & n2913 ) ;
  assign n6330 = n544 | n948 ;
  assign n6332 = n6331 ^ n6330 ^ n6206 ;
  assign n6333 = n6332 ^ n3282 ^ x12 ;
  assign n6327 = n4012 ^ n1266 ^ n908 ;
  assign n6328 = n192 | n6327 ;
  assign n6329 = n2999 | n6328 ;
  assign n6334 = n6333 ^ n6329 ^ 1'b0 ;
  assign n6336 = ( ~n608 & n1002 ) | ( ~n608 & n5811 ) | ( n1002 & n5811 ) ;
  assign n6335 = n2447 & n3135 ;
  assign n6337 = n6336 ^ n6335 ^ 1'b0 ;
  assign n6338 = n704 ^ n270 ^ 1'b0 ;
  assign n6339 = ~n1086 & n6164 ;
  assign n6340 = n6339 ^ n838 ^ 1'b0 ;
  assign n6341 = ( n4518 & n6338 ) | ( n4518 & n6340 ) | ( n6338 & n6340 ) ;
  assign n6342 = n4240 | n4423 ;
  assign n6344 = n2338 ^ x83 ^ 1'b0 ;
  assign n6343 = n776 ^ n738 ^ n454 ;
  assign n6345 = n6344 ^ n6343 ^ 1'b0 ;
  assign n6346 = ~n1889 & n3145 ;
  assign n6347 = n6346 ^ n3829 ^ 1'b0 ;
  assign n6348 = n6347 ^ n2433 ^ 1'b0 ;
  assign n6349 = n1060 & n6348 ;
  assign n6350 = n2062 | n6349 ;
  assign n6351 = n5064 ^ n986 ^ 1'b0 ;
  assign n6352 = ~n562 & n6351 ;
  assign n6353 = n6352 ^ n4778 ^ 1'b0 ;
  assign n6354 = n4181 & ~n6353 ;
  assign n6355 = n2134 ^ n770 ^ 1'b0 ;
  assign n6356 = x37 | n3375 ;
  assign n6357 = n6355 & ~n6356 ;
  assign n6358 = ~n1834 & n2365 ;
  assign n6359 = ( n2760 & n3874 ) | ( n2760 & ~n6358 ) | ( n3874 & ~n6358 ) ;
  assign n6360 = n4121 ^ n1769 ^ n1643 ;
  assign n6361 = n4339 ^ n1796 ^ 1'b0 ;
  assign n6362 = ( n4138 & ~n4156 ) | ( n4138 & n6361 ) | ( ~n4156 & n6361 ) ;
  assign n6363 = ( n1466 & ~n2240 ) | ( n1466 & n3798 ) | ( ~n2240 & n3798 ) ;
  assign n6364 = n1051 & ~n6363 ;
  assign n6365 = ~n1833 & n3050 ;
  assign n6366 = n3895 & n6365 ;
  assign n6367 = ~n903 & n4296 ;
  assign n6368 = n6367 ^ n3349 ^ 1'b0 ;
  assign n6369 = n6368 ^ n3105 ^ 1'b0 ;
  assign n6370 = n5810 | n6369 ;
  assign n6371 = n6366 | n6370 ;
  assign n6372 = n6364 & ~n6371 ;
  assign n6373 = n6372 ^ n1829 ^ 1'b0 ;
  assign n6374 = n1713 ^ n1490 ^ 1'b0 ;
  assign n6375 = n6374 ^ n4897 ^ 1'b0 ;
  assign n6376 = n3934 ^ x65 ^ 1'b0 ;
  assign n6377 = n6376 ^ n865 ^ 1'b0 ;
  assign n6378 = n2597 | n6377 ;
  assign n6379 = ( n1638 & ~n1666 ) | ( n1638 & n6378 ) | ( ~n1666 & n6378 ) ;
  assign n6380 = ( n4730 & ~n6375 ) | ( n4730 & n6379 ) | ( ~n6375 & n6379 ) ;
  assign n6381 = n4733 ^ n2112 ^ 1'b0 ;
  assign n6382 = x100 & n6381 ;
  assign n6383 = n2195 | n4476 ;
  assign n6384 = n6383 ^ n5375 ^ 1'b0 ;
  assign n6385 = n1086 & ~n2336 ;
  assign n6386 = ( n1194 & n6384 ) | ( n1194 & n6385 ) | ( n6384 & n6385 ) ;
  assign n6387 = n5397 ^ n1767 ^ n1246 ;
  assign n6388 = ( n755 & n3514 ) | ( n755 & n6387 ) | ( n3514 & n6387 ) ;
  assign n6389 = ~n1385 & n1689 ;
  assign n6390 = ~n6388 & n6389 ;
  assign n6391 = ( ~n6382 & n6386 ) | ( ~n6382 & n6390 ) | ( n6386 & n6390 ) ;
  assign n6392 = n6391 ^ x55 ^ 1'b0 ;
  assign n6393 = n6392 ^ n487 ^ n178 ;
  assign n6394 = ~n1137 & n2308 ;
  assign n6395 = n6393 & n6394 ;
  assign n6396 = n6395 ^ n3998 ^ 1'b0 ;
  assign n6397 = n2681 & n5890 ;
  assign n6398 = ~n773 & n6397 ;
  assign n6399 = n6398 ^ n441 ^ 1'b0 ;
  assign n6400 = ~n2326 & n4075 ;
  assign n6401 = ~n2430 & n6400 ;
  assign n6406 = ( n2165 & ~n2652 ) | ( n2165 & n4778 ) | ( ~n2652 & n4778 ) ;
  assign n6402 = n4221 ^ n2573 ^ n2131 ;
  assign n6403 = ( n1562 & n4517 ) | ( n1562 & n6402 ) | ( n4517 & n6402 ) ;
  assign n6404 = n2709 | n6403 ;
  assign n6405 = n6404 ^ n4699 ^ 1'b0 ;
  assign n6407 = n6406 ^ n6405 ^ 1'b0 ;
  assign n6408 = n5275 & n6407 ;
  assign n6409 = n4073 ^ n3729 ^ 1'b0 ;
  assign n6410 = n6409 ^ n5563 ^ x41 ;
  assign n6411 = n6410 ^ n2296 ^ 1'b0 ;
  assign n6412 = n2587 & ~n6411 ;
  assign n6413 = n2363 ^ n1597 ^ n401 ;
  assign n6414 = n6413 ^ n838 ^ 1'b0 ;
  assign n6415 = ( n1772 & ~n4991 ) | ( n1772 & n6414 ) | ( ~n4991 & n6414 ) ;
  assign n6416 = ( n180 & ~n1274 ) | ( n180 & n2917 ) | ( ~n1274 & n2917 ) ;
  assign n6417 = ( n1896 & ~n2674 ) | ( n1896 & n6416 ) | ( ~n2674 & n6416 ) ;
  assign n6418 = n5418 ^ n1415 ^ n204 ;
  assign n6419 = ( n2232 & n5415 ) | ( n2232 & ~n5963 ) | ( n5415 & ~n5963 ) ;
  assign n6420 = n4341 ^ n3613 ^ 1'b0 ;
  assign n6421 = n1256 ^ n318 ^ n146 ;
  assign n6422 = ( n2095 & n4792 ) | ( n2095 & ~n6421 ) | ( n4792 & ~n6421 ) ;
  assign n6423 = ~n1242 & n1627 ;
  assign n6424 = n6423 ^ n2205 ^ 1'b0 ;
  assign n6425 = ( n3168 & n5837 ) | ( n3168 & ~n6424 ) | ( n5837 & ~n6424 ) ;
  assign n6426 = n1149 & ~n5053 ;
  assign n6427 = n6426 ^ n3347 ^ 1'b0 ;
  assign n6428 = n2317 | n6427 ;
  assign n6430 = x53 & ~n1769 ;
  assign n6431 = n327 & n6430 ;
  assign n6432 = n6431 ^ n306 ^ 1'b0 ;
  assign n6429 = n3709 | n3883 ;
  assign n6433 = n6432 ^ n6429 ^ 1'b0 ;
  assign n6435 = n2487 & ~n2931 ;
  assign n6436 = n6435 ^ n787 ^ 1'b0 ;
  assign n6434 = n3382 ^ n1837 ^ 1'b0 ;
  assign n6437 = n6436 ^ n6434 ^ n3892 ;
  assign n6438 = n1096 ^ n689 ^ n620 ;
  assign n6439 = n3473 ^ n987 ^ 1'b0 ;
  assign n6440 = ( x30 & n768 ) | ( x30 & n5749 ) | ( n768 & n5749 ) ;
  assign n6441 = n6440 ^ n1153 ^ 1'b0 ;
  assign n6442 = n661 & n6441 ;
  assign n6443 = n3555 ^ n1770 ^ n1290 ;
  assign n6444 = n2638 & ~n3266 ;
  assign n6445 = n6443 & n6444 ;
  assign n6446 = ( n696 & n2101 ) | ( n696 & n3417 ) | ( n2101 & n3417 ) ;
  assign n6447 = n6446 ^ n738 ^ x86 ;
  assign n6449 = n1943 ^ n1113 ^ n506 ;
  assign n6450 = ~n5386 & n6449 ;
  assign n6448 = n2962 ^ n1969 ^ 1'b0 ;
  assign n6451 = n6450 ^ n6448 ^ n6416 ;
  assign n6452 = n6308 ^ n4493 ^ n2189 ;
  assign n6453 = n2422 & ~n6452 ;
  assign n6454 = n2217 ^ n1263 ^ 1'b0 ;
  assign n6455 = n5434 ^ n2805 ^ 1'b0 ;
  assign n6456 = n2515 ^ n1592 ^ n1252 ;
  assign n6457 = ~n4299 & n6456 ;
  assign n6458 = n6457 ^ n1837 ^ n1211 ;
  assign n6459 = ( n6454 & n6455 ) | ( n6454 & ~n6458 ) | ( n6455 & ~n6458 ) ;
  assign n6460 = n2440 ^ n1896 ^ 1'b0 ;
  assign n6461 = n5440 & n6460 ;
  assign n6462 = n6461 ^ n4034 ^ n2855 ;
  assign n6463 = n3715 ^ n1246 ^ 1'b0 ;
  assign n6465 = n889 & ~n3046 ;
  assign n6466 = n2992 & n6465 ;
  assign n6467 = n2981 ^ n2325 ^ n1699 ;
  assign n6468 = n129 & ~n6467 ;
  assign n6469 = n6466 & n6468 ;
  assign n6470 = n4710 | n6469 ;
  assign n6471 = n4527 & ~n6470 ;
  assign n6464 = n2141 & n4491 ;
  assign n6472 = n6471 ^ n6464 ^ 1'b0 ;
  assign n6479 = n6332 ^ n5054 ^ n3831 ;
  assign n6478 = n2493 | n3543 ;
  assign n6480 = n6479 ^ n6478 ^ 1'b0 ;
  assign n6481 = n4359 | n6480 ;
  assign n6482 = ( ~n1996 & n2970 ) | ( ~n1996 & n6481 ) | ( n2970 & n6481 ) ;
  assign n6473 = n1092 ^ x42 ^ 1'b0 ;
  assign n6474 = n6473 ^ n797 ^ 1'b0 ;
  assign n6475 = n455 & n6474 ;
  assign n6476 = n1038 & n6475 ;
  assign n6477 = n6476 ^ n1460 ^ 1'b0 ;
  assign n6483 = n6482 ^ n6477 ^ n3433 ;
  assign n6484 = ( n1808 & n1820 ) | ( n1808 & ~n2059 ) | ( n1820 & ~n2059 ) ;
  assign n6485 = ( n1547 & n2261 ) | ( n1547 & n3982 ) | ( n2261 & n3982 ) ;
  assign n6486 = n3349 & ~n6485 ;
  assign n6487 = n6484 & n6486 ;
  assign n6488 = n6487 ^ n2404 ^ 1'b0 ;
  assign n6494 = ( ~n1816 & n4611 ) | ( ~n1816 & n4828 ) | ( n4611 & n4828 ) ;
  assign n6495 = n6494 ^ n965 ^ 1'b0 ;
  assign n6492 = n363 | n2112 ;
  assign n6491 = ( x56 & ~n3049 ) | ( x56 & n4841 ) | ( ~n3049 & n4841 ) ;
  assign n6493 = n6492 ^ n6491 ^ n845 ;
  assign n6489 = n153 & n1925 ;
  assign n6490 = n4052 | n6489 ;
  assign n6496 = n6495 ^ n6493 ^ n6490 ;
  assign n6498 = n1579 ^ n538 ^ 1'b0 ;
  assign n6499 = n6498 ^ n3097 ^ 1'b0 ;
  assign n6500 = ~n4169 & n6499 ;
  assign n6497 = n3489 ^ x112 ^ 1'b0 ;
  assign n6501 = n6500 ^ n6497 ^ n227 ;
  assign n6506 = n1989 & ~n2156 ;
  assign n6507 = n6506 ^ n4100 ^ n1848 ;
  assign n6502 = ( x112 & n797 ) | ( x112 & ~n2248 ) | ( n797 & ~n2248 ) ;
  assign n6503 = n6502 ^ n955 ^ x70 ;
  assign n6504 = ~n383 & n6503 ;
  assign n6505 = n999 & n6504 ;
  assign n6508 = n6507 ^ n6505 ^ 1'b0 ;
  assign n6509 = n734 & ~n2072 ;
  assign n6510 = ~n3386 & n6509 ;
  assign n6511 = n3409 ^ n2934 ^ n1839 ;
  assign n6512 = n6511 ^ n664 ^ n511 ;
  assign n6514 = n874 | n1013 ;
  assign n6515 = n6514 ^ n2684 ^ 1'b0 ;
  assign n6513 = n2698 ^ n2290 ^ 1'b0 ;
  assign n6516 = n6515 ^ n6513 ^ n4108 ;
  assign n6517 = ~n6512 & n6516 ;
  assign n6518 = n6517 ^ n1834 ^ 1'b0 ;
  assign n6519 = n4220 | n6401 ;
  assign n6520 = n5512 ^ n3200 ^ x17 ;
  assign n6521 = n1363 | n2518 ;
  assign n6522 = n6521 ^ n725 ^ 1'b0 ;
  assign n6523 = n6522 ^ n2660 ^ 1'b0 ;
  assign n6524 = n3569 ^ n875 ^ n411 ;
  assign n6525 = n6524 ^ n4578 ^ 1'b0 ;
  assign n6529 = n3694 ^ n3072 ^ n1253 ;
  assign n6530 = n6529 ^ n3792 ^ n1726 ;
  assign n6531 = n903 ^ n744 ^ 1'b0 ;
  assign n6532 = n6530 | n6531 ;
  assign n6526 = n3013 ^ n679 ^ 1'b0 ;
  assign n6527 = n1146 | n6526 ;
  assign n6528 = ( ~n274 & n2819 ) | ( ~n274 & n6527 ) | ( n2819 & n6527 ) ;
  assign n6533 = n6532 ^ n6528 ^ 1'b0 ;
  assign n6534 = ( n280 & ~n3595 ) | ( n280 & n4190 ) | ( ~n3595 & n4190 ) ;
  assign n6535 = n6534 ^ n346 ^ 1'b0 ;
  assign n6540 = n2569 & n4650 ;
  assign n6541 = ~n4356 & n6540 ;
  assign n6536 = ~n2355 & n5493 ;
  assign n6537 = ~n5493 & n6536 ;
  assign n6538 = n1078 & n5172 ;
  assign n6539 = n6537 & n6538 ;
  assign n6542 = n6541 ^ n6539 ^ n540 ;
  assign n6543 = n1244 & ~n3161 ;
  assign n6544 = ~n991 & n6543 ;
  assign n6545 = n6544 ^ n4774 ^ 1'b0 ;
  assign n6546 = n6545 ^ n6084 ^ n333 ;
  assign n6547 = ( n2513 & ~n2794 ) | ( n2513 & n6546 ) | ( ~n2794 & n6546 ) ;
  assign n6548 = ~n1804 & n4647 ;
  assign n6549 = ( ~n241 & n6547 ) | ( ~n241 & n6548 ) | ( n6547 & n6548 ) ;
  assign n6554 = n2127 ^ n1802 ^ n287 ;
  assign n6550 = n4090 & ~n4836 ;
  assign n6551 = ~n4158 & n6550 ;
  assign n6552 = ~n577 & n1490 ;
  assign n6553 = n6551 & n6552 ;
  assign n6555 = n6554 ^ n6553 ^ n5717 ;
  assign n6556 = ~n1754 & n6555 ;
  assign n6557 = n6556 ^ n751 ^ 1'b0 ;
  assign n6558 = n3450 & ~n6557 ;
  assign n6559 = n3459 ^ n3069 ^ n824 ;
  assign n6560 = n6559 ^ n6366 ^ 1'b0 ;
  assign n6561 = n6558 & ~n6560 ;
  assign n6562 = n1355 | n5919 ;
  assign n6563 = n807 & ~n6562 ;
  assign n6564 = ~n6561 & n6563 ;
  assign n6565 = n673 | n1129 ;
  assign n6566 = ( n533 & ~n2072 ) | ( n533 & n6565 ) | ( ~n2072 & n6565 ) ;
  assign n6567 = n247 | n6566 ;
  assign n6568 = n2537 | n6567 ;
  assign n6569 = n5171 ^ n719 ^ 1'b0 ;
  assign n6570 = n1537 ^ n535 ^ 1'b0 ;
  assign n6571 = ( n1254 & ~n6050 ) | ( n1254 & n6570 ) | ( ~n6050 & n6570 ) ;
  assign n6574 = n184 | n1819 ;
  assign n6575 = x43 | n6574 ;
  assign n6576 = ( n1468 & ~n2693 ) | ( n1468 & n6575 ) | ( ~n2693 & n6575 ) ;
  assign n6572 = n4233 ^ n935 ^ n158 ;
  assign n6573 = n3668 & n6572 ;
  assign n6577 = n6576 ^ n6573 ^ 1'b0 ;
  assign n6578 = n6577 ^ n3966 ^ 1'b0 ;
  assign n6579 = n5437 ^ n4600 ^ n2582 ;
  assign n6580 = n6579 ^ n3903 ^ 1'b0 ;
  assign n6581 = n6248 ^ n4180 ^ n3144 ;
  assign n6582 = n6581 ^ n4783 ^ 1'b0 ;
  assign n6586 = ( n889 & ~n1254 ) | ( n889 & n2143 ) | ( ~n1254 & n2143 ) ;
  assign n6584 = ~n338 & n4020 ;
  assign n6585 = n6584 ^ n1084 ^ 1'b0 ;
  assign n6583 = ( n2631 & ~n2885 ) | ( n2631 & n3174 ) | ( ~n2885 & n3174 ) ;
  assign n6587 = n6586 ^ n6585 ^ n6583 ;
  assign n6588 = n2298 ^ n1702 ^ n1484 ;
  assign n6589 = n1944 | n6588 ;
  assign n6590 = n5471 & ~n6589 ;
  assign n6591 = n1583 ^ x31 ^ 1'b0 ;
  assign n6592 = n6591 ^ n5928 ^ n5163 ;
  assign n6593 = n6590 | n6592 ;
  assign n6594 = n5121 ^ n3081 ^ n1515 ;
  assign n6595 = n6594 ^ n2723 ^ 1'b0 ;
  assign n6596 = n3945 & ~n6595 ;
  assign n6597 = n6596 ^ n1068 ^ 1'b0 ;
  assign n6598 = n5122 | n6597 ;
  assign n6599 = n538 & n6546 ;
  assign n6600 = ( n528 & n2445 ) | ( n528 & n6599 ) | ( n2445 & n6599 ) ;
  assign n6606 = n994 ^ x100 ^ 1'b0 ;
  assign n6607 = n439 | n6606 ;
  assign n6603 = n1341 ^ n1193 ^ 1'b0 ;
  assign n6604 = ~n352 & n6603 ;
  assign n6605 = n6604 ^ n1078 ^ n549 ;
  assign n6608 = n6607 ^ n6605 ^ 1'b0 ;
  assign n6609 = n516 & n6608 ;
  assign n6601 = n2377 ^ n786 ^ 1'b0 ;
  assign n6602 = ~n3681 & n6601 ;
  assign n6610 = n6609 ^ n6602 ^ 1'b0 ;
  assign n6611 = ~n6600 & n6610 ;
  assign n6612 = n1623 & n6611 ;
  assign n6613 = n6598 & n6612 ;
  assign n6614 = ( n1713 & n2763 ) | ( n1713 & ~n4197 ) | ( n2763 & ~n4197 ) ;
  assign n6619 = n485 | n1543 ;
  assign n6620 = n3221 | n6079 ;
  assign n6621 = n6620 ^ n3411 ^ 1'b0 ;
  assign n6622 = n6619 | n6621 ;
  assign n6615 = n943 & n3630 ;
  assign n6616 = n5627 & n6615 ;
  assign n6617 = n4226 & n6616 ;
  assign n6618 = n599 & n6617 ;
  assign n6623 = n6622 ^ n6618 ^ 1'b0 ;
  assign n6624 = n6623 ^ n3124 ^ 1'b0 ;
  assign n6625 = n2587 | n4347 ;
  assign n6626 = n1083 & ~n6140 ;
  assign n6627 = n6626 ^ n6479 ^ 1'b0 ;
  assign n6628 = n2688 & ~n3311 ;
  assign n6629 = n6628 ^ n4120 ^ 1'b0 ;
  assign n6630 = n1954 ^ n1882 ^ 1'b0 ;
  assign n6631 = n168 & ~n5323 ;
  assign n6632 = n6631 ^ n3188 ^ 1'b0 ;
  assign n6633 = n2322 & ~n4681 ;
  assign n6634 = n1404 & n5842 ;
  assign n6635 = ~n3998 & n6634 ;
  assign n6636 = n6635 ^ n4450 ^ n3052 ;
  assign n6637 = n6636 ^ n3382 ^ n396 ;
  assign n6638 = ~n331 & n1120 ;
  assign n6639 = ~x67 & n6638 ;
  assign n6640 = ( ~n5390 & n6332 ) | ( ~n5390 & n6639 ) | ( n6332 & n6639 ) ;
  assign n6641 = ~n6637 & n6640 ;
  assign n6642 = n2913 & ~n6605 ;
  assign n6643 = n2788 & ~n3971 ;
  assign n6644 = n6643 ^ n1912 ^ 1'b0 ;
  assign n6645 = n2652 & ~n6644 ;
  assign n6646 = ~n6642 & n6645 ;
  assign n6647 = n6646 ^ n4732 ^ 1'b0 ;
  assign n6648 = n3463 ^ n1226 ^ 1'b0 ;
  assign n6649 = ~n5014 & n6648 ;
  assign n6650 = n3674 & n6649 ;
  assign n6651 = n6650 ^ n2131 ^ 1'b0 ;
  assign n6652 = n3374 ^ n2239 ^ n1246 ;
  assign n6653 = ( n525 & n4227 ) | ( n525 & ~n6652 ) | ( n4227 & ~n6652 ) ;
  assign n6654 = n4120 ^ n2836 ^ 1'b0 ;
  assign n6655 = n6654 ^ n4673 ^ n4415 ;
  assign n6656 = n4415 ^ n3326 ^ n894 ;
  assign n6657 = n4318 & ~n6656 ;
  assign n6661 = n6224 ^ n211 ^ 1'b0 ;
  assign n6662 = n3698 & n6661 ;
  assign n6658 = n1409 & n6528 ;
  assign n6659 = n6658 ^ n3349 ^ 1'b0 ;
  assign n6660 = ~n1940 & n6659 ;
  assign n6663 = n6662 ^ n6660 ^ 1'b0 ;
  assign n6664 = ~n1013 & n3253 ;
  assign n6665 = n6664 ^ n3258 ^ 1'b0 ;
  assign n6666 = n1898 & ~n6665 ;
  assign n6667 = n949 & ~n2748 ;
  assign n6668 = n2673 & n6667 ;
  assign n6669 = ( ~n3473 & n4101 ) | ( ~n3473 & n4660 ) | ( n4101 & n4660 ) ;
  assign n6670 = ( n3286 & n6668 ) | ( n3286 & n6669 ) | ( n6668 & n6669 ) ;
  assign n6671 = n2372 | n6670 ;
  assign n6672 = n689 | n6671 ;
  assign n6673 = ( n1761 & n6071 ) | ( n1761 & ~n6672 ) | ( n6071 & ~n6672 ) ;
  assign n6674 = n870 ^ x47 ^ 1'b0 ;
  assign n6675 = ( n580 & ~n1348 ) | ( n580 & n3776 ) | ( ~n1348 & n3776 ) ;
  assign n6676 = n6675 ^ n5788 ^ n3273 ;
  assign n6677 = ( ~x73 & n5065 ) | ( ~x73 & n6676 ) | ( n5065 & n6676 ) ;
  assign n6678 = n719 ^ n675 ^ 1'b0 ;
  assign n6679 = n6678 ^ n5120 ^ n264 ;
  assign n6680 = n608 & ~n1756 ;
  assign n6681 = n6680 ^ n293 ^ 1'b0 ;
  assign n6682 = n2061 | n2214 ;
  assign n6683 = n6682 ^ n478 ^ 1'b0 ;
  assign n6684 = n6683 ^ n2636 ^ n2190 ;
  assign n6685 = n6684 ^ n4135 ^ 1'b0 ;
  assign n6686 = n3134 ^ n1131 ^ 1'b0 ;
  assign n6687 = n3799 | n6686 ;
  assign n6688 = ~n265 & n4679 ;
  assign n6689 = n6688 ^ n2228 ^ 1'b0 ;
  assign n6690 = ( n449 & ~n1803 ) | ( n449 & n6233 ) | ( ~n1803 & n6233 ) ;
  assign n6691 = ~n3273 & n6690 ;
  assign n6692 = n6691 ^ n370 ^ 1'b0 ;
  assign n6693 = n6527 ^ n456 ^ 1'b0 ;
  assign n6694 = ~n6692 & n6693 ;
  assign n6695 = n6694 ^ n3076 ^ n1877 ;
  assign n6701 = n1062 ^ n851 ^ x40 ;
  assign n6696 = n184 | n471 ;
  assign n6697 = n2172 | n6696 ;
  assign n6698 = n2263 & n6697 ;
  assign n6699 = n6698 ^ n1789 ^ 1'b0 ;
  assign n6700 = n6699 ^ n5441 ^ n323 ;
  assign n6702 = n6701 ^ n6700 ^ n5281 ;
  assign n6703 = n4469 ^ n3403 ^ n604 ;
  assign n6704 = n5823 | n6703 ;
  assign n6705 = n5729 & n6704 ;
  assign n6706 = ( n725 & n1616 ) | ( n725 & ~n4561 ) | ( n1616 & ~n4561 ) ;
  assign n6707 = ( ~n890 & n1056 ) | ( ~n890 & n4703 ) | ( n1056 & n4703 ) ;
  assign n6708 = n6707 ^ n3120 ^ 1'b0 ;
  assign n6709 = n5172 & n6708 ;
  assign n6714 = n1543 ^ n1104 ^ 1'b0 ;
  assign n6710 = n5928 ^ n3133 ^ n1199 ;
  assign n6711 = ( n370 & ~n559 ) | ( n370 & n6534 ) | ( ~n559 & n6534 ) ;
  assign n6712 = ~n1132 & n6711 ;
  assign n6713 = ~n6710 & n6712 ;
  assign n6715 = n6714 ^ n6713 ^ 1'b0 ;
  assign n6716 = n3688 & ~n6345 ;
  assign n6717 = n6715 & n6716 ;
  assign n6718 = n4569 & ~n5215 ;
  assign n6719 = n6718 ^ x13 ^ 1'b0 ;
  assign n6720 = n1912 & ~n2377 ;
  assign n6721 = n6720 ^ n6215 ^ 1'b0 ;
  assign n6722 = n6256 ^ n2166 ^ n339 ;
  assign n6723 = n3476 | n4972 ;
  assign n6724 = n367 | n2766 ;
  assign n6725 = n6724 ^ n971 ^ 1'b0 ;
  assign n6726 = n6725 ^ n3521 ^ n1738 ;
  assign n6727 = n6726 ^ n554 ^ 1'b0 ;
  assign n6728 = n2460 | n6727 ;
  assign n6729 = n6728 ^ n6611 ^ 1'b0 ;
  assign n6730 = n2494 | n6729 ;
  assign n6731 = n6730 ^ n2129 ^ 1'b0 ;
  assign n6732 = ( ~n4179 & n4313 ) | ( ~n4179 & n6731 ) | ( n4313 & n6731 ) ;
  assign n6733 = n3772 & ~n5166 ;
  assign n6734 = n6392 ^ n2959 ^ 1'b0 ;
  assign n6735 = n6390 ^ n269 ^ 1'b0 ;
  assign n6736 = n3002 & n6735 ;
  assign n6737 = n6736 ^ n4594 ^ n3588 ;
  assign n6738 = n6734 & ~n6737 ;
  assign n6739 = n6738 ^ n3956 ^ 1'b0 ;
  assign n6740 = n2331 ^ n246 ^ 1'b0 ;
  assign n6741 = n6740 ^ n2060 ^ 1'b0 ;
  assign n6742 = x119 & ~n6741 ;
  assign n6743 = n1872 & ~n3047 ;
  assign n6744 = n4952 ^ n2631 ^ 1'b0 ;
  assign n6745 = ~n2356 & n3927 ;
  assign n6746 = n6745 ^ n3477 ^ 1'b0 ;
  assign n6747 = n1535 | n6746 ;
  assign n6748 = n6155 & ~n6747 ;
  assign n6749 = n6528 ^ n1400 ^ 1'b0 ;
  assign n6750 = n3174 & ~n3498 ;
  assign n6751 = n262 | n2889 ;
  assign n6752 = ( ~n4622 & n6750 ) | ( ~n4622 & n6751 ) | ( n6750 & n6751 ) ;
  assign n6753 = ~n885 & n2994 ;
  assign n6754 = n2914 & n6753 ;
  assign n6755 = ( ~n296 & n708 ) | ( ~n296 & n4073 ) | ( n708 & n4073 ) ;
  assign n6756 = ~n6754 & n6755 ;
  assign n6757 = n6756 ^ n4529 ^ 1'b0 ;
  assign n6758 = n5729 & ~n6757 ;
  assign n6759 = ~n296 & n383 ;
  assign n6760 = n6759 ^ n4327 ^ n2707 ;
  assign n6761 = ( n204 & ~n2623 ) | ( n204 & n6760 ) | ( ~n2623 & n6760 ) ;
  assign n6762 = n3220 | n6331 ;
  assign n6763 = n1872 & ~n6762 ;
  assign n6764 = n6050 | n6763 ;
  assign n6765 = n6761 | n6764 ;
  assign n6766 = n2872 & n6765 ;
  assign n6767 = ~n4185 & n6766 ;
  assign n6768 = ~n1240 & n1663 ;
  assign n6769 = ( n954 & n1482 ) | ( n954 & ~n6768 ) | ( n1482 & ~n6768 ) ;
  assign n6770 = n1767 & ~n2521 ;
  assign n6771 = n1728 | n6770 ;
  assign n6772 = n6771 ^ n2340 ^ 1'b0 ;
  assign n6773 = n723 ^ n668 ^ 1'b0 ;
  assign n6774 = n6772 | n6773 ;
  assign n6775 = n1762 ^ n500 ^ 1'b0 ;
  assign n6776 = n3672 ^ n851 ^ 1'b0 ;
  assign n6777 = n5367 | n6776 ;
  assign n6779 = ~n2014 & n2993 ;
  assign n6778 = ~n3856 & n4945 ;
  assign n6780 = n6779 ^ n6778 ^ 1'b0 ;
  assign n6781 = n6780 ^ n4232 ^ n867 ;
  assign n6782 = n6777 | n6781 ;
  assign n6783 = n2025 & ~n6782 ;
  assign n6784 = ( n381 & n6775 ) | ( n381 & n6783 ) | ( n6775 & n6783 ) ;
  assign n6785 = n1063 ^ n514 ^ 1'b0 ;
  assign n6786 = n3951 ^ n1498 ^ 1'b0 ;
  assign n6787 = ( n2969 & n4010 ) | ( n2969 & ~n6786 ) | ( n4010 & ~n6786 ) ;
  assign n6788 = n6785 & n6787 ;
  assign n6789 = ~n1688 & n6788 ;
  assign n6790 = n171 ^ x51 ^ 1'b0 ;
  assign n6791 = n5182 | n6790 ;
  assign n6792 = n1143 & ~n1838 ;
  assign n6793 = n6792 ^ n550 ^ 1'b0 ;
  assign n6794 = x66 & ~n1519 ;
  assign n6795 = ~n6336 & n6794 ;
  assign n6796 = n6793 & n6795 ;
  assign n6797 = n1830 ^ n219 ^ 1'b0 ;
  assign n6798 = n6797 ^ n1799 ^ 1'b0 ;
  assign n6799 = ~n1333 & n6798 ;
  assign n6800 = n6799 ^ n2794 ^ n2701 ;
  assign n6801 = n6800 ^ n4164 ^ 1'b0 ;
  assign n6802 = n6796 | n6801 ;
  assign n6803 = n266 & n2738 ;
  assign n6804 = n6803 ^ n1126 ^ 1'b0 ;
  assign n6805 = n657 & n3049 ;
  assign n6806 = ~n4592 & n6805 ;
  assign n6807 = n6806 ^ n3639 ^ 1'b0 ;
  assign n6808 = n6807 ^ n4858 ^ 1'b0 ;
  assign n6809 = n5890 ^ n3067 ^ n596 ;
  assign n6810 = n1056 ^ n680 ^ 1'b0 ;
  assign n6811 = ~n2869 & n6810 ;
  assign n6812 = n6811 ^ n483 ^ 1'b0 ;
  assign n6813 = n6809 & ~n6812 ;
  assign n6814 = n6030 ^ n2368 ^ n737 ;
  assign n6815 = n3440 & n6814 ;
  assign n6816 = n3086 & ~n3972 ;
  assign n6817 = ( n396 & n2639 ) | ( n396 & ~n6816 ) | ( n2639 & ~n6816 ) ;
  assign n6818 = n2798 ^ n2608 ^ n466 ;
  assign n6819 = n6449 | n6818 ;
  assign n6820 = n2579 ^ n1394 ^ 1'b0 ;
  assign n6821 = n2115 | n6820 ;
  assign n6822 = n2313 & ~n6821 ;
  assign n6823 = ( n842 & n5982 ) | ( n842 & n6822 ) | ( n5982 & n6822 ) ;
  assign n6824 = n6823 ^ n6233 ^ n3259 ;
  assign n6825 = ( n4907 & n6819 ) | ( n4907 & n6824 ) | ( n6819 & n6824 ) ;
  assign n6828 = ( n432 & n5570 ) | ( n432 & ~n5873 ) | ( n5570 & ~n5873 ) ;
  assign n6829 = x43 & n6828 ;
  assign n6830 = n6829 ^ n2550 ^ 1'b0 ;
  assign n6826 = n1485 ^ n1360 ^ 1'b0 ;
  assign n6827 = n1513 | n6826 ;
  assign n6831 = n6830 ^ n6827 ^ 1'b0 ;
  assign n6832 = n454 | n4534 ;
  assign n6833 = n5211 | n6832 ;
  assign n6834 = n3612 & n6833 ;
  assign n6835 = n5762 ^ n4357 ^ n2511 ;
  assign n6836 = n5290 ^ n3246 ^ 1'b0 ;
  assign n6837 = n6835 & n6836 ;
  assign n6838 = n5476 ^ n4636 ^ n1691 ;
  assign n6839 = n6838 ^ n6164 ^ n1071 ;
  assign n6840 = n5549 ^ n3711 ^ 1'b0 ;
  assign n6841 = ~n1855 & n6840 ;
  assign n6842 = n6841 ^ n554 ^ 1'b0 ;
  assign n6843 = ( ~n3108 & n3451 ) | ( ~n3108 & n5332 ) | ( n3451 & n5332 ) ;
  assign n6844 = n4506 ^ n1094 ^ 1'b0 ;
  assign n6845 = ~n1071 & n6844 ;
  assign n6846 = n1017 | n3851 ;
  assign n6847 = n6845 | n6846 ;
  assign n6848 = ~n6513 & n6847 ;
  assign n6849 = ( n1611 & n4579 ) | ( n1611 & ~n6848 ) | ( n4579 & ~n6848 ) ;
  assign n6850 = n3510 & ~n4838 ;
  assign n6851 = ~n1426 & n6850 ;
  assign n6857 = x102 & ~n1184 ;
  assign n6858 = n746 & n6857 ;
  assign n6855 = n5353 ^ n520 ^ 1'b0 ;
  assign n6856 = n194 & n6855 ;
  assign n6859 = n6858 ^ n6856 ^ n4955 ;
  assign n6860 = n3485 | n6859 ;
  assign n6852 = n1256 | n1426 ;
  assign n6853 = n1034 | n6852 ;
  assign n6854 = n4553 & n6853 ;
  assign n6861 = n6860 ^ n6854 ^ 1'b0 ;
  assign n6862 = n1104 & ~n4655 ;
  assign n6863 = n501 & ~n4832 ;
  assign n6864 = n4217 & n6863 ;
  assign n6865 = n955 & ~n6864 ;
  assign n6866 = n6865 ^ n2717 ^ 1'b0 ;
  assign n6867 = n5991 | n6866 ;
  assign n6868 = n6862 | n6867 ;
  assign n6869 = n3331 | n6868 ;
  assign n6870 = n6325 ^ n2131 ^ n739 ;
  assign n6871 = n5052 ^ n1646 ^ 1'b0 ;
  assign n6872 = n2913 & ~n5241 ;
  assign n6873 = ~n2102 & n6872 ;
  assign n6874 = n6871 | n6873 ;
  assign n6875 = n1397 & ~n6874 ;
  assign n6879 = ( ~n613 & n2561 ) | ( ~n613 & n4183 ) | ( n2561 & n4183 ) ;
  assign n6880 = n541 & ~n6879 ;
  assign n6881 = ~n2749 & n6880 ;
  assign n6876 = n2387 & ~n3154 ;
  assign n6877 = n6876 ^ n1223 ^ 1'b0 ;
  assign n6878 = ( ~n1160 & n1348 ) | ( ~n1160 & n6877 ) | ( n1348 & n6877 ) ;
  assign n6882 = n6881 ^ n6878 ^ n1558 ;
  assign n6883 = ( n1448 & ~n1972 ) | ( n1448 & n3065 ) | ( ~n1972 & n3065 ) ;
  assign n6884 = n3564 ^ n2228 ^ 1'b0 ;
  assign n6885 = n2372 ^ x94 ^ 1'b0 ;
  assign n6886 = n6884 & ~n6885 ;
  assign n6887 = n4758 & n6886 ;
  assign n6888 = n6887 ^ n2887 ^ 1'b0 ;
  assign n6891 = n2586 ^ n1628 ^ n1551 ;
  assign n6892 = ~n2296 & n6891 ;
  assign n6893 = n6892 ^ n2166 ^ 1'b0 ;
  assign n6889 = n3242 ^ n1639 ^ n1543 ;
  assign n6890 = n6889 ^ n6206 ^ n4371 ;
  assign n6894 = n6893 ^ n6890 ^ 1'b0 ;
  assign n6895 = n531 & ~n3664 ;
  assign n6896 = n6895 ^ n4137 ^ 1'b0 ;
  assign n6897 = n6896 ^ n487 ^ 1'b0 ;
  assign n6898 = n2618 & n6897 ;
  assign n6899 = n6545 & n6898 ;
  assign n6901 = n3468 ^ n2996 ^ n2378 ;
  assign n6900 = x21 & n6294 ;
  assign n6902 = n6901 ^ n6900 ^ 1'b0 ;
  assign n6903 = ( ~n1013 & n3562 ) | ( ~n1013 & n4934 ) | ( n3562 & n4934 ) ;
  assign n6904 = n4133 | n6903 ;
  assign n6905 = n3461 | n6904 ;
  assign n6906 = n5522 ^ n3524 ^ n1547 ;
  assign n6907 = n6668 ^ n3383 ^ 1'b0 ;
  assign n6908 = n1968 ^ n905 ^ n601 ;
  assign n6910 = n2737 ^ n2571 ^ 1'b0 ;
  assign n6909 = n4827 ^ n3140 ^ 1'b0 ;
  assign n6911 = n6910 ^ n6909 ^ n3194 ;
  assign n6912 = n5643 ^ n5002 ^ 1'b0 ;
  assign n6913 = n859 & n928 ;
  assign n6914 = ~n449 & n6913 ;
  assign n6915 = n2874 | n6914 ;
  assign n6916 = n6915 ^ n1306 ^ 1'b0 ;
  assign n6917 = n739 | n4987 ;
  assign n6918 = n6917 ^ n5615 ^ 1'b0 ;
  assign n6919 = n4671 & ~n6918 ;
  assign n6920 = n4774 ^ n274 ^ 1'b0 ;
  assign n6921 = n6447 & ~n6920 ;
  assign n6922 = n5676 ^ n4363 ^ n2372 ;
  assign n6923 = n5172 ^ n2835 ^ 1'b0 ;
  assign n6924 = ~n314 & n1357 ;
  assign n6925 = n821 ^ n654 ^ 1'b0 ;
  assign n6926 = n3897 | n6925 ;
  assign n6927 = ( n192 & n6811 ) | ( n192 & n6926 ) | ( n6811 & n6926 ) ;
  assign n6928 = ~n318 & n5343 ;
  assign n6929 = n6927 & n6928 ;
  assign n6930 = n5332 | n6875 ;
  assign n6931 = ~n826 & n4536 ;
  assign n6932 = ( n2921 & ~n5492 ) | ( n2921 & n6931 ) | ( ~n5492 & n6931 ) ;
  assign n6933 = x96 & ~n1184 ;
  assign n6934 = n1184 & n6933 ;
  assign n6935 = n6934 ^ n631 ^ n214 ;
  assign n6936 = n4466 ^ n2543 ^ 1'b0 ;
  assign n6937 = ( n5655 & n6935 ) | ( n5655 & ~n6936 ) | ( n6935 & ~n6936 ) ;
  assign n6938 = n238 | n2663 ;
  assign n6939 = ~n1111 & n6938 ;
  assign n6940 = n6939 ^ n4081 ^ 1'b0 ;
  assign n6941 = n1682 | n6524 ;
  assign n6942 = n6941 ^ n4257 ^ 1'b0 ;
  assign n6943 = x110 & ~n6942 ;
  assign n6944 = ~n3637 & n5993 ;
  assign n6945 = n6944 ^ n5760 ^ 1'b0 ;
  assign n6946 = ( n348 & n1397 ) | ( n348 & ~n6945 ) | ( n1397 & ~n6945 ) ;
  assign n6947 = n5702 ^ n1946 ^ 1'b0 ;
  assign n6948 = n6860 ^ n1846 ^ 1'b0 ;
  assign n6949 = n5041 | n6948 ;
  assign n6950 = n6949 ^ n1833 ^ 1'b0 ;
  assign n6951 = n3634 & ~n4030 ;
  assign n6952 = n2346 | n6951 ;
  assign n6953 = ( n605 & n848 ) | ( n605 & ~n1505 ) | ( n848 & ~n1505 ) ;
  assign n6954 = n6953 ^ n4699 ^ n349 ;
  assign n6955 = n6322 ^ n4627 ^ n1597 ;
  assign n6956 = n6598 ^ n3267 ^ n2663 ;
  assign n6957 = ( n1425 & ~n5590 ) | ( n1425 & n6956 ) | ( ~n5590 & n6956 ) ;
  assign n6960 = ( n2705 & ~n3124 ) | ( n2705 & n5672 ) | ( ~n3124 & n5672 ) ;
  assign n6958 = ( n243 & n334 ) | ( n243 & ~n3059 ) | ( n334 & ~n3059 ) ;
  assign n6959 = n6958 ^ n4261 ^ n1816 ;
  assign n6961 = n6960 ^ n6959 ^ n6216 ;
  assign n6962 = ( n1235 & n4525 ) | ( n1235 & ~n6961 ) | ( n4525 & ~n6961 ) ;
  assign n6963 = n4226 ^ n3761 ^ n1327 ;
  assign n6964 = n6963 ^ n2152 ^ 1'b0 ;
  assign n6965 = n2459 ^ n253 ^ 1'b0 ;
  assign n6966 = ( n2564 & n4699 ) | ( n2564 & n6965 ) | ( n4699 & n6965 ) ;
  assign n6967 = n2194 ^ x35 ^ 1'b0 ;
  assign n6968 = n1986 ^ n1559 ^ n230 ;
  assign n6969 = ( n2884 & n6967 ) | ( n2884 & n6968 ) | ( n6967 & n6968 ) ;
  assign n6970 = ( ~n1916 & n4821 ) | ( ~n1916 & n6969 ) | ( n4821 & n6969 ) ;
  assign n6971 = n4972 ^ n3253 ^ 1'b0 ;
  assign n6972 = n1661 | n2585 ;
  assign n6973 = n958 ^ x74 ^ 1'b0 ;
  assign n6974 = n967 | n6973 ;
  assign n6975 = ( n5454 & n6972 ) | ( n5454 & n6974 ) | ( n6972 & n6974 ) ;
  assign n6976 = ( n1913 & ~n4144 ) | ( n1913 & n6975 ) | ( ~n4144 & n6975 ) ;
  assign n6977 = ( n1134 & n1550 ) | ( n1134 & n4635 ) | ( n1550 & n4635 ) ;
  assign n6978 = ~n1634 & n2619 ;
  assign n6979 = n3772 & n6978 ;
  assign n6980 = n6332 ^ n5811 ^ 1'b0 ;
  assign n6981 = n6979 | n6980 ;
  assign n6982 = ~n3398 & n5582 ;
  assign n6983 = ~n3409 & n5287 ;
  assign n6984 = n6983 ^ n2296 ^ 1'b0 ;
  assign n6985 = ( n6981 & n6982 ) | ( n6981 & ~n6984 ) | ( n6982 & ~n6984 ) ;
  assign n6986 = n5013 ^ n3207 ^ n2879 ;
  assign n6987 = x93 & ~n6129 ;
  assign n6988 = n2701 ^ n2454 ^ n851 ;
  assign n6989 = n6988 ^ n5181 ^ n2490 ;
  assign n6990 = n5787 ^ n2285 ^ 1'b0 ;
  assign n6991 = ( n4000 & ~n6989 ) | ( n4000 & n6990 ) | ( ~n6989 & n6990 ) ;
  assign n6993 = n4089 ^ n2401 ^ n2239 ;
  assign n6992 = n1837 & ~n2065 ;
  assign n6994 = n6993 ^ n6992 ^ 1'b0 ;
  assign n6995 = n6994 ^ n3304 ^ n1466 ;
  assign n6996 = n1599 & ~n6995 ;
  assign n6997 = n6996 ^ n1206 ^ 1'b0 ;
  assign n7004 = n4747 & ~n5468 ;
  assign n7005 = n7004 ^ n3378 ^ 1'b0 ;
  assign n7006 = ( n586 & ~n1223 ) | ( n586 & n7005 ) | ( ~n1223 & n7005 ) ;
  assign n6998 = n141 & n4290 ;
  assign n6999 = n6998 ^ n619 ^ 1'b0 ;
  assign n7000 = n6999 ^ n973 ^ 1'b0 ;
  assign n7001 = n5206 ^ n1819 ^ 1'b0 ;
  assign n7002 = n4864 & ~n7001 ;
  assign n7003 = ( n1942 & n7000 ) | ( n1942 & ~n7002 ) | ( n7000 & ~n7002 ) ;
  assign n7007 = n7006 ^ n7003 ^ n2706 ;
  assign n7008 = n7007 ^ n6635 ^ n519 ;
  assign n7009 = n4354 ^ n3513 ^ n1830 ;
  assign n7010 = n5229 ^ n2401 ^ 1'b0 ;
  assign n7011 = n6030 & n7010 ;
  assign n7012 = n4733 ^ n1952 ^ 1'b0 ;
  assign n7013 = n1422 ^ n1420 ^ 1'b0 ;
  assign n7014 = n1196 & ~n7013 ;
  assign n7015 = ( ~n2955 & n3990 ) | ( ~n2955 & n7014 ) | ( n3990 & n7014 ) ;
  assign n7016 = ~n3670 & n7015 ;
  assign n7017 = n1072 & ~n2522 ;
  assign n7018 = n7017 ^ n3606 ^ 1'b0 ;
  assign n7019 = ( ~n3252 & n5753 ) | ( ~n3252 & n7018 ) | ( n5753 & n7018 ) ;
  assign n7020 = n7016 & ~n7019 ;
  assign n7021 = n7012 & n7020 ;
  assign n7022 = ( n1820 & ~n2025 ) | ( n1820 & n3648 ) | ( ~n2025 & n3648 ) ;
  assign n7023 = ~n1302 & n4331 ;
  assign n7024 = n3091 & n7023 ;
  assign n7025 = n7024 ^ n1739 ^ n822 ;
  assign n7026 = ( n2322 & n5048 ) | ( n2322 & ~n7025 ) | ( n5048 & ~n7025 ) ;
  assign n7027 = n7026 ^ n6171 ^ 1'b0 ;
  assign n7028 = ~n7022 & n7027 ;
  assign n7029 = ~n1036 & n7028 ;
  assign n7030 = ~n5405 & n7029 ;
  assign n7031 = n164 & ~n7030 ;
  assign n7032 = n3312 ^ n2254 ^ 1'b0 ;
  assign n7033 = n5948 ^ n2994 ^ 1'b0 ;
  assign n7034 = ( n5270 & ~n7032 ) | ( n5270 & n7033 ) | ( ~n7032 & n7033 ) ;
  assign n7035 = n7034 ^ n4489 ^ 1'b0 ;
  assign n7036 = n2537 & n2542 ;
  assign n7037 = n6439 ^ n2116 ^ 1'b0 ;
  assign n7038 = n2223 & ~n7037 ;
  assign n7039 = n460 | n2450 ;
  assign n7040 = ( n2703 & n3524 ) | ( n2703 & n7039 ) | ( n3524 & n7039 ) ;
  assign n7041 = ( ~n293 & n5468 ) | ( ~n293 & n7040 ) | ( n5468 & n7040 ) ;
  assign n7042 = n2121 | n2246 ;
  assign n7043 = ~n5387 & n7042 ;
  assign n7044 = n7043 ^ n4525 ^ 1'b0 ;
  assign n7045 = n3582 ^ n2707 ^ n774 ;
  assign n7046 = n2859 | n3482 ;
  assign n7047 = n1065 | n7046 ;
  assign n7048 = ( n227 & n3028 ) | ( n227 & ~n7047 ) | ( n3028 & ~n7047 ) ;
  assign n7049 = n4976 ^ n4857 ^ n3390 ;
  assign n7050 = n7049 ^ n4109 ^ n3654 ;
  assign n7051 = ( n6761 & ~n7048 ) | ( n6761 & n7050 ) | ( ~n7048 & n7050 ) ;
  assign n7052 = n3719 ^ n1022 ^ 1'b0 ;
  assign n7053 = n831 ^ n800 ^ 1'b0 ;
  assign n7054 = ~n7052 & n7053 ;
  assign n7055 = n3262 ^ n817 ^ 1'b0 ;
  assign n7056 = n7054 & ~n7055 ;
  assign n7057 = ( n3696 & ~n3968 ) | ( n3696 & n5051 ) | ( ~n3968 & n5051 ) ;
  assign n7059 = n862 & ~n1915 ;
  assign n7060 = n7059 ^ x107 ^ 1'b0 ;
  assign n7058 = n2634 & n5218 ;
  assign n7061 = n7060 ^ n7058 ^ 1'b0 ;
  assign n7063 = n5980 ^ n1270 ^ 1'b0 ;
  assign n7064 = n421 & n7063 ;
  assign n7062 = x4 & n5234 ;
  assign n7065 = n7064 ^ n7062 ^ 1'b0 ;
  assign n7066 = ~n2778 & n7065 ;
  assign n7071 = ~n901 & n1877 ;
  assign n7068 = ( n1575 & n2222 ) | ( n1575 & n2818 ) | ( n2222 & n2818 ) ;
  assign n7069 = n7068 ^ n4199 ^ 1'b0 ;
  assign n7070 = n1653 & ~n7069 ;
  assign n7067 = n3688 ^ n3580 ^ 1'b0 ;
  assign n7072 = n7071 ^ n7070 ^ n7067 ;
  assign n7074 = n3515 ^ n2198 ^ 1'b0 ;
  assign n7073 = ~n2974 & n5341 ;
  assign n7075 = n7074 ^ n7073 ^ 1'b0 ;
  assign n7076 = n5935 ^ n5000 ^ 1'b0 ;
  assign n7077 = n321 & ~n7076 ;
  assign n7078 = n7077 ^ n1199 ^ 1'b0 ;
  assign n7079 = n3049 & ~n7078 ;
  assign n7082 = n4092 ^ n2424 ^ n693 ;
  assign n7080 = n1025 & ~n5364 ;
  assign n7081 = x32 & n7080 ;
  assign n7083 = n7082 ^ n7081 ^ n2842 ;
  assign n7085 = x60 & n3581 ;
  assign n7084 = x94 & ~n1928 ;
  assign n7086 = n7085 ^ n7084 ^ 1'b0 ;
  assign n7087 = ~n2862 & n6330 ;
  assign n7088 = n7087 ^ n885 ^ 1'b0 ;
  assign n7089 = n4775 ^ n2605 ^ 1'b0 ;
  assign n7090 = n7089 ^ n364 ^ x105 ;
  assign n7091 = n5762 ^ n5760 ^ 1'b0 ;
  assign n7092 = n2802 | n3476 ;
  assign n7093 = ( n4239 & n5086 ) | ( n4239 & n7092 ) | ( n5086 & n7092 ) ;
  assign n7094 = n6224 ^ n3610 ^ 1'b0 ;
  assign n7095 = n7094 ^ n771 ^ 1'b0 ;
  assign n7096 = n5120 | n7015 ;
  assign n7097 = n470 & ~n569 ;
  assign n7098 = ~n4377 & n7097 ;
  assign n7099 = n7098 ^ n1761 ^ n826 ;
  assign n7101 = n842 & n1420 ;
  assign n7102 = n7101 ^ n1754 ^ 1'b0 ;
  assign n7103 = n7102 ^ n2458 ^ n2114 ;
  assign n7100 = ( n888 & n2692 ) | ( n888 & n4984 ) | ( n2692 & n4984 ) ;
  assign n7104 = n7103 ^ n7100 ^ n4960 ;
  assign n7106 = n2491 & ~n3598 ;
  assign n7107 = n3558 & n7106 ;
  assign n7105 = n4910 ^ n1570 ^ n272 ;
  assign n7108 = n7107 ^ n7105 ^ 1'b0 ;
  assign n7109 = n7108 ^ n2417 ^ 1'b0 ;
  assign n7110 = n141 & n3312 ;
  assign n7113 = n6586 ^ n1389 ^ n1027 ;
  assign n7114 = n302 & ~n7113 ;
  assign n7115 = ~n771 & n7114 ;
  assign n7111 = n374 & ~n3476 ;
  assign n7112 = n7111 ^ n3832 ^ 1'b0 ;
  assign n7116 = n7115 ^ n7112 ^ n3971 ;
  assign n7117 = n7110 | n7116 ;
  assign n7118 = x93 | n548 ;
  assign n7121 = n6517 ^ n6218 ^ n549 ;
  assign n7119 = ~n2824 & n2978 ;
  assign n7120 = n3964 & ~n7119 ;
  assign n7122 = n7121 ^ n7120 ^ 1'b0 ;
  assign n7123 = n7122 ^ n4719 ^ n4236 ;
  assign n7124 = n6945 ^ n4094 ^ 1'b0 ;
  assign n7125 = n4290 | n5052 ;
  assign n7126 = n292 & n1590 ;
  assign n7127 = n7126 ^ n173 ^ 1'b0 ;
  assign n7128 = n7127 ^ n6786 ^ n137 ;
  assign n7129 = n3482 ^ n2211 ^ 1'b0 ;
  assign n7130 = n7129 ^ n6196 ^ 1'b0 ;
  assign n7131 = ~n562 & n1488 ;
  assign n7132 = ~n5218 & n7131 ;
  assign n7133 = n1468 & ~n2914 ;
  assign n7134 = n7133 ^ n3874 ^ 1'b0 ;
  assign n7135 = n7132 & ~n7134 ;
  assign n7137 = n2172 ^ n601 ^ 1'b0 ;
  assign n7138 = n2749 & ~n7137 ;
  assign n7136 = n3628 ^ n859 ^ n141 ;
  assign n7139 = n7138 ^ n7136 ^ 1'b0 ;
  assign n7140 = n1176 & ~n7139 ;
  assign n7148 = n2101 ^ n222 ^ 1'b0 ;
  assign n7147 = n1176 & n2251 ;
  assign n7149 = n7148 ^ n7147 ^ 1'b0 ;
  assign n7144 = n3162 ^ n2465 ^ 1'b0 ;
  assign n7145 = n3367 & n7144 ;
  assign n7141 = x15 & x88 ;
  assign n7142 = n299 & n7141 ;
  assign n7143 = n3239 & n7142 ;
  assign n7146 = n7145 ^ n7143 ^ n2077 ;
  assign n7150 = n7149 ^ n7146 ^ n6193 ;
  assign n7151 = n4727 & ~n5012 ;
  assign n7152 = n7151 ^ n4567 ^ 1'b0 ;
  assign n7153 = n6146 & ~n7152 ;
  assign n7154 = ( x73 & ~x98 ) | ( x73 & n7153 ) | ( ~x98 & n7153 ) ;
  assign n7157 = n1781 & ~n5495 ;
  assign n7155 = n540 & ~n2614 ;
  assign n7156 = ( n2387 & n5822 ) | ( n2387 & n7155 ) | ( n5822 & n7155 ) ;
  assign n7158 = n7157 ^ n7156 ^ n1754 ;
  assign n7160 = ~n4544 & n6010 ;
  assign n7161 = ~n2281 & n7160 ;
  assign n7162 = n7161 ^ n3033 ^ 1'b0 ;
  assign n7159 = n6317 ^ n5296 ^ 1'b0 ;
  assign n7163 = n7162 ^ n7159 ^ n3624 ;
  assign n7164 = n477 & ~n5759 ;
  assign n7165 = n7164 ^ n2199 ^ 1'b0 ;
  assign n7166 = n2324 & n4443 ;
  assign n7167 = n7166 ^ n4907 ^ 1'b0 ;
  assign n7168 = ( ~n1406 & n5396 ) | ( ~n1406 & n7068 ) | ( n5396 & n7068 ) ;
  assign n7169 = ( x102 & n721 ) | ( x102 & n1689 ) | ( n721 & n1689 ) ;
  assign n7174 = n1488 ^ n850 ^ x115 ;
  assign n7173 = n250 | n347 ;
  assign n7175 = n7174 ^ n7173 ^ 1'b0 ;
  assign n7176 = ( n4390 & ~n5736 ) | ( n4390 & n7175 ) | ( ~n5736 & n7175 ) ;
  assign n7170 = ~n497 & n2998 ;
  assign n7171 = ~n691 & n7170 ;
  assign n7172 = n7171 ^ n5318 ^ 1'b0 ;
  assign n7177 = n7176 ^ n7172 ^ n4907 ;
  assign n7178 = ( ~n505 & n4747 ) | ( ~n505 & n6281 ) | ( n4747 & n6281 ) ;
  assign n7179 = ~n381 & n771 ;
  assign n7180 = ~n285 & n7179 ;
  assign n7181 = n3438 & ~n7180 ;
  assign n7182 = ~n3926 & n7181 ;
  assign n7183 = n6802 ^ n810 ^ x59 ;
  assign n7184 = ~n1862 & n3666 ;
  assign n7185 = n7183 & n7184 ;
  assign n7187 = n3291 & ~n4182 ;
  assign n7188 = n7187 ^ n2381 ^ 1'b0 ;
  assign n7189 = n7188 ^ n5054 ^ n4939 ;
  assign n7186 = n3735 ^ n3546 ^ n1699 ;
  assign n7190 = n7189 ^ n7186 ^ 1'b0 ;
  assign n7191 = n7190 ^ n4152 ^ 1'b0 ;
  assign n7192 = ( n1836 & n3609 ) | ( n1836 & ~n4871 ) | ( n3609 & ~n4871 ) ;
  assign n7193 = ~n1172 & n4717 ;
  assign n7194 = n2958 & ~n7193 ;
  assign n7195 = n7194 ^ n5340 ^ 1'b0 ;
  assign n7196 = n3200 & n7195 ;
  assign n7197 = n7192 & n7196 ;
  assign n7199 = n1673 & n4949 ;
  assign n7200 = n7199 ^ n4859 ^ n4407 ;
  assign n7198 = ~n2315 & n6393 ;
  assign n7201 = n7200 ^ n7198 ^ n2929 ;
  assign n7202 = ~n4550 & n7176 ;
  assign n7203 = n2017 & n7202 ;
  assign n7204 = n3483 ^ n3378 ^ 1'b0 ;
  assign n7205 = n7204 ^ n4740 ^ 1'b0 ;
  assign n7206 = ( n5243 & n7203 ) | ( n5243 & ~n7205 ) | ( n7203 & ~n7205 ) ;
  assign n7207 = ~n1131 & n1830 ;
  assign n7208 = ( n2389 & n5522 ) | ( n2389 & ~n7207 ) | ( n5522 & ~n7207 ) ;
  assign n7209 = ( n3363 & ~n5956 ) | ( n3363 & n7208 ) | ( ~n5956 & n7208 ) ;
  assign n7210 = ~n6192 & n7209 ;
  assign n7211 = n7210 ^ n1764 ^ 1'b0 ;
  assign n7212 = n739 & ~n1687 ;
  assign n7213 = n7212 ^ n5084 ^ 1'b0 ;
  assign n7214 = n7213 ^ n7028 ^ n3961 ;
  assign n7215 = ( x88 & n953 ) | ( x88 & n6364 ) | ( n953 & n6364 ) ;
  assign n7216 = ( n5949 & n6347 ) | ( n5949 & n6432 ) | ( n6347 & n6432 ) ;
  assign n7218 = ( n1206 & n2124 ) | ( n1206 & n3260 ) | ( n2124 & n3260 ) ;
  assign n7217 = n595 & n1229 ;
  assign n7219 = n7218 ^ n7217 ^ 1'b0 ;
  assign n7220 = n7219 ^ n2129 ^ 1'b0 ;
  assign n7221 = ( ~x45 & n270 ) | ( ~x45 & n7220 ) | ( n270 & n7220 ) ;
  assign n7222 = n5588 ^ n2434 ^ 1'b0 ;
  assign n7223 = ~n5176 & n7222 ;
  assign n7224 = n6793 ^ n6374 ^ 1'b0 ;
  assign n7225 = n7224 ^ n4635 ^ n379 ;
  assign n7226 = n7225 ^ n5982 ^ n2160 ;
  assign n7227 = n3325 ^ n1625 ^ 1'b0 ;
  assign n7228 = n7227 ^ n3532 ^ n1914 ;
  assign n7229 = ( n3723 & n6040 ) | ( n3723 & n7228 ) | ( n6040 & n7228 ) ;
  assign n7230 = n2745 ^ n2542 ^ 1'b0 ;
  assign n7231 = n1977 ^ n1468 ^ 1'b0 ;
  assign n7232 = n7230 & n7231 ;
  assign n7233 = ( n6086 & n6723 ) | ( n6086 & n7232 ) | ( n6723 & n7232 ) ;
  assign n7235 = x111 & ~n3640 ;
  assign n7236 = n4828 & n7235 ;
  assign n7234 = n6529 ^ n5021 ^ 1'b0 ;
  assign n7237 = n7236 ^ n7234 ^ n1229 ;
  assign n7238 = n7237 ^ n4554 ^ n2199 ;
  assign n7239 = n1860 ^ n1407 ^ n1357 ;
  assign n7240 = n7239 ^ n2319 ^ n921 ;
  assign n7241 = ( n574 & ~n987 ) | ( n574 & n2328 ) | ( ~n987 & n2328 ) ;
  assign n7242 = n7241 ^ n1621 ^ n232 ;
  assign n7243 = ~n2140 & n4010 ;
  assign n7244 = ( n283 & n3274 ) | ( n283 & ~n7243 ) | ( n3274 & ~n7243 ) ;
  assign n7245 = n7244 ^ x98 ^ 1'b0 ;
  assign n7246 = n7242 & n7245 ;
  assign n7247 = ( n835 & ~n1080 ) | ( n835 & n4307 ) | ( ~n1080 & n4307 ) ;
  assign n7248 = n5632 ^ n2322 ^ 1'b0 ;
  assign n7249 = ~n5917 & n7248 ;
  assign n7250 = n1383 & n2919 ;
  assign n7251 = n7250 ^ n6910 ^ 1'b0 ;
  assign n7252 = ~n4613 & n7251 ;
  assign n7253 = ~n4538 & n7252 ;
  assign n7254 = n1862 & n7253 ;
  assign n7255 = n802 | n3207 ;
  assign n7256 = n7255 ^ n3257 ^ 1'b0 ;
  assign n7257 = n7256 ^ n6893 ^ x94 ;
  assign n7258 = x126 & ~n1107 ;
  assign n7259 = ~x74 & n7258 ;
  assign n7260 = n7242 & ~n7259 ;
  assign n7261 = n620 & n7260 ;
  assign n7262 = n7261 ^ n4781 ^ n1369 ;
  assign n7263 = n7262 ^ n5584 ^ 1'b0 ;
  assign n7264 = n576 | n2114 ;
  assign n7265 = n211 & ~n7264 ;
  assign n7266 = n1448 & ~n6703 ;
  assign n7267 = ( n1046 & ~n2373 ) | ( n1046 & n2834 ) | ( ~n2373 & n2834 ) ;
  assign n7268 = n7267 ^ n5940 ^ n4181 ;
  assign n7269 = ( ~n4316 & n5387 ) | ( ~n4316 & n6328 ) | ( n5387 & n6328 ) ;
  assign n7270 = n5629 ^ n2145 ^ n477 ;
  assign n7271 = ( n5944 & ~n6780 ) | ( n5944 & n7270 ) | ( ~n6780 & n7270 ) ;
  assign n7272 = n1221 & ~n5160 ;
  assign n7273 = n7271 & n7272 ;
  assign n7274 = n2965 | n5339 ;
  assign n7275 = n7274 ^ n2815 ^ 1'b0 ;
  assign n7276 = ~n2086 & n2101 ;
  assign n7277 = n7275 & n7276 ;
  assign n7278 = n4101 ^ n2275 ^ n348 ;
  assign n7279 = n2796 & ~n7278 ;
  assign n7280 = n7241 ^ n7214 ^ 1'b0 ;
  assign n7281 = n6651 ^ n1282 ^ 1'b0 ;
  assign n7282 = n4925 & ~n7281 ;
  assign n7283 = n1384 | n1493 ;
  assign n7284 = n7283 ^ n1088 ^ 1'b0 ;
  assign n7285 = ( n2285 & ~n4815 ) | ( n2285 & n6151 ) | ( ~n4815 & n6151 ) ;
  assign n7286 = ( n6755 & ~n7284 ) | ( n6755 & n7285 ) | ( ~n7284 & n7285 ) ;
  assign n7287 = n4701 | n6412 ;
  assign n7288 = n2422 | n6448 ;
  assign n7289 = n1275 | n7288 ;
  assign n7290 = ~n623 & n1178 ;
  assign n7291 = ~n5110 & n7290 ;
  assign n7293 = ( n1556 & n2227 ) | ( n1556 & ~n3027 ) | ( n2227 & ~n3027 ) ;
  assign n7292 = ( n1294 & n2739 ) | ( n1294 & n3062 ) | ( n2739 & n3062 ) ;
  assign n7294 = n7293 ^ n7292 ^ n5719 ;
  assign n7298 = n607 & ~n4602 ;
  assign n7299 = n243 & n7298 ;
  assign n7295 = n1103 & n3763 ;
  assign n7296 = n7295 ^ n3473 ^ 1'b0 ;
  assign n7297 = n7125 & ~n7296 ;
  assign n7300 = n7299 ^ n7297 ^ 1'b0 ;
  assign n7301 = n2222 & ~n7300 ;
  assign n7302 = x59 & ~n1613 ;
  assign n7303 = ~n3087 & n7302 ;
  assign n7304 = ( n4792 & ~n5302 ) | ( n4792 & n7303 ) | ( ~n5302 & n7303 ) ;
  assign n7305 = n7304 ^ n5332 ^ 1'b0 ;
  assign n7306 = ( ~n1794 & n7052 ) | ( ~n1794 & n7237 ) | ( n7052 & n7237 ) ;
  assign n7307 = ( x49 & n7305 ) | ( x49 & n7306 ) | ( n7305 & n7306 ) ;
  assign n7308 = n1791 ^ n1715 ^ n1019 ;
  assign n7309 = n7308 ^ n6273 ^ n6180 ;
  assign n7314 = n4179 ^ n3355 ^ 1'b0 ;
  assign n7312 = n985 & ~n1877 ;
  assign n7313 = ~n170 & n7312 ;
  assign n7310 = n3711 & ~n4046 ;
  assign n7311 = n7310 ^ n4837 ^ 1'b0 ;
  assign n7315 = n7314 ^ n7313 ^ n7311 ;
  assign n7316 = x117 & n525 ;
  assign n7317 = n7316 ^ n1434 ^ 1'b0 ;
  assign n7318 = n7317 ^ n3563 ^ n2289 ;
  assign n7319 = n7318 ^ n3332 ^ n691 ;
  assign n7320 = n4231 & ~n7319 ;
  assign n7321 = n171 & n1065 ;
  assign n7322 = ~n1492 & n7321 ;
  assign n7323 = ( x77 & ~n3303 ) | ( x77 & n7299 ) | ( ~n3303 & n7299 ) ;
  assign n7324 = n7323 ^ n2043 ^ n1534 ;
  assign n7325 = n7324 ^ n4013 ^ n3389 ;
  assign n7326 = ( n670 & ~n7322 ) | ( n670 & n7325 ) | ( ~n7322 & n7325 ) ;
  assign n7327 = ( n6310 & ~n6438 ) | ( n6310 & n7326 ) | ( ~n6438 & n7326 ) ;
  assign n7328 = n1077 | n4256 ;
  assign n7330 = n5302 ^ n575 ^ n304 ;
  assign n7329 = n1711 & n6388 ;
  assign n7331 = n7330 ^ n7329 ^ 1'b0 ;
  assign n7332 = ~n2029 & n3299 ;
  assign n7333 = n6959 & n7332 ;
  assign n7334 = n4013 & n5341 ;
  assign n7335 = n7334 ^ n5127 ^ n134 ;
  assign n7336 = n2900 ^ n295 ^ 1'b0 ;
  assign n7337 = n571 & ~n7336 ;
  assign n7338 = ( ~n3744 & n7335 ) | ( ~n3744 & n7337 ) | ( n7335 & n7337 ) ;
  assign n7339 = n5936 ^ n3573 ^ n2472 ;
  assign n7340 = n3453 ^ x59 ^ 1'b0 ;
  assign n7341 = n3905 & ~n7340 ;
  assign n7342 = n7341 ^ n1146 ^ 1'b0 ;
  assign n7343 = ( ~n4396 & n7339 ) | ( ~n4396 & n7342 ) | ( n7339 & n7342 ) ;
  assign n7344 = n3840 ^ n3704 ^ 1'b0 ;
  assign n7345 = ~n667 & n3616 ;
  assign n7346 = n7345 ^ n4192 ^ 1'b0 ;
  assign n7347 = x48 & n7346 ;
  assign n7348 = ( n2274 & n7344 ) | ( n2274 & n7347 ) | ( n7344 & n7347 ) ;
  assign n7349 = n3436 ^ n2715 ^ n1774 ;
  assign n7350 = n3563 | n7349 ;
  assign n7351 = n7350 ^ n1798 ^ 1'b0 ;
  assign n7352 = n2042 ^ n1346 ^ 1'b0 ;
  assign n7353 = n4541 | n7352 ;
  assign n7354 = n7353 ^ n4488 ^ n1818 ;
  assign n7355 = n2336 ^ n1185 ^ 1'b0 ;
  assign n7356 = ~n2404 & n5549 ;
  assign n7357 = n2515 & n7356 ;
  assign n7358 = n7357 ^ x79 ^ 1'b0 ;
  assign n7359 = n1927 & n4936 ;
  assign n7360 = ~n787 & n7359 ;
  assign n7361 = ( n7355 & n7358 ) | ( n7355 & ~n7360 ) | ( n7358 & ~n7360 ) ;
  assign n7362 = ( n884 & ~n1329 ) | ( n884 & n5131 ) | ( ~n1329 & n5131 ) ;
  assign n7363 = n2375 & ~n2730 ;
  assign n7364 = n7363 ^ n4036 ^ 1'b0 ;
  assign n7365 = n1872 ^ n1057 ^ n550 ;
  assign n7366 = ( n2787 & ~n6402 ) | ( n2787 & n7365 ) | ( ~n6402 & n7365 ) ;
  assign n7367 = n5608 | n7366 ;
  assign n7368 = n6769 ^ n6701 ^ n6534 ;
  assign n7370 = ( n1598 & n1897 ) | ( n1598 & n7228 ) | ( n1897 & n7228 ) ;
  assign n7369 = ( n3952 & n5062 ) | ( n3952 & n6151 ) | ( n5062 & n6151 ) ;
  assign n7371 = n7370 ^ n7369 ^ 1'b0 ;
  assign n7372 = ~n7368 & n7371 ;
  assign n7373 = ( n1057 & n1789 ) | ( n1057 & n2320 ) | ( n1789 & n2320 ) ;
  assign n7374 = ( n2878 & ~n3974 ) | ( n2878 & n7373 ) | ( ~n3974 & n7373 ) ;
  assign n7375 = ( n2906 & n3913 ) | ( n2906 & n5742 ) | ( n3913 & n5742 ) ;
  assign n7376 = ( n4635 & n5572 ) | ( n4635 & ~n7375 ) | ( n5572 & ~n7375 ) ;
  assign n7377 = n7374 & ~n7376 ;
  assign n7378 = ~n3449 & n3547 ;
  assign n7380 = ( ~n1022 & n1598 ) | ( ~n1022 & n6384 ) | ( n1598 & n6384 ) ;
  assign n7379 = n1530 & ~n5071 ;
  assign n7381 = n7380 ^ n7379 ^ n6412 ;
  assign n7382 = ~n7378 & n7381 ;
  assign n7383 = n3045 | n5036 ;
  assign n7384 = n1083 & n1095 ;
  assign n7385 = n394 & n5727 ;
  assign n7386 = n7385 ^ n6986 ^ 1'b0 ;
  assign n7387 = n1774 | n7386 ;
  assign n7388 = n4042 & n5381 ;
  assign n7389 = ~n2673 & n3692 ;
  assign n7390 = n7389 ^ n390 ^ 1'b0 ;
  assign n7391 = ~n7388 & n7390 ;
  assign n7392 = n7391 ^ n3238 ^ 1'b0 ;
  assign n7393 = n7230 ^ n1493 ^ 1'b0 ;
  assign n7394 = n7392 | n7393 ;
  assign n7395 = n1724 & ~n2819 ;
  assign n7396 = n7395 ^ n3484 ^ n3315 ;
  assign n7397 = n3416 ^ n1980 ^ n1146 ;
  assign n7398 = n3221 & n7397 ;
  assign n7399 = n2776 & ~n7398 ;
  assign n7401 = n3124 | n6524 ;
  assign n7402 = ( n5507 & ~n6759 ) | ( n5507 & n7401 ) | ( ~n6759 & n7401 ) ;
  assign n7400 = n1276 & ~n5692 ;
  assign n7403 = n7402 ^ n7400 ^ n1993 ;
  assign n7404 = n3718 ^ n3158 ^ 1'b0 ;
  assign n7405 = n5455 ^ n2059 ^ 1'b0 ;
  assign n7406 = n1018 | n7405 ;
  assign n7407 = ( ~n4582 & n4800 ) | ( ~n4582 & n7406 ) | ( n4800 & n7406 ) ;
  assign n7408 = n3420 & n4176 ;
  assign n7409 = n7407 & n7408 ;
  assign n7410 = n7409 ^ n2746 ^ 1'b0 ;
  assign n7411 = n7410 ^ n2985 ^ 1'b0 ;
  assign n7412 = n4443 ^ n2692 ^ 1'b0 ;
  assign n7418 = n5616 ^ n791 ^ 1'b0 ;
  assign n7419 = ( n4096 & ~n6210 ) | ( n4096 & n7418 ) | ( ~n6210 & n7418 ) ;
  assign n7420 = n4440 ^ n241 ^ 1'b0 ;
  assign n7421 = ~n7419 & n7420 ;
  assign n7413 = n3025 & n6151 ;
  assign n7414 = n7251 ^ n1000 ^ 1'b0 ;
  assign n7415 = n7413 | n7414 ;
  assign n7416 = n7415 ^ n2863 ^ 1'b0 ;
  assign n7417 = ~n7026 & n7416 ;
  assign n7422 = n7421 ^ n7417 ^ n3701 ;
  assign n7423 = ( ~n4208 & n7412 ) | ( ~n4208 & n7422 ) | ( n7412 & n7422 ) ;
  assign n7424 = ( n7404 & ~n7411 ) | ( n7404 & n7423 ) | ( ~n7411 & n7423 ) ;
  assign n7425 = ( n872 & ~n2036 ) | ( n872 & n3750 ) | ( ~n2036 & n3750 ) ;
  assign n7426 = ( n691 & n2285 ) | ( n691 & ~n4897 ) | ( n2285 & ~n4897 ) ;
  assign n7427 = n3579 & n7426 ;
  assign n7428 = n6714 & ~n7427 ;
  assign n7429 = n7425 & n7428 ;
  assign n7430 = ~n3666 & n4902 ;
  assign n7433 = n1984 ^ n379 ^ 1'b0 ;
  assign n7431 = n2657 ^ n2174 ^ 1'b0 ;
  assign n7432 = ~n649 & n7431 ;
  assign n7434 = n7433 ^ n7432 ^ 1'b0 ;
  assign n7435 = ~n7430 & n7434 ;
  assign n7436 = ~n2903 & n7435 ;
  assign n7437 = ~n1290 & n2541 ;
  assign n7438 = n298 & n477 ;
  assign n7439 = ~n298 & n7438 ;
  assign n7440 = n7439 ^ n5154 ^ 1'b0 ;
  assign n7451 = n260 & n1507 ;
  assign n7449 = n7042 ^ n3732 ^ 1'b0 ;
  assign n7441 = n227 & ~n2254 ;
  assign n7442 = n7441 ^ n3130 ^ n1326 ;
  assign n7445 = ~n344 & n2760 ;
  assign n7446 = n7445 ^ n808 ^ 1'b0 ;
  assign n7443 = ~n1608 & n4290 ;
  assign n7444 = ~n1074 & n7443 ;
  assign n7447 = n7446 ^ n7444 ^ 1'b0 ;
  assign n7448 = n7442 | n7447 ;
  assign n7450 = n7449 ^ n7448 ^ 1'b0 ;
  assign n7452 = n7451 ^ n7450 ^ 1'b0 ;
  assign n7453 = ~n7440 & n7452 ;
  assign n7454 = n6304 ^ n3010 ^ 1'b0 ;
  assign n7455 = ~n4421 & n7454 ;
  assign n7456 = ( n855 & n6699 ) | ( n855 & n7455 ) | ( n6699 & n7455 ) ;
  assign n7457 = ~x37 & n1310 ;
  assign n7458 = n7456 & n7457 ;
  assign n7459 = ~n1745 & n3691 ;
  assign n7460 = n1976 & ~n2401 ;
  assign n7461 = ( n1176 & n7459 ) | ( n1176 & ~n7460 ) | ( n7459 & ~n7460 ) ;
  assign n7462 = n6125 ^ x126 ^ 1'b0 ;
  assign n7463 = n3784 ^ x10 ^ 1'b0 ;
  assign n7464 = n7462 & n7463 ;
  assign n7465 = n2619 ^ n1851 ^ 1'b0 ;
  assign n7466 = n7465 ^ n6111 ^ n3130 ;
  assign n7467 = n1605 & n7466 ;
  assign n7468 = n3020 ^ n174 ^ 1'b0 ;
  assign n7469 = ( n202 & n1413 ) | ( n202 & n4085 ) | ( n1413 & n4085 ) ;
  assign n7470 = ~n1053 & n7469 ;
  assign n7471 = ~x58 & n4356 ;
  assign n7472 = n4772 ^ n1314 ^ x23 ;
  assign n7473 = n7355 ^ n5443 ^ n144 ;
  assign n7474 = n7472 | n7473 ;
  assign n7475 = n7474 ^ n2834 ^ 1'b0 ;
  assign n7476 = n6040 ^ n2292 ^ n1176 ;
  assign n7477 = n915 ^ n878 ^ 1'b0 ;
  assign n7478 = n7477 ^ n897 ^ 1'b0 ;
  assign n7480 = n174 & n2251 ;
  assign n7481 = n7480 ^ n539 ^ 1'b0 ;
  assign n7482 = n2251 ^ n483 ^ n232 ;
  assign n7483 = ( n2927 & n7481 ) | ( n2927 & n7482 ) | ( n7481 & n7482 ) ;
  assign n7484 = ( n1028 & n2553 ) | ( n1028 & n4966 ) | ( n2553 & n4966 ) ;
  assign n7485 = n1078 & ~n7484 ;
  assign n7486 = n7485 ^ n3005 ^ 1'b0 ;
  assign n7487 = ~n2918 & n7486 ;
  assign n7488 = ( n3502 & ~n7483 ) | ( n3502 & n7487 ) | ( ~n7483 & n7487 ) ;
  assign n7479 = n4728 | n6751 ;
  assign n7489 = n7488 ^ n7479 ^ 1'b0 ;
  assign n7490 = n7489 ^ n4973 ^ 1'b0 ;
  assign n7491 = ~n2079 & n2272 ;
  assign n7492 = n7491 ^ n3691 ^ n1861 ;
  assign n7493 = ~n613 & n7492 ;
  assign n7494 = n7493 ^ n3324 ^ 1'b0 ;
  assign n7495 = n7494 ^ n838 ^ 1'b0 ;
  assign n7496 = n1702 & n7495 ;
  assign n7497 = n4574 | n7496 ;
  assign n7498 = n5386 ^ n5068 ^ n2758 ;
  assign n7503 = n5858 ^ n2860 ^ 1'b0 ;
  assign n7499 = n2179 ^ n1013 ^ n171 ;
  assign n7500 = ~n250 & n7499 ;
  assign n7501 = n5894 & n7500 ;
  assign n7502 = n5621 | n7501 ;
  assign n7504 = n7503 ^ n7502 ^ 1'b0 ;
  assign n7505 = n7504 ^ n4033 ^ 1'b0 ;
  assign n7506 = ~n6971 & n7505 ;
  assign n7507 = ~n612 & n2468 ;
  assign n7508 = ( n2324 & n2908 ) | ( n2324 & n7507 ) | ( n2908 & n7507 ) ;
  assign n7509 = n605 & n2503 ;
  assign n7510 = ( x43 & n541 ) | ( x43 & n3774 ) | ( n541 & n3774 ) ;
  assign n7511 = ~n7509 & n7510 ;
  assign n7512 = n2425 & n7511 ;
  assign n7513 = n5924 & ~n7512 ;
  assign n7514 = n7513 ^ n5672 ^ 1'b0 ;
  assign n7515 = ~n7508 & n7514 ;
  assign n7516 = n7481 ^ n4234 ^ n1333 ;
  assign n7517 = ~n921 & n2760 ;
  assign n7518 = n4689 & n7517 ;
  assign n7519 = n2606 & ~n7518 ;
  assign n7520 = n6475 ^ n3217 ^ n1769 ;
  assign n7521 = n5023 | n7520 ;
  assign n7522 = n5071 ^ n1537 ^ 1'b0 ;
  assign n7523 = n491 & n7522 ;
  assign n7532 = ( n1521 & ~n2572 ) | ( n1521 & n3592 ) | ( ~n2572 & n3592 ) ;
  assign n7528 = n4942 ^ n2781 ^ n2111 ;
  assign n7529 = n2063 & ~n7528 ;
  assign n7530 = n6725 & n7529 ;
  assign n7524 = ( n1211 & n1323 ) | ( n1211 & ~n2058 ) | ( n1323 & ~n2058 ) ;
  assign n7525 = n1597 & n3943 ;
  assign n7526 = n7525 ^ n2113 ^ 1'b0 ;
  assign n7527 = ~n7524 & n7526 ;
  assign n7531 = n7530 ^ n7527 ^ 1'b0 ;
  assign n7533 = n7532 ^ n7531 ^ 1'b0 ;
  assign n7534 = n7523 & ~n7533 ;
  assign n7538 = n1143 & n4571 ;
  assign n7539 = n7538 ^ n1568 ^ 1'b0 ;
  assign n7540 = n7539 ^ n1487 ^ n1450 ;
  assign n7541 = n3872 & ~n5667 ;
  assign n7542 = n7540 & n7541 ;
  assign n7535 = n2776 ^ x13 ^ 1'b0 ;
  assign n7536 = n3524 & n7535 ;
  assign n7537 = n4867 & n7536 ;
  assign n7543 = n7542 ^ n7537 ^ 1'b0 ;
  assign n7544 = n7251 ^ n3881 ^ 1'b0 ;
  assign n7545 = n4750 & n7544 ;
  assign n7559 = n888 & n2660 ;
  assign n7554 = n679 & n2150 ;
  assign n7555 = ~n2536 & n7554 ;
  assign n7556 = ( n752 & n5040 ) | ( n752 & n5655 ) | ( n5040 & n5655 ) ;
  assign n7557 = n350 & ~n7556 ;
  assign n7558 = n7555 & n7557 ;
  assign n7560 = n7559 ^ n7558 ^ n927 ;
  assign n7549 = ~n531 & n1548 ;
  assign n7550 = n7549 ^ n2205 ^ 1'b0 ;
  assign n7548 = n566 | n7339 ;
  assign n7551 = n7550 ^ n7548 ^ 1'b0 ;
  assign n7552 = n7551 ^ n7413 ^ 1'b0 ;
  assign n7553 = ~n248 & n7552 ;
  assign n7546 = n4675 & ~n7332 ;
  assign n7547 = n7546 ^ n1022 ^ 1'b0 ;
  assign n7561 = n7560 ^ n7553 ^ n7547 ;
  assign n7562 = n3799 ^ n477 ^ n394 ;
  assign n7563 = n1762 ^ n1159 ^ n485 ;
  assign n7567 = n940 | n4201 ;
  assign n7568 = n7567 ^ n3861 ^ 1'b0 ;
  assign n7564 = n573 ^ x125 ^ 1'b0 ;
  assign n7565 = n1490 & ~n7564 ;
  assign n7566 = ~n675 & n7565 ;
  assign n7569 = n7568 ^ n7566 ^ n7385 ;
  assign n7571 = n6382 ^ n2641 ^ 1'b0 ;
  assign n7570 = n4216 | n6370 ;
  assign n7572 = n7571 ^ n7570 ^ 1'b0 ;
  assign n7573 = n5811 ^ n2242 ^ 1'b0 ;
  assign n7574 = n7572 & n7573 ;
  assign n7575 = n7574 ^ n3629 ^ 1'b0 ;
  assign n7576 = n7575 ^ n7197 ^ n2944 ;
  assign n7577 = n6480 ^ n2380 ^ 1'b0 ;
  assign n7578 = n5110 & n7577 ;
  assign n7579 = ( ~n1686 & n5726 ) | ( ~n1686 & n7578 ) | ( n5726 & n7578 ) ;
  assign n7580 = n4049 ^ n1944 ^ 1'b0 ;
  assign n7581 = n3393 | n7580 ;
  assign n7582 = n7579 & ~n7581 ;
  assign n7583 = ~n200 & n310 ;
  assign n7584 = n7583 ^ n6562 ^ 1'b0 ;
  assign n7585 = n7584 ^ n4183 ^ x21 ;
  assign n7587 = ~n2244 & n2324 ;
  assign n7588 = n7587 ^ n4269 ^ 1'b0 ;
  assign n7586 = ( n149 & ~n451 ) | ( n149 & n5443 ) | ( ~n451 & n5443 ) ;
  assign n7589 = n7588 ^ n7586 ^ 1'b0 ;
  assign n7590 = n1850 & n6359 ;
  assign n7591 = n7590 ^ n2956 ^ 1'b0 ;
  assign n7592 = n594 & ~n1193 ;
  assign n7593 = ~n169 & n7592 ;
  assign n7594 = n3484 & n6835 ;
  assign n7595 = ( n1467 & n1772 ) | ( n1467 & n7594 ) | ( n1772 & n7594 ) ;
  assign n7596 = n7088 ^ n1745 ^ 1'b0 ;
  assign n7597 = n6101 ^ n3727 ^ 1'b0 ;
  assign n7598 = n7415 | n7597 ;
  assign n7599 = n7598 ^ n3244 ^ 1'b0 ;
  assign n7600 = n2200 ^ n1759 ^ 1'b0 ;
  assign n7601 = ( n1188 & ~n1366 ) | ( n1188 & n7600 ) | ( ~n1366 & n7600 ) ;
  assign n7602 = ( n1138 & ~n6226 ) | ( n1138 & n7594 ) | ( ~n6226 & n7594 ) ;
  assign n7603 = n7602 ^ n6755 ^ 1'b0 ;
  assign n7604 = n7601 & ~n7603 ;
  assign n7605 = ( n1317 & n3176 ) | ( n1317 & n4630 ) | ( n3176 & n4630 ) ;
  assign n7606 = n2328 | n3616 ;
  assign n7607 = n7606 ^ n2599 ^ 1'b0 ;
  assign n7608 = ~n2511 & n7607 ;
  assign n7610 = n2262 ^ n445 ^ 1'b0 ;
  assign n7611 = n7407 | n7610 ;
  assign n7609 = n1538 & ~n2440 ;
  assign n7612 = n7611 ^ n7609 ^ 1'b0 ;
  assign n7613 = n388 & ~n2975 ;
  assign n7614 = n3888 ^ n1460 ^ 1'b0 ;
  assign n7615 = n7613 | n7614 ;
  assign n7616 = n7615 ^ n3409 ^ 1'b0 ;
  assign n7617 = n7616 ^ n5801 ^ n294 ;
  assign n7618 = n2058 & n3542 ;
  assign n7619 = n7618 ^ n3801 ^ n1618 ;
  assign n7620 = ~n1934 & n3607 ;
  assign n7621 = n7620 ^ n3340 ^ 1'b0 ;
  assign n7622 = n7621 ^ n2733 ^ n509 ;
  assign n7623 = n2111 ^ n267 ^ 1'b0 ;
  assign n7624 = n4320 & n7623 ;
  assign n7625 = ( ~n3956 & n6466 ) | ( ~n3956 & n7624 ) | ( n6466 & n7624 ) ;
  assign n7626 = n7625 ^ n2067 ^ n1053 ;
  assign n7627 = ~n3202 & n7626 ;
  assign n7628 = n4181 & ~n7627 ;
  assign n7629 = n2737 | n5032 ;
  assign n7630 = ( n1230 & n4791 ) | ( n1230 & ~n7629 ) | ( n4791 & ~n7629 ) ;
  assign n7631 = n885 ^ n298 ^ 1'b0 ;
  assign n7632 = n3073 | n7631 ;
  assign n7633 = n5228 & ~n7632 ;
  assign n7634 = n7269 ^ n2038 ^ n456 ;
  assign n7638 = n1666 & n1777 ;
  assign n7639 = n7638 ^ n1422 ^ 1'b0 ;
  assign n7640 = n636 & ~n7639 ;
  assign n7641 = n7113 ^ n2870 ^ n1030 ;
  assign n7642 = ~n7640 & n7641 ;
  assign n7643 = n2921 & n7642 ;
  assign n7635 = n1867 & n3075 ;
  assign n7636 = n1829 & n3059 ;
  assign n7637 = ~n7635 & n7636 ;
  assign n7644 = n7643 ^ n7637 ^ 1'b0 ;
  assign n7647 = n2101 ^ n1134 ^ 1'b0 ;
  assign n7648 = ~n861 & n7647 ;
  assign n7649 = ~n794 & n7648 ;
  assign n7650 = n7649 ^ n3888 ^ n1700 ;
  assign n7645 = n4118 & ~n4576 ;
  assign n7646 = ~n4224 & n7645 ;
  assign n7651 = n7650 ^ n7646 ^ 1'b0 ;
  assign n7652 = x91 & n7651 ;
  assign n7653 = n5562 ^ n2832 ^ 1'b0 ;
  assign n7654 = n5503 & n7653 ;
  assign n7655 = n208 & n7654 ;
  assign n7656 = n4374 ^ n1400 ^ 1'b0 ;
  assign n7657 = ~n5387 & n7656 ;
  assign n7658 = ~n7655 & n7657 ;
  assign n7659 = n5328 & n7658 ;
  assign n7660 = ( ~n2884 & n3102 ) | ( ~n2884 & n4704 ) | ( n3102 & n4704 ) ;
  assign n7661 = n7660 ^ n3025 ^ n182 ;
  assign n7662 = n1994 | n7661 ;
  assign n7663 = n1108 | n7662 ;
  assign n7664 = n7663 ^ n5472 ^ 1'b0 ;
  assign n7665 = n5873 ^ n2934 ^ 1'b0 ;
  assign n7666 = ( n655 & n2086 ) | ( n655 & ~n6886 ) | ( n2086 & ~n6886 ) ;
  assign n7667 = n2589 ^ n332 ^ 1'b0 ;
  assign n7668 = n1405 & n7667 ;
  assign n7669 = n7666 & n7668 ;
  assign n7670 = n7669 ^ n3533 ^ 1'b0 ;
  assign n7671 = n7417 & ~n7670 ;
  assign n7673 = n4642 ^ n2462 ^ 1'b0 ;
  assign n7674 = n2993 & n7673 ;
  assign n7675 = n1306 & n7674 ;
  assign n7672 = n2361 & ~n6281 ;
  assign n7676 = n7675 ^ n7672 ^ 1'b0 ;
  assign n7677 = n5420 ^ n608 ^ 1'b0 ;
  assign n7678 = n1821 & ~n7677 ;
  assign n7679 = n2743 & n7678 ;
  assign n7680 = ~x25 & n7584 ;
  assign n7681 = n810 | n1190 ;
  assign n7682 = n3134 & ~n7681 ;
  assign n7683 = n7682 ^ n1553 ^ 1'b0 ;
  assign n7684 = ~n3611 & n7243 ;
  assign n7685 = n7684 ^ n3971 ^ n305 ;
  assign n7687 = n285 & ~n1940 ;
  assign n7688 = ~n4587 & n7687 ;
  assign n7686 = n3402 & ~n4397 ;
  assign n7689 = n7688 ^ n7686 ^ 1'b0 ;
  assign n7690 = x6 & n2532 ;
  assign n7691 = n7503 & n7690 ;
  assign n7692 = n7691 ^ n2243 ^ 1'b0 ;
  assign n7693 = ~n4990 & n7669 ;
  assign n7694 = ~n3612 & n4912 ;
  assign n7695 = n7694 ^ n333 ^ 1'b0 ;
  assign n7698 = n4807 ^ n982 ^ n646 ;
  assign n7696 = n1793 ^ n1154 ^ 1'b0 ;
  assign n7697 = ~n2436 & n7696 ;
  assign n7699 = n7698 ^ n7697 ^ 1'b0 ;
  assign n7700 = ~n2354 & n7699 ;
  assign n7701 = n7700 ^ n3134 ^ n557 ;
  assign n7702 = ~n5455 & n7701 ;
  assign n7703 = x0 & ~n2870 ;
  assign n7704 = n7703 ^ n6639 ^ 1'b0 ;
  assign n7705 = ( n1256 & n5238 ) | ( n1256 & n7704 ) | ( n5238 & n7704 ) ;
  assign n7706 = n6845 ^ n3200 ^ n1611 ;
  assign n7707 = ( ~n7702 & n7705 ) | ( ~n7702 & n7706 ) | ( n7705 & n7706 ) ;
  assign n7708 = ( n5521 & ~n7695 ) | ( n5521 & n7707 ) | ( ~n7695 & n7707 ) ;
  assign n7709 = n3096 | n7349 ;
  assign n7710 = n7709 ^ n363 ^ 1'b0 ;
  assign n7711 = ( n3256 & n5230 ) | ( n3256 & n7710 ) | ( n5230 & n7710 ) ;
  assign n7712 = n3945 ^ n2898 ^ n2222 ;
  assign n7713 = n6930 & n7712 ;
  assign n7714 = n7713 ^ n5600 ^ 1'b0 ;
  assign n7718 = n5764 & ~n6104 ;
  assign n7719 = n5521 & n7718 ;
  assign n7720 = ( ~n2466 & n3126 ) | ( ~n2466 & n4974 ) | ( n3126 & n4974 ) ;
  assign n7721 = ( n3573 & n7719 ) | ( n3573 & n7720 ) | ( n7719 & n7720 ) ;
  assign n7715 = n1462 & n6940 ;
  assign n7716 = n7715 ^ n5836 ^ 1'b0 ;
  assign n7717 = n7716 ^ n2443 ^ n732 ;
  assign n7722 = n7721 ^ n7717 ^ n6918 ;
  assign n7723 = n589 & n1429 ;
  assign n7724 = n1943 & n7723 ;
  assign n7725 = n3451 ^ n3003 ^ 1'b0 ;
  assign n7726 = n2310 ^ n1641 ^ 1'b0 ;
  assign n7727 = n7726 ^ n6393 ^ n852 ;
  assign n7729 = x116 & ~n565 ;
  assign n7730 = n7729 ^ n2377 ^ n2198 ;
  assign n7728 = n624 & n3237 ;
  assign n7731 = n7730 ^ n7728 ^ 1'b0 ;
  assign n7732 = n7731 ^ n7113 ^ 1'b0 ;
  assign n7733 = n7732 ^ n6566 ^ n5756 ;
  assign n7734 = n7733 ^ n6291 ^ n4002 ;
  assign n7737 = n3171 ^ n1013 ^ n171 ;
  assign n7738 = ( n2770 & ~n3042 ) | ( n2770 & n7737 ) | ( ~n3042 & n7737 ) ;
  assign n7739 = ( n1482 & n1513 ) | ( n1482 & n7738 ) | ( n1513 & n7738 ) ;
  assign n7740 = ( n2421 & n5144 ) | ( n2421 & ~n7739 ) | ( n5144 & ~n7739 ) ;
  assign n7735 = n4413 ^ n1901 ^ 1'b0 ;
  assign n7736 = n7628 & n7735 ;
  assign n7741 = n7740 ^ n7736 ^ 1'b0 ;
  assign n7743 = n3451 ^ n2688 ^ 1'b0 ;
  assign n7742 = ~n2487 & n5272 ;
  assign n7744 = n7743 ^ n7742 ^ n1745 ;
  assign n7745 = ~n2372 & n7239 ;
  assign n7746 = n230 & n7745 ;
  assign n7747 = n3087 & n7746 ;
  assign n7748 = n3254 ^ n2626 ^ n2239 ;
  assign n7749 = n6675 ^ n4857 ^ 1'b0 ;
  assign n7750 = n7748 & n7749 ;
  assign n7751 = ~n4010 & n7750 ;
  assign n7752 = ~n2632 & n6803 ;
  assign n7753 = x113 & n7752 ;
  assign n7759 = n6364 ^ n5690 ^ n1070 ;
  assign n7754 = n3144 & n6799 ;
  assign n7755 = n6012 ^ n4200 ^ 1'b0 ;
  assign n7756 = n5390 & n7755 ;
  assign n7757 = ( ~n6254 & n7754 ) | ( ~n6254 & n7756 ) | ( n7754 & n7756 ) ;
  assign n7758 = n3924 & n7757 ;
  assign n7760 = n7759 ^ n7758 ^ 1'b0 ;
  assign n7761 = n2408 & ~n6357 ;
  assign n7762 = n7761 ^ n1770 ^ 1'b0 ;
  assign n7763 = n2811 ^ n571 ^ n272 ;
  assign n7764 = n6924 & n7763 ;
  assign n7765 = ~n4818 & n7764 ;
  assign n7766 = ( x0 & n3862 ) | ( x0 & n5557 ) | ( n3862 & n5557 ) ;
  assign n7767 = n920 & n1420 ;
  assign n7768 = n7767 ^ n7204 ^ 1'b0 ;
  assign n7769 = n7768 ^ n4960 ^ 1'b0 ;
  assign n7772 = n1374 ^ x24 ^ 1'b0 ;
  assign n7770 = ( n468 & ~n815 ) | ( n468 & n4160 ) | ( ~n815 & n4160 ) ;
  assign n7771 = ~n1235 & n7770 ;
  assign n7773 = n7772 ^ n7771 ^ n3398 ;
  assign n7782 = n4536 ^ n3418 ^ n485 ;
  assign n7783 = ( ~n3459 & n7102 ) | ( ~n3459 & n7782 ) | ( n7102 & n7782 ) ;
  assign n7780 = n366 & ~n460 ;
  assign n7774 = n4717 ^ n2130 ^ x30 ;
  assign n7775 = n7774 ^ x67 ^ 1'b0 ;
  assign n7776 = n4252 & ~n7775 ;
  assign n7777 = n755 & n7776 ;
  assign n7778 = n7777 ^ n4605 ^ 1'b0 ;
  assign n7779 = n1923 & ~n7778 ;
  assign n7781 = n7780 ^ n7779 ^ n2151 ;
  assign n7784 = n7783 ^ n7781 ^ 1'b0 ;
  assign n7789 = n5629 ^ x19 ^ 1'b0 ;
  assign n7786 = ( n627 & ~n2687 ) | ( n627 & n3470 ) | ( ~n2687 & n3470 ) ;
  assign n7785 = ( ~n2433 & n4357 ) | ( ~n2433 & n4811 ) | ( n4357 & n4811 ) ;
  assign n7787 = n7786 ^ n7785 ^ 1'b0 ;
  assign n7788 = n5842 & ~n7787 ;
  assign n7790 = n7789 ^ n7788 ^ n3696 ;
  assign n7791 = n2934 & n3385 ;
  assign n7792 = n7791 ^ n3501 ^ x102 ;
  assign n7793 = ( x87 & ~n388 ) | ( x87 & n7792 ) | ( ~n388 & n7792 ) ;
  assign n7794 = ( n2522 & n2898 ) | ( n2522 & n2992 ) | ( n2898 & n2992 ) ;
  assign n7795 = n7794 ^ n3625 ^ n1883 ;
  assign n7796 = n2523 & ~n6575 ;
  assign n7797 = n2219 ^ n2010 ^ n1935 ;
  assign n7798 = ( n3580 & n7796 ) | ( n3580 & ~n7797 ) | ( n7796 & ~n7797 ) ;
  assign n7799 = n7795 | n7798 ;
  assign n7800 = n7793 | n7799 ;
  assign n7801 = ~n6853 & n7800 ;
  assign n7802 = n424 | n2303 ;
  assign n7803 = ~n4955 & n5064 ;
  assign n7804 = ~n7802 & n7803 ;
  assign n7805 = ( n894 & n3897 ) | ( n894 & n5062 ) | ( n3897 & n5062 ) ;
  assign n7806 = n5942 ^ n2985 ^ n1250 ;
  assign n7807 = ( n1394 & n3921 ) | ( n1394 & ~n7806 ) | ( n3921 & ~n7806 ) ;
  assign n7808 = ~n2542 & n5351 ;
  assign n7809 = ~n1814 & n7808 ;
  assign n7810 = n921 & ~n5052 ;
  assign n7811 = n7810 ^ x19 ^ 1'b0 ;
  assign n7812 = ~n2885 & n7811 ;
  assign n7813 = n7812 ^ n3200 ^ n2678 ;
  assign n7814 = ( x90 & ~n3766 ) | ( x90 & n7813 ) | ( ~n3766 & n7813 ) ;
  assign n7815 = ( n848 & ~n7809 ) | ( n848 & n7814 ) | ( ~n7809 & n7814 ) ;
  assign n7816 = n5962 ^ n1188 ^ 1'b0 ;
  assign n7817 = n7816 ^ n3653 ^ n3611 ;
  assign n7818 = n1028 & ~n6914 ;
  assign n7819 = n7818 ^ n1258 ^ 1'b0 ;
  assign n7820 = n4642 ^ n2360 ^ 1'b0 ;
  assign n7825 = ( ~n947 & n2870 ) | ( ~n947 & n3929 ) | ( n2870 & n3929 ) ;
  assign n7821 = n1764 & n3386 ;
  assign n7822 = n4012 & n7821 ;
  assign n7823 = n7822 ^ n2587 ^ 1'b0 ;
  assign n7824 = n2830 | n7823 ;
  assign n7826 = n7825 ^ n7824 ^ n270 ;
  assign n7832 = ( n1405 & n2511 ) | ( n1405 & n3341 ) | ( n2511 & n3341 ) ;
  assign n7831 = n210 | n3715 ;
  assign n7833 = n7832 ^ n7831 ^ 1'b0 ;
  assign n7834 = n7833 ^ n5498 ^ 1'b0 ;
  assign n7835 = n2204 | n7834 ;
  assign n7828 = n5511 ^ n2163 ^ n462 ;
  assign n7827 = n7200 ^ n4343 ^ n4260 ;
  assign n7829 = n7828 ^ n7827 ^ n5488 ;
  assign n7830 = n7088 & n7829 ;
  assign n7836 = n7835 ^ n7830 ^ n5318 ;
  assign n7837 = n3489 | n4469 ;
  assign n7838 = n797 & ~n7837 ;
  assign n7839 = ( n464 & n1288 ) | ( n464 & ~n1783 ) | ( n1288 & ~n1783 ) ;
  assign n7840 = n7839 ^ n2668 ^ x19 ;
  assign n7841 = n2921 | n7840 ;
  assign n7842 = n7841 ^ n3567 ^ 1'b0 ;
  assign n7843 = n5665 ^ n920 ^ 1'b0 ;
  assign n7844 = ( n7838 & ~n7842 ) | ( n7838 & n7843 ) | ( ~n7842 & n7843 ) ;
  assign n7845 = n7844 ^ n3971 ^ n724 ;
  assign n7846 = ~n3069 & n4660 ;
  assign n7847 = n2071 | n5718 ;
  assign n7848 = n7847 ^ n791 ^ 1'b0 ;
  assign n7853 = n2927 ^ n2748 ^ 1'b0 ;
  assign n7851 = n2311 & n4000 ;
  assign n7852 = n7851 ^ n5259 ^ 1'b0 ;
  assign n7849 = ~n413 & n4522 ;
  assign n7850 = ~x13 & n7849 ;
  assign n7854 = n7853 ^ n7852 ^ n7850 ;
  assign n7855 = ( n4216 & ~n7848 ) | ( n4216 & n7854 ) | ( ~n7848 & n7854 ) ;
  assign n7856 = n196 | n5164 ;
  assign n7857 = n1374 & ~n7856 ;
  assign n7858 = n7857 ^ n3934 ^ 1'b0 ;
  assign n7859 = n7855 & n7858 ;
  assign n7860 = n3277 ^ n2798 ^ 1'b0 ;
  assign n7861 = n7859 & n7860 ;
  assign n7862 = ~n1246 & n5573 ;
  assign n7863 = n5621 & n7862 ;
  assign n7864 = n1071 | n7863 ;
  assign n7865 = n169 & ~n2182 ;
  assign n7866 = n3394 | n7865 ;
  assign n7867 = n7866 ^ n4195 ^ 1'b0 ;
  assign n7868 = n6982 & ~n7867 ;
  assign n7869 = n6416 ^ n2418 ^ 1'b0 ;
  assign n7870 = n7869 ^ n3032 ^ 1'b0 ;
  assign n7871 = ~n2810 & n7870 ;
  assign n7872 = ~n3424 & n3853 ;
  assign n7873 = n3587 & n7872 ;
  assign n7877 = n3383 ^ n1743 ^ 1'b0 ;
  assign n7878 = n4750 & n7877 ;
  assign n7874 = n1591 ^ n829 ^ n392 ;
  assign n7875 = ( n2567 & ~n3651 ) | ( n2567 & n7874 ) | ( ~n3651 & n7874 ) ;
  assign n7876 = ( n1554 & n1695 ) | ( n1554 & ~n7875 ) | ( n1695 & ~n7875 ) ;
  assign n7879 = n7878 ^ n7876 ^ n2199 ;
  assign n7880 = ~n866 & n4528 ;
  assign n7881 = n2377 & n7880 ;
  assign n7885 = n7782 ^ n4200 ^ n1731 ;
  assign n7882 = n1334 ^ n680 ^ x41 ;
  assign n7883 = n2687 | n7882 ;
  assign n7884 = n4875 & ~n7883 ;
  assign n7886 = n7885 ^ n7884 ^ n747 ;
  assign n7887 = n6811 ^ n1407 ^ 1'b0 ;
  assign n7888 = ~n5507 & n7887 ;
  assign n7889 = n4294 & n7888 ;
  assign n7890 = n331 & ~n7889 ;
  assign n7896 = n3399 ^ n3258 ^ n979 ;
  assign n7893 = x44 & ~n265 ;
  assign n7894 = n7893 ^ n1349 ^ 1'b0 ;
  assign n7895 = x102 & n7894 ;
  assign n7897 = n7896 ^ n7895 ^ 1'b0 ;
  assign n7891 = ( n224 & ~n3692 ) | ( n224 & n7866 ) | ( ~n3692 & n7866 ) ;
  assign n7892 = n5231 & ~n7891 ;
  assign n7898 = n7897 ^ n7892 ^ 1'b0 ;
  assign n7899 = n3200 ^ n2926 ^ n915 ;
  assign n7900 = n6510 ^ n6507 ^ n3619 ;
  assign n7901 = n3919 ^ n2175 ^ 1'b0 ;
  assign n7902 = n4762 & n7901 ;
  assign n7903 = n7902 ^ n6012 ^ n4304 ;
  assign n7906 = n3179 | n5468 ;
  assign n7907 = n7906 ^ n5198 ^ 1'b0 ;
  assign n7904 = ~n320 & n1105 ;
  assign n7905 = n7904 ^ n5360 ^ 1'b0 ;
  assign n7908 = n7907 ^ n7905 ^ 1'b0 ;
  assign n7909 = n6353 ^ n6180 ^ n4164 ;
  assign n7913 = ( n1569 & n2426 ) | ( n1569 & n4247 ) | ( n2426 & n4247 ) ;
  assign n7911 = n6066 ^ n304 ^ 1'b0 ;
  assign n7912 = ( n1964 & n2511 ) | ( n1964 & ~n7911 ) | ( n2511 & ~n7911 ) ;
  assign n7910 = ~n2418 & n6856 ;
  assign n7914 = n7913 ^ n7912 ^ n7910 ;
  assign n7915 = ~n7909 & n7914 ;
  assign n7916 = n6314 & n7915 ;
  assign n7918 = n4059 ^ n1422 ^ 1'b0 ;
  assign n7917 = n7840 ^ n2036 ^ 1'b0 ;
  assign n7919 = n7918 ^ n7917 ^ n3121 ;
  assign n7920 = n5298 & n5398 ;
  assign n7921 = n3801 ^ x114 ^ 1'b0 ;
  assign n7922 = n5764 ^ n2018 ^ 1'b0 ;
  assign n7923 = ~n1601 & n7922 ;
  assign n7924 = ( n2385 & ~n7921 ) | ( n2385 & n7923 ) | ( ~n7921 & n7923 ) ;
  assign n7929 = ( n1547 & n1986 ) | ( n1547 & n4123 ) | ( n1986 & n4123 ) ;
  assign n7925 = n2918 | n3257 ;
  assign n7926 = n1028 | n7925 ;
  assign n7927 = n2592 & n7926 ;
  assign n7928 = n7927 ^ n3096 ^ 1'b0 ;
  assign n7930 = n7929 ^ n7928 ^ 1'b0 ;
  assign n7931 = ( x9 & ~n675 ) | ( x9 & n1061 ) | ( ~n675 & n1061 ) ;
  assign n7932 = n4302 ^ n512 ^ 1'b0 ;
  assign n7933 = ( n3177 & n7931 ) | ( n3177 & ~n7932 ) | ( n7931 & ~n7932 ) ;
  assign n7934 = ( n3415 & n3642 ) | ( n3415 & ~n6811 ) | ( n3642 & ~n6811 ) ;
  assign n7935 = ( ~n443 & n6602 ) | ( ~n443 & n7934 ) | ( n6602 & n7934 ) ;
  assign n7936 = ~n171 & n6961 ;
  assign n7937 = n7270 | n7936 ;
  assign n7938 = n3293 | n7937 ;
  assign n7939 = x108 & n5513 ;
  assign n7942 = n1912 ^ n1226 ^ n1067 ;
  assign n7940 = ( n237 & n1084 ) | ( n237 & n4097 ) | ( n1084 & n4097 ) ;
  assign n7941 = n7940 ^ n368 ^ 1'b0 ;
  assign n7943 = n7942 ^ n7941 ^ n2623 ;
  assign n7944 = n2199 & ~n7943 ;
  assign n7945 = n7944 ^ n401 ^ 1'b0 ;
  assign n7946 = ( n601 & ~n1251 ) | ( n601 & n7945 ) | ( ~n1251 & n7945 ) ;
  assign n7947 = ( n6214 & n6920 ) | ( n6214 & ~n7822 ) | ( n6920 & ~n7822 ) ;
  assign n7948 = n2878 & ~n6092 ;
  assign n7949 = n3721 ^ n2007 ^ n452 ;
  assign n7950 = n5935 ^ x5 ^ 1'b0 ;
  assign n7951 = n5493 & ~n7950 ;
  assign n7952 = n7951 ^ n1355 ^ n796 ;
  assign n7953 = n850 | n7952 ;
  assign n7954 = n7949 | n7953 ;
  assign n7955 = ~n4048 & n7954 ;
  assign n7956 = ( n1861 & ~n3254 ) | ( n1861 & n7955 ) | ( ~n3254 & n7955 ) ;
  assign n7957 = ( ~n647 & n7948 ) | ( ~n647 & n7956 ) | ( n7948 & n7956 ) ;
  assign n7958 = n3653 ^ n2959 ^ 1'b0 ;
  assign n7959 = n7472 ^ n4534 ^ n2072 ;
  assign n7960 = n7959 ^ n7731 ^ x123 ;
  assign n7961 = ( n5023 & ~n7958 ) | ( n5023 & n7960 ) | ( ~n7958 & n7960 ) ;
  assign n7962 = n7806 ^ n3893 ^ 1'b0 ;
  assign n7963 = n7238 & n7962 ;
  assign n7966 = n1067 ^ n985 ^ 1'b0 ;
  assign n7967 = x59 & ~n1059 ;
  assign n7968 = ~n7966 & n7967 ;
  assign n7964 = ~n1714 & n1952 ;
  assign n7965 = n7964 ^ n5567 ^ 1'b0 ;
  assign n7969 = n7968 ^ n7965 ^ n4713 ;
  assign n7970 = n1077 ^ n727 ^ 1'b0 ;
  assign n7971 = n7969 & ~n7970 ;
  assign n7972 = x90 | n7528 ;
  assign n7973 = n2917 ^ n1783 ^ 1'b0 ;
  assign n7974 = n2705 & ~n7973 ;
  assign n7975 = ~n3607 & n7974 ;
  assign n7976 = ~n7972 & n7975 ;
  assign n7980 = n501 & ~n547 ;
  assign n7981 = n7980 ^ n331 ^ 1'b0 ;
  assign n7982 = n5873 & ~n7981 ;
  assign n7977 = n1349 ^ n318 ^ 1'b0 ;
  assign n7978 = ~n2567 & n7977 ;
  assign n7979 = ( n3688 & ~n7355 ) | ( n3688 & n7978 ) | ( ~n7355 & n7978 ) ;
  assign n7983 = n7982 ^ n7979 ^ n3358 ;
  assign n7984 = n7695 ^ n3562 ^ x19 ;
  assign n7985 = n2337 ^ n2227 ^ n946 ;
  assign n7986 = n3749 | n7985 ;
  assign n7987 = n7986 ^ n1211 ^ 1'b0 ;
  assign n7995 = n1501 & n6235 ;
  assign n7993 = n5391 ^ n4157 ^ 1'b0 ;
  assign n7988 = n589 ^ n474 ^ n259 ;
  assign n7989 = n474 & n5274 ;
  assign n7990 = n7989 ^ n4073 ^ 1'b0 ;
  assign n7991 = n4323 & n7990 ;
  assign n7992 = ~n7988 & n7991 ;
  assign n7994 = n7993 ^ n7992 ^ n5421 ;
  assign n7996 = n7995 ^ n7994 ^ 1'b0 ;
  assign n7997 = n1907 | n7996 ;
  assign n7998 = n1455 ^ n958 ^ 1'b0 ;
  assign n7999 = n3732 | n7998 ;
  assign n8000 = ~n2985 & n6813 ;
  assign n8001 = n2835 & ~n5131 ;
  assign n8002 = n8001 ^ n5659 ^ 1'b0 ;
  assign n8003 = ( ~n3784 & n5973 ) | ( ~n3784 & n8002 ) | ( n5973 & n8002 ) ;
  assign n8004 = n4008 ^ n2608 ^ 1'b0 ;
  assign n8005 = n6301 ^ n2178 ^ 1'b0 ;
  assign n8007 = n7344 & ~n7388 ;
  assign n8008 = n8007 ^ n2951 ^ 1'b0 ;
  assign n8006 = n5145 | n7167 ;
  assign n8009 = n8008 ^ n8006 ^ n2564 ;
  assign n8010 = n4569 ^ n4103 ^ n3375 ;
  assign n8011 = n5338 | n8010 ;
  assign n8012 = n4699 ^ n4252 ^ n2418 ;
  assign n8013 = n3888 | n6985 ;
  assign n8014 = n1332 | n8013 ;
  assign n8015 = n3718 ^ n2264 ^ n1804 ;
  assign n8016 = n3206 & n7523 ;
  assign n8017 = n6546 & n8016 ;
  assign n8018 = ( n6053 & n7797 ) | ( n6053 & n8017 ) | ( n7797 & n8017 ) ;
  assign n8019 = n8018 ^ n807 ^ n693 ;
  assign n8020 = n1125 & n2563 ;
  assign n8021 = n1822 & ~n8020 ;
  assign n8022 = n2951 & n8021 ;
  assign n8023 = n5606 ^ x126 ^ 1'b0 ;
  assign n8024 = ( n5249 & n7942 ) | ( n5249 & ~n8023 ) | ( n7942 & ~n8023 ) ;
  assign n8025 = n572 & n824 ;
  assign n8026 = n7483 ^ n6085 ^ 1'b0 ;
  assign n8035 = n3429 ^ n1523 ^ n1462 ;
  assign n8036 = n3396 & n8035 ;
  assign n8037 = ~n3926 & n8036 ;
  assign n8038 = ~n3227 & n8037 ;
  assign n8039 = n8038 ^ n1519 ^ 1'b0 ;
  assign n8031 = n4201 ^ n523 ^ 1'b0 ;
  assign n8032 = n8031 ^ n4742 ^ n2360 ;
  assign n8028 = n2724 ^ n1966 ^ n1883 ;
  assign n8027 = n3762 & n4733 ;
  assign n8029 = n8028 ^ n8027 ^ 1'b0 ;
  assign n8030 = n5076 | n8029 ;
  assign n8033 = n8032 ^ n8030 ^ 1'b0 ;
  assign n8034 = n550 | n8033 ;
  assign n8040 = n8039 ^ n8034 ^ 1'b0 ;
  assign n8041 = ~n903 & n2522 ;
  assign n8042 = n781 & n2822 ;
  assign n8043 = ( n5888 & ~n5948 ) | ( n5888 & n8042 ) | ( ~n5948 & n8042 ) ;
  assign n8044 = ~n8041 & n8043 ;
  assign n8045 = n5334 & n8044 ;
  assign n8046 = n1697 | n6136 ;
  assign n8047 = n364 & n4296 ;
  assign n8048 = n8047 ^ n4224 ^ n2752 ;
  assign n8049 = n2945 ^ n2067 ^ n692 ;
  assign n8050 = n2536 & n8049 ;
  assign n8051 = n866 & n8050 ;
  assign n8052 = n8051 ^ n5220 ^ n2153 ;
  assign n8053 = ~n4299 & n7840 ;
  assign n8054 = ( n174 & n1342 ) | ( n174 & ~n8053 ) | ( n1342 & ~n8053 ) ;
  assign n8055 = ( ~n2154 & n5117 ) | ( ~n2154 & n8054 ) | ( n5117 & n8054 ) ;
  assign n8056 = ( ~n230 & n4133 ) | ( ~n230 & n5445 ) | ( n4133 & n5445 ) ;
  assign n8057 = n1646 & n6016 ;
  assign n8058 = n8057 ^ n5449 ^ 1'b0 ;
  assign n8059 = n3597 ^ n2732 ^ n1201 ;
  assign n8060 = n2163 & ~n8059 ;
  assign n8061 = n8060 ^ n6796 ^ 1'b0 ;
  assign n8062 = ( ~n1027 & n8058 ) | ( ~n1027 & n8061 ) | ( n8058 & n8061 ) ;
  assign n8063 = n2749 & n6750 ;
  assign n8064 = ~n2444 & n8063 ;
  assign n8065 = x111 & ~n3848 ;
  assign n8066 = n2553 ^ n692 ^ 1'b0 ;
  assign n8067 = ( n2469 & n8065 ) | ( n2469 & n8066 ) | ( n8065 & n8066 ) ;
  assign n8068 = ( n2161 & n7555 ) | ( n2161 & ~n8067 ) | ( n7555 & ~n8067 ) ;
  assign n8069 = n3764 ^ n826 ^ x70 ;
  assign n8070 = ~n1262 & n2348 ;
  assign n8071 = n8070 ^ n527 ^ 1'b0 ;
  assign n8072 = n3772 | n8071 ;
  assign n8073 = n8072 ^ n6728 ^ 1'b0 ;
  assign n8076 = ( n295 & ~n1575 ) | ( n295 & n1704 ) | ( ~n1575 & n1704 ) ;
  assign n8077 = n8076 ^ n2931 ^ 1'b0 ;
  assign n8078 = n8077 ^ n5458 ^ n4064 ;
  assign n8074 = n655 & n2968 ;
  assign n8075 = ( n6995 & n7666 ) | ( n6995 & n8074 ) | ( n7666 & n8074 ) ;
  assign n8079 = n8078 ^ n8075 ^ 1'b0 ;
  assign n8080 = ( n8069 & ~n8073 ) | ( n8069 & n8079 ) | ( ~n8073 & n8079 ) ;
  assign n8081 = n8080 ^ n7914 ^ n1619 ;
  assign n8082 = n3556 & n8081 ;
  assign n8083 = n8082 ^ n1691 ^ 1'b0 ;
  assign n8084 = n2813 ^ n2640 ^ 1'b0 ;
  assign n8085 = n3123 ^ n3031 ^ 1'b0 ;
  assign n8086 = n8084 | n8085 ;
  assign n8087 = n7042 ^ n4354 ^ 1'b0 ;
  assign n8088 = n5788 | n8087 ;
  assign n8089 = n4349 ^ n559 ^ 1'b0 ;
  assign n8090 = ~n474 & n8089 ;
  assign n8091 = ~n4259 & n8090 ;
  assign n8092 = n8091 ^ n5151 ^ 1'b0 ;
  assign n8093 = n4703 ^ n1898 ^ 1'b0 ;
  assign n8094 = n2498 & ~n4362 ;
  assign n8095 = ~n8093 & n8094 ;
  assign n8102 = n6309 ^ n2959 ^ n1976 ;
  assign n8103 = n8102 ^ n6951 ^ n3407 ;
  assign n8101 = n2365 ^ n708 ^ n508 ;
  assign n8096 = n2271 & n2726 ;
  assign n8097 = n8096 ^ x99 ^ 1'b0 ;
  assign n8098 = n6896 & ~n8097 ;
  assign n8099 = n8098 ^ n3904 ^ 1'b0 ;
  assign n8100 = n8099 ^ n3715 ^ n2592 ;
  assign n8104 = n8103 ^ n8101 ^ n8100 ;
  assign n8105 = n8104 ^ n6697 ^ 1'b0 ;
  assign n8107 = n2438 | n3307 ;
  assign n8108 = n8107 ^ n4165 ^ 1'b0 ;
  assign n8106 = n6297 ^ n3699 ^ 1'b0 ;
  assign n8109 = n8108 ^ n8106 ^ n2757 ;
  assign n8110 = n1808 & n8109 ;
  assign n8111 = n608 & n2693 ;
  assign n8112 = n2008 & n8111 ;
  assign n8113 = n3845 & n8112 ;
  assign n8114 = n802 ^ n506 ^ n462 ;
  assign n8115 = n8113 | n8114 ;
  assign n8116 = n6287 ^ n6029 ^ n3467 ;
  assign n8117 = n2590 | n5936 ;
  assign n8118 = n1441 | n2298 ;
  assign n8119 = n8117 | n8118 ;
  assign n8120 = n8119 ^ n2098 ^ 1'b0 ;
  assign n8121 = n8116 & n8120 ;
  assign n8122 = ~n1427 & n8121 ;
  assign n8123 = n8122 ^ n626 ^ 1'b0 ;
  assign n8124 = n139 & ~n5618 ;
  assign n8125 = n287 & n5909 ;
  assign n8126 = ~n266 & n8125 ;
  assign n8127 = n6779 ^ n4182 ^ 1'b0 ;
  assign n8128 = n8126 | n8127 ;
  assign n8129 = n7817 | n8112 ;
  assign n8131 = ( n1051 & n2744 ) | ( n1051 & ~n2856 ) | ( n2744 & ~n2856 ) ;
  assign n8130 = ( ~n3254 & n4941 ) | ( ~n3254 & n6326 ) | ( n4941 & n6326 ) ;
  assign n8132 = n8131 ^ n8130 ^ 1'b0 ;
  assign n8133 = n549 & ~n7239 ;
  assign n8134 = ( n1645 & n3351 ) | ( n1645 & n8133 ) | ( n3351 & n8133 ) ;
  assign n8135 = x18 & ~n4203 ;
  assign n8136 = n2473 & ~n8135 ;
  assign n8137 = n8134 & n8136 ;
  assign n8138 = n4160 ^ n3304 ^ 1'b0 ;
  assign n8139 = n3838 & ~n8138 ;
  assign n8140 = n8139 ^ n7214 ^ n4653 ;
  assign n8142 = n3468 | n3504 ;
  assign n8141 = n4470 ^ n1426 ^ x75 ;
  assign n8143 = n8142 ^ n8141 ^ n2670 ;
  assign n8144 = n1754 | n8143 ;
  assign n8145 = n4373 | n8144 ;
  assign n8146 = ~n533 & n5997 ;
  assign n8147 = n2838 & ~n5570 ;
  assign n8148 = n8147 ^ n214 ^ 1'b0 ;
  assign n8149 = n8148 ^ n3980 ^ n1485 ;
  assign n8153 = x7 & ~n770 ;
  assign n8154 = x37 & n8153 ;
  assign n8155 = n8154 ^ n3790 ^ n2522 ;
  assign n8150 = n848 | n4094 ;
  assign n8151 = n8150 ^ n6605 ^ 1'b0 ;
  assign n8152 = n8151 ^ n5746 ^ n2122 ;
  assign n8156 = n8155 ^ n8152 ^ n2840 ;
  assign n8157 = n6336 ^ n6266 ^ n3686 ;
  assign n8158 = ( n2177 & n2465 ) | ( n2177 & ~n6853 ) | ( n2465 & ~n6853 ) ;
  assign n8159 = n8158 ^ n1105 ^ 1'b0 ;
  assign n8160 = n2623 & ~n6639 ;
  assign n8161 = ( n1097 & ~n4279 ) | ( n1097 & n6858 ) | ( ~n4279 & n6858 ) ;
  assign n8162 = n2082 | n2141 ;
  assign n8163 = n8162 ^ n7891 ^ n6828 ;
  assign n8164 = n8163 ^ n6794 ^ n6654 ;
  assign n8165 = n4302 & ~n4327 ;
  assign n8166 = n8165 ^ n2659 ^ 1'b0 ;
  assign n8167 = ~n1897 & n8166 ;
  assign n8168 = n8164 & n8167 ;
  assign n8169 = n1718 | n4598 ;
  assign n8170 = n8169 ^ n1688 ^ 1'b0 ;
  assign n8171 = n3896 & ~n4113 ;
  assign n8172 = ~n851 & n8171 ;
  assign n8173 = ( n2366 & n8170 ) | ( n2366 & n8172 ) | ( n8170 & n8172 ) ;
  assign n8174 = n7018 ^ n984 ^ 1'b0 ;
  assign n8175 = n8173 | n8174 ;
  assign n8176 = n2624 ^ n821 ^ 1'b0 ;
  assign n8177 = ~n7270 & n8176 ;
  assign n8178 = n5473 & n6168 ;
  assign n8179 = n1243 & n1629 ;
  assign n8180 = ( ~n2590 & n8178 ) | ( ~n2590 & n8179 ) | ( n8178 & n8179 ) ;
  assign n8181 = ( ~n1410 & n2557 ) | ( ~n1410 & n4524 ) | ( n2557 & n4524 ) ;
  assign n8182 = n3503 & n6016 ;
  assign n8183 = n1211 & ~n6624 ;
  assign n8184 = n3121 ^ n267 ^ 1'b0 ;
  assign n8185 = n3267 | n8184 ;
  assign n8186 = x19 & n2292 ;
  assign n8187 = n8185 & n8186 ;
  assign n8188 = n219 | n1972 ;
  assign n8189 = n8188 ^ n1279 ^ 1'b0 ;
  assign n8190 = n2483 & n8189 ;
  assign n8191 = n8190 ^ n2790 ^ 1'b0 ;
  assign n8192 = n4313 ^ n1314 ^ n871 ;
  assign n8193 = n5129 | n8192 ;
  assign n8194 = n871 ^ x121 ^ 1'b0 ;
  assign n8195 = n2452 & n3597 ;
  assign n8196 = n8195 ^ n370 ^ 1'b0 ;
  assign n8197 = ~n613 & n1058 ;
  assign n8198 = n8196 & n8197 ;
  assign n8199 = ( ~n4623 & n5225 ) | ( ~n4623 & n8198 ) | ( n5225 & n8198 ) ;
  assign n8200 = n8199 ^ n2352 ^ n1852 ;
  assign n8201 = ( n7933 & ~n8194 ) | ( n7933 & n8200 ) | ( ~n8194 & n8200 ) ;
  assign n8202 = ( n2874 & ~n6131 ) | ( n2874 & n6151 ) | ( ~n6131 & n6151 ) ;
  assign n8203 = n8202 ^ n3935 ^ n2915 ;
  assign n8204 = n186 | n3364 ;
  assign n8205 = n2693 | n8204 ;
  assign n8206 = ( n798 & n4346 ) | ( n798 & ~n8205 ) | ( n4346 & ~n8205 ) ;
  assign n8207 = ( n1175 & n4175 ) | ( n1175 & n8206 ) | ( n4175 & n8206 ) ;
  assign n8208 = n7727 ^ n4493 ^ n3986 ;
  assign n8209 = n5872 ^ n4520 ^ 1'b0 ;
  assign n8210 = n6046 & n8209 ;
  assign n8211 = n3631 ^ n898 ^ 1'b0 ;
  assign n8214 = n3703 ^ n491 ^ 1'b0 ;
  assign n8215 = x26 | n8214 ;
  assign n8212 = n899 & ~n4800 ;
  assign n8213 = n2682 | n8212 ;
  assign n8216 = n8215 ^ n8213 ^ 1'b0 ;
  assign n8217 = ( n1143 & ~n3063 ) | ( n1143 & n6073 ) | ( ~n3063 & n6073 ) ;
  assign n8218 = ~n3189 & n7738 ;
  assign n8219 = ~n5519 & n8218 ;
  assign n8225 = n2860 ^ n2515 ^ 1'b0 ;
  assign n8226 = n136 & n8225 ;
  assign n8227 = n8226 ^ n1266 ^ 1'b0 ;
  assign n8228 = n1242 | n2324 ;
  assign n8229 = ( n659 & ~n8227 ) | ( n659 & n8228 ) | ( ~n8227 & n8228 ) ;
  assign n8221 = ~n497 & n781 ;
  assign n8222 = n8221 ^ n1846 ^ 1'b0 ;
  assign n8220 = ( n1065 & n2093 ) | ( n1065 & ~n3237 ) | ( n2093 & ~n3237 ) ;
  assign n8223 = n8222 ^ n8220 ^ n4998 ;
  assign n8224 = ( n481 & n1762 ) | ( n481 & n8223 ) | ( n1762 & n8223 ) ;
  assign n8230 = n8229 ^ n8224 ^ 1'b0 ;
  assign n8231 = n858 & n8230 ;
  assign n8232 = n1164 & n3377 ;
  assign n8233 = n612 & n6126 ;
  assign n8234 = ( ~n3642 & n3988 ) | ( ~n3642 & n7193 ) | ( n3988 & n7193 ) ;
  assign n8235 = ( n837 & n2932 ) | ( n837 & ~n8234 ) | ( n2932 & ~n8234 ) ;
  assign n8236 = n1564 & ~n4376 ;
  assign n8237 = n8236 ^ n6296 ^ 1'b0 ;
  assign n8238 = n4180 ^ n934 ^ 1'b0 ;
  assign n8239 = n8238 ^ n7757 ^ 1'b0 ;
  assign n8240 = n2199 ^ n1784 ^ 1'b0 ;
  assign n8241 = n4391 | n7695 ;
  assign n8242 = n8240 | n8241 ;
  assign n8243 = ( ~n219 & n4022 ) | ( ~n219 & n4882 ) | ( n4022 & n4882 ) ;
  assign n8244 = n3741 & ~n4693 ;
  assign n8245 = n8243 & n8244 ;
  assign n8246 = n2457 & ~n4313 ;
  assign n8247 = ~n580 & n8246 ;
  assign n8248 = n4594 ^ n3158 ^ 1'b0 ;
  assign n8249 = ~n3020 & n8248 ;
  assign n8250 = ( ~n4201 & n5052 ) | ( ~n4201 & n8249 ) | ( n5052 & n8249 ) ;
  assign n8251 = n6306 | n8250 ;
  assign n8252 = n8251 ^ n7743 ^ 1'b0 ;
  assign n8253 = n5005 | n8252 ;
  assign n8254 = ( n598 & ~n2425 ) | ( n598 & n8253 ) | ( ~n2425 & n8253 ) ;
  assign n8255 = ( n415 & n1302 ) | ( n415 & n2855 ) | ( n1302 & n2855 ) ;
  assign n8256 = n8255 ^ n1326 ^ 1'b0 ;
  assign n8257 = n7918 ^ n1518 ^ 1'b0 ;
  assign n8258 = n556 | n8257 ;
  assign n8259 = n8258 ^ n5522 ^ 1'b0 ;
  assign n8260 = ~n8256 & n8259 ;
  assign n8261 = n8260 ^ n1454 ^ 1'b0 ;
  assign n8262 = n4430 & ~n6494 ;
  assign n8263 = n1339 & n8262 ;
  assign n8264 = ~n535 & n8263 ;
  assign n8265 = n754 ^ x116 ^ 1'b0 ;
  assign n8266 = n2163 & n8265 ;
  assign n8267 = n8264 & n8266 ;
  assign n8268 = n4807 ^ n1490 ^ 1'b0 ;
  assign n8269 = ~n4541 & n8268 ;
  assign n8270 = n6739 ^ n4862 ^ 1'b0 ;
  assign n8271 = ( n1481 & n5373 ) | ( n1481 & n7701 ) | ( n5373 & n7701 ) ;
  assign n8272 = n6016 ^ n4859 ^ n3437 ;
  assign n8273 = n8272 ^ n5550 ^ n1736 ;
  assign n8274 = n8273 ^ n1852 ^ n972 ;
  assign n8275 = n415 & n3099 ;
  assign n8276 = ( ~n1541 & n8274 ) | ( ~n1541 & n8275 ) | ( n8274 & n8275 ) ;
  assign n8277 = ( n1916 & ~n7640 ) | ( n1916 & n8276 ) | ( ~n7640 & n8276 ) ;
  assign n8282 = n655 & n734 ;
  assign n8283 = n8282 ^ n3617 ^ n650 ;
  assign n8278 = n2631 ^ n2232 ^ 1'b0 ;
  assign n8279 = n1302 | n8278 ;
  assign n8280 = n8279 ^ n1244 ^ 1'b0 ;
  assign n8281 = ~x59 & n8280 ;
  assign n8284 = n8283 ^ n8281 ^ 1'b0 ;
  assign n8285 = n5414 ^ n1283 ^ 1'b0 ;
  assign n8286 = ~n1384 & n8285 ;
  assign n8288 = n4711 ^ n4401 ^ n1617 ;
  assign n8287 = n2751 ^ n1810 ^ n637 ;
  assign n8289 = n8288 ^ n8287 ^ n2048 ;
  assign n8290 = n1759 & ~n7459 ;
  assign n8291 = ( n3431 & n8289 ) | ( n3431 & n8290 ) | ( n8289 & n8290 ) ;
  assign n8292 = n6374 ^ n3389 ^ 1'b0 ;
  assign n8293 = ~n742 & n8292 ;
  assign n8294 = n3640 & n8293 ;
  assign n8295 = ( n272 & n4539 ) | ( n272 & n8294 ) | ( n4539 & n8294 ) ;
  assign n8300 = n5161 ^ n1515 ^ 1'b0 ;
  assign n8301 = n1818 & ~n8300 ;
  assign n8296 = n4791 & ~n7180 ;
  assign n8297 = ~n531 & n5748 ;
  assign n8298 = n8297 ^ n2402 ^ n2296 ;
  assign n8299 = n8296 & ~n8298 ;
  assign n8302 = n8301 ^ n8299 ^ 1'b0 ;
  assign n8303 = n5600 ^ n1515 ^ 1'b0 ;
  assign n8304 = n7379 ^ n262 ^ 1'b0 ;
  assign n8305 = ~n5040 & n8304 ;
  assign n8306 = ( n1490 & n3283 ) | ( n1490 & ~n8305 ) | ( n3283 & ~n8305 ) ;
  assign n8308 = ~n2116 & n2329 ;
  assign n8307 = n222 & ~n3384 ;
  assign n8309 = n8308 ^ n8307 ^ 1'b0 ;
  assign n8310 = n1765 | n3509 ;
  assign n8311 = ( n3688 & ~n8240 ) | ( n3688 & n8310 ) | ( ~n8240 & n8310 ) ;
  assign n8312 = ( n680 & n6366 ) | ( n680 & n8311 ) | ( n6366 & n8311 ) ;
  assign n8314 = n5739 ^ n1038 ^ n141 ;
  assign n8315 = n2170 | n8314 ;
  assign n8316 = n143 | n8315 ;
  assign n8313 = ~n5889 & n6059 ;
  assign n8317 = n8316 ^ n8313 ^ 1'b0 ;
  assign n8318 = n1162 & ~n5430 ;
  assign n8319 = n3346 & ~n4127 ;
  assign n8320 = n5723 & n8319 ;
  assign n8321 = n2660 & ~n8320 ;
  assign n8322 = n8318 & n8321 ;
  assign n8326 = n2504 & ~n5181 ;
  assign n8323 = n5400 ^ n4157 ^ n4067 ;
  assign n8324 = n8323 ^ n5051 ^ n985 ;
  assign n8325 = ~n3389 & n8324 ;
  assign n8327 = n8326 ^ n8325 ^ 1'b0 ;
  assign n8328 = n2027 | n3071 ;
  assign n8329 = n6226 ^ n2509 ^ n1048 ;
  assign n8330 = n8329 ^ n4825 ^ 1'b0 ;
  assign n8331 = n2687 ^ n2499 ^ n1754 ;
  assign n8332 = n6008 & ~n8331 ;
  assign n8333 = ~n2487 & n8332 ;
  assign n8335 = n1171 | n1514 ;
  assign n8336 = n6559 | n8335 ;
  assign n8334 = n8215 ^ n2315 ^ n230 ;
  assign n8337 = n8336 ^ n8334 ^ n4921 ;
  assign n8338 = n4703 & ~n7518 ;
  assign n8339 = n4588 & ~n8288 ;
  assign n8340 = n4949 ^ n4457 ^ n3369 ;
  assign n8341 = n2243 & ~n8340 ;
  assign n8342 = n4099 ^ n2009 ^ n984 ;
  assign n8343 = n6658 ^ n182 ^ 1'b0 ;
  assign n8344 = n7924 ^ n7515 ^ 1'b0 ;
  assign n8345 = n1110 ^ n915 ^ 1'b0 ;
  assign n8346 = n3691 & ~n8345 ;
  assign n8347 = n7735 & n8346 ;
  assign n8348 = ~n8049 & n8347 ;
  assign n8349 = n6191 ^ n3649 ^ 1'b0 ;
  assign n8353 = ~n514 & n2273 ;
  assign n8354 = n8353 ^ n2090 ^ 1'b0 ;
  assign n8350 = n7838 ^ n3982 ^ n3670 ;
  assign n8351 = ( ~n245 & n2903 ) | ( ~n245 & n3536 ) | ( n2903 & n3536 ) ;
  assign n8352 = ( n3934 & n8350 ) | ( n3934 & n8351 ) | ( n8350 & n8351 ) ;
  assign n8355 = n8354 ^ n8352 ^ n555 ;
  assign n8356 = n2369 & ~n6136 ;
  assign n8357 = n806 & n8356 ;
  assign n8358 = n3778 & ~n8043 ;
  assign n8359 = n8358 ^ n883 ^ 1'b0 ;
  assign n8360 = n8359 ^ n8064 ^ n620 ;
  assign n8361 = n4107 ^ n3688 ^ 1'b0 ;
  assign n8362 = n8361 ^ n4602 ^ 1'b0 ;
  assign n8363 = x122 & ~n2113 ;
  assign n8364 = n2104 & n8363 ;
  assign n8365 = n1250 & n1283 ;
  assign n8366 = n7449 ^ n3685 ^ n1770 ;
  assign n8367 = n891 & ~n2438 ;
  assign n8368 = n8366 & n8367 ;
  assign n8369 = ( n1571 & n3609 ) | ( n1571 & n8368 ) | ( n3609 & n8368 ) ;
  assign n8370 = n5076 ^ n2451 ^ n2056 ;
  assign n8371 = n8370 ^ n1449 ^ 1'b0 ;
  assign n8372 = n8371 ^ n1034 ^ 1'b0 ;
  assign n8373 = n2000 & ~n8071 ;
  assign n8374 = n8373 ^ n1044 ^ 1'b0 ;
  assign n8375 = n4841 ^ n4406 ^ 1'b0 ;
  assign n8376 = ~n4689 & n8375 ;
  assign n8377 = ~n8374 & n8376 ;
  assign n8378 = n2018 & n7639 ;
  assign n8379 = n8378 ^ n636 ^ 1'b0 ;
  assign n8380 = ( n525 & ~n3260 ) | ( n525 & n8379 ) | ( ~n3260 & n8379 ) ;
  assign n8382 = n2359 & ~n5963 ;
  assign n8381 = ( n2401 & n2730 ) | ( n2401 & ~n3144 ) | ( n2730 & ~n3144 ) ;
  assign n8383 = n8382 ^ n8381 ^ n5101 ;
  assign n8384 = n6151 | n6312 ;
  assign n8385 = n5102 | n8384 ;
  assign n8386 = ~n307 & n8249 ;
  assign n8387 = ~n5689 & n8386 ;
  assign n8388 = n8387 ^ n872 ^ 1'b0 ;
  assign n8389 = ~n3479 & n3561 ;
  assign n8390 = ~n7775 & n8389 ;
  assign n8391 = n531 & ~n8390 ;
  assign n8392 = n8391 ^ n5807 ^ 1'b0 ;
  assign n8395 = n3703 ^ n897 ^ 1'b0 ;
  assign n8396 = n1150 & ~n8395 ;
  assign n8393 = n2948 ^ n2794 ^ n2061 ;
  assign n8394 = ( n2891 & n6532 ) | ( n2891 & n8393 ) | ( n6532 & n8393 ) ;
  assign n8397 = n8396 ^ n8394 ^ n3418 ;
  assign n8399 = n4492 ^ n2871 ^ 1'b0 ;
  assign n8398 = n1624 | n6600 ;
  assign n8400 = n8399 ^ n8398 ^ 1'b0 ;
  assign n8401 = n751 & n8400 ;
  assign n8402 = n8401 ^ n1688 ^ 1'b0 ;
  assign n8403 = ~n8397 & n8402 ;
  assign n8404 = ( n6590 & ~n8392 ) | ( n6590 & n8403 ) | ( ~n8392 & n8403 ) ;
  assign n8405 = n7705 ^ n1671 ^ 1'b0 ;
  assign n8407 = n3489 ^ x35 ^ 1'b0 ;
  assign n8406 = n7494 ^ n1585 ^ 1'b0 ;
  assign n8408 = n8407 ^ n8406 ^ 1'b0 ;
  assign n8409 = n826 & ~n4131 ;
  assign n8410 = n3715 & n8409 ;
  assign n8411 = n1321 ^ x115 ^ 1'b0 ;
  assign n8412 = ( n2102 & n8410 ) | ( n2102 & ~n8411 ) | ( n8410 & ~n8411 ) ;
  assign n8413 = n652 & n7304 ;
  assign n8414 = ( n567 & n4443 ) | ( n567 & n8275 ) | ( n4443 & n8275 ) ;
  assign n8415 = n8413 | n8414 ;
  assign n8416 = n1258 & ~n3215 ;
  assign n8417 = ( n1178 & n7842 ) | ( n1178 & n8416 ) | ( n7842 & n8416 ) ;
  assign n8418 = ~n8415 & n8417 ;
  assign n8419 = n8418 ^ n6086 ^ 1'b0 ;
  assign n8420 = n912 & ~n3637 ;
  assign n8421 = n5633 & n8420 ;
  assign n8423 = n4802 ^ x3 ^ 1'b0 ;
  assign n8424 = n1538 & n3218 ;
  assign n8425 = ~n6443 & n8424 ;
  assign n8426 = ~n8423 & n8425 ;
  assign n8422 = ( ~n1573 & n1935 ) | ( ~n1573 & n4854 ) | ( n1935 & n4854 ) ;
  assign n8427 = n8426 ^ n8422 ^ n2356 ;
  assign n8428 = n4587 & ~n8427 ;
  assign n8429 = n8428 ^ n1535 ^ 1'b0 ;
  assign n8430 = n6137 & n8429 ;
  assign n8431 = ( n3885 & n4403 ) | ( n3885 & ~n4423 ) | ( n4403 & ~n4423 ) ;
  assign n8432 = n1165 & n3895 ;
  assign n8433 = ( x99 & ~n8309 ) | ( x99 & n8432 ) | ( ~n8309 & n8432 ) ;
  assign n8434 = n7812 ^ n3311 ^ 1'b0 ;
  assign n8435 = n7033 ^ n243 ^ 1'b0 ;
  assign n8436 = n7998 & n8435 ;
  assign n8437 = n8436 ^ n7785 ^ n4198 ;
  assign n8438 = n6697 ^ n1598 ^ 1'b0 ;
  assign n8444 = n3979 & n4063 ;
  assign n8439 = n239 ^ n149 ^ 1'b0 ;
  assign n8441 = ( ~n3047 & n4754 ) | ( ~n3047 & n8170 ) | ( n4754 & n8170 ) ;
  assign n8440 = ( n1359 & ~n6621 ) | ( n1359 & n7366 ) | ( ~n6621 & n7366 ) ;
  assign n8442 = n8441 ^ n8440 ^ n4376 ;
  assign n8443 = n8439 & ~n8442 ;
  assign n8445 = n8444 ^ n8443 ^ 1'b0 ;
  assign n8449 = n1586 & ~n2211 ;
  assign n8450 = n338 & n8449 ;
  assign n8448 = ~n3018 & n5697 ;
  assign n8451 = n8450 ^ n8448 ^ 1'b0 ;
  assign n8452 = n2328 | n8451 ;
  assign n8447 = n6304 & n6517 ;
  assign n8446 = n7731 ^ n7423 ^ n2242 ;
  assign n8453 = n8452 ^ n8447 ^ n8446 ;
  assign n8454 = n2598 ^ n1454 ^ x106 ;
  assign n8455 = n4261 ^ n3633 ^ n2536 ;
  assign n8456 = ( n5418 & n8454 ) | ( n5418 & ~n8455 ) | ( n8454 & ~n8455 ) ;
  assign n8457 = n1986 | n2876 ;
  assign n8458 = ( ~n3656 & n7604 ) | ( ~n3656 & n8457 ) | ( n7604 & n8457 ) ;
  assign n8459 = n2662 | n5746 ;
  assign n8460 = n8459 ^ n4087 ^ 1'b0 ;
  assign n8461 = ( n357 & n2334 ) | ( n357 & n8460 ) | ( n2334 & n8460 ) ;
  assign n8462 = n6133 ^ n3766 ^ 1'b0 ;
  assign n8463 = n3642 ^ n1117 ^ 1'b0 ;
  assign n8464 = n1468 & ~n8463 ;
  assign n8465 = n849 | n3587 ;
  assign n8466 = n8464 | n8465 ;
  assign n8471 = n5014 ^ n4221 ^ n797 ;
  assign n8469 = n724 | n2378 ;
  assign n8467 = n2191 & n5347 ;
  assign n8468 = n8467 ^ n2632 ^ 1'b0 ;
  assign n8470 = n8469 ^ n8468 ^ 1'b0 ;
  assign n8472 = n8471 ^ n8470 ^ n4644 ;
  assign n8473 = n4899 & n6038 ;
  assign n8474 = n997 ^ n901 ^ 1'b0 ;
  assign n8475 = ( n885 & n1217 ) | ( n885 & n3413 ) | ( n1217 & n3413 ) ;
  assign n8476 = n8475 ^ n3345 ^ 1'b0 ;
  assign n8477 = ( n490 & n1769 ) | ( n490 & n8476 ) | ( n1769 & n8476 ) ;
  assign n8478 = ( n930 & ~n8474 ) | ( n930 & n8477 ) | ( ~n8474 & n8477 ) ;
  assign n8479 = n817 & n8478 ;
  assign n8480 = ( n3154 & n8473 ) | ( n3154 & n8479 ) | ( n8473 & n8479 ) ;
  assign n8481 = n2654 ^ n1320 ^ 1'b0 ;
  assign n8482 = n692 | n8481 ;
  assign n8483 = ~n3137 & n8482 ;
  assign n8484 = n2895 & ~n6781 ;
  assign n8485 = n8484 ^ n5655 ^ 1'b0 ;
  assign n8486 = n912 & n3738 ;
  assign n8487 = n8486 ^ n3850 ^ 1'b0 ;
  assign n8488 = ~n5714 & n7855 ;
  assign n8489 = n8487 & n8488 ;
  assign n8490 = ( n375 & n1060 ) | ( n375 & n5248 ) | ( n1060 & n5248 ) ;
  assign n8491 = n8490 ^ n2151 ^ 1'b0 ;
  assign n8492 = ~n6065 & n8491 ;
  assign n8493 = n8492 ^ n4367 ^ n1517 ;
  assign n8494 = n8493 ^ n3869 ^ n2621 ;
  assign n8495 = n239 & ~n3869 ;
  assign n8496 = n1339 & n7236 ;
  assign n8497 = ~n1229 & n2098 ;
  assign n8498 = n3306 & ~n8497 ;
  assign n8499 = n8496 & n8498 ;
  assign n8500 = ( n6714 & ~n6780 ) | ( n6714 & n8499 ) | ( ~n6780 & n8499 ) ;
  assign n8501 = n1447 & ~n5525 ;
  assign n8502 = n2206 & n8113 ;
  assign n8503 = n8502 ^ n5773 ^ 1'b0 ;
  assign n8504 = n2644 ^ n599 ^ 1'b0 ;
  assign n8505 = n4179 & ~n8504 ;
  assign n8506 = n8505 ^ n5093 ^ n188 ;
  assign n8507 = ~n2400 & n8506 ;
  assign n8518 = n209 & n3211 ;
  assign n8519 = ~n2232 & n8518 ;
  assign n8508 = n5530 ^ n4611 ^ n964 ;
  assign n8509 = n1139 & n2781 ;
  assign n8510 = n8509 ^ n2277 ^ 1'b0 ;
  assign n8511 = ~n831 & n8510 ;
  assign n8512 = n915 & n8511 ;
  assign n8513 = n1541 & n4976 ;
  assign n8514 = n3772 & n8513 ;
  assign n8515 = n8514 ^ x7 ^ 1'b0 ;
  assign n8516 = n8512 | n8515 ;
  assign n8517 = ( n1564 & n8508 ) | ( n1564 & ~n8516 ) | ( n8508 & ~n8516 ) ;
  assign n8520 = n8519 ^ n8517 ^ 1'b0 ;
  assign n8521 = ( n3719 & ~n4094 ) | ( n3719 & n8041 ) | ( ~n4094 & n8041 ) ;
  assign n8522 = n7026 ^ n1886 ^ 1'b0 ;
  assign n8523 = ( n260 & ~n570 ) | ( n260 & n8522 ) | ( ~n570 & n8522 ) ;
  assign n8524 = n1704 | n4546 ;
  assign n8525 = n8524 ^ n4356 ^ 1'b0 ;
  assign n8526 = n1287 & n5286 ;
  assign n8527 = ~n8525 & n8526 ;
  assign n8528 = n3795 ^ n2883 ^ n462 ;
  assign n8529 = n8528 ^ n6382 ^ n4605 ;
  assign n8530 = n8529 ^ n6838 ^ n3321 ;
  assign n8531 = n8396 ^ n7256 ^ 1'b0 ;
  assign n8532 = x108 & ~n8531 ;
  assign n8537 = n2340 & ~n7110 ;
  assign n8538 = ~n5209 & n8537 ;
  assign n8533 = n2029 ^ n457 ^ 1'b0 ;
  assign n8534 = ~n3770 & n8533 ;
  assign n8535 = n3197 | n8534 ;
  assign n8536 = n8535 ^ n6164 ^ n5030 ;
  assign n8539 = n8538 ^ n8536 ^ n7344 ;
  assign n8540 = n1339 & n4417 ;
  assign n8541 = ~n5764 & n8540 ;
  assign n8542 = n6311 | n8541 ;
  assign n8543 = n7100 & n8542 ;
  assign n8544 = n7889 ^ n5492 ^ 1'b0 ;
  assign n8545 = n306 | n3686 ;
  assign n8546 = n5298 ^ n3262 ^ 1'b0 ;
  assign n8547 = n6150 ^ n1405 ^ 1'b0 ;
  assign n8548 = n8546 & ~n8547 ;
  assign n8549 = ~n1590 & n8548 ;
  assign n8550 = ( n4166 & n8545 ) | ( n4166 & n8549 ) | ( n8545 & n8549 ) ;
  assign n8551 = n968 ^ n826 ^ 1'b0 ;
  assign n8552 = ~n1715 & n8551 ;
  assign n8553 = n8552 ^ n4014 ^ 1'b0 ;
  assign n8554 = n7929 | n8553 ;
  assign n8555 = ( n3178 & ~n5122 ) | ( n3178 & n8554 ) | ( ~n5122 & n8554 ) ;
  assign n8556 = n8555 ^ n4370 ^ 1'b0 ;
  assign n8557 = n1279 & n8556 ;
  assign n8558 = n8557 ^ n6105 ^ n3881 ;
  assign n8563 = n5597 ^ n1756 ^ 1'b0 ;
  assign n8564 = n8563 ^ n3200 ^ n2309 ;
  assign n8559 = n2375 & ~n2789 ;
  assign n8560 = n8559 ^ n1511 ^ 1'b0 ;
  assign n8561 = ( ~n3378 & n6118 ) | ( ~n3378 & n8560 ) | ( n6118 & n8560 ) ;
  assign n8562 = n8561 ^ n1011 ^ 1'b0 ;
  assign n8565 = n8564 ^ n8562 ^ n3592 ;
  assign n8566 = x120 & ~n1460 ;
  assign n8567 = n5370 ^ n3700 ^ n1366 ;
  assign n8568 = ( n737 & n8566 ) | ( n737 & n8567 ) | ( n8566 & n8567 ) ;
  assign n8569 = n2101 & n8330 ;
  assign n8570 = n8569 ^ n7200 ^ 1'b0 ;
  assign n8571 = n2400 & ~n2847 ;
  assign n8572 = n2095 ^ x31 ^ 1'b0 ;
  assign n8573 = ~n1316 & n8049 ;
  assign n8574 = ( n8571 & n8572 ) | ( n8571 & ~n8573 ) | ( n8572 & ~n8573 ) ;
  assign n8575 = ( n2092 & n3894 ) | ( n2092 & ~n6954 ) | ( n3894 & ~n6954 ) ;
  assign n8576 = n365 & ~n1741 ;
  assign n8577 = n6207 ^ n2701 ^ n813 ;
  assign n8578 = ( n8414 & n8576 ) | ( n8414 & ~n8577 ) | ( n8576 & ~n8577 ) ;
  assign n8579 = n6635 ^ n3365 ^ n2003 ;
  assign n8580 = ( n5353 & n7795 ) | ( n5353 & n8579 ) | ( n7795 & n8579 ) ;
  assign n8581 = ( n3971 & n8253 ) | ( n3971 & ~n8580 ) | ( n8253 & ~n8580 ) ;
  assign n8582 = n7457 ^ n3191 ^ 1'b0 ;
  assign n8583 = n8582 ^ n7373 ^ 1'b0 ;
  assign n8584 = n1944 ^ n1588 ^ 1'b0 ;
  assign n8585 = n182 | n7096 ;
  assign n8586 = n8585 ^ n3722 ^ 1'b0 ;
  assign n8587 = ( n612 & n8584 ) | ( n612 & n8586 ) | ( n8584 & n8586 ) ;
  assign n8590 = ( n2377 & n2417 ) | ( n2377 & n5615 ) | ( n2417 & n5615 ) ;
  assign n8588 = ( n984 & n3718 ) | ( n984 & n4390 ) | ( n3718 & n4390 ) ;
  assign n8589 = n8588 ^ n6838 ^ n6670 ;
  assign n8591 = n8590 ^ n8589 ^ 1'b0 ;
  assign n8592 = n2770 ^ n2007 ^ 1'b0 ;
  assign n8593 = n8592 ^ n2423 ^ n1622 ;
  assign n8594 = ~n2715 & n6241 ;
  assign n8595 = ~n7756 & n8594 ;
  assign n8596 = n1290 ^ n1206 ^ n552 ;
  assign n8597 = n8596 ^ n3051 ^ 1'b0 ;
  assign n8598 = n8597 ^ n8134 ^ n7987 ;
  assign n8599 = n3998 ^ n2681 ^ 1'b0 ;
  assign n8600 = ~n1063 & n8599 ;
  assign n8601 = n8600 ^ n1876 ^ 1'b0 ;
  assign n8602 = n5870 ^ x117 ^ 1'b0 ;
  assign n8603 = ~n3939 & n8602 ;
  assign n8604 = n8603 ^ n2072 ^ 1'b0 ;
  assign n8605 = n8601 | n8604 ;
  assign n8606 = n7024 ^ n296 ^ 1'b0 ;
  assign n8607 = ~n2346 & n4645 ;
  assign n8608 = n8606 & n8607 ;
  assign n8609 = n4167 ^ x120 ^ 1'b0 ;
  assign n8610 = n7145 | n8277 ;
  assign n8611 = n5121 ^ n563 ^ n447 ;
  assign n8612 = n216 & n8611 ;
  assign n8613 = n6821 & n8612 ;
  assign n8614 = n2036 & n7481 ;
  assign n8615 = n8614 ^ n1184 ^ 1'b0 ;
  assign n8616 = n8615 ^ n7698 ^ 1'b0 ;
  assign n8617 = n2764 & ~n8100 ;
  assign n8618 = ~n8616 & n8617 ;
  assign n8619 = n7853 ^ n2475 ^ n831 ;
  assign n8623 = n1590 & n1730 ;
  assign n8621 = ( ~n218 & n228 ) | ( ~n218 & n641 ) | ( n228 & n641 ) ;
  assign n8620 = ~n2179 & n5386 ;
  assign n8622 = n8621 ^ n8620 ^ n6368 ;
  assign n8624 = n8623 ^ n8622 ^ n3134 ;
  assign n8625 = n689 ^ x18 ^ 1'b0 ;
  assign n8626 = n771 & n8625 ;
  assign n8627 = n1718 ^ n1137 ^ 1'b0 ;
  assign n8628 = n2842 & n8627 ;
  assign n8629 = n2017 & n8628 ;
  assign n8630 = ( n1212 & n1654 ) | ( n1212 & ~n8629 ) | ( n1654 & ~n8629 ) ;
  assign n8631 = n8305 & ~n8630 ;
  assign n8632 = n8631 ^ n2532 ^ 1'b0 ;
  assign n8633 = n3314 & ~n3827 ;
  assign n8634 = n8633 ^ n4361 ^ 1'b0 ;
  assign n8635 = n620 | n8634 ;
  assign n8636 = n8632 | n8635 ;
  assign n8637 = n8636 ^ n6111 ^ 1'b0 ;
  assign n8638 = ( n5124 & ~n8626 ) | ( n5124 & n8637 ) | ( ~n8626 & n8637 ) ;
  assign n8639 = n1326 & n7735 ;
  assign n8640 = n8638 & n8639 ;
  assign n8641 = n8640 ^ n4107 ^ n4048 ;
  assign n8642 = ~n4175 & n8641 ;
  assign n8643 = n8642 ^ n989 ^ 1'b0 ;
  assign n8644 = ( ~n2422 & n7724 ) | ( ~n2422 & n8643 ) | ( n7724 & n8643 ) ;
  assign n8645 = n1797 ^ n1533 ^ n1496 ;
  assign n8646 = n8645 ^ n3722 ^ 1'b0 ;
  assign n8647 = n218 | n8646 ;
  assign n8648 = n390 & n7432 ;
  assign n8649 = n1804 & ~n2704 ;
  assign n8650 = n348 & ~n8649 ;
  assign n8652 = n4766 & n7578 ;
  assign n8653 = ~n2334 & n8652 ;
  assign n8651 = n5118 ^ n2036 ^ n670 ;
  assign n8654 = n8653 ^ n8651 ^ n4957 ;
  assign n8655 = n4227 ^ n4182 ^ n349 ;
  assign n8656 = n8655 ^ n7198 ^ n4374 ;
  assign n8657 = ( n4597 & n4792 ) | ( n4597 & ~n6416 ) | ( n4792 & ~n6416 ) ;
  assign n8658 = ( ~n4127 & n7719 ) | ( ~n4127 & n8482 ) | ( n7719 & n8482 ) ;
  assign n8659 = n3288 ^ n2470 ^ 1'b0 ;
  assign n8660 = ~n3569 & n8659 ;
  assign n8661 = n8660 ^ n6446 ^ n1740 ;
  assign n8662 = ( n486 & ~n1192 ) | ( n486 & n4370 ) | ( ~n1192 & n4370 ) ;
  assign n8663 = n5159 & n8662 ;
  assign n8664 = ~n149 & n8663 ;
  assign n8665 = ( n2177 & ~n8661 ) | ( n2177 & n8664 ) | ( ~n8661 & n8664 ) ;
  assign n8666 = n7367 ^ n3095 ^ 1'b0 ;
  assign n8667 = ( n761 & n1301 ) | ( n761 & n1525 ) | ( n1301 & n1525 ) ;
  assign n8668 = x112 | n3774 ;
  assign n8669 = n1466 | n8668 ;
  assign n8670 = ( n5865 & n6891 ) | ( n5865 & n8669 ) | ( n6891 & n8669 ) ;
  assign n8671 = n3190 ^ n908 ^ 1'b0 ;
  assign n8672 = n1446 & ~n8671 ;
  assign n8673 = n2400 & ~n8672 ;
  assign n8674 = n3036 & ~n3790 ;
  assign n8675 = ( ~n837 & n7741 ) | ( ~n837 & n8080 ) | ( n7741 & n8080 ) ;
  assign n8677 = n1721 | n4137 ;
  assign n8676 = ( ~n838 & n2007 ) | ( ~n838 & n2205 ) | ( n2007 & n2205 ) ;
  assign n8678 = n8677 ^ n8676 ^ n1419 ;
  assign n8679 = n321 & n8678 ;
  assign n8680 = n8675 & ~n8679 ;
  assign n8681 = n6756 ^ n5801 ^ 1'b0 ;
  assign n8682 = ~n6243 & n7469 ;
  assign n8687 = ( x20 & n4322 ) | ( x20 & ~n5016 ) | ( n4322 & ~n5016 ) ;
  assign n8683 = n4703 ^ n3346 ^ n151 ;
  assign n8684 = n3649 & n7954 ;
  assign n8685 = n8683 & n8684 ;
  assign n8686 = n3146 & n8685 ;
  assign n8688 = n8687 ^ n8686 ^ 1'b0 ;
  assign n8691 = n565 | n2738 ;
  assign n8692 = ( n3864 & ~n5463 ) | ( n3864 & n8691 ) | ( ~n5463 & n8691 ) ;
  assign n8689 = n2808 & n8101 ;
  assign n8690 = ~n3712 & n8689 ;
  assign n8693 = n8692 ^ n8690 ^ 1'b0 ;
  assign n8694 = ( n2072 & n2419 ) | ( n2072 & ~n4208 ) | ( n2419 & ~n4208 ) ;
  assign n8695 = n6466 ^ n5028 ^ n3389 ;
  assign n8700 = ~n2004 & n5657 ;
  assign n8701 = n8700 ^ n7819 ^ 1'b0 ;
  assign n8696 = x43 & n781 ;
  assign n8697 = n260 & n8696 ;
  assign n8698 = n3645 | n8697 ;
  assign n8699 = n4136 & ~n8698 ;
  assign n8702 = n8701 ^ n8699 ^ 1'b0 ;
  assign n8703 = n8695 | n8702 ;
  assign n8704 = n8694 | n8703 ;
  assign n8705 = ( n1201 & n3108 ) | ( n1201 & ~n3904 ) | ( n3108 & ~n3904 ) ;
  assign n8706 = n1484 & n8705 ;
  assign n8707 = n8706 ^ n2968 ^ 1'b0 ;
  assign n8708 = ( ~n7104 & n7402 ) | ( ~n7104 & n8707 ) | ( n7402 & n8707 ) ;
  assign n8709 = n266 & n8708 ;
  assign n8710 = n8709 ^ n6611 ^ 1'b0 ;
  assign n8711 = n5377 ^ n796 ^ n294 ;
  assign n8712 = n6301 ^ n4429 ^ 1'b0 ;
  assign n8713 = n751 & n8712 ;
  assign n8714 = n8713 ^ n4752 ^ 1'b0 ;
  assign n8715 = n8711 & ~n8714 ;
  assign n8716 = n8715 ^ n8129 ^ 1'b0 ;
  assign n8717 = ~n2339 & n2415 ;
  assign n8718 = n8192 & n8717 ;
  assign n8719 = n1687 | n8718 ;
  assign n8720 = n7781 ^ n6471 ^ 1'b0 ;
  assign n8721 = ( x47 & n1547 ) | ( x47 & n5432 ) | ( n1547 & n5432 ) ;
  assign n8722 = x59 & ~n7152 ;
  assign n8723 = ( ~n5390 & n8721 ) | ( ~n5390 & n8722 ) | ( n8721 & n8722 ) ;
  assign n8724 = n1256 & ~n2296 ;
  assign n8725 = n2079 | n7613 ;
  assign n8726 = n8724 | n8725 ;
  assign n8727 = n6517 ^ n1887 ^ 1'b0 ;
  assign n8728 = n7425 ^ n3808 ^ 1'b0 ;
  assign n8729 = ~n4005 & n8728 ;
  assign n8730 = ( n1632 & ~n4887 ) | ( n1632 & n8729 ) | ( ~n4887 & n8729 ) ;
  assign n8731 = n8730 ^ n5268 ^ 1'b0 ;
  assign n8732 = n3459 ^ n620 ^ 1'b0 ;
  assign n8733 = ~n8731 & n8732 ;
  assign n8734 = ( ~n2595 & n6842 ) | ( ~n2595 & n8733 ) | ( n6842 & n8733 ) ;
  assign n8735 = ( n4758 & ~n4962 ) | ( n4758 & n5875 ) | ( ~n4962 & n5875 ) ;
  assign n8736 = n8735 ^ n6135 ^ n721 ;
  assign n8743 = n232 | n1258 ;
  assign n8744 = n8743 ^ n4030 ^ 1'b0 ;
  assign n8737 = n4955 ^ n3207 ^ 1'b0 ;
  assign n8738 = n4192 & n8737 ;
  assign n8739 = n3950 & ~n4784 ;
  assign n8740 = ~x81 & n8739 ;
  assign n8741 = n8738 & ~n8740 ;
  assign n8742 = n8741 ^ n2292 ^ 1'b0 ;
  assign n8745 = n8744 ^ n8742 ^ 1'b0 ;
  assign n8746 = ~x32 & n3691 ;
  assign n8747 = n4194 ^ n2705 ^ n492 ;
  assign n8748 = ( n2650 & ~n4712 ) | ( n2650 & n8747 ) | ( ~n4712 & n8747 ) ;
  assign n8749 = ( n381 & n8746 ) | ( n381 & ~n8748 ) | ( n8746 & ~n8748 ) ;
  assign n8750 = n8745 | n8749 ;
  assign n8754 = n1762 | n2704 ;
  assign n8753 = n2060 ^ n2035 ^ 1'b0 ;
  assign n8751 = n6247 ^ n4164 ^ 1'b0 ;
  assign n8752 = n2254 & ~n8751 ;
  assign n8755 = n8754 ^ n8753 ^ n8752 ;
  assign n8756 = n8755 ^ n1994 ^ 1'b0 ;
  assign n8757 = ~n2409 & n4163 ;
  assign n8758 = n8757 ^ n211 ^ 1'b0 ;
  assign n8759 = n1390 ^ n1123 ^ n776 ;
  assign n8760 = n8759 ^ n7337 ^ n806 ;
  assign n8761 = n1400 | n3121 ;
  assign n8762 = n1202 & ~n8761 ;
  assign n8763 = n3565 & ~n8762 ;
  assign n8764 = n7174 | n8763 ;
  assign n8765 = n2280 | n8764 ;
  assign n8766 = n8760 | n8765 ;
  assign n8767 = n6361 ^ n4110 ^ 1'b0 ;
  assign n8768 = n2375 ^ n182 ^ 1'b0 ;
  assign n8769 = n1611 & ~n4394 ;
  assign n8770 = n8769 ^ x60 ^ 1'b0 ;
  assign n8771 = n3247 ^ n238 ^ 1'b0 ;
  assign n8772 = ~n6110 & n8771 ;
  assign n8773 = ( n2406 & n7234 ) | ( n2406 & n8772 ) | ( n7234 & n8772 ) ;
  assign n8774 = ( n7524 & ~n7978 ) | ( n7524 & n8773 ) | ( ~n7978 & n8773 ) ;
  assign n8775 = n6488 ^ n2339 ^ 1'b0 ;
  assign n8776 = n8775 ^ n8747 ^ n3160 ;
  assign n8777 = n2219 ^ n872 ^ 1'b0 ;
  assign n8778 = n4300 & ~n6119 ;
  assign n8779 = n4376 & n8778 ;
  assign n8780 = n8779 ^ n644 ^ n408 ;
  assign n8781 = n2383 & ~n8780 ;
  assign n8782 = n8777 & n8781 ;
  assign n8783 = n1686 & ~n8782 ;
  assign n8784 = n8783 ^ n5529 ^ 1'b0 ;
  assign n8785 = n8329 ^ n6416 ^ n5216 ;
  assign n8786 = ( n1327 & n4389 ) | ( n1327 & ~n8785 ) | ( n4389 & ~n8785 ) ;
  assign n8787 = ( n483 & n2058 ) | ( n483 & ~n4772 ) | ( n2058 & ~n4772 ) ;
  assign n8788 = ~n2931 & n3940 ;
  assign n8789 = ~n8787 & n8788 ;
  assign n8792 = n1959 & ~n3831 ;
  assign n8793 = n2211 & n8792 ;
  assign n8794 = n4457 ^ n2035 ^ 1'b0 ;
  assign n8795 = ~n8793 & n8794 ;
  assign n8790 = n3894 ^ n1654 ^ 1'b0 ;
  assign n8791 = ~n7792 & n8790 ;
  assign n8796 = n8795 ^ n8791 ^ n5519 ;
  assign n8797 = ~n783 & n7519 ;
  assign n8798 = n8409 & n8797 ;
  assign n8799 = n1429 & n8113 ;
  assign n8800 = n6336 & n8799 ;
  assign n8803 = n5712 ^ n3840 ^ n3489 ;
  assign n8801 = n3552 ^ n511 ^ n236 ;
  assign n8802 = ( ~n2010 & n4747 ) | ( ~n2010 & n8801 ) | ( n4747 & n8801 ) ;
  assign n8804 = n8803 ^ n8802 ^ 1'b0 ;
  assign n8805 = ~n8800 & n8804 ;
  assign n8806 = ~n7113 & n8805 ;
  assign n8807 = n8806 ^ n6143 ^ 1'b0 ;
  assign n8808 = ( n4647 & ~n6670 ) | ( n4647 & n7136 ) | ( ~n6670 & n7136 ) ;
  assign n8809 = n7998 ^ n7721 ^ n1299 ;
  assign n8810 = ~n5920 & n7482 ;
  assign n8811 = ( n628 & n6273 ) | ( n628 & ~n7614 ) | ( n6273 & ~n7614 ) ;
  assign n8812 = n5984 ^ n3443 ^ 1'b0 ;
  assign n8813 = n2698 & n8812 ;
  assign n8814 = ~n3519 & n8813 ;
  assign n8815 = n3721 ^ n1666 ^ x113 ;
  assign n8816 = ( n3587 & n3694 ) | ( n3587 & ~n8815 ) | ( n3694 & ~n8815 ) ;
  assign n8817 = n7262 ^ n758 ^ 1'b0 ;
  assign n8818 = n3139 & ~n8817 ;
  assign n8820 = ( n2896 & n5480 ) | ( n2896 & n7555 ) | ( n5480 & n7555 ) ;
  assign n8819 = n2279 & ~n7702 ;
  assign n8821 = n8820 ^ n8819 ^ 1'b0 ;
  assign n8823 = n3133 ^ n2650 ^ 1'b0 ;
  assign n8824 = ( n8308 & n8759 ) | ( n8308 & n8823 ) | ( n8759 & n8823 ) ;
  assign n8825 = n8824 ^ n3793 ^ n604 ;
  assign n8822 = n5278 ^ n4017 ^ n583 ;
  assign n8826 = n8825 ^ n8822 ^ 1'b0 ;
  assign n8827 = n4090 ^ n1756 ^ n156 ;
  assign n8828 = n3188 | n8827 ;
  assign n8829 = ( n160 & n1818 ) | ( n160 & n3164 ) | ( n1818 & n3164 ) ;
  assign n8830 = n8829 ^ n1852 ^ n567 ;
  assign n8831 = n1834 & ~n1870 ;
  assign n8832 = n2157 & n8831 ;
  assign n8833 = ( ~n8828 & n8830 ) | ( ~n8828 & n8832 ) | ( n8830 & n8832 ) ;
  assign n8836 = n3378 ^ n3286 ^ n1146 ;
  assign n8834 = n2974 | n6443 ;
  assign n8835 = n8451 | n8834 ;
  assign n8837 = n8836 ^ n8835 ^ n2518 ;
  assign n8838 = x66 | n1342 ;
  assign n8839 = n3503 & n8838 ;
  assign n8840 = n6577 ^ n4234 ^ 1'b0 ;
  assign n8841 = n8839 | n8840 ;
  assign n8842 = n1828 & ~n4931 ;
  assign n8843 = n5766 & n8842 ;
  assign n8844 = n5745 & ~n7499 ;
  assign n8845 = n8844 ^ n4313 ^ n3106 ;
  assign n8846 = n7542 ^ n4165 ^ n1396 ;
  assign n8847 = n7794 & n7804 ;
  assign n8848 = n3688 & n6098 ;
  assign n8849 = ~n7089 & n8848 ;
  assign n8850 = ~n1537 & n2624 ;
  assign n8851 = ~n5069 & n8850 ;
  assign n8852 = n8851 ^ n2326 ^ 1'b0 ;
  assign n8853 = n180 & n8852 ;
  assign n8854 = n8853 ^ n6621 ^ n6309 ;
  assign n8855 = ( n3373 & n4094 ) | ( n3373 & n5428 ) | ( n4094 & n5428 ) ;
  assign n8856 = n2396 ^ n1419 ^ n807 ;
  assign n8857 = x54 & ~n8856 ;
  assign n8858 = n8857 ^ n8446 ^ 1'b0 ;
  assign n8859 = ( n627 & n1763 ) | ( n627 & n1925 ) | ( n1763 & n1925 ) ;
  assign n8860 = n8859 ^ n1328 ^ 1'b0 ;
  assign n8861 = ~n262 & n8860 ;
  assign n8862 = n7337 ^ n6333 ^ 1'b0 ;
  assign n8863 = n7402 ^ n5319 ^ n1625 ;
  assign n8864 = n8206 ^ n4528 ^ n3424 ;
  assign n8865 = ( n701 & n1794 ) | ( n701 & ~n3626 ) | ( n1794 & ~n3626 ) ;
  assign n8866 = n3505 & ~n4408 ;
  assign n8867 = n8866 ^ n4147 ^ 1'b0 ;
  assign n8868 = ( ~n2678 & n8865 ) | ( ~n2678 & n8867 ) | ( n8865 & n8867 ) ;
  assign n8869 = n6669 ^ n508 ^ 1'b0 ;
  assign n8870 = n6122 ^ x52 ^ 1'b0 ;
  assign n8871 = n8869 & ~n8870 ;
  assign n8872 = n7614 ^ n1493 ^ 1'b0 ;
  assign n8873 = ( ~n2621 & n2713 ) | ( ~n2621 & n8872 ) | ( n2713 & n8872 ) ;
  assign n8874 = n8158 ^ n4914 ^ n3517 ;
  assign n8875 = n8357 ^ n2151 ^ 1'b0 ;
  assign n8876 = n8874 | n8875 ;
  assign n8877 = n2749 ^ n766 ^ 1'b0 ;
  assign n8878 = n307 & n8877 ;
  assign n8879 = n8878 ^ n3101 ^ 1'b0 ;
  assign n8883 = ( n266 & ~n2172 ) | ( n266 & n8397 ) | ( ~n2172 & n8397 ) ;
  assign n8880 = n1986 & n2308 ;
  assign n8881 = ~n188 & n8880 ;
  assign n8882 = n8881 ^ n4090 ^ 1'b0 ;
  assign n8884 = n8883 ^ n8882 ^ n2061 ;
  assign n8885 = ( ~n508 & n3221 ) | ( ~n508 & n4982 ) | ( n3221 & n4982 ) ;
  assign n8886 = x113 & ~n8885 ;
  assign n8887 = n6213 & n8886 ;
  assign n8888 = ( n3966 & n8288 ) | ( n3966 & ~n8887 ) | ( n8288 & ~n8887 ) ;
  assign n8889 = n8117 & ~n8888 ;
  assign n8890 = n8889 ^ n1089 ^ 1'b0 ;
  assign n8891 = n4472 ^ n577 ^ n472 ;
  assign n8892 = n2255 & ~n8891 ;
  assign n8893 = n8892 ^ n7794 ^ 1'b0 ;
  assign n8894 = n7227 ^ n7026 ^ n6590 ;
  assign n8895 = n2749 & ~n4124 ;
  assign n8896 = n8895 ^ n2545 ^ n199 ;
  assign n8897 = ~n4208 & n6256 ;
  assign n8898 = ~n1116 & n8897 ;
  assign n8899 = ( n970 & n3668 ) | ( n970 & n4008 ) | ( n3668 & n4008 ) ;
  assign n8900 = n1569 & ~n8899 ;
  assign n8901 = n8172 & n8900 ;
  assign n8902 = n3257 ^ n250 ^ 1'b0 ;
  assign n8903 = ~n7353 & n8902 ;
  assign n8904 = n5491 ^ n462 ^ n170 ;
  assign n8905 = n2757 ^ n1089 ^ 1'b0 ;
  assign n8906 = ~n7033 & n7830 ;
  assign n8907 = ~n6625 & n8906 ;
  assign n8908 = n7753 ^ n1460 ^ 1'b0 ;
  assign n8909 = n8908 ^ n6057 ^ x82 ;
  assign n8912 = n7370 ^ n6513 ^ n2994 ;
  assign n8910 = n4185 ^ n3477 ^ n1097 ;
  assign n8911 = n8910 ^ n3666 ^ 1'b0 ;
  assign n8913 = n8912 ^ n8911 ^ n4409 ;
  assign n8914 = ~n1046 & n8913 ;
  assign n8915 = ~n8326 & n8914 ;
  assign n8916 = n8915 ^ n915 ^ 1'b0 ;
  assign n8917 = n3780 | n3947 ;
  assign n8918 = n8917 ^ n673 ^ 1'b0 ;
  assign n8919 = ( n3321 & n7501 ) | ( n3321 & ~n8918 ) | ( n7501 & ~n8918 ) ;
  assign n8920 = n3357 | n4505 ;
  assign n8921 = n8920 ^ n8043 ^ n1002 ;
  assign n8922 = ( n794 & n6043 ) | ( n794 & n8921 ) | ( n6043 & n8921 ) ;
  assign n8923 = ( n4096 & ~n5295 ) | ( n4096 & n5973 ) | ( ~n5295 & n5973 ) ;
  assign n8924 = n8923 ^ n1084 ^ 1'b0 ;
  assign n8925 = n6769 | n8924 ;
  assign n8926 = n1164 & ~n2581 ;
  assign n8927 = n8851 ^ n4677 ^ n366 ;
  assign n8928 = n8927 ^ n3511 ^ n383 ;
  assign n8929 = ( n2780 & n3610 ) | ( n2780 & n8928 ) | ( n3610 & n8928 ) ;
  assign n8930 = n3436 ^ n2125 ^ 1'b0 ;
  assign n8931 = ~n2490 & n7252 ;
  assign n8932 = ( n3721 & ~n8782 ) | ( n3721 & n8931 ) | ( ~n8782 & n8931 ) ;
  assign n8933 = n4822 ^ n2001 ^ 1'b0 ;
  assign n8934 = ~n2156 & n8933 ;
  assign n8935 = x33 & n8934 ;
  assign n8936 = n659 & n8935 ;
  assign n8937 = n8723 ^ n2190 ^ 1'b0 ;
  assign n8938 = n4808 & ~n8937 ;
  assign n8939 = n7584 ^ n4115 ^ 1'b0 ;
  assign n8940 = n376 | n5099 ;
  assign n8941 = n7051 | n8940 ;
  assign n8942 = n596 & ~n2593 ;
  assign n8943 = n8942 ^ n831 ^ 1'b0 ;
  assign n8944 = n2434 & n8943 ;
  assign n8945 = x115 & ~n2085 ;
  assign n8946 = n8945 ^ n466 ^ 1'b0 ;
  assign n8947 = n143 & n7571 ;
  assign n8948 = ~n8946 & n8947 ;
  assign n8949 = n1053 | n2515 ;
  assign n8950 = n8949 ^ n535 ^ 1'b0 ;
  assign n8951 = ~n8012 & n8950 ;
  assign n8953 = n5332 ^ n4332 ^ n2609 ;
  assign n8954 = n8953 ^ n6579 ^ n461 ;
  assign n8952 = n2051 | n2885 ;
  assign n8955 = n8954 ^ n8952 ^ 1'b0 ;
  assign n8956 = n761 ^ n255 ^ 1'b0 ;
  assign n8957 = ~n8691 & n8956 ;
  assign n8958 = n7218 ^ n4611 ^ n3681 ;
  assign n8959 = ( ~n1123 & n8523 ) | ( ~n1123 & n8958 ) | ( n8523 & n8958 ) ;
  assign n8960 = ( n405 & ~n2733 ) | ( n405 & n3386 ) | ( ~n2733 & n3386 ) ;
  assign n8961 = n1927 | n8960 ;
  assign n8962 = n1999 ^ n1426 ^ 1'b0 ;
  assign n8963 = n8962 ^ n5635 ^ n328 ;
  assign n8964 = n3950 ^ n253 ^ 1'b0 ;
  assign n8965 = ( n1054 & ~n2368 ) | ( n1054 & n6312 ) | ( ~n2368 & n6312 ) ;
  assign n8966 = n6576 ^ n3600 ^ x120 ;
  assign n8967 = n550 | n1553 ;
  assign n8968 = n3448 ^ n2845 ^ 1'b0 ;
  assign n8969 = n6082 & ~n8968 ;
  assign n8970 = ( n2779 & n8967 ) | ( n2779 & n8969 ) | ( n8967 & n8969 ) ;
  assign n8971 = n6783 ^ n2307 ^ 1'b0 ;
  assign n8972 = n8970 & n8971 ;
  assign n8973 = n8972 ^ n6963 ^ n2070 ;
  assign n8977 = n3152 & ~n6743 ;
  assign n8978 = n8977 ^ n2372 ^ 1'b0 ;
  assign n8974 = n3101 & n8576 ;
  assign n8975 = n8974 ^ x114 ^ 1'b0 ;
  assign n8976 = n4633 | n8975 ;
  assign n8979 = n8978 ^ n8976 ^ 1'b0 ;
  assign n8980 = ~n531 & n5928 ;
  assign n8981 = ~x109 & n8980 ;
  assign n8982 = ( n2036 & n2544 ) | ( n2036 & ~n3631 ) | ( n2544 & ~n3631 ) ;
  assign n8983 = n8981 | n8982 ;
  assign n8984 = n1020 & ~n8983 ;
  assign n8985 = n8251 | n8984 ;
  assign n8986 = n2424 | n5021 ;
  assign n8987 = n8986 ^ n3617 ^ 1'b0 ;
  assign n8988 = n8987 ^ n1796 ^ 1'b0 ;
  assign n8989 = n2598 | n4387 ;
  assign n8990 = n3772 & ~n8989 ;
  assign n8991 = n8990 ^ n1773 ^ n737 ;
  assign n8992 = n4567 ^ n1918 ^ x45 ;
  assign n8993 = ( n8988 & n8991 ) | ( n8988 & n8992 ) | ( n8991 & n8992 ) ;
  assign n8994 = n771 & ~n5566 ;
  assign n8995 = ~n8035 & n8994 ;
  assign n8996 = n1046 | n8995 ;
  assign n8997 = n8996 ^ n1388 ^ 1'b0 ;
  assign n8998 = n8997 ^ n2950 ^ 1'b0 ;
  assign n8999 = ~n8993 & n8998 ;
  assign n9005 = n551 | n4383 ;
  assign n9007 = n4094 ^ n295 ^ x122 ;
  assign n9006 = n238 | n1448 ;
  assign n9008 = n9007 ^ n9006 ^ 1'b0 ;
  assign n9009 = n9008 ^ n5729 ^ n2565 ;
  assign n9010 = n9009 ^ n1350 ^ 1'b0 ;
  assign n9011 = n9005 & ~n9010 ;
  assign n9001 = ( n981 & n1068 ) | ( n981 & n3083 ) | ( n1068 & n3083 ) ;
  assign n9000 = n7144 ^ n4808 ^ n1646 ;
  assign n9002 = n9001 ^ n9000 ^ n3301 ;
  assign n9003 = ( n2140 & n2913 ) | ( n2140 & n9002 ) | ( n2913 & n9002 ) ;
  assign n9004 = n1554 & n9003 ;
  assign n9012 = n9011 ^ n9004 ^ 1'b0 ;
  assign n9013 = ~n233 & n1922 ;
  assign n9014 = n9013 ^ n1576 ^ 1'b0 ;
  assign n9015 = n9014 ^ n2219 ^ 1'b0 ;
  assign n9016 = ( n1100 & n4286 ) | ( n1100 & ~n9015 ) | ( n4286 & ~n9015 ) ;
  assign n9017 = n9016 ^ n7432 ^ 1'b0 ;
  assign n9018 = ( ~n1466 & n3850 ) | ( ~n1466 & n7234 ) | ( n3850 & n7234 ) ;
  assign n9019 = n1343 ^ n1236 ^ 1'b0 ;
  assign n9020 = n9019 ^ n2513 ^ 1'b0 ;
  assign n9021 = n9018 | n9020 ;
  assign n9023 = n4561 ^ n2088 ^ 1'b0 ;
  assign n9024 = n9023 ^ n2355 ^ 1'b0 ;
  assign n9022 = n5808 ^ n4087 ^ n1628 ;
  assign n9025 = n9024 ^ n9022 ^ n6867 ;
  assign n9026 = ( n738 & ~n1907 ) | ( n738 & n6298 ) | ( ~n1907 & n6298 ) ;
  assign n9027 = n1453 ^ n840 ^ 1'b0 ;
  assign n9028 = n9026 & n9027 ;
  assign n9029 = ~n3482 & n5211 ;
  assign n9030 = ~n9028 & n9029 ;
  assign n9031 = ~n721 & n5036 ;
  assign n9032 = ~n5629 & n9031 ;
  assign n9033 = n2835 ^ n2401 ^ 1'b0 ;
  assign n9034 = n4378 ^ n469 ^ 1'b0 ;
  assign n9037 = n1797 & ~n3817 ;
  assign n9038 = n9037 ^ n6330 ^ 1'b0 ;
  assign n9039 = ( n4791 & n5902 ) | ( n4791 & n9038 ) | ( n5902 & n9038 ) ;
  assign n9035 = n1765 ^ n246 ^ 1'b0 ;
  assign n9036 = n9035 ^ n1496 ^ n1098 ;
  assign n9040 = n9039 ^ n9036 ^ n5472 ;
  assign n9041 = n6656 | n7695 ;
  assign n9042 = n2175 ^ n1573 ^ 1'b0 ;
  assign n9043 = n2337 | n5596 ;
  assign n9044 = n9042 & n9043 ;
  assign n9045 = ~n573 & n2859 ;
  assign n9046 = n9045 ^ n6768 ^ n2833 ;
  assign n9047 = n9046 ^ n3114 ^ n1927 ;
  assign n9048 = n9047 ^ n3335 ^ 1'b0 ;
  assign n9049 = n9048 ^ n6593 ^ n1171 ;
  assign n9050 = n7727 ^ n5385 ^ n3557 ;
  assign n9051 = ~n2122 & n7827 ;
  assign n9052 = n9051 ^ n8861 ^ 1'b0 ;
  assign n9053 = ~n3104 & n5364 ;
  assign n9054 = ( n1202 & n2686 ) | ( n1202 & n4201 ) | ( n2686 & n4201 ) ;
  assign n9055 = n7748 & ~n9054 ;
  assign n9056 = ~n687 & n9055 ;
  assign n9057 = n4141 & ~n9056 ;
  assign n9058 = ~n1686 & n9057 ;
  assign n9059 = n9053 & n9058 ;
  assign n9060 = n9059 ^ n4618 ^ 1'b0 ;
  assign n9061 = ( n6315 & ~n8039 ) | ( n6315 & n9060 ) | ( ~n8039 & n9060 ) ;
  assign n9062 = n2801 ^ n1736 ^ n1287 ;
  assign n9063 = n3290 & n6042 ;
  assign n9064 = n9063 ^ n7611 ^ n991 ;
  assign n9065 = n9064 ^ n8748 ^ 1'b0 ;
  assign n9066 = n9065 ^ n5216 ^ 1'b0 ;
  assign n9067 = ~n8194 & n9066 ;
  assign n9068 = n5904 | n7068 ;
  assign n9069 = n9068 ^ n5012 ^ 1'b0 ;
  assign n9070 = n7854 & ~n8272 ;
  assign n9071 = ~n1143 & n9070 ;
  assign n9072 = n2467 & ~n8202 ;
  assign n9073 = n9072 ^ n6233 ^ 1'b0 ;
  assign n9074 = n9073 ^ n162 ^ 1'b0 ;
  assign n9075 = ( n291 & n4747 ) | ( n291 & ~n6790 ) | ( n4747 & ~n6790 ) ;
  assign n9076 = n4700 ^ n2817 ^ 1'b0 ;
  assign n9077 = n9076 ^ n2625 ^ 1'b0 ;
  assign n9078 = n3831 | n7897 ;
  assign n9079 = n9025 & ~n9078 ;
  assign n9080 = n1442 | n4172 ;
  assign n9081 = n4774 & ~n9080 ;
  assign n9082 = n9081 ^ n5695 ^ n3046 ;
  assign n9083 = n9082 ^ n3134 ^ 1'b0 ;
  assign n9084 = n2971 | n9083 ;
  assign n9085 = n6344 | n9084 ;
  assign n9086 = n1568 & ~n9085 ;
  assign n9087 = ( ~n4127 & n5050 ) | ( ~n4127 & n7982 ) | ( n5050 & n7982 ) ;
  assign n9088 = n9087 ^ n1799 ^ n865 ;
  assign n9089 = n6419 ^ n6405 ^ n4310 ;
  assign n9090 = n691 & n5340 ;
  assign n9091 = ~n1110 & n9090 ;
  assign n9092 = n9091 ^ n3556 ^ 1'b0 ;
  assign n9093 = n9089 & n9092 ;
  assign n9094 = n1666 ^ n1075 ^ 1'b0 ;
  assign n9095 = n129 & ~n9094 ;
  assign n9096 = n5139 ^ n3965 ^ n1986 ;
  assign n9097 = n9096 ^ n8318 ^ 1'b0 ;
  assign n9103 = ( x127 & n291 ) | ( x127 & ~n1723 ) | ( n291 & ~n1723 ) ;
  assign n9098 = n4100 ^ n485 ^ 1'b0 ;
  assign n9099 = ~n2582 & n3135 ;
  assign n9100 = ~n754 & n9099 ;
  assign n9101 = ( ~n3146 & n9098 ) | ( ~n3146 & n9100 ) | ( n9098 & n9100 ) ;
  assign n9102 = n9101 ^ n3766 ^ 1'b0 ;
  assign n9104 = n9103 ^ n9102 ^ n912 ;
  assign n9105 = ( ~n3077 & n3903 ) | ( ~n3077 & n5897 ) | ( n3903 & n5897 ) ;
  assign n9106 = n2996 ^ n1555 ^ n973 ;
  assign n9107 = n1635 & n6583 ;
  assign n9108 = n3093 | n3722 ;
  assign n9109 = n9108 ^ n3840 ^ 1'b0 ;
  assign n9110 = n3220 | n5210 ;
  assign n9114 = ~n1827 & n1850 ;
  assign n9111 = n3169 ^ n1688 ^ x16 ;
  assign n9112 = n4094 | n9111 ;
  assign n9113 = n9112 ^ n7882 ^ 1'b0 ;
  assign n9115 = n9114 ^ n9113 ^ n1732 ;
  assign n9116 = n5088 ^ n1801 ^ n255 ;
  assign n9117 = ( n3710 & n8704 ) | ( n3710 & ~n9116 ) | ( n8704 & ~n9116 ) ;
  assign n9118 = n5355 ^ n3507 ^ 1'b0 ;
  assign n9119 = n8097 & n9118 ;
  assign n9122 = n1196 & ~n2494 ;
  assign n9123 = n9122 ^ n2713 ^ 1'b0 ;
  assign n9124 = n9123 ^ n1762 ^ 1'b0 ;
  assign n9125 = ~n7754 & n9124 ;
  assign n9120 = n7647 ^ n5289 ^ n3262 ;
  assign n9121 = ( n222 & ~n2065 ) | ( n222 & n9120 ) | ( ~n2065 & n9120 ) ;
  assign n9126 = n9125 ^ n9121 ^ n6866 ;
  assign n9131 = n1726 & ~n2730 ;
  assign n9132 = n5942 & n9131 ;
  assign n9133 = n6816 | n9132 ;
  assign n9134 = n9133 ^ n3611 ^ 1'b0 ;
  assign n9127 = n5126 ^ n4406 ^ n2770 ;
  assign n9128 = n6758 & n9127 ;
  assign n9129 = n9128 ^ n9059 ^ 1'b0 ;
  assign n9130 = n1188 & ~n9129 ;
  assign n9135 = n9134 ^ n9130 ^ 1'b0 ;
  assign n9136 = n7556 ^ n4096 ^ n1287 ;
  assign n9137 = n9136 ^ n3100 ^ 1'b0 ;
  assign n9138 = n7620 & n9137 ;
  assign n9139 = n4007 ^ n2518 ^ 1'b0 ;
  assign n9140 = n3847 | n5521 ;
  assign n9141 = n9139 | n9140 ;
  assign n9142 = n4468 | n4714 ;
  assign n9143 = n9142 ^ n7254 ^ n763 ;
  assign n9144 = n392 & n2793 ;
  assign n9145 = x57 & n2581 ;
  assign n9146 = n9145 ^ n2463 ^ n1456 ;
  assign n9147 = n1605 & n1658 ;
  assign n9148 = n9146 & ~n9147 ;
  assign n9149 = n9148 ^ n1870 ^ 1'b0 ;
  assign n9151 = n6803 ^ n676 ^ 1'b0 ;
  assign n9150 = n4802 & ~n7770 ;
  assign n9152 = n9151 ^ n9150 ^ 1'b0 ;
  assign n9153 = n4864 & ~n9152 ;
  assign n9154 = n9153 ^ n5590 ^ 1'b0 ;
  assign n9155 = n5008 ^ n2805 ^ n2019 ;
  assign n9156 = n8403 ^ n1394 ^ 1'b0 ;
  assign n9157 = n9155 & ~n9156 ;
  assign n9158 = n7719 ^ n4823 ^ n3979 ;
  assign n9159 = n9158 ^ n4807 ^ 1'b0 ;
  assign n9160 = n3580 ^ n1989 ^ n1000 ;
  assign n9161 = n8103 ^ n1980 ^ n899 ;
  assign n9162 = ~n5271 & n9161 ;
  assign n9163 = n9162 ^ n5120 ^ 1'b0 ;
  assign n9164 = ~n9160 & n9163 ;
  assign n9165 = n9164 ^ x6 ^ 1'b0 ;
  assign n9166 = n9165 ^ n3015 ^ 1'b0 ;
  assign n9167 = ( n1199 & n1301 ) | ( n1199 & n2320 ) | ( n1301 & n2320 ) ;
  assign n9168 = n7156 & ~n9167 ;
  assign n9169 = n464 & ~n5741 ;
  assign n9170 = n9169 ^ n2192 ^ 1'b0 ;
  assign n9171 = n8982 | n9170 ;
  assign n9172 = n6332 | n9171 ;
  assign n9173 = n9172 ^ n8365 ^ n2338 ;
  assign n9174 = n7115 ^ n6249 ^ 1'b0 ;
  assign n9175 = n9174 ^ n7832 ^ n7412 ;
  assign n9176 = n9175 ^ n5510 ^ n3858 ;
  assign n9177 = n5420 ^ n1840 ^ 1'b0 ;
  assign n9178 = n8393 ^ n8273 ^ n3816 ;
  assign n9179 = n7760 ^ n985 ^ 1'b0 ;
  assign n9180 = ( n3433 & n5386 ) | ( n3433 & n5552 ) | ( n5386 & n5552 ) ;
  assign n9181 = ( ~n4684 & n9179 ) | ( ~n4684 & n9180 ) | ( n9179 & n9180 ) ;
  assign n9182 = x20 & n1899 ;
  assign n9183 = n9182 ^ n6502 ^ 1'b0 ;
  assign n9184 = ~n6317 & n9158 ;
  assign n9185 = n1833 | n9184 ;
  assign n9186 = n9185 ^ n4036 ^ 1'b0 ;
  assign n9187 = n9183 & ~n9186 ;
  assign n9188 = n6450 | n9187 ;
  assign n9189 = n9188 ^ x113 ^ 1'b0 ;
  assign n9190 = n4025 ^ n3578 ^ n3011 ;
  assign n9191 = ~n6588 & n9190 ;
  assign n9192 = n1785 & n9191 ;
  assign n9193 = n3718 & ~n9192 ;
  assign n9194 = ( n2003 & n3390 ) | ( n2003 & ~n6045 ) | ( n3390 & ~n6045 ) ;
  assign n9195 = n3709 & n9194 ;
  assign n9196 = n9193 | n9195 ;
  assign n9197 = n9196 ^ n7525 ^ 1'b0 ;
  assign n9198 = n1178 & n3803 ;
  assign n9199 = ( ~n5441 & n9197 ) | ( ~n5441 & n9198 ) | ( n9197 & n9198 ) ;
  assign n9200 = n8330 ^ n5361 ^ n5079 ;
  assign n9201 = n6640 ^ n5008 ^ n378 ;
  assign n9202 = n1077 & n5289 ;
  assign n9203 = n2281 & n9202 ;
  assign n9204 = ~n764 & n8268 ;
  assign n9205 = n4827 & ~n8322 ;
  assign n9206 = ( n2165 & n4409 ) | ( n2165 & n6207 ) | ( n4409 & n6207 ) ;
  assign n9207 = ( ~n2060 & n2829 ) | ( ~n2060 & n2965 ) | ( n2829 & n2965 ) ;
  assign n9208 = n1786 | n6192 ;
  assign n9209 = n9208 ^ n2559 ^ 1'b0 ;
  assign n9210 = n9209 ^ n7335 ^ x79 ;
  assign n9211 = n930 & ~n3131 ;
  assign n9212 = x7 & ~n2399 ;
  assign n9213 = n9212 ^ n3288 ^ 1'b0 ;
  assign n9214 = ~n1086 & n5368 ;
  assign n9215 = n9214 ^ n7612 ^ 1'b0 ;
  assign n9216 = n1317 | n4882 ;
  assign n9217 = ( n2805 & n8374 ) | ( n2805 & n9216 ) | ( n8374 & n9216 ) ;
  assign n9223 = ( n1025 & n2157 ) | ( n1025 & ~n2360 ) | ( n2157 & ~n2360 ) ;
  assign n9218 = n4164 ^ n2457 ^ n2240 ;
  assign n9219 = x113 & n2365 ;
  assign n9220 = ~n1656 & n9219 ;
  assign n9221 = n6384 & ~n9220 ;
  assign n9222 = n9218 & n9221 ;
  assign n9224 = n9223 ^ n9222 ^ 1'b0 ;
  assign n9226 = n2853 ^ n2243 ^ n789 ;
  assign n9227 = ( ~n831 & n1080 ) | ( ~n831 & n9226 ) | ( n1080 & n9226 ) ;
  assign n9228 = n9227 ^ n5041 ^ 1'b0 ;
  assign n9225 = n3027 ^ n349 ^ 1'b0 ;
  assign n9229 = n9228 ^ n9225 ^ n1890 ;
  assign n9230 = n180 | n1545 ;
  assign n9231 = n3024 | n8441 ;
  assign n9232 = n1767 & ~n6969 ;
  assign n9233 = n9231 & n9232 ;
  assign n9234 = n2048 | n5631 ;
  assign n9235 = n9233 & ~n9234 ;
  assign n9236 = n2254 | n6891 ;
  assign n9237 = n9236 ^ n8007 ^ 1'b0 ;
  assign n9238 = n5822 ^ n1209 ^ 1'b0 ;
  assign n9239 = n3991 & n9238 ;
  assign n9240 = n9239 ^ n3267 ^ n1784 ;
  assign n9241 = ( ~n2483 & n2970 ) | ( ~n2483 & n4694 ) | ( n2970 & n4694 ) ;
  assign n9242 = n434 & n2838 ;
  assign n9243 = n9242 ^ n3162 ^ n1679 ;
  assign n9244 = ~n1215 & n9243 ;
  assign n9245 = n9244 ^ n1218 ^ 1'b0 ;
  assign n9246 = n2377 ^ n2162 ^ n1951 ;
  assign n9247 = ( n2631 & n9245 ) | ( n2631 & ~n9246 ) | ( n9245 & ~n9246 ) ;
  assign n9248 = x110 & ~n1448 ;
  assign n9249 = n9248 ^ n6314 ^ 1'b0 ;
  assign n9250 = n8065 | n9249 ;
  assign n9251 = n7806 ^ n2411 ^ 1'b0 ;
  assign n9252 = n8408 ^ n1204 ^ 1'b0 ;
  assign n9253 = n955 | n1523 ;
  assign n9254 = ~n4594 & n9253 ;
  assign n9255 = ~n2213 & n9254 ;
  assign n9256 = n4625 & n9255 ;
  assign n9257 = n9256 ^ n2917 ^ 1'b0 ;
  assign n9258 = ~n3617 & n4321 ;
  assign n9259 = ~n6985 & n9258 ;
  assign n9260 = n7988 ^ n5093 ^ 1'b0 ;
  assign n9261 = n8775 ^ n5606 ^ 1'b0 ;
  assign n9262 = ~n1509 & n2369 ;
  assign n9263 = n9262 ^ n8502 ^ 1'b0 ;
  assign n9264 = n9263 ^ n2738 ^ 1'b0 ;
  assign n9265 = ~n6244 & n9264 ;
  assign n9266 = n9265 ^ n2688 ^ 1'b0 ;
  assign n9267 = n9266 ^ n8121 ^ n1699 ;
  assign n9268 = n8596 ^ n7512 ^ n1485 ;
  assign n9269 = ( ~n547 & n822 ) | ( ~n547 & n2532 ) | ( n822 & n2532 ) ;
  assign n9270 = n4302 & n9269 ;
  assign n9271 = n9270 ^ n6674 ^ 1'b0 ;
  assign n9272 = ( ~n432 & n783 ) | ( ~n432 & n7187 ) | ( n783 & n7187 ) ;
  assign n9273 = n9272 ^ n4176 ^ 1'b0 ;
  assign n9274 = n7014 ^ n2101 ^ 1'b0 ;
  assign n9275 = ( n3075 & n3310 ) | ( n3075 & ~n9274 ) | ( n3310 & ~n9274 ) ;
  assign n9276 = n4297 & n7100 ;
  assign n9277 = n9276 ^ n3565 ^ 1'b0 ;
  assign n9278 = ~n2637 & n9277 ;
  assign n9279 = n1540 & n9278 ;
  assign n9280 = n9279 ^ n7659 ^ 1'b0 ;
  assign n9281 = n3540 & ~n6506 ;
  assign n9282 = ( ~n3355 & n7190 ) | ( ~n3355 & n9281 ) | ( n7190 & n9281 ) ;
  assign n9283 = n8237 ^ n2732 ^ 1'b0 ;
  assign n9284 = n3576 ^ n232 ^ 1'b0 ;
  assign n9285 = n6399 | n9284 ;
  assign n9286 = n9285 ^ n3274 ^ n256 ;
  assign n9287 = n1573 & n5848 ;
  assign n9288 = ( n257 & n2331 ) | ( n257 & n2581 ) | ( n2331 & n2581 ) ;
  assign n9289 = n1270 ^ x119 ^ 1'b0 ;
  assign n9290 = ~n9288 & n9289 ;
  assign n9291 = n6137 & n9290 ;
  assign n9292 = n9291 ^ n1639 ^ 1'b0 ;
  assign n9293 = n6043 ^ n2597 ^ 1'b0 ;
  assign n9294 = ~n3614 & n9293 ;
  assign n9295 = x79 & ~n733 ;
  assign n9296 = n9295 ^ n4086 ^ n3035 ;
  assign n9297 = ~n1342 & n2015 ;
  assign n9298 = n9297 ^ n7488 ^ 1'b0 ;
  assign n9299 = n9296 & ~n9298 ;
  assign n9300 = n5985 ^ x49 ^ 1'b0 ;
  assign n9301 = n5915 ^ n786 ^ 1'b0 ;
  assign n9302 = n2539 ^ n1534 ^ 1'b0 ;
  assign n9303 = n4867 ^ n4247 ^ n893 ;
  assign n9304 = ( n7003 & n8591 ) | ( n7003 & ~n9303 ) | ( n8591 & ~n9303 ) ;
  assign n9305 = ( ~n2163 & n7625 ) | ( ~n2163 & n9106 ) | ( n7625 & n9106 ) ;
  assign n9306 = n7072 ^ n4740 ^ n3488 ;
  assign n9307 = n6701 ^ n3877 ^ 1'b0 ;
  assign n9308 = n9307 ^ x127 ^ 1'b0 ;
  assign n9309 = n9308 ^ n7340 ^ n3548 ;
  assign n9310 = n636 & n1234 ;
  assign n9311 = ~n1217 & n3480 ;
  assign n9312 = n567 & n9311 ;
  assign n9313 = n7896 ^ n917 ^ 1'b0 ;
  assign n9314 = ~n9312 & n9313 ;
  assign n9315 = ( n7774 & ~n7882 ) | ( n7774 & n9314 ) | ( ~n7882 & n9314 ) ;
  assign n9316 = ( n7560 & n7776 ) | ( n7560 & n9315 ) | ( n7776 & n9315 ) ;
  assign n9317 = n1905 | n9316 ;
  assign n9318 = n6284 & ~n6541 ;
  assign n9319 = ~x59 & n9318 ;
  assign n9320 = n2782 & ~n9319 ;
  assign n9321 = ~n2334 & n9320 ;
  assign n9322 = n5605 ^ n4280 ^ n915 ;
  assign n9323 = n9322 ^ n1200 ^ 1'b0 ;
  assign n9324 = n6485 ^ n6316 ^ 1'b0 ;
  assign n9325 = n2101 & ~n4172 ;
  assign n9326 = ~n5762 & n9325 ;
  assign n9335 = n890 & n4466 ;
  assign n9334 = n6670 ^ n887 ^ 1'b0 ;
  assign n9327 = n605 | n2826 ;
  assign n9328 = n9327 ^ n3602 ^ 1'b0 ;
  assign n9329 = n9328 ^ n1410 ^ 1'b0 ;
  assign n9330 = n1623 & ~n9329 ;
  assign n9331 = n9330 ^ n3374 ^ n2127 ;
  assign n9332 = n2987 & n9331 ;
  assign n9333 = ~n5873 & n9332 ;
  assign n9336 = n9335 ^ n9334 ^ n9333 ;
  assign n9337 = n9336 ^ n8480 ^ 1'b0 ;
  assign n9338 = n9326 | n9337 ;
  assign n9339 = ( n997 & ~n9324 ) | ( n997 & n9338 ) | ( ~n9324 & n9338 ) ;
  assign n9341 = n2797 ^ x69 ^ 1'b0 ;
  assign n9342 = ~n3827 & n9341 ;
  assign n9343 = n8198 | n9342 ;
  assign n9340 = n4100 & ~n5247 ;
  assign n9344 = n9343 ^ n9340 ^ 1'b0 ;
  assign n9345 = n4029 ^ n447 ^ 1'b0 ;
  assign n9346 = n4039 & n9345 ;
  assign n9347 = n6527 ^ n4952 ^ 1'b0 ;
  assign n9348 = ~n1770 & n9347 ;
  assign n9349 = ( n550 & n9346 ) | ( n550 & n9348 ) | ( n9346 & n9348 ) ;
  assign n9353 = n2922 ^ n960 ^ 1'b0 ;
  assign n9354 = ~n3956 & n9353 ;
  assign n9350 = n4329 ^ n1759 ^ n1730 ;
  assign n9351 = n6196 ^ n1741 ^ n1343 ;
  assign n9352 = n9350 & ~n9351 ;
  assign n9355 = n9354 ^ n9352 ^ 1'b0 ;
  assign n9356 = ~n328 & n3178 ;
  assign n9357 = ( ~n5001 & n6409 ) | ( ~n5001 & n9356 ) | ( n6409 & n9356 ) ;
  assign n9358 = n6477 & n9357 ;
  assign n9359 = ~n756 & n9358 ;
  assign n9360 = n5584 ^ n3195 ^ n1781 ;
  assign n9361 = n2851 ^ n2472 ^ 1'b0 ;
  assign n9362 = n2175 & n3411 ;
  assign n9363 = n9194 ^ n7193 ^ n425 ;
  assign n9364 = x77 & ~n3534 ;
  assign n9365 = n9363 & ~n9364 ;
  assign n9366 = n9365 ^ n5545 ^ n949 ;
  assign n9367 = ~n1423 & n3712 ;
  assign n9368 = n442 & n9367 ;
  assign n9369 = n2514 | n9368 ;
  assign n9373 = n4530 ^ n3567 ^ 1'b0 ;
  assign n9371 = n4267 & ~n6196 ;
  assign n9372 = n9371 ^ n8308 ^ n2022 ;
  assign n9370 = n4464 & ~n8010 ;
  assign n9374 = n9373 ^ n9372 ^ n9370 ;
  assign n9375 = ( ~n822 & n9369 ) | ( ~n822 & n9374 ) | ( n9369 & n9374 ) ;
  assign n9376 = ~n517 & n8611 ;
  assign n9377 = ~n9375 & n9376 ;
  assign n9378 = ( n182 & n2449 ) | ( n182 & n2921 ) | ( n2449 & n2921 ) ;
  assign n9379 = n9378 ^ n1879 ^ 1'b0 ;
  assign n9380 = n2200 & n4525 ;
  assign n9381 = ~n8065 & n9380 ;
  assign n9382 = n8497 ^ n4133 ^ 1'b0 ;
  assign n9383 = ~n367 & n9382 ;
  assign n9384 = ( n982 & n2342 ) | ( n982 & ~n3154 ) | ( n2342 & ~n3154 ) ;
  assign n9385 = ( n5099 & ~n5304 ) | ( n5099 & n9384 ) | ( ~n5304 & n9384 ) ;
  assign n9387 = n5367 ^ n2422 ^ 1'b0 ;
  assign n9388 = n4078 & n9387 ;
  assign n9386 = n580 & ~n2048 ;
  assign n9389 = n9388 ^ n9386 ^ n141 ;
  assign n9390 = ( ~n1899 & n2792 ) | ( ~n1899 & n6456 ) | ( n2792 & n6456 ) ;
  assign n9391 = ( n2391 & n3405 ) | ( n2391 & ~n3557 ) | ( n3405 & ~n3557 ) ;
  assign n9392 = ~n9390 & n9391 ;
  assign n9393 = n5045 & n9392 ;
  assign n9394 = n599 | n9393 ;
  assign n9395 = n6327 ^ n2348 ^ 1'b0 ;
  assign n9396 = n4973 | n9395 ;
  assign n9397 = ( x59 & ~n9394 ) | ( x59 & n9396 ) | ( ~n9394 & n9396 ) ;
  assign n9398 = n4483 ^ n2293 ^ 1'b0 ;
  assign n9399 = n559 | n9398 ;
  assign n9400 = n7367 | n9399 ;
  assign n9401 = n1123 & n3043 ;
  assign n9402 = ~n1590 & n9401 ;
  assign n9403 = n2469 & ~n3932 ;
  assign n9404 = ( ~n6524 & n9402 ) | ( ~n6524 & n9403 ) | ( n9402 & n9403 ) ;
  assign n9405 = n5528 & n9404 ;
  assign n9406 = n5229 & n9405 ;
  assign n9407 = n1326 & n1808 ;
  assign n9408 = n9406 & n9407 ;
  assign n9409 = n7369 ^ n6454 ^ n171 ;
  assign n9410 = ~n5716 & n9409 ;
  assign n9411 = n9410 ^ n6621 ^ 1'b0 ;
  assign n9412 = n5069 ^ n793 ^ 1'b0 ;
  assign n9413 = x4 & n9412 ;
  assign n9414 = n3919 ^ n1339 ^ n804 ;
  assign n9417 = n5641 & ~n8450 ;
  assign n9418 = n9417 ^ n2253 ^ 1'b0 ;
  assign n9415 = n1067 ^ n294 ^ 1'b0 ;
  assign n9416 = n5431 & ~n9415 ;
  assign n9419 = n9418 ^ n9416 ^ n2863 ;
  assign n9420 = n9419 ^ n5389 ^ n2227 ;
  assign n9421 = n1733 ^ n205 ^ 1'b0 ;
  assign n9429 = n7324 ^ n5886 ^ n1797 ;
  assign n9422 = n1876 | n7192 ;
  assign n9423 = n1448 & ~n9422 ;
  assign n9424 = n321 & ~n1994 ;
  assign n9425 = n9423 & n9424 ;
  assign n9426 = n5772 & ~n9425 ;
  assign n9427 = ~n2134 & n9426 ;
  assign n9428 = n6800 | n9427 ;
  assign n9430 = n9429 ^ n9428 ^ 1'b0 ;
  assign n9431 = n2416 ^ n2228 ^ 1'b0 ;
  assign n9432 = n4242 ^ n544 ^ 1'b0 ;
  assign n9433 = n7600 | n9432 ;
  assign n9434 = ( ~n915 & n1521 ) | ( ~n915 & n5640 ) | ( n1521 & n5640 ) ;
  assign n9435 = ( n5510 & ~n6755 ) | ( n5510 & n9434 ) | ( ~n6755 & n9434 ) ;
  assign n9436 = n9435 ^ n2293 ^ 1'b0 ;
  assign n9437 = n6449 ^ n5937 ^ n2949 ;
  assign n9439 = n2543 ^ n2029 ^ n1001 ;
  assign n9438 = n413 | n5610 ;
  assign n9440 = n9439 ^ n9438 ^ 1'b0 ;
  assign n9441 = n1519 | n9440 ;
  assign n9442 = ~n1204 & n9111 ;
  assign n9443 = n9442 ^ n5766 ^ n2640 ;
  assign n9444 = n8510 ^ n456 ^ 1'b0 ;
  assign n9445 = n9443 & n9444 ;
  assign n9446 = ( n3867 & n6969 ) | ( n3867 & n9445 ) | ( n6969 & n9445 ) ;
  assign n9447 = n9446 ^ n2968 ^ 1'b0 ;
  assign n9448 = n3812 | n9447 ;
  assign n9449 = n6974 ^ n3947 ^ n399 ;
  assign n9450 = n8753 ^ n5610 ^ n1652 ;
  assign n9452 = n3639 & ~n9218 ;
  assign n9453 = n9452 ^ n4405 ^ 1'b0 ;
  assign n9451 = n6317 ^ n158 ^ 1'b0 ;
  assign n9454 = n9453 ^ n9451 ^ n6604 ;
  assign n9455 = ~n1638 & n3477 ;
  assign n9456 = n2402 ^ n1290 ^ n134 ;
  assign n9457 = n4807 ^ n3917 ^ 1'b0 ;
  assign n9458 = n9456 & ~n9457 ;
  assign n9459 = n3341 ^ n1707 ^ 1'b0 ;
  assign n9460 = ~n2493 & n9459 ;
  assign n9461 = n1553 & ~n2636 ;
  assign n9462 = n4394 & n9461 ;
  assign n9463 = n4653 ^ n2284 ^ 1'b0 ;
  assign n9464 = n9463 ^ n7243 ^ 1'b0 ;
  assign n9465 = x63 & n2573 ;
  assign n9466 = ( ~n9462 & n9464 ) | ( ~n9462 & n9465 ) | ( n9464 & n9465 ) ;
  assign n9467 = n4656 & n8490 ;
  assign n9468 = ~n3047 & n9467 ;
  assign n9469 = n2490 | n9468 ;
  assign n9470 = n2632 | n5355 ;
  assign n9471 = n8838 ^ n856 ^ 1'b0 ;
  assign n9472 = n9471 ^ n1433 ^ 1'b0 ;
  assign n9473 = ( ~n372 & n2088 ) | ( ~n372 & n2927 ) | ( n2088 & n2927 ) ;
  assign n9474 = n2342 & ~n4285 ;
  assign n9475 = n9473 & n9474 ;
  assign n9476 = n9475 ^ n3737 ^ 1'b0 ;
  assign n9477 = n9472 | n9476 ;
  assign n9478 = n1089 & n9477 ;
  assign n9479 = n7333 & ~n9478 ;
  assign n9480 = ( n610 & ~n855 ) | ( n610 & n5765 ) | ( ~n855 & n5765 ) ;
  assign n9481 = n2691 ^ n1921 ^ 1'b0 ;
  assign n9482 = ~n5791 & n9481 ;
  assign n9483 = n6086 ^ n4007 ^ 1'b0 ;
  assign n9484 = ( n6274 & n9482 ) | ( n6274 & ~n9483 ) | ( n9482 & ~n9483 ) ;
  assign n9489 = n1435 | n6206 ;
  assign n9485 = n4259 ^ n1571 ^ 1'b0 ;
  assign n9486 = ( n2522 & n3351 ) | ( n2522 & ~n9485 ) | ( n3351 & ~n9485 ) ;
  assign n9487 = n4408 | n9486 ;
  assign n9488 = n5101 & ~n9487 ;
  assign n9490 = n9489 ^ n9488 ^ 1'b0 ;
  assign n9491 = n8932 & ~n9490 ;
  assign n9492 = ( ~n4127 & n4597 ) | ( ~n4127 & n6103 ) | ( n4597 & n6103 ) ;
  assign n9493 = n7954 & ~n9492 ;
  assign n9494 = ( n4046 & n5355 ) | ( n4046 & ~n8923 ) | ( n5355 & ~n8923 ) ;
  assign n9496 = n5002 ^ n3175 ^ 1'b0 ;
  assign n9497 = ~n1096 & n9496 ;
  assign n9498 = ~n2007 & n9497 ;
  assign n9499 = n9498 ^ n5201 ^ 1'b0 ;
  assign n9495 = n2584 & ~n6319 ;
  assign n9500 = n9499 ^ n9495 ^ n3946 ;
  assign n9501 = n972 & ~n4339 ;
  assign n9502 = n9501 ^ n652 ^ 1'b0 ;
  assign n9503 = n8237 | n9502 ;
  assign n9504 = n9503 ^ n8499 ^ 1'b0 ;
  assign n9511 = ( n597 & n1986 ) | ( n597 & ~n3042 ) | ( n1986 & ~n3042 ) ;
  assign n9512 = n2322 | n9511 ;
  assign n9505 = n5021 ^ n1840 ^ 1'b0 ;
  assign n9506 = n6103 ^ n2242 ^ n770 ;
  assign n9507 = n5598 & ~n9506 ;
  assign n9508 = n9507 ^ n2774 ^ n1131 ;
  assign n9509 = n9508 ^ n7066 ^ n4987 ;
  assign n9510 = n9505 | n9509 ;
  assign n9513 = n9512 ^ n9510 ^ 1'b0 ;
  assign n9514 = n6993 ^ n383 ^ 1'b0 ;
  assign n9515 = n1043 & n2202 ;
  assign n9516 = n9515 ^ n9442 ^ 1'b0 ;
  assign n9517 = ~n9514 & n9516 ;
  assign n9518 = n4390 & n9517 ;
  assign n9519 = n5418 & ~n7430 ;
  assign n9520 = n9519 ^ n8291 ^ 1'b0 ;
  assign n9521 = n4384 ^ n1670 ^ 1'b0 ;
  assign n9522 = n956 ^ n408 ^ 1'b0 ;
  assign n9523 = n9522 ^ n1635 ^ 1'b0 ;
  assign n9524 = ~n808 & n9523 ;
  assign n9525 = ~n2863 & n5371 ;
  assign n9526 = n4195 & n9525 ;
  assign n9527 = n947 & ~n2077 ;
  assign n9528 = n9527 ^ x22 ^ 1'b0 ;
  assign n9529 = n5512 ^ n1942 ^ n1464 ;
  assign n9530 = n4875 & ~n7132 ;
  assign n9531 = n9529 & n9530 ;
  assign n9532 = n9531 ^ n752 ^ 1'b0 ;
  assign n9533 = n1697 | n9532 ;
  assign n9534 = n5832 ^ n5476 ^ n3766 ;
  assign n9535 = n911 | n4814 ;
  assign n9536 = n9534 | n9535 ;
  assign n9537 = n2811 | n6065 ;
  assign n9538 = ~n3068 & n9537 ;
  assign n9539 = ~n9536 & n9538 ;
  assign n9540 = n9539 ^ n4120 ^ 1'b0 ;
  assign n9541 = ~n9533 & n9540 ;
  assign n9542 = ~n1580 & n4867 ;
  assign n9543 = n9542 ^ n8664 ^ 1'b0 ;
  assign n9544 = ( n9528 & ~n9541 ) | ( n9528 & n9543 ) | ( ~n9541 & n9543 ) ;
  assign n9547 = n4090 & n9463 ;
  assign n9545 = ( n2093 & n2181 ) | ( n2093 & ~n3842 ) | ( n2181 & ~n3842 ) ;
  assign n9546 = n9545 ^ n7559 ^ 1'b0 ;
  assign n9548 = n9547 ^ n9546 ^ x103 ;
  assign n9549 = x61 & n932 ;
  assign n9550 = ~n5533 & n9549 ;
  assign n9552 = ~n983 & n2953 ;
  assign n9553 = n6853 & n9552 ;
  assign n9551 = n5326 & ~n5905 ;
  assign n9554 = n9553 ^ n9551 ^ n3670 ;
  assign n9557 = n2528 | n4700 ;
  assign n9558 = n9557 ^ n4365 ^ 1'b0 ;
  assign n9555 = n3232 ^ n1924 ^ 1'b0 ;
  assign n9556 = n7056 & ~n9555 ;
  assign n9559 = n9558 ^ n9556 ^ n643 ;
  assign n9560 = n1753 ^ n1498 ^ 1'b0 ;
  assign n9561 = n7467 & n9560 ;
  assign n9562 = n1773 ^ n1534 ^ 1'b0 ;
  assign n9563 = n4391 & ~n9562 ;
  assign n9564 = n1072 & ~n1145 ;
  assign n9565 = n9563 & n9564 ;
  assign n9566 = ( x38 & n1929 ) | ( x38 & ~n8441 ) | ( n1929 & ~n8441 ) ;
  assign n9569 = n5610 ^ n2595 ^ n1959 ;
  assign n9567 = n1019 ^ n520 ^ 1'b0 ;
  assign n9568 = n7719 | n9567 ;
  assign n9570 = n9569 ^ n9568 ^ 1'b0 ;
  assign n9571 = ~n3224 & n9570 ;
  assign n9573 = n7199 ^ n451 ^ 1'b0 ;
  assign n9572 = n793 & n6358 ;
  assign n9574 = n9573 ^ n9572 ^ 1'b0 ;
  assign n9575 = ~n1481 & n9574 ;
  assign n9576 = n9575 ^ n5675 ^ 1'b0 ;
  assign n9577 = n9470 & ~n9576 ;
  assign n9578 = n1996 | n8196 ;
  assign n9579 = n2932 & n6528 ;
  assign n9580 = ~n2112 & n9579 ;
  assign n9581 = n1138 | n9580 ;
  assign n9582 = n9581 ^ n6046 ^ 1'b0 ;
  assign n9583 = n947 & ~n994 ;
  assign n9584 = ~n364 & n9583 ;
  assign n9585 = ( ~n1838 & n5260 ) | ( ~n1838 & n9584 ) | ( n5260 & n9584 ) ;
  assign n9586 = n1798 & n9585 ;
  assign n9587 = ~n6027 & n9586 ;
  assign n9588 = n9587 ^ n3386 ^ 1'b0 ;
  assign n9589 = n4187 & n5683 ;
  assign n9590 = n6481 & ~n7256 ;
  assign n9591 = n2202 & n9590 ;
  assign n9592 = n6571 & ~n9591 ;
  assign n9593 = n9592 ^ n5760 ^ 1'b0 ;
  assign n9600 = n272 & n2854 ;
  assign n9601 = n5418 & ~n9600 ;
  assign n9602 = n1290 | n9601 ;
  assign n9596 = n2655 & n3658 ;
  assign n9597 = n9596 ^ n4880 ^ 1'b0 ;
  assign n9594 = n1671 & n3288 ;
  assign n9595 = ~n9170 & n9594 ;
  assign n9598 = n9597 ^ n9595 ^ n411 ;
  assign n9599 = n4527 | n9598 ;
  assign n9603 = n9602 ^ n9599 ^ 1'b0 ;
  assign n9604 = n5314 ^ n2947 ^ 1'b0 ;
  assign n9605 = n2756 & ~n9604 ;
  assign n9606 = n5339 | n8755 ;
  assign n9607 = n6206 | n9606 ;
  assign n9608 = n9607 ^ n3926 ^ n2219 ;
  assign n9609 = n3008 ^ n1676 ^ 1'b0 ;
  assign n9610 = n9609 ^ n2601 ^ 1'b0 ;
  assign n9611 = n3646 & n9610 ;
  assign n9612 = ( ~n9605 & n9608 ) | ( ~n9605 & n9611 ) | ( n9608 & n9611 ) ;
  assign n9613 = n4882 & ~n5220 ;
  assign n9614 = n4703 | n9613 ;
  assign n9616 = n3639 & n7978 ;
  assign n9617 = ~n7009 & n9616 ;
  assign n9615 = ( ~n1555 & n3527 ) | ( ~n1555 & n7536 ) | ( n3527 & n7536 ) ;
  assign n9618 = n9617 ^ n9615 ^ 1'b0 ;
  assign n9619 = n2304 | n2424 ;
  assign n9620 = n2152 | n9619 ;
  assign n9621 = n9620 ^ n1188 ^ 1'b0 ;
  assign n9622 = n8112 | n9621 ;
  assign n9623 = n4062 ^ n1070 ^ 1'b0 ;
  assign n9624 = n9622 | n9623 ;
  assign n9625 = n1328 & ~n4094 ;
  assign n9626 = ~n8215 & n9625 ;
  assign n9627 = n5886 ^ n1411 ^ 1'b0 ;
  assign n9628 = ( n4844 & n6150 ) | ( n4844 & n9627 ) | ( n6150 & n9627 ) ;
  assign n9629 = n6416 & ~n9628 ;
  assign n9630 = ~n2724 & n9629 ;
  assign n9631 = n7461 & ~n9630 ;
  assign n9632 = n9626 & n9631 ;
  assign n9633 = n6004 ^ n4436 ^ 1'b0 ;
  assign n9634 = n4405 | n9633 ;
  assign n9635 = n7071 ^ n2735 ^ 1'b0 ;
  assign n9636 = n9229 & ~n9635 ;
  assign n9637 = n9636 ^ n3829 ^ 1'b0 ;
  assign n9638 = ( n7789 & ~n8558 ) | ( n7789 & n8620 ) | ( ~n8558 & n8620 ) ;
  assign n9642 = n7064 & n8669 ;
  assign n9643 = n1855 & n9642 ;
  assign n9644 = n5128 | n9643 ;
  assign n9639 = n2294 & ~n2320 ;
  assign n9640 = n8545 | n9639 ;
  assign n9641 = n4765 | n9640 ;
  assign n9645 = n9644 ^ n9641 ^ 1'b0 ;
  assign n9646 = ~n473 & n2882 ;
  assign n9647 = n9646 ^ n2154 ^ 1'b0 ;
  assign n9648 = ~n2934 & n9647 ;
  assign n9649 = n4784 | n5870 ;
  assign n9650 = n619 & n2177 ;
  assign n9651 = ~n646 & n9650 ;
  assign n9652 = n9123 & ~n9651 ;
  assign n9653 = ~n9649 & n9652 ;
  assign n9663 = n4164 & ~n5170 ;
  assign n9664 = n9663 ^ n8490 ^ 1'b0 ;
  assign n9660 = n3740 ^ n2766 ^ n2491 ;
  assign n9661 = ( n259 & n1339 ) | ( n259 & ~n9660 ) | ( n1339 & ~n9660 ) ;
  assign n9662 = ( n773 & n924 ) | ( n773 & ~n9661 ) | ( n924 & ~n9661 ) ;
  assign n9665 = n9664 ^ n9662 ^ n9241 ;
  assign n9654 = ( n1934 & n4163 ) | ( n1934 & ~n6790 ) | ( n4163 & ~n6790 ) ;
  assign n9655 = n5276 | n9654 ;
  assign n9656 = n2831 | n9655 ;
  assign n9657 = n9656 ^ n623 ^ 1'b0 ;
  assign n9658 = n9657 ^ n8632 ^ 1'b0 ;
  assign n9659 = n5102 & ~n9658 ;
  assign n9666 = n9665 ^ n9659 ^ 1'b0 ;
  assign n9668 = n9639 ^ n3473 ^ 1'b0 ;
  assign n9669 = n3857 & ~n9668 ;
  assign n9670 = ( n5425 & ~n6833 ) | ( n5425 & n9669 ) | ( ~n6833 & n9669 ) ;
  assign n9671 = ~n4598 & n5666 ;
  assign n9672 = n1932 & n9671 ;
  assign n9673 = n1205 & n2453 ;
  assign n9674 = ( n1773 & n6338 ) | ( n1773 & n9673 ) | ( n6338 & n9673 ) ;
  assign n9675 = n9672 & ~n9674 ;
  assign n9676 = n9675 ^ n5544 ^ 1'b0 ;
  assign n9677 = n9670 | n9676 ;
  assign n9667 = n7686 & n8067 ;
  assign n9678 = n9677 ^ n9667 ^ 1'b0 ;
  assign n9679 = n5166 ^ n1599 ^ x98 ;
  assign n9680 = n9679 ^ n5325 ^ 1'b0 ;
  assign n9681 = n2623 & ~n9680 ;
  assign n9682 = n624 & ~n7259 ;
  assign n9683 = n9682 ^ n7136 ^ 1'b0 ;
  assign n9684 = n2058 & n9683 ;
  assign n9685 = n9684 ^ n4877 ^ 1'b0 ;
  assign n9686 = n887 & ~n9685 ;
  assign n9687 = n3614 & n9686 ;
  assign n9688 = n9687 ^ n7743 ^ 1'b0 ;
  assign n9689 = n8224 | n9688 ;
  assign n9690 = n3393 ^ n1731 ^ 1'b0 ;
  assign n9691 = ( n1978 & ~n3410 ) | ( n1978 & n9690 ) | ( ~n3410 & n9690 ) ;
  assign n9692 = n9691 ^ n1018 ^ 1'b0 ;
  assign n9693 = ~n1751 & n9692 ;
  assign n9694 = n4474 & n9693 ;
  assign n9695 = n6283 & n9694 ;
  assign n9696 = ~n6649 & n9695 ;
  assign n9697 = n7270 ^ n4634 ^ 1'b0 ;
  assign n9698 = ~n1877 & n9697 ;
  assign n9699 = n8765 ^ n8692 ^ n4566 ;
  assign n9700 = n9698 & ~n9699 ;
  assign n9701 = n1329 ^ n308 ^ 1'b0 ;
  assign n9702 = n9673 | n9701 ;
  assign n9703 = n2779 ^ n1939 ^ 1'b0 ;
  assign n9704 = n4022 & ~n9703 ;
  assign n9705 = ( ~n1699 & n9702 ) | ( ~n1699 & n9704 ) | ( n9702 & n9704 ) ;
  assign n9706 = ~n218 & n8298 ;
  assign n9707 = ~n5362 & n9706 ;
  assign n9708 = n6454 & n9707 ;
  assign n9709 = n9708 ^ n8712 ^ 1'b0 ;
  assign n9710 = n833 & n9709 ;
  assign n9711 = n8059 ^ n3004 ^ n1654 ;
  assign n9712 = n260 & ~n1939 ;
  assign n9713 = n3532 & n9712 ;
  assign n9714 = n9534 | n9713 ;
  assign n9715 = n4852 ^ n4440 ^ n1538 ;
  assign n9716 = n9715 ^ n5681 ^ n4772 ;
  assign n9717 = n5500 & ~n9716 ;
  assign n9718 = n6749 | n9717 ;
  assign n9719 = n627 & ~n9718 ;
  assign n9720 = n7932 & ~n9719 ;
  assign n9721 = ~n5262 & n9720 ;
  assign n9722 = n9721 ^ n1200 ^ n917 ;
  assign n9723 = n798 | n9722 ;
  assign n9724 = n7719 ^ x59 ^ 1'b0 ;
  assign n9725 = n4625 | n9724 ;
  assign n9732 = n2971 & ~n9508 ;
  assign n9733 = n7319 & n9732 ;
  assign n9726 = n3763 ^ n1800 ^ n710 ;
  assign n9727 = n6881 ^ n5302 ^ 1'b0 ;
  assign n9728 = n9726 & ~n9727 ;
  assign n9729 = ( n143 & ~n1718 ) | ( n143 & n8318 ) | ( ~n1718 & n8318 ) ;
  assign n9730 = n9729 ^ n3413 ^ 1'b0 ;
  assign n9731 = n9728 & n9730 ;
  assign n9734 = n9733 ^ n9731 ^ 1'b0 ;
  assign n9735 = ~n3136 & n4482 ;
  assign n9736 = n9735 ^ n5942 ^ 1'b0 ;
  assign n9737 = n466 & ~n9736 ;
  assign n9738 = n7919 ^ n6185 ^ 1'b0 ;
  assign n9739 = ~n7955 & n9738 ;
  assign n9741 = n4483 ^ n2490 ^ 1'b0 ;
  assign n9742 = ~n2244 & n9741 ;
  assign n9743 = n9742 ^ n1137 ^ 1'b0 ;
  assign n9744 = ~n248 & n9743 ;
  assign n9740 = n2799 ^ n796 ^ 1'b0 ;
  assign n9745 = n9744 ^ n9740 ^ 1'b0 ;
  assign n9751 = n2179 ^ n402 ^ 1'b0 ;
  assign n9747 = n6891 ^ x101 ^ 1'b0 ;
  assign n9748 = n3470 | n9747 ;
  assign n9746 = n383 & ~n1779 ;
  assign n9749 = n9748 ^ n9746 ^ n3433 ;
  assign n9750 = ~n6824 & n9749 ;
  assign n9752 = n9751 ^ n9750 ^ 1'b0 ;
  assign n9753 = x42 & n8372 ;
  assign n9754 = n9752 & n9753 ;
  assign n9757 = ( n1087 & ~n1246 ) | ( n1087 & n1551 ) | ( ~n1246 & n1551 ) ;
  assign n9755 = n4390 ^ n827 ^ 1'b0 ;
  assign n9756 = n4723 & ~n9755 ;
  assign n9758 = n9757 ^ n9756 ^ 1'b0 ;
  assign n9760 = ~n331 & n1818 ;
  assign n9761 = ~n1382 & n9760 ;
  assign n9759 = n971 | n3178 ;
  assign n9762 = n9761 ^ n9759 ^ 1'b0 ;
  assign n9763 = n227 | n9762 ;
  assign n9764 = n9763 ^ n9615 ^ 1'b0 ;
  assign n9765 = n8916 ^ n1846 ^ 1'b0 ;
  assign n9766 = ( n1117 & n3555 ) | ( n1117 & n7015 ) | ( n3555 & n7015 ) ;
  assign n9767 = ( x96 & n5156 ) | ( x96 & n9766 ) | ( n5156 & n9766 ) ;
  assign n9768 = n9767 ^ n7019 ^ n5233 ;
  assign n9769 = n6617 ^ n3955 ^ 1'b0 ;
  assign n9770 = n2175 & ~n9769 ;
  assign n9771 = n8757 ^ n5991 ^ n2981 ;
  assign n9775 = n1990 ^ n857 ^ 1'b0 ;
  assign n9776 = n9775 ^ n5505 ^ 1'b0 ;
  assign n9777 = n1339 & n9776 ;
  assign n9772 = ~n3175 & n3596 ;
  assign n9773 = ~n4606 & n9772 ;
  assign n9774 = n3940 & ~n9773 ;
  assign n9778 = n9777 ^ n9774 ^ 1'b0 ;
  assign n9779 = n9778 ^ n689 ^ 1'b0 ;
  assign n9780 = n5717 & n9779 ;
  assign n9781 = n8820 ^ n7589 ^ n6198 ;
  assign n9782 = n4200 ^ n1494 ^ 1'b0 ;
  assign n9783 = n7988 ^ n1683 ^ 1'b0 ;
  assign n9784 = ~n1458 & n9783 ;
  assign n9785 = n9784 ^ n8454 ^ 1'b0 ;
  assign n9786 = n5673 & n9785 ;
  assign n9787 = n9782 & n9786 ;
  assign n9788 = n141 | n2008 ;
  assign n9789 = n9788 ^ n234 ^ 1'b0 ;
  assign n9790 = n9789 ^ n7494 ^ n3972 ;
  assign n9791 = n9437 ^ n1056 ^ 1'b0 ;
  assign n9792 = n7451 & ~n9791 ;
  assign n9793 = n6453 ^ n4238 ^ 1'b0 ;
  assign n9794 = x54 & n2823 ;
  assign n9795 = ~n2434 & n9794 ;
  assign n9796 = n8060 ^ n2929 ^ 1'b0 ;
  assign n9797 = ~n3654 & n9796 ;
  assign n9801 = ( n1954 & ~n2537 ) | ( n1954 & n4602 ) | ( ~n2537 & n4602 ) ;
  assign n9802 = n366 & n5022 ;
  assign n9803 = ~n894 & n9802 ;
  assign n9804 = ~n5932 & n9803 ;
  assign n9805 = n6989 ^ n3390 ^ n2967 ;
  assign n9806 = ( n8394 & n9804 ) | ( n8394 & n9805 ) | ( n9804 & n9805 ) ;
  assign n9807 = ~n9801 & n9806 ;
  assign n9808 = n9807 ^ n7048 ^ 1'b0 ;
  assign n9798 = n560 | n4329 ;
  assign n9799 = n7132 & ~n9798 ;
  assign n9800 = n2247 & n9799 ;
  assign n9809 = n9808 ^ n9800 ^ 1'b0 ;
  assign n9810 = n5596 ^ n2530 ^ x85 ;
  assign n9811 = n9190 ^ n1433 ^ 1'b0 ;
  assign n9812 = n2036 & ~n4394 ;
  assign n9813 = n9811 & n9812 ;
  assign n9814 = ~n2573 & n9813 ;
  assign n9815 = ( n2131 & ~n4711 ) | ( n2131 & n9419 ) | ( ~n4711 & n9419 ) ;
  assign n9816 = ( n4135 & ~n9814 ) | ( n4135 & n9815 ) | ( ~n9814 & n9815 ) ;
  assign n9817 = n875 ^ n155 ^ 1'b0 ;
  assign n9818 = n4774 ^ n4090 ^ 1'b0 ;
  assign n9819 = ~n9817 & n9818 ;
  assign n9820 = n7840 & n9819 ;
  assign n9821 = n9820 ^ n4230 ^ 1'b0 ;
  assign n9822 = ~n401 & n9821 ;
  assign n9823 = n7968 ^ n5454 ^ n2339 ;
  assign n9824 = n2235 ^ n1969 ^ n558 ;
  assign n9825 = n3646 & n9824 ;
  assign n9826 = n9810 & n9825 ;
  assign n9827 = ( n477 & n831 ) | ( n477 & n5421 ) | ( n831 & n5421 ) ;
  assign n9828 = ( n2165 & n2338 ) | ( n2165 & n4885 ) | ( n2338 & n4885 ) ;
  assign n9829 = ( n6530 & n9827 ) | ( n6530 & ~n9828 ) | ( n9827 & ~n9828 ) ;
  assign n9830 = n5308 & ~n9829 ;
  assign n9831 = n3628 | n7012 ;
  assign n9832 = n2897 | n9831 ;
  assign n9833 = n6623 & n9832 ;
  assign n9834 = n3648 & n9833 ;
  assign n9838 = ( n2262 & n3626 ) | ( n2262 & ~n4822 ) | ( n3626 & ~n4822 ) ;
  assign n9835 = n3585 ^ n2265 ^ n1861 ;
  assign n9836 = n9835 ^ n4728 ^ 1'b0 ;
  assign n9837 = n4445 & ~n9836 ;
  assign n9839 = n9838 ^ n9837 ^ n6561 ;
  assign n9840 = n3501 & n7794 ;
  assign n9841 = ~n2762 & n9840 ;
  assign n9842 = n4642 ^ n2165 ^ n1069 ;
  assign n9843 = ( ~n4039 & n9841 ) | ( ~n4039 & n9842 ) | ( n9841 & n9842 ) ;
  assign n9844 = n6250 ^ n3572 ^ 1'b0 ;
  assign n9845 = ~n6197 & n9844 ;
  assign n9846 = n4663 ^ n2303 ^ 1'b0 ;
  assign n9847 = n5083 ^ n592 ^ 1'b0 ;
  assign n9848 = ~n9846 & n9847 ;
  assign n9849 = ( ~n4407 & n9845 ) | ( ~n4407 & n9848 ) | ( n9845 & n9848 ) ;
  assign n9850 = ( n5929 & ~n7591 ) | ( n5929 & n9849 ) | ( ~n7591 & n9849 ) ;
  assign n9851 = n7103 & n9850 ;
  assign n9852 = n2348 & n9851 ;
  assign n9853 = n9852 ^ n4488 ^ 1'b0 ;
  assign n9854 = n2462 | n8289 ;
  assign n9855 = n6211 | n9854 ;
  assign n9856 = n3303 ^ n2302 ^ 1'b0 ;
  assign n9857 = n1579 & ~n9856 ;
  assign n9858 = ~n6502 & n9857 ;
  assign n9859 = n9858 ^ n1796 ^ 1'b0 ;
  assign n9860 = n7014 ^ n1671 ^ n1640 ;
  assign n9861 = ~n9859 & n9860 ;
  assign n9862 = n9861 ^ n4705 ^ 1'b0 ;
  assign n9863 = n9855 & n9862 ;
  assign n9864 = n241 | n514 ;
  assign n9865 = n9864 ^ n2978 ^ 1'b0 ;
  assign n9868 = n1120 & ~n2459 ;
  assign n9869 = n2668 & n9868 ;
  assign n9866 = n3133 ^ n308 ^ 1'b0 ;
  assign n9867 = n4208 & n9866 ;
  assign n9870 = n9869 ^ n9867 ^ 1'b0 ;
  assign n9871 = ( ~n1813 & n4944 ) | ( ~n1813 & n9870 ) | ( n4944 & n9870 ) ;
  assign n9872 = n6988 ^ n3820 ^ 1'b0 ;
  assign n9873 = n3011 | n9872 ;
  assign n9874 = n9873 ^ n9648 ^ 1'b0 ;
  assign n9875 = ~n1460 & n9874 ;
  assign n9876 = n3646 ^ n1973 ^ n299 ;
  assign n9877 = n3293 ^ n307 ^ 1'b0 ;
  assign n9878 = n6872 & ~n9877 ;
  assign n9879 = n9878 ^ n7941 ^ 1'b0 ;
  assign n9880 = n356 & ~n9879 ;
  assign n9881 = n9880 ^ n2688 ^ 1'b0 ;
  assign n9882 = n9881 ^ n3697 ^ 1'b0 ;
  assign n9883 = n9876 & ~n9882 ;
  assign n9884 = n6824 ^ n5154 ^ n4516 ;
  assign n9885 = ( ~n540 & n3475 ) | ( ~n540 & n6137 ) | ( n3475 & n6137 ) ;
  assign n9886 = ~n1451 & n2698 ;
  assign n9887 = ~n4583 & n9886 ;
  assign n9888 = n9887 ^ n9246 ^ n4103 ;
  assign n9889 = n6858 ^ n5700 ^ n497 ;
  assign n9890 = ( n5614 & n9192 ) | ( n5614 & n9889 ) | ( n9192 & n9889 ) ;
  assign n9891 = n7183 ^ n6059 ^ 1'b0 ;
  assign n9892 = ~n7373 & n9891 ;
  assign n9893 = n149 | n2296 ;
  assign n9894 = n9893 ^ n6151 ^ 1'b0 ;
  assign n9895 = ~n4266 & n7402 ;
  assign n9896 = n9894 & n9895 ;
  assign n9897 = n9896 ^ n2272 ^ 1'b0 ;
  assign n9898 = n2820 & n9897 ;
  assign n9899 = n8031 ^ n1268 ^ n1196 ;
  assign n9900 = n5629 & n9899 ;
  assign n9901 = ~n9898 & n9900 ;
  assign n9902 = ~n1701 & n4283 ;
  assign n9903 = n5381 & n9902 ;
  assign n9904 = n9903 ^ n7842 ^ 1'b0 ;
  assign n9905 = n9904 ^ n5795 ^ 1'b0 ;
  assign n9906 = ( n3015 & ~n4202 ) | ( n3015 & n9905 ) | ( ~n4202 & n9905 ) ;
  assign n9907 = ( n7489 & n9901 ) | ( n7489 & n9906 ) | ( n9901 & n9906 ) ;
  assign n9909 = n8552 ^ x109 ^ 1'b0 ;
  assign n9908 = n4192 & n5325 ;
  assign n9910 = n9909 ^ n9908 ^ 1'b0 ;
  assign n9911 = n269 & n9186 ;
  assign n9912 = n9910 | n9911 ;
  assign n9916 = n3396 & ~n8076 ;
  assign n9913 = n4013 & ~n6502 ;
  assign n9914 = ~n5875 & n9913 ;
  assign n9915 = n9073 & n9914 ;
  assign n9917 = n9916 ^ n9915 ^ 1'b0 ;
  assign n9922 = n5625 ^ n4222 ^ 1'b0 ;
  assign n9918 = n6953 ^ n3028 ^ n2889 ;
  assign n9919 = ( x24 & n4114 ) | ( x24 & ~n9918 ) | ( n4114 & ~n9918 ) ;
  assign n9920 = n9919 ^ n2415 ^ 1'b0 ;
  assign n9921 = n9920 ^ n9277 ^ n8173 ;
  assign n9923 = n9922 ^ n9921 ^ n4296 ;
  assign n9924 = n7143 ^ n2571 ^ 1'b0 ;
  assign n9927 = ~n2516 & n4379 ;
  assign n9925 = n1431 | n8076 ;
  assign n9926 = n9925 ^ n5121 ^ x115 ;
  assign n9928 = n9927 ^ n9926 ^ n4686 ;
  assign n9929 = n9928 ^ n136 ^ 1'b0 ;
  assign n9930 = n1368 ^ n322 ^ 1'b0 ;
  assign n9931 = ~n1073 & n9930 ;
  assign n9932 = n3883 | n9931 ;
  assign n9933 = n4949 ^ n302 ^ 1'b0 ;
  assign n9934 = n3264 & n9933 ;
  assign n9935 = n9934 ^ n222 ^ 1'b0 ;
  assign n9936 = n857 & ~n3035 ;
  assign n9937 = n9936 ^ n3832 ^ n1114 ;
  assign n9938 = n9937 ^ n9562 ^ n3249 ;
  assign n9939 = n4377 & n6639 ;
  assign n9940 = ( n9935 & ~n9938 ) | ( n9935 & n9939 ) | ( ~n9938 & n9939 ) ;
  assign n9941 = n8215 ^ n1280 ^ x13 ;
  assign n9942 = n9941 ^ n8800 ^ n1258 ;
  assign n9943 = n5265 ^ n2122 ^ 1'b0 ;
  assign n9944 = x113 | n6841 ;
  assign n9945 = n9944 ^ n3220 ^ n2214 ;
  assign n9946 = n2601 ^ n2227 ^ 1'b0 ;
  assign n9947 = ~n4787 & n9946 ;
  assign n9948 = n9945 & n9947 ;
  assign n9955 = ( n202 & ~n1009 ) | ( n202 & n1545 ) | ( ~n1009 & n1545 ) ;
  assign n9949 = ( ~n3904 & n7446 ) | ( ~n3904 & n7840 ) | ( n7446 & n7840 ) ;
  assign n9950 = ~n4772 & n7565 ;
  assign n9951 = n1780 & n9950 ;
  assign n9952 = n1707 | n9951 ;
  assign n9953 = n9952 ^ n4470 ^ 1'b0 ;
  assign n9954 = n9949 | n9953 ;
  assign n9956 = n9955 ^ n9954 ^ n9531 ;
  assign n9957 = ( n905 & ~n1343 ) | ( n905 & n3523 ) | ( ~n1343 & n3523 ) ;
  assign n9958 = ( n897 & n3065 ) | ( n897 & n9957 ) | ( n3065 & n9957 ) ;
  assign n9959 = n9958 ^ n8730 ^ n789 ;
  assign n9961 = n1966 ^ n1499 ^ 1'b0 ;
  assign n9962 = n1686 & ~n9961 ;
  assign n9963 = n9962 ^ n7088 ^ n2579 ;
  assign n9960 = n9045 ^ n7832 ^ n7251 ;
  assign n9964 = n9963 ^ n9960 ^ n2473 ;
  assign n9965 = n4233 ^ n2489 ^ n2029 ;
  assign n9966 = n7028 | n9965 ;
  assign n9967 = ( n1616 & ~n3067 ) | ( n1616 & n4677 ) | ( ~n3067 & n4677 ) ;
  assign n9968 = n9967 ^ x96 ^ 1'b0 ;
  assign n9969 = n5451 ^ n5113 ^ 1'b0 ;
  assign n9970 = n7026 ^ n6717 ^ n2051 ;
  assign n9971 = n6994 ^ n4665 ^ 1'b0 ;
  assign n9972 = n9971 ^ n7824 ^ n487 ;
  assign n9973 = n9972 ^ n7418 ^ 1'b0 ;
  assign n9974 = n1114 | n9973 ;
  assign n9975 = n9974 ^ n5280 ^ 1'b0 ;
  assign n9976 = ~n6185 & n9975 ;
  assign n9977 = n9976 ^ n6004 ^ n373 ;
  assign n9978 = n9977 ^ n4877 ^ 1'b0 ;
  assign n9979 = ~n1399 & n9978 ;
  assign n9980 = n4106 & n4306 ;
  assign n9981 = n9980 ^ n800 ^ 1'b0 ;
  assign n9982 = n1114 | n9981 ;
  assign n9983 = n4881 ^ n1389 ^ 1'b0 ;
  assign n9984 = n5445 | n9983 ;
  assign n9985 = n787 | n9984 ;
  assign n9986 = n1170 & n1339 ;
  assign n9987 = ( n5529 & n7215 ) | ( n5529 & n9986 ) | ( n7215 & n9986 ) ;
  assign n9988 = n3303 ^ n3070 ^ n2055 ;
  assign n9989 = n1378 & n9988 ;
  assign n9993 = n8588 ^ n7094 ^ 1'b0 ;
  assign n9990 = n7505 & ~n9427 ;
  assign n9991 = n5580 & n9990 ;
  assign n9992 = n7085 & ~n9991 ;
  assign n9994 = n9993 ^ n9992 ^ 1'b0 ;
  assign n9995 = n1490 & ~n4585 ;
  assign n9996 = n1585 & n8320 ;
  assign n9997 = n6218 ^ n3753 ^ n3276 ;
  assign n9998 = ( n3634 & n9842 ) | ( n3634 & ~n9997 ) | ( n9842 & ~n9997 ) ;
  assign n9999 = n1658 ^ x108 ^ 1'b0 ;
  assign n10000 = n5840 ^ n2962 ^ 1'b0 ;
  assign n10001 = ( n887 & n9999 ) | ( n887 & n10000 ) | ( n9999 & n10000 ) ;
  assign n10002 = ~n3677 & n10001 ;
  assign n10003 = ( n1086 & n1400 ) | ( n1086 & n4409 ) | ( n1400 & n4409 ) ;
  assign n10004 = n2772 & ~n10003 ;
  assign n10005 = ( n2262 & n4049 ) | ( n2262 & n10004 ) | ( n4049 & n10004 ) ;
  assign n10006 = n5228 ^ n4843 ^ 1'b0 ;
  assign n10007 = n7913 & n10006 ;
  assign n10008 = n266 & ~n5872 ;
  assign n10009 = ~n10007 & n10008 ;
  assign n10010 = n10009 ^ n251 ^ 1'b0 ;
  assign n10011 = ~n1230 & n10010 ;
  assign n10012 = ( ~n4430 & n6580 ) | ( ~n4430 & n9390 ) | ( n6580 & n9390 ) ;
  assign n10013 = n10011 & n10012 ;
  assign n10014 = n3749 & ~n7820 ;
  assign n10027 = ( n164 & n237 ) | ( n164 & n1067 ) | ( n237 & n1067 ) ;
  assign n10028 = n5791 ^ n2955 ^ 1'b0 ;
  assign n10029 = ~n10027 & n10028 ;
  assign n10030 = ( n5529 & ~n6629 ) | ( n5529 & n10029 ) | ( ~n6629 & n10029 ) ;
  assign n10015 = n4320 ^ n2587 ^ 1'b0 ;
  assign n10016 = n136 & ~n10015 ;
  assign n10017 = ( ~n551 & n8475 ) | ( ~n551 & n10016 ) | ( n8475 & n10016 ) ;
  assign n10018 = n1006 | n9664 ;
  assign n10019 = n1371 & ~n2898 ;
  assign n10020 = n4552 ^ n3304 ^ n1327 ;
  assign n10021 = n5034 & n10020 ;
  assign n10022 = ~n4238 & n10021 ;
  assign n10023 = n1246 & ~n10022 ;
  assign n10024 = ( n541 & ~n2573 ) | ( n541 & n10023 ) | ( ~n2573 & n10023 ) ;
  assign n10025 = n10019 & n10024 ;
  assign n10026 = ( n10017 & ~n10018 ) | ( n10017 & n10025 ) | ( ~n10018 & n10025 ) ;
  assign n10031 = n10030 ^ n10026 ^ n5569 ;
  assign n10032 = ( n3001 & n3579 ) | ( n3001 & n6730 ) | ( n3579 & n6730 ) ;
  assign n10042 = n9045 ^ n8753 ^ n7794 ;
  assign n10035 = n522 & n3597 ;
  assign n10036 = ~n1935 & n10035 ;
  assign n10037 = n7167 ^ n3051 ^ 1'b0 ;
  assign n10038 = n2389 & ~n10037 ;
  assign n10039 = n10038 ^ n2728 ^ 1'b0 ;
  assign n10040 = ~n10036 & n10039 ;
  assign n10041 = ~n3974 & n10040 ;
  assign n10043 = n10042 ^ n10041 ^ 1'b0 ;
  assign n10033 = n8268 ^ n3123 ^ n147 ;
  assign n10034 = n2200 & ~n10033 ;
  assign n10044 = n10043 ^ n10034 ^ 1'b0 ;
  assign n10045 = n3054 & ~n4761 ;
  assign n10046 = n296 | n615 ;
  assign n10047 = n10046 ^ x120 ^ 1'b0 ;
  assign n10048 = ( n676 & n760 ) | ( n676 & n1057 ) | ( n760 & n1057 ) ;
  assign n10049 = n10048 ^ n3929 ^ n1607 ;
  assign n10050 = ( n9017 & n10047 ) | ( n9017 & n10049 ) | ( n10047 & n10049 ) ;
  assign n10051 = n1476 & n2734 ;
  assign n10052 = n5308 & ~n10051 ;
  assign n10053 = n6477 ^ n1514 ^ 1'b0 ;
  assign n10054 = n3507 ^ n1999 ^ n774 ;
  assign n10055 = n2069 & ~n3424 ;
  assign n10056 = n10055 ^ n2638 ^ 1'b0 ;
  assign n10057 = n10056 ^ n5210 ^ n888 ;
  assign n10058 = n3323 & n10057 ;
  assign n10059 = n10058 ^ n558 ^ 1'b0 ;
  assign n10060 = n10054 & n10059 ;
  assign n10061 = ~n2869 & n10060 ;
  assign n10062 = n10061 ^ n8561 ^ 1'b0 ;
  assign n10063 = n10062 ^ n5853 ^ 1'b0 ;
  assign n10064 = n10053 | n10063 ;
  assign n10066 = n3959 & ~n7130 ;
  assign n10065 = n9675 ^ n6406 ^ 1'b0 ;
  assign n10067 = n10066 ^ n10065 ^ n4880 ;
  assign n10068 = ( ~n1861 & n4450 ) | ( ~n1861 & n6273 ) | ( n4450 & n6273 ) ;
  assign n10069 = ( n3499 & n8242 ) | ( n3499 & ~n10068 ) | ( n8242 & ~n10068 ) ;
  assign n10070 = n9058 ^ n4115 ^ 1'b0 ;
  assign n10071 = n10069 | n10070 ;
  assign n10072 = n807 & ~n2425 ;
  assign n10073 = n10072 ^ n1600 ^ 1'b0 ;
  assign n10074 = n9475 ^ n7526 ^ n3394 ;
  assign n10075 = n10074 ^ n5129 ^ n800 ;
  assign n10076 = n2491 | n8782 ;
  assign n10077 = ( n369 & n3742 ) | ( n369 & ~n5206 ) | ( n3742 & ~n5206 ) ;
  assign n10078 = ~n5041 & n5211 ;
  assign n10079 = n10078 ^ n3600 ^ 1'b0 ;
  assign n10080 = n10079 ^ n4647 ^ 1'b0 ;
  assign n10081 = n6787 & n10080 ;
  assign n10082 = n791 & n10081 ;
  assign n10083 = ~n289 & n2420 ;
  assign n10084 = n804 & n10083 ;
  assign n10087 = ~n5713 & n5729 ;
  assign n10085 = ( n1899 & n5643 ) | ( n1899 & ~n7710 ) | ( n5643 & ~n7710 ) ;
  assign n10086 = n6984 & n10085 ;
  assign n10088 = n10087 ^ n10086 ^ 1'b0 ;
  assign n10089 = n10084 | n10088 ;
  assign n10090 = n7930 & ~n10089 ;
  assign n10091 = n180 & n3325 ;
  assign n10092 = n1250 & n10091 ;
  assign n10093 = n1360 & ~n4198 ;
  assign n10094 = n10093 ^ n6835 ^ 1'b0 ;
  assign n10095 = n6987 & n10094 ;
  assign n10096 = ( n5436 & n10092 ) | ( n5436 & ~n10095 ) | ( n10092 & ~n10095 ) ;
  assign n10097 = n1238 | n1282 ;
  assign n10098 = n1230 & ~n10097 ;
  assign n10099 = n10098 ^ n4781 ^ 1'b0 ;
  assign n10100 = n10099 ^ n2565 ^ 1'b0 ;
  assign n10101 = n8865 ^ n5016 ^ 1'b0 ;
  assign n10102 = n3671 & ~n4083 ;
  assign n10103 = n10102 ^ n3420 ^ 1'b0 ;
  assign n10104 = ( n1426 & ~n6150 ) | ( n1426 & n7613 ) | ( ~n6150 & n7613 ) ;
  assign n10105 = n10104 ^ n7832 ^ 1'b0 ;
  assign n10106 = ( n10101 & n10103 ) | ( n10101 & n10105 ) | ( n10103 & n10105 ) ;
  assign n10107 = n5323 ^ n168 ^ 1'b0 ;
  assign n10108 = n2177 & ~n10107 ;
  assign n10109 = n10108 ^ n9341 ^ 1'b0 ;
  assign n10110 = n10109 ^ n5362 ^ 1'b0 ;
  assign n10111 = n1279 & ~n10110 ;
  assign n10112 = n10111 ^ n2363 ^ 1'b0 ;
  assign n10113 = n5304 ^ n305 ^ 1'b0 ;
  assign n10114 = n9269 & ~n10113 ;
  assign n10115 = n1219 | n5408 ;
  assign n10116 = n10115 ^ n1363 ^ 1'b0 ;
  assign n10117 = ( ~n6551 & n7682 ) | ( ~n6551 & n10116 ) | ( n7682 & n10116 ) ;
  assign n10118 = ( n2458 & n2615 ) | ( n2458 & n4578 ) | ( n2615 & n4578 ) ;
  assign n10119 = n4576 | n10118 ;
  assign n10120 = n5345 & ~n10119 ;
  assign n10121 = n6948 ^ n2129 ^ 1'b0 ;
  assign n10122 = ( n5713 & ~n6953 ) | ( n5713 & n10121 ) | ( ~n6953 & n10121 ) ;
  assign n10123 = n6153 & n10122 ;
  assign n10124 = n10123 ^ n2766 ^ n1575 ;
  assign n10128 = n8997 ^ n5780 ^ 1'b0 ;
  assign n10125 = n646 | n3374 ;
  assign n10126 = n10125 ^ n5311 ^ 1'b0 ;
  assign n10127 = n1769 | n10126 ;
  assign n10129 = n10128 ^ n10127 ^ n3734 ;
  assign n10130 = ~n2859 & n7432 ;
  assign n10131 = ( n1545 & n3947 ) | ( n1545 & n8458 ) | ( n3947 & n8458 ) ;
  assign n10132 = n1287 ^ n994 ^ 1'b0 ;
  assign n10133 = n1861 ^ n162 ^ 1'b0 ;
  assign n10134 = n2544 | n10133 ;
  assign n10135 = n10134 ^ n9716 ^ 1'b0 ;
  assign n10136 = ( x61 & n4030 ) | ( x61 & ~n4418 ) | ( n4030 & ~n4418 ) ;
  assign n10137 = ~n4006 & n6963 ;
  assign n10138 = n10137 ^ n4574 ^ n1645 ;
  assign n10139 = n9649 ^ n9620 ^ n318 ;
  assign n10140 = n2460 ^ n1804 ^ x21 ;
  assign n10141 = n5909 ^ n5521 ^ n4778 ;
  assign n10142 = ~n10140 & n10141 ;
  assign n10143 = ~n9106 & n10142 ;
  assign n10144 = n9464 & n10143 ;
  assign n10145 = n3921 ^ n2923 ^ 1'b0 ;
  assign n10146 = n9664 ^ n4066 ^ 1'b0 ;
  assign n10147 = n8801 | n10146 ;
  assign n10148 = n2319 & ~n2465 ;
  assign n10149 = n8954 ^ n5093 ^ 1'b0 ;
  assign n10150 = ( n9513 & n10148 ) | ( n9513 & ~n10149 ) | ( n10148 & ~n10149 ) ;
  assign n10156 = n5543 ^ n2732 ^ 1'b0 ;
  assign n10154 = n4944 ^ n2763 ^ 1'b0 ;
  assign n10155 = n1219 | n10154 ;
  assign n10157 = n10156 ^ n10155 ^ 1'b0 ;
  assign n10151 = n4322 | n9773 ;
  assign n10152 = n5967 | n10151 ;
  assign n10153 = ~n372 & n10152 ;
  assign n10158 = n10157 ^ n10153 ^ n8979 ;
  assign n10159 = ( n1410 & n1894 ) | ( n1410 & n2153 ) | ( n1894 & n2153 ) ;
  assign n10160 = n10159 ^ n3895 ^ n388 ;
  assign n10161 = n10160 ^ n5872 ^ n567 ;
  assign n10162 = n10161 ^ n4717 ^ n1217 ;
  assign n10163 = n7999 & ~n9079 ;
  assign n10164 = ~n10162 & n10163 ;
  assign n10165 = ~n3527 & n8454 ;
  assign n10166 = n1018 ^ n972 ^ n819 ;
  assign n10167 = n10166 ^ n4002 ^ 1'b0 ;
  assign n10168 = ~n2317 & n10167 ;
  assign n10169 = ( n5644 & n10165 ) | ( n5644 & ~n10168 ) | ( n10165 & ~n10168 ) ;
  assign n10176 = ( n467 & n1574 ) | ( n467 & ~n7812 ) | ( n1574 & ~n7812 ) ;
  assign n10171 = ~n1240 & n4162 ;
  assign n10172 = n10171 ^ n3332 ^ 1'b0 ;
  assign n10173 = n2036 & ~n10172 ;
  assign n10174 = ~n1850 & n10173 ;
  assign n10170 = n1984 | n9442 ;
  assign n10175 = n10174 ^ n10170 ^ 1'b0 ;
  assign n10177 = n10176 ^ n10175 ^ n2232 ;
  assign n10178 = n2044 & ~n4237 ;
  assign n10179 = n413 & ~n7611 ;
  assign n10180 = ( x52 & ~n3074 ) | ( x52 & n4745 ) | ( ~n3074 & n4745 ) ;
  assign n10181 = ~n6092 & n10180 ;
  assign n10182 = ( n2895 & n6233 ) | ( n2895 & n10181 ) | ( n6233 & n10181 ) ;
  assign n10183 = ( n3406 & n10179 ) | ( n3406 & n10182 ) | ( n10179 & n10182 ) ;
  assign n10184 = ~n7487 & n10183 ;
  assign n10185 = n9965 ^ n4192 ^ 1'b0 ;
  assign n10186 = n4932 ^ n3551 ^ n3504 ;
  assign n10187 = ~n8704 & n9876 ;
  assign n10188 = x7 & ~n10187 ;
  assign n10189 = n10188 ^ n314 ^ 1'b0 ;
  assign n10190 = ( n3489 & n7141 ) | ( n3489 & n7711 ) | ( n7141 & n7711 ) ;
  assign n10191 = n10190 ^ n4081 ^ 1'b0 ;
  assign n10194 = n2865 | n3354 ;
  assign n10195 = n10194 ^ n1801 ^ 1'b0 ;
  assign n10193 = n2569 & n4270 ;
  assign n10192 = n2267 ^ n401 ^ n305 ;
  assign n10196 = n10195 ^ n10193 ^ n10192 ;
  assign n10197 = n10196 ^ n3698 ^ n1202 ;
  assign n10198 = n2377 | n5913 ;
  assign n10199 = n5925 | n10198 ;
  assign n10200 = n8036 ^ n3398 ^ 1'b0 ;
  assign n10201 = n10200 ^ n5817 ^ 1'b0 ;
  assign n10202 = n2539 & n10201 ;
  assign n10203 = n10202 ^ n8830 ^ 1'b0 ;
  assign n10204 = n7917 & ~n7959 ;
  assign n10205 = n3293 | n10204 ;
  assign n10206 = n6410 ^ n6095 ^ n3842 ;
  assign n10207 = ~n6217 & n10206 ;
  assign n10208 = n5929 ^ n5639 ^ 1'b0 ;
  assign n10209 = n8196 | n10208 ;
  assign n10210 = n3169 ^ n2709 ^ 1'b0 ;
  assign n10211 = n2522 | n10210 ;
  assign n10212 = n4230 & ~n10211 ;
  assign n10213 = n9820 | n10212 ;
  assign n10214 = n1993 ^ n1867 ^ n1683 ;
  assign n10215 = ~n1015 & n4627 ;
  assign n10216 = ~n10214 & n10215 ;
  assign n10217 = n8836 ^ n971 ^ 1'b0 ;
  assign n10218 = n10216 | n10217 ;
  assign n10219 = n1802 ^ n1025 ^ 1'b0 ;
  assign n10220 = n831 | n10219 ;
  assign n10221 = n10218 & n10220 ;
  assign n10222 = ~n8081 & n10221 ;
  assign n10223 = n3228 ^ n1345 ^ 1'b0 ;
  assign n10224 = n4329 & ~n10223 ;
  assign n10225 = ( n2897 & ~n4089 ) | ( n2897 & n9626 ) | ( ~n4089 & n9626 ) ;
  assign n10226 = n468 | n10225 ;
  assign n10227 = n10224 | n10226 ;
  assign n10228 = n6705 | n6851 ;
  assign n10229 = n10228 ^ n9272 ^ 1'b0 ;
  assign n10230 = n7629 ^ n6616 ^ 1'b0 ;
  assign n10231 = n5607 ^ n1860 ^ n1143 ;
  assign n10232 = n10231 ^ n7639 ^ n5689 ;
  assign n10234 = ( n2149 & n2423 ) | ( n2149 & n7064 ) | ( n2423 & n7064 ) ;
  assign n10233 = n2036 & n5326 ;
  assign n10235 = n10234 ^ n10233 ^ 1'b0 ;
  assign n10236 = n3379 & ~n10235 ;
  assign n10237 = ( ~n4624 & n6889 ) | ( ~n4624 & n7024 ) | ( n6889 & n7024 ) ;
  assign n10238 = n1252 | n7682 ;
  assign n10239 = n1693 & n3420 ;
  assign n10240 = n3424 ^ n1978 ^ n486 ;
  assign n10241 = n10240 ^ n9151 ^ 1'b0 ;
  assign n10242 = n6196 & n10241 ;
  assign n10243 = n10242 ^ n1387 ^ 1'b0 ;
  assign n10244 = n10239 & n10243 ;
  assign n10246 = n272 | n7806 ;
  assign n10247 = n10246 ^ n3582 ^ 1'b0 ;
  assign n10248 = ( n260 & n466 ) | ( n260 & n10247 ) | ( n466 & n10247 ) ;
  assign n10249 = ~n1190 & n10248 ;
  assign n10245 = ~n5041 & n7866 ;
  assign n10250 = n10249 ^ n10245 ^ 1'b0 ;
  assign n10251 = ( n1178 & n6946 ) | ( n1178 & n10250 ) | ( n6946 & n10250 ) ;
  assign n10253 = ( n1283 & ~n3784 ) | ( n1283 & n7355 ) | ( ~n3784 & n7355 ) ;
  assign n10254 = ~n4199 & n10253 ;
  assign n10255 = n10254 ^ x115 ^ 1'b0 ;
  assign n10256 = n10255 ^ n6101 ^ 1'b0 ;
  assign n10252 = ~n5316 & n9955 ;
  assign n10257 = n10256 ^ n10252 ^ n5171 ;
  assign n10263 = n2870 ^ n2618 ^ n1799 ;
  assign n10264 = n1915 | n10263 ;
  assign n10258 = n5414 ^ n1837 ^ 1'b0 ;
  assign n10259 = n10258 ^ n2388 ^ 1'b0 ;
  assign n10260 = n10259 ^ n8042 ^ n1043 ;
  assign n10261 = n10260 ^ n153 ^ 1'b0 ;
  assign n10262 = ~n1316 & n10261 ;
  assign n10265 = n10264 ^ n10262 ^ 1'b0 ;
  assign n10266 = n3319 ^ n2823 ^ n1301 ;
  assign n10267 = n10266 ^ n3560 ^ n478 ;
  assign n10268 = ~n5445 & n9777 ;
  assign n10269 = n10268 ^ n2098 ^ 1'b0 ;
  assign n10270 = n5336 ^ n916 ^ n664 ;
  assign n10271 = n10270 ^ n3573 ^ n1632 ;
  assign n10275 = n7141 ^ n3565 ^ 1'b0 ;
  assign n10272 = n3548 ^ n940 ^ 1'b0 ;
  assign n10273 = n10272 ^ n3410 ^ n2524 ;
  assign n10274 = n2140 & ~n10273 ;
  assign n10276 = n10275 ^ n10274 ^ 1'b0 ;
  assign n10277 = ~n10271 & n10276 ;
  assign n10278 = ( ~n2738 & n7068 ) | ( ~n2738 & n8238 ) | ( n7068 & n8238 ) ;
  assign n10279 = n8323 & n8534 ;
  assign n10280 = n522 & n1920 ;
  assign n10281 = ( ~n3242 & n5094 ) | ( ~n3242 & n6172 ) | ( n5094 & n6172 ) ;
  assign n10282 = n7909 ^ n4735 ^ 1'b0 ;
  assign n10283 = n9714 ^ n3744 ^ n1922 ;
  assign n10284 = n1600 & ~n1710 ;
  assign n10285 = n2067 & n4162 ;
  assign n10286 = n10285 ^ n7523 ^ n2334 ;
  assign n10289 = n2220 ^ n1405 ^ n696 ;
  assign n10290 = ( ~n2764 & n4163 ) | ( ~n2764 & n10289 ) | ( n4163 & n10289 ) ;
  assign n10291 = n10290 ^ n1076 ^ 1'b0 ;
  assign n10287 = n2660 & n7232 ;
  assign n10288 = ~n5629 & n10287 ;
  assign n10292 = n10291 ^ n10288 ^ 1'b0 ;
  assign n10293 = ~n10286 & n10292 ;
  assign n10294 = n171 & n1385 ;
  assign n10295 = n10294 ^ n2469 ^ 1'b0 ;
  assign n10296 = n2079 | n4948 ;
  assign n10297 = n10295 & ~n10296 ;
  assign n10298 = ~n2110 & n9799 ;
  assign n10299 = ~x54 & n10298 ;
  assign n10300 = ( n9698 & n10297 ) | ( n9698 & ~n10299 ) | ( n10297 & ~n10299 ) ;
  assign n10301 = n9608 ^ n6668 ^ n6347 ;
  assign n10302 = ~n2978 & n5962 ;
  assign n10303 = n3636 ^ n452 ^ 1'b0 ;
  assign n10304 = ~n1037 & n10303 ;
  assign n10308 = ( ~n1011 & n3128 ) | ( ~n1011 & n5982 ) | ( n3128 & n5982 ) ;
  assign n10305 = ~n1586 & n4849 ;
  assign n10306 = ~n5493 & n10305 ;
  assign n10307 = n4837 & ~n10306 ;
  assign n10309 = n10308 ^ n10307 ^ 1'b0 ;
  assign n10310 = n641 | n5224 ;
  assign n10311 = n4957 | n10310 ;
  assign n10312 = n10311 ^ x1 ^ 1'b0 ;
  assign n10313 = n10309 & n10312 ;
  assign n10314 = n8225 ^ n6585 ^ 1'b0 ;
  assign n10315 = n10314 ^ n9106 ^ n4336 ;
  assign n10316 = n1308 & ~n7721 ;
  assign n10320 = n4094 ^ n3204 ^ 1'b0 ;
  assign n10317 = n3326 & n5454 ;
  assign n10318 = n8662 ^ n5900 ^ n232 ;
  assign n10319 = n10317 | n10318 ;
  assign n10321 = n10320 ^ n10319 ^ 1'b0 ;
  assign n10322 = n5654 & n10321 ;
  assign n10323 = n8008 & ~n10322 ;
  assign n10324 = ~n1126 & n10323 ;
  assign n10325 = n6486 & ~n6957 ;
  assign n10326 = n10325 ^ n4510 ^ 1'b0 ;
  assign n10327 = ( n4506 & n4642 ) | ( n4506 & ~n7838 ) | ( n4642 & ~n7838 ) ;
  assign n10328 = n7455 & n10327 ;
  assign n10329 = n10328 ^ n1656 ^ 1'b0 ;
  assign n10330 = x50 & ~n10329 ;
  assign n10331 = n10330 ^ n9266 ^ n4921 ;
  assign n10332 = ~n4497 & n10331 ;
  assign n10333 = n3333 & ~n4814 ;
  assign n10334 = x1 | n6353 ;
  assign n10335 = n5225 | n10334 ;
  assign n10336 = n10335 ^ n3498 ^ 1'b0 ;
  assign n10337 = ( n2417 & n4830 ) | ( n2417 & ~n10336 ) | ( n4830 & ~n10336 ) ;
  assign n10338 = n4462 ^ n980 ^ 1'b0 ;
  assign n10339 = n3355 | n10338 ;
  assign n10340 = n4214 | n7155 ;
  assign n10341 = n4125 | n10340 ;
  assign n10343 = n7791 ^ n4021 ^ 1'b0 ;
  assign n10342 = ( ~n1096 & n6148 ) | ( ~n1096 & n6604 ) | ( n6148 & n6604 ) ;
  assign n10344 = n10343 ^ n10342 ^ 1'b0 ;
  assign n10345 = n10341 & ~n10344 ;
  assign n10351 = n3314 ^ n2107 ^ 1'b0 ;
  assign n10348 = ~n4597 & n8336 ;
  assign n10347 = n255 & ~n3100 ;
  assign n10349 = n10348 ^ n10347 ^ 1'b0 ;
  assign n10350 = n10349 ^ x30 ^ 1'b0 ;
  assign n10346 = n4199 ^ n1092 ^ 1'b0 ;
  assign n10352 = n10351 ^ n10350 ^ n10346 ;
  assign n10353 = ( n1019 & ~n2858 ) | ( n1019 & n3484 ) | ( ~n2858 & n3484 ) ;
  assign n10354 = n10353 ^ n6562 ^ n5630 ;
  assign n10355 = n3124 & ~n7053 ;
  assign n10356 = n10354 & n10355 ;
  assign n10357 = n5711 & n10356 ;
  assign n10358 = n449 & n2756 ;
  assign n10359 = n3956 & n10358 ;
  assign n10360 = n5480 | n10359 ;
  assign n10361 = ( ~n4100 & n10357 ) | ( ~n4100 & n10360 ) | ( n10357 & n10360 ) ;
  assign n10362 = n1800 ^ n917 ^ 1'b0 ;
  assign n10363 = n4742 ^ n2497 ^ 1'b0 ;
  assign n10364 = n357 & ~n10363 ;
  assign n10365 = ~n2104 & n8065 ;
  assign n10366 = ~n10364 & n10365 ;
  assign n10367 = ~n466 & n2756 ;
  assign n10368 = ~n2022 & n10367 ;
  assign n10373 = n1785 ^ n1572 ^ n699 ;
  assign n10374 = ( n486 & ~n2036 ) | ( n486 & n10373 ) | ( ~n2036 & n10373 ) ;
  assign n10369 = n2179 ^ n1204 ^ 1'b0 ;
  assign n10370 = n5616 | n10369 ;
  assign n10371 = n4543 ^ n505 ^ 1'b0 ;
  assign n10372 = ~n10370 & n10371 ;
  assign n10375 = n10374 ^ n10372 ^ 1'b0 ;
  assign n10376 = n10368 | n10375 ;
  assign n10377 = n2906 & ~n10376 ;
  assign n10378 = ~n4415 & n10377 ;
  assign n10379 = n8234 ^ n2652 ^ n1034 ;
  assign n10381 = n156 & n3443 ;
  assign n10382 = n10381 ^ n6368 ^ 1'b0 ;
  assign n10380 = n10125 ^ n8943 ^ n6451 ;
  assign n10383 = n10382 ^ n10380 ^ 1'b0 ;
  assign n10384 = n3354 & ~n10383 ;
  assign n10385 = n4987 ^ n3213 ^ 1'b0 ;
  assign n10386 = ~n798 & n10385 ;
  assign n10387 = n7623 ^ n3964 ^ 1'b0 ;
  assign n10388 = n339 & n10387 ;
  assign n10389 = ~n10386 & n10388 ;
  assign n10390 = n10384 | n10389 ;
  assign n10391 = n9475 ^ n9090 ^ n2211 ;
  assign n10392 = n10391 ^ n6862 ^ n3314 ;
  assign n10393 = n10392 ^ n6022 ^ n5730 ;
  assign n10394 = n182 & n4706 ;
  assign n10395 = ( n2027 & n8301 ) | ( n2027 & ~n10394 ) | ( n8301 & ~n10394 ) ;
  assign n10396 = n5436 & ~n10395 ;
  assign n10397 = n7071 ^ n3829 ^ 1'b0 ;
  assign n10398 = n4696 & ~n10397 ;
  assign n10399 = ~n7110 & n10398 ;
  assign n10400 = n10399 ^ x86 ^ 1'b0 ;
  assign n10401 = n10400 ^ n552 ^ 1'b0 ;
  assign n10402 = n964 & n5605 ;
  assign n10403 = n5799 ^ n2621 ^ 1'b0 ;
  assign n10404 = n8552 & ~n10403 ;
  assign n10405 = n9482 ^ n5353 ^ 1'b0 ;
  assign n10406 = n6879 ^ n6829 ^ n1357 ;
  assign n10407 = ( n464 & n1555 ) | ( n464 & n3207 ) | ( n1555 & n3207 ) ;
  assign n10408 = n5044 | n10407 ;
  assign n10409 = n10408 ^ n4722 ^ 1'b0 ;
  assign n10410 = ~n10406 & n10409 ;
  assign n10411 = ( ~n919 & n3437 ) | ( ~n919 & n8746 ) | ( n3437 & n8746 ) ;
  assign n10412 = ( n285 & ~n6920 ) | ( n285 & n10411 ) | ( ~n6920 & n10411 ) ;
  assign n10413 = n10412 ^ n8563 ^ 1'b0 ;
  assign n10414 = n2335 ^ n643 ^ x67 ;
  assign n10415 = n8827 & ~n9063 ;
  assign n10416 = ( n2662 & ~n10414 ) | ( n2662 & n10415 ) | ( ~n10414 & n10415 ) ;
  assign n10417 = n10191 ^ n3826 ^ n1668 ;
  assign n10418 = n2788 & n5630 ;
  assign n10419 = n318 & n3640 ;
  assign n10420 = ( n3471 & n3660 ) | ( n3471 & ~n10419 ) | ( n3660 & ~n10419 ) ;
  assign n10421 = n10420 ^ n8439 ^ 1'b0 ;
  assign n10422 = ~n8024 & n10421 ;
  assign n10423 = n10422 ^ n5179 ^ 1'b0 ;
  assign n10424 = n10418 & n10423 ;
  assign n10430 = ~n4058 & n9962 ;
  assign n10431 = ~n5371 & n10430 ;
  assign n10432 = n10431 ^ n9363 ^ n2722 ;
  assign n10425 = n5502 ^ n1159 ^ n497 ;
  assign n10426 = ( ~n516 & n4752 ) | ( ~n516 & n6085 ) | ( n4752 & n6085 ) ;
  assign n10427 = n10426 ^ n1321 ^ n708 ;
  assign n10428 = ( ~n6092 & n10425 ) | ( ~n6092 & n10427 ) | ( n10425 & n10427 ) ;
  assign n10429 = ~n5227 & n10428 ;
  assign n10433 = n10432 ^ n10429 ^ 1'b0 ;
  assign n10434 = n10433 ^ n6781 ^ 1'b0 ;
  assign n10435 = ( n2757 & ~n7002 ) | ( n2757 & n10434 ) | ( ~n7002 & n10434 ) ;
  assign n10436 = ( n4619 & ~n5154 ) | ( n4619 & n5866 ) | ( ~n5154 & n5866 ) ;
  assign n10437 = ~n5338 & n8305 ;
  assign n10439 = ( x64 & ~n1791 ) | ( x64 & n9660 ) | ( ~n1791 & n9660 ) ;
  assign n10438 = x88 & ~n6390 ;
  assign n10440 = n10439 ^ n10438 ^ 1'b0 ;
  assign n10441 = n10440 ^ n7388 ^ 1'b0 ;
  assign n10442 = n10023 | n10441 ;
  assign n10443 = ( n967 & n3473 ) | ( n967 & ~n4952 ) | ( n3473 & ~n4952 ) ;
  assign n10444 = n10443 ^ n7374 ^ 1'b0 ;
  assign n10445 = n920 & n10444 ;
  assign n10447 = ( n935 & n4133 ) | ( n935 & ~n6103 ) | ( n4133 & ~n6103 ) ;
  assign n10448 = n10447 ^ n6190 ^ n2901 ;
  assign n10446 = n1996 & ~n5334 ;
  assign n10449 = n10448 ^ n10446 ^ 1'b0 ;
  assign n10450 = ( ~n6153 & n8638 ) | ( ~n6153 & n10449 ) | ( n8638 & n10449 ) ;
  assign n10451 = ( n3293 & ~n5472 ) | ( n3293 & n10216 ) | ( ~n5472 & n10216 ) ;
  assign n10452 = ( ~n4741 & n5898 ) | ( ~n4741 & n10451 ) | ( n5898 & n10451 ) ;
  assign n10453 = ~n10450 & n10452 ;
  assign n10454 = n10445 & n10453 ;
  assign n10455 = ~n2424 & n4305 ;
  assign n10456 = n1090 & n10455 ;
  assign n10457 = n7326 | n10456 ;
  assign n10458 = n1387 & ~n1809 ;
  assign n10459 = ( n685 & n5041 ) | ( n685 & n5071 ) | ( n5041 & n5071 ) ;
  assign n10460 = n10459 ^ n4080 ^ n2642 ;
  assign n10461 = n7536 ^ n477 ^ 1'b0 ;
  assign n10462 = n10460 & n10461 ;
  assign n10463 = n5096 & ~n10462 ;
  assign n10464 = n2561 | n2682 ;
  assign n10465 = n10463 & ~n10464 ;
  assign n10466 = ( ~n6221 & n10458 ) | ( ~n6221 & n10465 ) | ( n10458 & n10465 ) ;
  assign n10467 = ( x47 & ~n1456 ) | ( x47 & n3416 ) | ( ~n1456 & n3416 ) ;
  assign n10468 = n3382 ^ n1828 ^ 1'b0 ;
  assign n10469 = n10467 | n10468 ;
  assign n10470 = n3001 & ~n10469 ;
  assign n10471 = n10470 ^ n5425 ^ 1'b0 ;
  assign n10472 = n7994 & ~n8466 ;
  assign n10473 = ~n738 & n1581 ;
  assign n10474 = ~n209 & n10473 ;
  assign n10475 = n10474 ^ n784 ^ x28 ;
  assign n10476 = n10475 ^ n5018 ^ n2944 ;
  assign n10477 = n2884 ^ n851 ^ n739 ;
  assign n10478 = n10477 ^ n257 ^ 1'b0 ;
  assign n10479 = n7729 ^ n4177 ^ 1'b0 ;
  assign n10480 = ~n8214 & n10479 ;
  assign n10481 = ~n5839 & n10480 ;
  assign n10482 = n2097 & n10481 ;
  assign n10483 = n7340 & n10482 ;
  assign n10484 = n9045 ^ n7353 ^ 1'b0 ;
  assign n10485 = ~n7219 & n10484 ;
  assign n10486 = ( n3815 & n9522 ) | ( n3815 & n10485 ) | ( n9522 & n10485 ) ;
  assign n10493 = ~n2207 & n8867 ;
  assign n10494 = n4509 & n10493 ;
  assign n10492 = n5561 & ~n8020 ;
  assign n10487 = n170 & ~n9691 ;
  assign n10488 = n1692 & n10487 ;
  assign n10489 = n1397 & n5909 ;
  assign n10490 = n10489 ^ x123 ^ 1'b0 ;
  assign n10491 = ~n10488 & n10490 ;
  assign n10495 = n10494 ^ n10492 ^ n10491 ;
  assign n10498 = n7200 ^ n5516 ^ 1'b0 ;
  assign n10499 = n6803 | n10498 ;
  assign n10496 = ~n4142 & n4217 ;
  assign n10497 = n10496 ^ n10193 ^ 1'b0 ;
  assign n10500 = n10499 ^ n10497 ^ n2140 ;
  assign n10501 = ~n6790 & n10500 ;
  assign n10502 = n1023 & ~n2195 ;
  assign n10503 = n10502 ^ n775 ^ 1'b0 ;
  assign n10504 = n10503 ^ n1493 ^ n270 ;
  assign n10505 = x16 & n4052 ;
  assign n10506 = n10505 ^ n6896 ^ 1'b0 ;
  assign n10507 = n862 & ~n1588 ;
  assign n10508 = n10506 & n10507 ;
  assign n10509 = n10508 ^ n194 ^ 1'b0 ;
  assign n10510 = n6498 & n10509 ;
  assign n10511 = n10510 ^ n523 ^ 1'b0 ;
  assign n10512 = n4194 & ~n10511 ;
  assign n10513 = n1692 ^ x126 ^ 1'b0 ;
  assign n10514 = ( ~n1223 & n10481 ) | ( ~n1223 & n10513 ) | ( n10481 & n10513 ) ;
  assign n10515 = n460 | n10514 ;
  assign n10516 = ( n1244 & n1385 ) | ( n1244 & n5822 ) | ( n1385 & n5822 ) ;
  assign n10517 = n10516 ^ n6668 ^ n2018 ;
  assign n10518 = ( n3315 & ~n10056 ) | ( n3315 & n10317 ) | ( ~n10056 & n10317 ) ;
  assign n10519 = ~n3661 & n10518 ;
  assign n10520 = n10519 ^ n5143 ^ 1'b0 ;
  assign n10521 = n10517 | n10520 ;
  assign n10522 = n4857 ^ n3238 ^ 1'b0 ;
  assign n10523 = ( x65 & n1223 ) | ( x65 & ~n3605 ) | ( n1223 & ~n3605 ) ;
  assign n10524 = n4477 & n8896 ;
  assign n10525 = ~n897 & n1041 ;
  assign n10526 = n1912 & n3290 ;
  assign n10527 = n10526 ^ n4280 ^ 1'b0 ;
  assign n10528 = n8007 | n10527 ;
  assign n10529 = n9506 ^ n1032 ^ 1'b0 ;
  assign n10530 = n2098 & ~n2499 ;
  assign n10531 = n10529 & n10530 ;
  assign n10532 = n10528 & n10531 ;
  assign n10533 = n1229 & ~n2965 ;
  assign n10534 = n10533 ^ n955 ^ 1'b0 ;
  assign n10535 = n2887 | n10534 ;
  assign n10538 = ( n1234 & n5665 ) | ( n1234 & n8151 ) | ( n5665 & n8151 ) ;
  assign n10536 = n4613 ^ n1986 ^ n283 ;
  assign n10537 = ( x103 & n3566 ) | ( x103 & ~n10536 ) | ( n3566 & ~n10536 ) ;
  assign n10539 = n10538 ^ n10537 ^ 1'b0 ;
  assign n10540 = n10539 ^ n357 ^ 1'b0 ;
  assign n10541 = n8298 & n10540 ;
  assign n10542 = ( n3806 & n10535 ) | ( n3806 & n10541 ) | ( n10535 & n10541 ) ;
  assign n10543 = n4144 ^ n919 ^ 1'b0 ;
  assign n10544 = n10543 ^ n3459 ^ 1'b0 ;
  assign n10545 = n6674 ^ n1454 ^ n331 ;
  assign n10546 = n6750 ^ n3035 ^ 1'b0 ;
  assign n10547 = n10299 | n10546 ;
  assign n10548 = n10545 & n10547 ;
  assign n10549 = ( ~n1849 & n5336 ) | ( ~n1849 & n6306 ) | ( n5336 & n6306 ) ;
  assign n10550 = n3475 & n10549 ;
  assign n10551 = n3401 & n10550 ;
  assign n10552 = n586 & ~n10551 ;
  assign n10553 = n7076 | n8475 ;
  assign n10554 = n3639 ^ n3471 ^ n3378 ;
  assign n10555 = n1769 & n5082 ;
  assign n10556 = ( n4180 & ~n10554 ) | ( n4180 & n10555 ) | ( ~n10554 & n10555 ) ;
  assign n10557 = ~n3666 & n8250 ;
  assign n10558 = n3401 ^ n3174 ^ 1'b0 ;
  assign n10559 = n8129 | n10558 ;
  assign n10560 = n10557 & ~n10559 ;
  assign n10561 = n958 ^ n925 ^ 1'b0 ;
  assign n10562 = n8293 & n10561 ;
  assign n10563 = n10562 ^ n3432 ^ 1'b0 ;
  assign n10564 = ~n3051 & n10563 ;
  assign n10565 = n2675 & ~n10564 ;
  assign n10566 = ( ~n1274 & n6144 ) | ( ~n1274 & n10565 ) | ( n6144 & n10565 ) ;
  assign n10567 = n9866 ^ n4905 ^ x59 ;
  assign n10568 = n3975 & ~n4484 ;
  assign n10569 = n2735 | n2748 ;
  assign n10570 = n8333 | n9002 ;
  assign n10571 = n633 & ~n7219 ;
  assign n10572 = n2914 | n10571 ;
  assign n10573 = n9673 ^ n4792 ^ n4413 ;
  assign n10574 = n7654 ^ n3990 ^ 1'b0 ;
  assign n10575 = n6843 & ~n10574 ;
  assign n10576 = n9177 & n10575 ;
  assign n10577 = n10576 ^ n4566 ^ 1'b0 ;
  assign n10578 = n8417 ^ n4075 ^ n3256 ;
  assign n10579 = n6640 ^ n5276 ^ 1'b0 ;
  assign n10580 = ~n3324 & n10579 ;
  assign n10581 = n151 & ~n10580 ;
  assign n10582 = n10463 & n10581 ;
  assign n10589 = n2823 & n9605 ;
  assign n10590 = n2720 & n10589 ;
  assign n10585 = ( ~n191 & n1067 ) | ( ~n191 & n4772 ) | ( n1067 & n4772 ) ;
  assign n10586 = n10585 ^ n7528 ^ n7520 ;
  assign n10583 = n6231 ^ n2929 ^ 1'b0 ;
  assign n10584 = n7043 & ~n10583 ;
  assign n10587 = n10586 ^ n10584 ^ n7306 ;
  assign n10588 = ~n7956 & n10587 ;
  assign n10591 = n10590 ^ n10588 ^ 1'b0 ;
  assign n10592 = n3749 ^ n1771 ^ n1025 ;
  assign n10593 = n10592 ^ n620 ^ 1'b0 ;
  assign n10594 = n10593 ^ n5270 ^ 1'b0 ;
  assign n10596 = n1615 ^ n1198 ^ x57 ;
  assign n10597 = ( n5453 & ~n10419 ) | ( n5453 & n10596 ) | ( ~n10419 & n10596 ) ;
  assign n10595 = n2408 & n10093 ;
  assign n10598 = n10597 ^ n10595 ^ n6685 ;
  assign n10601 = n6324 ^ n4063 ^ n2466 ;
  assign n10599 = ~n3734 & n9733 ;
  assign n10600 = n10599 ^ n4854 ^ n302 ;
  assign n10602 = n10601 ^ n10600 ^ 1'b0 ;
  assign n10603 = n6184 ^ n1464 ^ 1'b0 ;
  assign n10604 = n10602 & n10603 ;
  assign n10605 = ( n807 & n1006 ) | ( n807 & ~n1345 ) | ( n1006 & ~n1345 ) ;
  assign n10606 = n512 & n10605 ;
  assign n10607 = n10606 ^ n646 ^ 1'b0 ;
  assign n10608 = n8519 ^ x42 ^ 1'b0 ;
  assign n10609 = n4914 & ~n10608 ;
  assign n10610 = n10607 | n10609 ;
  assign n10611 = ( x11 & n1289 ) | ( x11 & ~n2463 ) | ( n1289 & ~n2463 ) ;
  assign n10612 = ~n1946 & n10611 ;
  assign n10613 = n9015 & n10612 ;
  assign n10614 = n10613 ^ n8314 ^ 1'b0 ;
  assign n10615 = n10610 & n10614 ;
  assign n10616 = ~n316 & n2744 ;
  assign n10617 = n10616 ^ n6252 ^ n938 ;
  assign n10618 = n4096 ^ n456 ^ 1'b0 ;
  assign n10619 = ~n1939 & n10618 ;
  assign n10620 = ~n6459 & n10619 ;
  assign n10621 = n10620 ^ n7284 ^ 1'b0 ;
  assign n10623 = n5455 ^ n3975 ^ n3186 ;
  assign n10624 = n10623 ^ n5507 ^ n511 ;
  assign n10622 = n7096 ^ n6794 ^ 1'b0 ;
  assign n10625 = n10624 ^ n10622 ^ n2631 ;
  assign n10626 = n7200 & n10625 ;
  assign n10627 = n9023 ^ n6793 ^ n4181 ;
  assign n10628 = n6085 | n10627 ;
  assign n10629 = n2926 | n10628 ;
  assign n10630 = n10629 ^ n6440 ^ 1'b0 ;
  assign n10631 = n10626 & n10630 ;
  assign n10632 = ( ~n6230 & n9845 ) | ( ~n6230 & n10242 ) | ( n9845 & n10242 ) ;
  assign n10634 = ~n6466 & n7233 ;
  assign n10633 = n5272 & ~n8253 ;
  assign n10635 = n10634 ^ n10633 ^ 1'b0 ;
  assign n10636 = n1268 ^ n319 ^ 1'b0 ;
  assign n10637 = n10636 ^ n3620 ^ n878 ;
  assign n10638 = n10637 ^ n9000 ^ 1'b0 ;
  assign n10639 = n3271 | n7754 ;
  assign n10640 = n8074 | n10639 ;
  assign n10641 = n10640 ^ n5771 ^ 1'b0 ;
  assign n10642 = n2060 ^ n1942 ^ 1'b0 ;
  assign n10643 = ( n3778 & n4684 ) | ( n3778 & n10642 ) | ( n4684 & n10642 ) ;
  assign n10644 = n541 & ~n4807 ;
  assign n10645 = n4432 & n10644 ;
  assign n10646 = n10645 ^ n3197 ^ 1'b0 ;
  assign n10647 = ~n573 & n10646 ;
  assign n10648 = ( n3768 & ~n10643 ) | ( n3768 & n10647 ) | ( ~n10643 & n10647 ) ;
  assign n10649 = n3059 & n5332 ;
  assign n10650 = ~n2145 & n10649 ;
  assign n10651 = n10650 ^ n6067 ^ 1'b0 ;
  assign n10652 = n10360 ^ n6989 ^ n4018 ;
  assign n10653 = n10607 ^ n5801 ^ 1'b0 ;
  assign n10654 = n334 & ~n10653 ;
  assign n10655 = ( n1509 & ~n3923 ) | ( n1509 & n10654 ) | ( ~n3923 & n10654 ) ;
  assign n10656 = n3507 ^ n2212 ^ 1'b0 ;
  assign n10657 = x51 & ~n6814 ;
  assign n10658 = n3402 ^ n2756 ^ 1'b0 ;
  assign n10659 = n9748 | n10658 ;
  assign n10660 = ( ~n1409 & n3872 ) | ( ~n1409 & n4593 ) | ( n3872 & n4593 ) ;
  assign n10661 = n1641 & ~n5633 ;
  assign n10662 = n10661 ^ n6180 ^ 1'b0 ;
  assign n10663 = n1767 ^ n390 ^ 1'b0 ;
  assign n10664 = ( ~n416 & n983 ) | ( ~n416 & n10663 ) | ( n983 & n10663 ) ;
  assign n10665 = ( n8762 & n9098 ) | ( n8762 & n10214 ) | ( n9098 & n10214 ) ;
  assign n10673 = n619 & ~n5326 ;
  assign n10674 = n1769 & n10673 ;
  assign n10666 = n2406 & n3968 ;
  assign n10667 = n10666 ^ n1649 ^ 1'b0 ;
  assign n10668 = n10667 ^ n2498 ^ 1'b0 ;
  assign n10669 = n2363 & ~n3178 ;
  assign n10670 = n10427 & n10669 ;
  assign n10671 = n10373 | n10670 ;
  assign n10672 = n10668 & ~n10671 ;
  assign n10675 = n10674 ^ n10672 ^ 1'b0 ;
  assign n10676 = ~n10665 & n10675 ;
  assign n10677 = n1253 | n2090 ;
  assign n10678 = n8577 | n10677 ;
  assign n10679 = n5786 & n10678 ;
  assign n10680 = n533 | n3273 ;
  assign n10681 = n2235 | n10680 ;
  assign n10682 = ~x120 & n10681 ;
  assign n10683 = ~n8748 & n10682 ;
  assign n10684 = n10683 ^ n4743 ^ n2047 ;
  assign n10685 = ( n474 & n1400 ) | ( n474 & ~n6520 ) | ( n1400 & ~n6520 ) ;
  assign n10686 = n6739 ^ n2225 ^ 1'b0 ;
  assign n10689 = n266 | n4825 ;
  assign n10687 = n2342 & n4240 ;
  assign n10688 = ~n8995 & n10687 ;
  assign n10690 = n10689 ^ n10688 ^ 1'b0 ;
  assign n10691 = ~n9495 & n9870 ;
  assign n10692 = n10691 ^ n4978 ^ 1'b0 ;
  assign n10693 = n4020 ^ n2521 ^ 1'b0 ;
  assign n10694 = n1009 & ~n3602 ;
  assign n10695 = n10693 & n10694 ;
  assign n10696 = ~n2347 & n7842 ;
  assign n10697 = ~n1572 & n2369 ;
  assign n10698 = ~n2348 & n10697 ;
  assign n10699 = n9231 ^ n2732 ^ n1754 ;
  assign n10700 = n10699 ^ n6609 ^ n4710 ;
  assign n10701 = n10700 ^ n5382 ^ n1537 ;
  assign n10702 = ~n10698 & n10701 ;
  assign n10703 = n4343 & n10702 ;
  assign n10704 = n6206 ^ n2116 ^ n1962 ;
  assign n10705 = n10704 ^ n6409 ^ 1'b0 ;
  assign n10706 = n10443 & n10705 ;
  assign n10707 = ( n3503 & ~n6787 ) | ( n3503 & n10706 ) | ( ~n6787 & n10706 ) ;
  assign n10708 = n4212 & ~n10707 ;
  assign n10709 = n10708 ^ n5748 ^ n4641 ;
  assign n10710 = n9274 ^ n6172 ^ 1'b0 ;
  assign n10715 = n1622 & n4761 ;
  assign n10716 = ( ~n327 & n8658 ) | ( ~n327 & n10715 ) | ( n8658 & n10715 ) ;
  assign n10711 = n8451 ^ n851 ^ 1'b0 ;
  assign n10712 = n4371 & ~n10711 ;
  assign n10713 = n10712 ^ n319 ^ 1'b0 ;
  assign n10714 = ( n1732 & n6831 ) | ( n1732 & ~n10713 ) | ( n6831 & ~n10713 ) ;
  assign n10717 = n10716 ^ n10714 ^ n4138 ;
  assign n10718 = n4059 & n4897 ;
  assign n10719 = n756 ^ n550 ^ x83 ;
  assign n10720 = n10719 ^ n8224 ^ n714 ;
  assign n10721 = n10720 ^ n5025 ^ n3838 ;
  assign n10722 = ( ~n4594 & n9801 ) | ( ~n4594 & n10414 ) | ( n9801 & n10414 ) ;
  assign n10723 = n2235 & ~n10722 ;
  assign n10724 = ~n6649 & n10723 ;
  assign n10725 = n10721 | n10724 ;
  assign n10726 = n10725 ^ n8408 ^ 1'b0 ;
  assign n10727 = ~n3488 & n4254 ;
  assign n10728 = n9446 | n10450 ;
  assign n10729 = n2929 & ~n10728 ;
  assign n10730 = ( ~n547 & n5906 ) | ( ~n547 & n8995 ) | ( n5906 & n8995 ) ;
  assign n10731 = ~n3073 & n10730 ;
  assign n10732 = ( n3111 & n5924 ) | ( n3111 & ~n10731 ) | ( n5924 & ~n10731 ) ;
  assign n10733 = n10732 ^ n2157 ^ n1769 ;
  assign n10734 = n4686 ^ n2914 ^ 1'b0 ;
  assign n10735 = ~n1653 & n4904 ;
  assign n10736 = n2036 & ~n10735 ;
  assign n10737 = n10373 ^ n6261 ^ 1'b0 ;
  assign n10738 = n4530 & ~n10737 ;
  assign n10739 = n6121 ^ n3161 ^ 1'b0 ;
  assign n10740 = ~n10177 & n10739 ;
  assign n10741 = n4715 ^ n2567 ^ 1'b0 ;
  assign n10742 = ~n2211 & n10741 ;
  assign n10743 = n3964 & n10742 ;
  assign n10744 = n6026 & n10743 ;
  assign n10745 = n10744 ^ n4546 ^ n2865 ;
  assign n10746 = n10346 ^ n266 ^ 1'b0 ;
  assign n10747 = ~n993 & n10527 ;
  assign n10748 = ~n8240 & n10747 ;
  assign n10749 = ( n1072 & n2207 ) | ( n1072 & n3829 ) | ( n2207 & n3829 ) ;
  assign n10750 = ( n169 & n3621 ) | ( n169 & n10749 ) | ( n3621 & n10749 ) ;
  assign n10751 = ( n549 & n3578 ) | ( n549 & n6344 ) | ( n3578 & n6344 ) ;
  assign n10752 = ( ~n1157 & n9714 ) | ( ~n1157 & n10751 ) | ( n9714 & n10751 ) ;
  assign n10753 = n5430 | n5695 ;
  assign n10754 = n10575 ^ n4306 ^ n2704 ;
  assign n10755 = n2450 & n9770 ;
  assign n10756 = n10755 ^ n6886 ^ 1'b0 ;
  assign n10757 = n5654 & ~n10756 ;
  assign n10758 = n3167 & n4342 ;
  assign n10759 = n10758 ^ n8375 ^ 1'b0 ;
  assign n10760 = ( ~n2476 & n3904 ) | ( ~n2476 & n4190 ) | ( n3904 & n4190 ) ;
  assign n10761 = ( n361 & ~n4862 ) | ( n361 & n10760 ) | ( ~n4862 & n10760 ) ;
  assign n10762 = n10761 ^ n1829 ^ 1'b0 ;
  assign n10763 = n10762 ^ n1379 ^ n378 ;
  assign n10771 = ( n2569 & ~n2863 ) | ( n2569 & n3951 ) | ( ~n2863 & n3951 ) ;
  assign n10764 = n6186 ^ n4107 ^ n1568 ;
  assign n10765 = ( ~n617 & n3844 ) | ( ~n617 & n5259 ) | ( n3844 & n5259 ) ;
  assign n10766 = n5680 | n10765 ;
  assign n10767 = n4039 | n10766 ;
  assign n10768 = n10767 ^ n6226 ^ 1'b0 ;
  assign n10769 = n3838 | n10768 ;
  assign n10770 = ( n7119 & n10764 ) | ( n7119 & n10769 ) | ( n10764 & n10769 ) ;
  assign n10772 = n10771 ^ n10770 ^ 1'b0 ;
  assign n10773 = n10763 & ~n10772 ;
  assign n10774 = n3062 & ~n10773 ;
  assign n10781 = ( ~n4101 & n5309 ) | ( ~n4101 & n5453 ) | ( n5309 & n5453 ) ;
  assign n10775 = n859 & ~n4006 ;
  assign n10776 = ~n5817 & n10775 ;
  assign n10777 = n8545 ^ n2926 ^ x71 ;
  assign n10778 = n1816 & n2724 ;
  assign n10779 = ~n10777 & n10778 ;
  assign n10780 = ( n2918 & n10776 ) | ( n2918 & ~n10779 ) | ( n10776 & ~n10779 ) ;
  assign n10782 = n10781 ^ n10780 ^ n5441 ;
  assign n10783 = n4489 ^ n1153 ^ 1'b0 ;
  assign n10784 = ~n2899 & n10783 ;
  assign n10785 = ( ~n149 & n549 ) | ( ~n149 & n707 ) | ( n549 & n707 ) ;
  assign n10786 = n4939 & n10785 ;
  assign n10787 = n10786 ^ n4440 ^ 1'b0 ;
  assign n10788 = n5801 & n6424 ;
  assign n10789 = ( n537 & n10787 ) | ( n537 & n10788 ) | ( n10787 & n10788 ) ;
  assign n10790 = ~n4459 & n8586 ;
  assign n10791 = ( n8808 & n10789 ) | ( n8808 & n10790 ) | ( n10789 & n10790 ) ;
  assign n10792 = ( n4228 & ~n9621 ) | ( n4228 & n9846 ) | ( ~n9621 & n9846 ) ;
  assign n10793 = n3482 | n4176 ;
  assign n10794 = n2013 | n10793 ;
  assign n10795 = n10792 & n10794 ;
  assign n10796 = ( n131 & n5906 ) | ( n131 & n10795 ) | ( n5906 & n10795 ) ;
  assign n10797 = n4964 & n10796 ;
  assign n10798 = n8240 ^ n1921 ^ 1'b0 ;
  assign n10803 = ( ~n652 & n2727 ) | ( ~n652 & n8265 ) | ( n2727 & n8265 ) ;
  assign n10799 = n1733 ^ n1040 ^ 1'b0 ;
  assign n10800 = ( n3440 & n7572 ) | ( n3440 & n10799 ) | ( n7572 & n10799 ) ;
  assign n10801 = ~n4872 & n10800 ;
  assign n10802 = n6215 & n10801 ;
  assign n10804 = n10803 ^ n10802 ^ 1'b0 ;
  assign n10806 = ( n2445 & ~n4732 ) | ( n2445 & n9620 ) | ( ~n4732 & n9620 ) ;
  assign n10807 = n10806 ^ n4812 ^ 1'b0 ;
  assign n10805 = ~n1317 & n3750 ;
  assign n10808 = n10807 ^ n10805 ^ 1'b0 ;
  assign n10809 = n10808 ^ n9499 ^ 1'b0 ;
  assign n10810 = n516 & n629 ;
  assign n10811 = ~n2646 & n10810 ;
  assign n10812 = n10811 ^ n1955 ^ n756 ;
  assign n10813 = n6327 ^ n5625 ^ 1'b0 ;
  assign n10814 = ~n10812 & n10813 ;
  assign n10815 = n3897 | n4902 ;
  assign n10816 = n10815 ^ n8469 ^ n7071 ;
  assign n10817 = n2647 & n4684 ;
  assign n10818 = n8340 ^ n7075 ^ 1'b0 ;
  assign n10819 = n10817 & n10818 ;
  assign n10820 = ~n1128 & n2194 ;
  assign n10821 = n4089 ^ n3223 ^ n461 ;
  assign n10822 = ( n260 & n635 ) | ( n260 & ~n4856 ) | ( n635 & ~n4856 ) ;
  assign n10823 = n1527 & n6951 ;
  assign n10824 = ~n5915 & n10823 ;
  assign n10825 = ( n4169 & n10822 ) | ( n4169 & n10824 ) | ( n10822 & n10824 ) ;
  assign n10826 = n10825 ^ n9954 ^ n1616 ;
  assign n10827 = ~n1915 & n10826 ;
  assign n10828 = ( ~n2472 & n6170 ) | ( ~n2472 & n10827 ) | ( n6170 & n10827 ) ;
  assign n10829 = n8636 ^ n6926 ^ n4792 ;
  assign n10831 = ( n2036 & ~n2370 ) | ( n2036 & n6668 ) | ( ~n2370 & n6668 ) ;
  assign n10830 = n357 | n3706 ;
  assign n10832 = n10831 ^ n10830 ^ n8214 ;
  assign n10833 = ( ~n4046 & n8287 ) | ( ~n4046 & n10832 ) | ( n8287 & n10832 ) ;
  assign n10834 = ~n5148 & n5293 ;
  assign n10835 = n10834 ^ n8346 ^ n4436 ;
  assign n10837 = n5603 ^ n3550 ^ n1883 ;
  assign n10836 = n3862 ^ n3797 ^ n1145 ;
  assign n10838 = n10837 ^ n10836 ^ n2805 ;
  assign n10843 = n8370 ^ n1318 ^ n154 ;
  assign n10840 = ( n508 & ~n1038 ) | ( n508 & n3095 ) | ( ~n1038 & n3095 ) ;
  assign n10841 = n989 & n10840 ;
  assign n10842 = n2242 & n10841 ;
  assign n10839 = n5935 ^ n1736 ^ n1697 ;
  assign n10844 = n10843 ^ n10842 ^ n10839 ;
  assign n10845 = n10838 & n10844 ;
  assign n10846 = x112 | n471 ;
  assign n10847 = n10141 & n10846 ;
  assign n10848 = ( x24 & ~n3258 ) | ( x24 & n5578 ) | ( ~n3258 & n5578 ) ;
  assign n10849 = n7259 ^ n1693 ^ 1'b0 ;
  assign n10850 = n4774 | n10849 ;
  assign n10851 = n10850 ^ n4032 ^ 1'b0 ;
  assign n10852 = n1266 & n10851 ;
  assign n10853 = ~n10848 & n10852 ;
  assign n10854 = n8495 | n10853 ;
  assign n10855 = n5309 ^ n636 ^ 1'b0 ;
  assign n10856 = n7682 ^ n5001 ^ n1968 ;
  assign n10857 = ( n2262 & ~n2794 ) | ( n2262 & n10856 ) | ( ~n2794 & n10856 ) ;
  assign n10858 = n10857 ^ n2903 ^ n1971 ;
  assign n10863 = n9123 ^ n8793 ^ 1'b0 ;
  assign n10859 = n6936 ^ n4887 ^ 1'b0 ;
  assign n10860 = n501 & n10859 ;
  assign n10861 = n9518 ^ n2970 ^ 1'b0 ;
  assign n10862 = n10860 & n10861 ;
  assign n10864 = n10863 ^ n10862 ^ n1979 ;
  assign n10867 = ( ~n316 & n562 ) | ( ~n316 & n1289 ) | ( n562 & n1289 ) ;
  assign n10868 = n8316 & ~n10867 ;
  assign n10869 = n10868 ^ n2502 ^ 1'b0 ;
  assign n10870 = n10869 ^ n3098 ^ 1'b0 ;
  assign n10871 = n5977 & ~n10870 ;
  assign n10865 = n3822 & ~n5101 ;
  assign n10866 = n9042 & n10865 ;
  assign n10872 = n10871 ^ n10866 ^ n4246 ;
  assign n10873 = n4535 & ~n8601 ;
  assign n10874 = ~x32 & n10873 ;
  assign n10875 = n10874 ^ n7604 ^ 1'b0 ;
  assign n10876 = n227 | n10875 ;
  assign n10877 = n10872 & n10876 ;
  assign n10878 = n10877 ^ n8303 ^ 1'b0 ;
  assign n10881 = ( ~n523 & n1751 ) | ( ~n523 & n2896 ) | ( n1751 & n2896 ) ;
  assign n10879 = n849 | n2372 ;
  assign n10880 = n5159 | n10879 ;
  assign n10882 = n10881 ^ n10880 ^ n3735 ;
  assign n10883 = ( n2579 & ~n8824 ) | ( n2579 & n9161 ) | ( ~n8824 & n9161 ) ;
  assign n10884 = ( n6701 & n7326 ) | ( n6701 & n10883 ) | ( n7326 & n10883 ) ;
  assign n10885 = n10884 ^ n5753 ^ 1'b0 ;
  assign n10886 = n4050 | n10885 ;
  assign n10887 = ( ~n2646 & n4323 ) | ( ~n2646 & n8018 ) | ( n4323 & n8018 ) ;
  assign n10888 = n4684 & ~n10887 ;
  assign n10889 = ( n3149 & n3217 ) | ( n3149 & ~n8957 ) | ( n3217 & ~n8957 ) ;
  assign n10890 = n10889 ^ n2001 ^ n739 ;
  assign n10891 = n9331 ^ n4200 ^ 1'b0 ;
  assign n10892 = n5488 & ~n6351 ;
  assign n10893 = n5460 & ~n7251 ;
  assign n10894 = n7889 ^ n3220 ^ 1'b0 ;
  assign n10895 = n2280 ^ n893 ^ 1'b0 ;
  assign n10896 = n10895 ^ n6216 ^ n2953 ;
  assign n10897 = n2660 ^ n613 ^ 1'b0 ;
  assign n10898 = n742 | n10897 ;
  assign n10899 = n3950 & ~n10898 ;
  assign n10900 = ~n3869 & n10899 ;
  assign n10901 = n10900 ^ n1041 ^ 1'b0 ;
  assign n10902 = n1051 & ~n10901 ;
  assign n10903 = n10902 ^ n4160 ^ 1'b0 ;
  assign n10904 = n3777 ^ n1332 ^ 1'b0 ;
  assign n10905 = ~n2153 & n10904 ;
  assign n10906 = n10905 ^ n5806 ^ 1'b0 ;
  assign n10908 = n6607 ^ n1415 ^ 1'b0 ;
  assign n10907 = n4391 | n8237 ;
  assign n10909 = n10908 ^ n10907 ^ 1'b0 ;
  assign n10910 = n7349 ^ n1068 ^ n306 ;
  assign n10917 = n2283 & ~n2786 ;
  assign n10918 = n10917 ^ n10159 ^ n8967 ;
  assign n10911 = ( ~n454 & n601 ) | ( ~n454 & n4216 ) | ( n601 & n4216 ) ;
  assign n10912 = ~n1932 & n4415 ;
  assign n10913 = n10912 ^ n2205 ^ 1'b0 ;
  assign n10914 = n4961 ^ n2834 ^ 1'b0 ;
  assign n10915 = n10913 | n10914 ;
  assign n10916 = n10911 | n10915 ;
  assign n10919 = n10918 ^ n10916 ^ 1'b0 ;
  assign n10920 = n10910 & ~n10919 ;
  assign n10921 = ~n5572 & n7330 ;
  assign n10922 = n5005 ^ n2038 ^ 1'b0 ;
  assign n10923 = n7189 ^ n1718 ^ 1'b0 ;
  assign n10924 = n10923 ^ n3046 ^ 1'b0 ;
  assign n10925 = ~n2951 & n7599 ;
  assign n10926 = n4441 ^ n3980 ^ n1928 ;
  assign n10927 = n10926 ^ n2352 ^ 1'b0 ;
  assign n10928 = ~n5580 & n10927 ;
  assign n10929 = ~n8824 & n10928 ;
  assign n10930 = n1832 & n10929 ;
  assign n10931 = n10547 ^ n9509 ^ n6443 ;
  assign n10932 = ~n2430 & n5453 ;
  assign n10933 = n10932 ^ n1406 ^ 1'b0 ;
  assign n10934 = n10933 ^ n551 ^ 1'b0 ;
  assign n10935 = n10934 ^ n2567 ^ 1'b0 ;
  assign n10936 = ( n5971 & n10326 ) | ( n5971 & n10935 ) | ( n10326 & n10935 ) ;
  assign n10937 = ~n7824 & n7998 ;
  assign n10938 = n6410 & n10937 ;
  assign n10939 = n200 | n3735 ;
  assign n10940 = n1215 & ~n10939 ;
  assign n10941 = ~n2688 & n2776 ;
  assign n10942 = n5053 & n10941 ;
  assign n10943 = n10942 ^ n5521 ^ 1'b0 ;
  assign n10944 = ~n6140 & n10943 ;
  assign n10945 = ( ~n802 & n10940 ) | ( ~n802 & n10944 ) | ( n10940 & n10944 ) ;
  assign n10946 = ( n431 & ~n10938 ) | ( n431 & n10945 ) | ( ~n10938 & n10945 ) ;
  assign n10947 = n10946 ^ n3948 ^ n1837 ;
  assign n10948 = n3973 ^ n1697 ^ 1'b0 ;
  assign n10949 = n5554 ^ n3206 ^ n283 ;
  assign n10950 = ( n2113 & ~n2428 ) | ( n2113 & n10949 ) | ( ~n2428 & n10949 ) ;
  assign n10951 = n10105 ^ n9889 ^ n1710 ;
  assign n10952 = n10951 ^ n9810 ^ 1'b0 ;
  assign n10953 = n10950 | n10952 ;
  assign n10954 = ~n1797 & n3865 ;
  assign n10955 = ( n5721 & n7919 ) | ( n5721 & n10954 ) | ( n7919 & n10954 ) ;
  assign n10956 = n571 & n1658 ;
  assign n10957 = n10956 ^ n592 ^ 1'b0 ;
  assign n10958 = n10957 ^ n5440 ^ 1'b0 ;
  assign n10959 = ~n9553 & n10958 ;
  assign n10960 = ( n844 & n10955 ) | ( n844 & ~n10959 ) | ( n10955 & ~n10959 ) ;
  assign n10961 = ( n1445 & n1568 ) | ( n1445 & n3286 ) | ( n1568 & n3286 ) ;
  assign n10962 = n6760 & ~n10961 ;
  assign n10963 = ( n2043 & n8344 ) | ( n2043 & n10962 ) | ( n8344 & n10962 ) ;
  assign n10964 = ~n348 & n3118 ;
  assign n10965 = ~n10311 & n10964 ;
  assign n10966 = n1341 & n3813 ;
  assign n10967 = n10966 ^ n6424 ^ 1'b0 ;
  assign n10968 = n5778 ^ n1785 ^ 1'b0 ;
  assign n10969 = n3511 ^ n3247 ^ 1'b0 ;
  assign n10970 = ~n7909 & n10969 ;
  assign n10971 = n596 & ~n10970 ;
  assign n10972 = n3752 ^ n958 ^ 1'b0 ;
  assign n10973 = ~n9160 & n10972 ;
  assign n10974 = n4251 & n8812 ;
  assign n10975 = n10974 ^ n1515 ^ 1'b0 ;
  assign n10976 = ( n149 & ~n565 ) | ( n149 & n2077 ) | ( ~n565 & n2077 ) ;
  assign n10977 = n10976 ^ n3570 ^ n3347 ;
  assign n10978 = ( n2424 & n4266 ) | ( n2424 & n10977 ) | ( n4266 & n10977 ) ;
  assign n10979 = ~n478 & n3964 ;
  assign n10980 = ~n2025 & n10979 ;
  assign n10981 = n10980 ^ n7726 ^ 1'b0 ;
  assign n10983 = n3162 ^ n747 ^ n641 ;
  assign n10982 = ( n1810 & ~n3413 ) | ( n1810 & n7318 ) | ( ~n3413 & n7318 ) ;
  assign n10984 = n10983 ^ n10982 ^ 1'b0 ;
  assign n10985 = ( n8990 & ~n10981 ) | ( n8990 & n10984 ) | ( ~n10981 & n10984 ) ;
  assign n10986 = ( n2101 & ~n6099 ) | ( n2101 & n10985 ) | ( ~n6099 & n10985 ) ;
  assign n10987 = n7407 & ~n9455 ;
  assign n10991 = n3551 ^ n2011 ^ n1339 ;
  assign n10988 = x36 ^ x20 ^ 1'b0 ;
  assign n10989 = n2278 & n10988 ;
  assign n10990 = n10989 ^ n3976 ^ n386 ;
  assign n10992 = n10991 ^ n10990 ^ n10875 ;
  assign n10994 = n2862 ^ n431 ^ 1'b0 ;
  assign n10995 = n1103 & ~n10994 ;
  assign n10996 = n10995 ^ n1282 ^ 1'b0 ;
  assign n10997 = n6575 & ~n10996 ;
  assign n10993 = n8692 ^ n2495 ^ n2493 ;
  assign n10998 = n10997 ^ n10993 ^ 1'b0 ;
  assign n10999 = n10998 ^ n9883 ^ n519 ;
  assign n11000 = n8336 ^ n155 ^ 1'b0 ;
  assign n11001 = n6962 | n7898 ;
  assign n11002 = n894 | n11001 ;
  assign n11003 = n5021 ^ n318 ^ 1'b0 ;
  assign n11004 = n4356 & n11003 ;
  assign n11005 = ~n8805 & n11004 ;
  assign n11006 = ( n608 & ~n7903 ) | ( n608 & n10042 ) | ( ~n7903 & n10042 ) ;
  assign n11007 = x92 & n3191 ;
  assign n11008 = ~n605 & n11007 ;
  assign n11009 = ( n1143 & n5167 ) | ( n1143 & n11008 ) | ( n5167 & n11008 ) ;
  assign n11010 = ~n3870 & n11009 ;
  assign n11011 = n11010 ^ n7738 ^ n7691 ;
  assign n11012 = n5169 & n5728 ;
  assign n11013 = n11011 & ~n11012 ;
  assign n11014 = ~n8874 & n11013 ;
  assign n11015 = ~n3337 & n8314 ;
  assign n11016 = n11015 ^ n1668 ^ 1'b0 ;
  assign n11017 = ( n239 & n845 ) | ( n239 & ~n4364 ) | ( n845 & ~n4364 ) ;
  assign n11018 = n11017 ^ n6334 ^ 1'b0 ;
  assign n11019 = ( n4124 & n5635 ) | ( n4124 & n6800 ) | ( n5635 & n6800 ) ;
  assign n11020 = ~n4183 & n8113 ;
  assign n11021 = n11020 ^ n2523 ^ 1'b0 ;
  assign n11022 = n11021 ^ n3752 ^ 1'b0 ;
  assign n11025 = n10558 ^ n8620 ^ 1'b0 ;
  assign n11026 = ~n1037 & n11025 ;
  assign n11027 = n11026 ^ n2153 ^ 1'b0 ;
  assign n11028 = n8836 ^ n1104 ^ 1'b0 ;
  assign n11029 = n11028 ^ n2557 ^ 1'b0 ;
  assign n11030 = n11027 & n11029 ;
  assign n11023 = ( n194 & ~n844 ) | ( n194 & n3207 ) | ( ~n844 & n3207 ) ;
  assign n11024 = n3010 & n11023 ;
  assign n11031 = n11030 ^ n11024 ^ 1'b0 ;
  assign n11032 = n7835 ^ n4195 ^ n3214 ;
  assign n11033 = n881 & n11032 ;
  assign n11034 = n11031 & n11033 ;
  assign n11035 = n8007 | n11034 ;
  assign n11036 = n3244 | n11035 ;
  assign n11037 = ~n9165 & n10785 ;
  assign n11038 = n3842 & ~n5492 ;
  assign n11039 = ( n777 & ~n838 ) | ( n777 & n6416 ) | ( ~n838 & n6416 ) ;
  assign n11040 = n6021 & ~n11039 ;
  assign n11041 = n11038 & ~n11040 ;
  assign n11042 = n11041 ^ n9733 ^ 1'b0 ;
  assign n11043 = n8967 ^ n3274 ^ 1'b0 ;
  assign n11044 = ( n569 & n4877 ) | ( n569 & ~n8002 ) | ( n4877 & ~n8002 ) ;
  assign n11045 = n2447 ^ n1220 ^ 1'b0 ;
  assign n11046 = ( x74 & n6958 ) | ( x74 & n9084 ) | ( n6958 & n9084 ) ;
  assign n11050 = n6475 ^ n3421 ^ x112 ;
  assign n11049 = n477 & n500 ;
  assign n11051 = n11050 ^ n11049 ^ n4769 ;
  assign n11052 = n10895 ^ n4294 ^ n1679 ;
  assign n11053 = ( ~n1073 & n3509 ) | ( ~n1073 & n11052 ) | ( n3509 & n11052 ) ;
  assign n11054 = n11053 ^ n6958 ^ 1'b0 ;
  assign n11055 = ~n11051 & n11054 ;
  assign n11056 = n11055 ^ n4125 ^ 1'b0 ;
  assign n11047 = n10321 ^ n9701 ^ n9630 ;
  assign n11048 = n10267 & ~n11047 ;
  assign n11057 = n11056 ^ n11048 ^ 1'b0 ;
  assign n11059 = n877 & n7794 ;
  assign n11058 = n4708 & ~n4873 ;
  assign n11060 = n11059 ^ n11058 ^ 1'b0 ;
  assign n11061 = n3554 | n3938 ;
  assign n11062 = n6145 ^ n1492 ^ n165 ;
  assign n11063 = n754 & ~n11062 ;
  assign n11064 = n11063 ^ n2255 ^ 1'b0 ;
  assign n11065 = ( ~n2896 & n3774 ) | ( ~n2896 & n7832 ) | ( n3774 & n7832 ) ;
  assign n11067 = n7233 ^ n1390 ^ 1'b0 ;
  assign n11068 = ~n3100 & n10558 ;
  assign n11069 = n11068 ^ n5257 ^ 1'b0 ;
  assign n11070 = n11067 & ~n11069 ;
  assign n11066 = ~n5810 & n8161 ;
  assign n11071 = n11070 ^ n11066 ^ 1'b0 ;
  assign n11072 = n11071 ^ n1590 ^ 1'b0 ;
  assign n11073 = ( n3631 & ~n7498 ) | ( n3631 & n11072 ) | ( ~n7498 & n11072 ) ;
  assign n11074 = n7259 ^ n7075 ^ 1'b0 ;
  assign n11075 = n11074 ^ n1687 ^ 1'b0 ;
  assign n11076 = n1377 & ~n9092 ;
  assign n11077 = n3600 & n11076 ;
  assign n11078 = n7172 ^ n3287 ^ 1'b0 ;
  assign n11079 = n5474 ^ n2578 ^ n1084 ;
  assign n11080 = n4023 & ~n10255 ;
  assign n11085 = n1083 & ~n4625 ;
  assign n11086 = n543 & n11085 ;
  assign n11087 = ( n833 & n2910 ) | ( n833 & n11086 ) | ( n2910 & n11086 ) ;
  assign n11081 = n989 & n2279 ;
  assign n11082 = ~n269 & n11081 ;
  assign n11083 = ( n1385 & ~n10658 ) | ( n1385 & n11082 ) | ( ~n10658 & n11082 ) ;
  assign n11084 = n11083 ^ n6382 ^ 1'b0 ;
  assign n11088 = n11087 ^ n11084 ^ n2219 ;
  assign n11089 = n1018 | n5975 ;
  assign n11090 = n11089 ^ n9546 ^ 1'b0 ;
  assign n11091 = ~n1447 & n5679 ;
  assign n11092 = ~n5272 & n11091 ;
  assign n11093 = n11092 ^ n4639 ^ 1'b0 ;
  assign n11094 = ( n1741 & n7819 ) | ( n1741 & n11093 ) | ( n7819 & n11093 ) ;
  assign n11095 = n1480 | n6114 ;
  assign n11096 = n11094 | n11095 ;
  assign n11098 = n4463 ^ n573 ^ n392 ;
  assign n11097 = n6960 ^ n1275 ^ 1'b0 ;
  assign n11099 = n11098 ^ n11097 ^ n1019 ;
  assign n11100 = ~n4174 & n5676 ;
  assign n11101 = n11100 ^ n5151 ^ n4857 ;
  assign n11102 = n5290 & n11101 ;
  assign n11104 = ( ~n1914 & n4576 ) | ( ~n1914 & n4593 ) | ( n4576 & n4593 ) ;
  assign n11103 = n1104 & ~n7952 ;
  assign n11105 = n11104 ^ n11103 ^ 1'b0 ;
  assign n11106 = ~n8170 & n11105 ;
  assign n11107 = n11106 ^ n11080 ^ 1'b0 ;
  assign n11108 = n4385 ^ n2536 ^ n1339 ;
  assign n11109 = n8281 & ~n11108 ;
  assign n11110 = ( n921 & ~n951 ) | ( n921 & n11109 ) | ( ~n951 & n11109 ) ;
  assign n11111 = n1017 | n7530 ;
  assign n11112 = n500 | n11111 ;
  assign n11113 = n4177 & n11112 ;
  assign n11114 = ~x60 & n11113 ;
  assign n11115 = ( n4712 & n10554 ) | ( n4712 & ~n11114 ) | ( n10554 & ~n11114 ) ;
  assign n11116 = n11115 ^ n8388 ^ 1'b0 ;
  assign n11117 = x62 & n11116 ;
  assign n11118 = n11117 ^ n679 ^ 1'b0 ;
  assign n11119 = n8069 ^ n4048 ^ 1'b0 ;
  assign n11120 = ( ~n372 & n1882 ) | ( ~n372 & n5280 ) | ( n1882 & n5280 ) ;
  assign n11121 = n1447 & ~n7508 ;
  assign n11122 = n11120 & n11121 ;
  assign n11123 = n10600 ^ n2219 ^ 1'b0 ;
  assign n11124 = n171 & ~n11123 ;
  assign n11125 = ~x17 & n8681 ;
  assign n11126 = n425 | n527 ;
  assign n11127 = n2296 ^ n219 ^ 1'b0 ;
  assign n11128 = n3671 & ~n11127 ;
  assign n11129 = ( ~n2177 & n4837 ) | ( ~n2177 & n11128 ) | ( n4837 & n11128 ) ;
  assign n11130 = n5608 ^ n2624 ^ n752 ;
  assign n11131 = ( ~n954 & n6138 ) | ( ~n954 & n6524 ) | ( n6138 & n6524 ) ;
  assign n11132 = n11131 ^ n1460 ^ 1'b0 ;
  assign n11133 = n2505 & ~n11132 ;
  assign n11135 = ( ~n589 & n1434 ) | ( ~n589 & n4626 ) | ( n1434 & n4626 ) ;
  assign n11134 = ~n5762 & n5792 ;
  assign n11136 = n11135 ^ n11134 ^ n6614 ;
  assign n11137 = ( n8640 & n9475 ) | ( n8640 & n9698 ) | ( n9475 & n9698 ) ;
  assign n11138 = ~n826 & n5170 ;
  assign n11139 = n11138 ^ n6569 ^ 1'b0 ;
  assign n11140 = n10016 & n11139 ;
  assign n11141 = ~n11137 & n11140 ;
  assign n11142 = n11141 ^ n2682 ^ 1'b0 ;
  assign n11143 = n687 & n2895 ;
  assign n11144 = ~n8192 & n11143 ;
  assign n11145 = n11144 ^ x114 ^ 1'b0 ;
  assign n11146 = n793 & ~n11145 ;
  assign n11147 = n11146 ^ n7813 ^ 1'b0 ;
  assign n11148 = ( n250 & ~n366 ) | ( n250 & n11147 ) | ( ~n366 & n11147 ) ;
  assign n11152 = ( ~n675 & n2418 ) | ( ~n675 & n5478 ) | ( n2418 & n5478 ) ;
  assign n11149 = n1476 & ~n6541 ;
  assign n11150 = ~n5206 & n11149 ;
  assign n11151 = n11150 ^ n6114 ^ 1'b0 ;
  assign n11153 = n11152 ^ n11151 ^ 1'b0 ;
  assign n11154 = ( n481 & n1687 ) | ( n481 & ~n8318 ) | ( n1687 & ~n8318 ) ;
  assign n11155 = ( n1382 & n9160 ) | ( n1382 & n11154 ) | ( n9160 & n11154 ) ;
  assign n11156 = n9976 & n11155 ;
  assign n11157 = n5291 & n11156 ;
  assign n11159 = x32 | n9160 ;
  assign n11158 = ~n4320 & n5762 ;
  assign n11160 = n11159 ^ n11158 ^ 1'b0 ;
  assign n11161 = n4878 ^ n474 ^ 1'b0 ;
  assign n11162 = n11160 | n11161 ;
  assign n11163 = n7806 & ~n10414 ;
  assign n11164 = ~n3527 & n11163 ;
  assign n11165 = n390 & n974 ;
  assign n11166 = n11164 & n11165 ;
  assign n11167 = n3557 ^ n1954 ^ 1'b0 ;
  assign n11168 = ~n2450 & n11167 ;
  assign n11169 = ( n8949 & n10247 ) | ( n8949 & ~n11168 ) | ( n10247 & ~n11168 ) ;
  assign n11170 = ( n7368 & n11166 ) | ( n7368 & n11169 ) | ( n11166 & n11169 ) ;
  assign n11171 = ~n3409 & n7805 ;
  assign n11172 = n9767 ^ n4550 ^ 1'b0 ;
  assign n11173 = n4238 & ~n11172 ;
  assign n11175 = n5440 ^ x54 ^ 1'b0 ;
  assign n11176 = ~n1076 & n11175 ;
  assign n11177 = n11176 ^ n993 ^ 1'b0 ;
  assign n11178 = x80 & ~n11177 ;
  assign n11174 = n9059 & ~n9344 ;
  assign n11179 = n11178 ^ n11174 ^ 1'b0 ;
  assign n11180 = n4341 & ~n7491 ;
  assign n11181 = ~n5030 & n5301 ;
  assign n11182 = ( ~n3070 & n10592 ) | ( ~n3070 & n11181 ) | ( n10592 & n11181 ) ;
  assign n11183 = n4221 ^ n528 ^ n171 ;
  assign n11184 = n11183 ^ n2738 ^ n1338 ;
  assign n11185 = ( n1682 & n2547 ) | ( n1682 & n11184 ) | ( n2547 & n11184 ) ;
  assign n11186 = ( n7334 & n9894 ) | ( n7334 & n11185 ) | ( n9894 & n11185 ) ;
  assign n11187 = n4156 ^ n1096 ^ 1'b0 ;
  assign n11188 = n4231 ^ n576 ^ 1'b0 ;
  assign n11189 = ( ~n10494 & n11187 ) | ( ~n10494 & n11188 ) | ( n11187 & n11188 ) ;
  assign n11190 = n1600 | n5284 ;
  assign n11195 = n863 & ~n4616 ;
  assign n11191 = ( ~x23 & n1992 ) | ( ~x23 & n2681 ) | ( n1992 & n2681 ) ;
  assign n11192 = ( n7455 & ~n10636 ) | ( n7455 & n11191 ) | ( ~n10636 & n11191 ) ;
  assign n11193 = ~n744 & n11192 ;
  assign n11194 = n5322 & ~n11193 ;
  assign n11196 = n11195 ^ n11194 ^ 1'b0 ;
  assign n11197 = ( n6557 & ~n11190 ) | ( n6557 & n11196 ) | ( ~n11190 & n11196 ) ;
  assign n11198 = n159 | n192 ;
  assign n11199 = ( ~n3750 & n7388 ) | ( ~n3750 & n11198 ) | ( n7388 & n11198 ) ;
  assign n11200 = ~n11198 & n11199 ;
  assign n11201 = n4365 & n11200 ;
  assign n11202 = n1446 & ~n4344 ;
  assign n11203 = n7110 ^ n608 ^ n560 ;
  assign n11204 = n8825 | n11203 ;
  assign n11205 = n11202 | n11204 ;
  assign n11206 = n4087 & ~n6116 ;
  assign n11207 = n6710 & n11206 ;
  assign n11211 = ( ~n773 & n3857 ) | ( ~n773 & n5023 ) | ( n3857 & n5023 ) ;
  assign n11212 = n11211 ^ n6371 ^ n2613 ;
  assign n11213 = n11212 ^ n6787 ^ n6769 ;
  assign n11208 = x22 | n3566 ;
  assign n11209 = ( n1327 & n1940 ) | ( n1327 & ~n3781 ) | ( n1940 & ~n3781 ) ;
  assign n11210 = ( ~n492 & n11208 ) | ( ~n492 & n11209 ) | ( n11208 & n11209 ) ;
  assign n11214 = n11213 ^ n11210 ^ n4279 ;
  assign n11215 = n3483 ^ n2734 ^ n2641 ;
  assign n11216 = n11215 ^ n6831 ^ n796 ;
  assign n11217 = n10524 ^ n7536 ^ 1'b0 ;
  assign n11218 = n938 & ~n4057 ;
  assign n11219 = n570 & n11218 ;
  assign n11220 = n11219 ^ n5068 ^ n1638 ;
  assign n11221 = n11220 ^ n5283 ^ n3106 ;
  assign n11222 = n10558 ^ n3582 ^ n3547 ;
  assign n11223 = n11222 ^ n1464 ^ 1'b0 ;
  assign n11224 = n9152 ^ n5685 ^ 1'b0 ;
  assign n11225 = n11223 & ~n11224 ;
  assign n11226 = ~n474 & n8251 ;
  assign n11227 = n11226 ^ n7323 ^ n4505 ;
  assign n11228 = n7156 ^ n2832 ^ 1'b0 ;
  assign n11229 = n5325 & n11228 ;
  assign n11230 = n4797 & n11229 ;
  assign n11231 = n11230 ^ n7375 ^ 1'b0 ;
  assign n11232 = ~n9335 & n9824 ;
  assign n11233 = n2365 & ~n5539 ;
  assign n11234 = n11233 ^ n9813 ^ 1'b0 ;
  assign n11235 = n11234 ^ n8757 ^ 1'b0 ;
  assign n11236 = n10698 ^ n1611 ^ 1'b0 ;
  assign n11237 = n10678 | n11236 ;
  assign n11246 = n6086 ^ n3483 ^ n1444 ;
  assign n11238 = n9507 ^ n5865 ^ n4525 ;
  assign n11241 = n6273 ^ n5056 ^ n4832 ;
  assign n11242 = n11241 ^ n714 ^ 1'b0 ;
  assign n11243 = n470 & n11242 ;
  assign n11239 = ( ~n1238 & n1682 ) | ( ~n1238 & n10329 ) | ( n1682 & n10329 ) ;
  assign n11240 = n11239 ^ n2228 ^ 1'b0 ;
  assign n11244 = n11243 ^ n11240 ^ 1'b0 ;
  assign n11245 = n11238 & ~n11244 ;
  assign n11247 = n11246 ^ n11245 ^ n6823 ;
  assign n11250 = n8596 ^ n6454 ^ 1'b0 ;
  assign n11248 = n10002 ^ n337 ^ 1'b0 ;
  assign n11249 = n5956 & ~n11248 ;
  assign n11251 = n11250 ^ n11249 ^ 1'b0 ;
  assign n11252 = n3020 ^ n1363 ^ 1'b0 ;
  assign n11253 = n7812 & n11252 ;
  assign n11254 = n1285 & n1743 ;
  assign n11255 = ~n11253 & n11254 ;
  assign n11256 = n605 ^ x121 ^ 1'b0 ;
  assign n11257 = ~n5622 & n11256 ;
  assign n11258 = ( n2989 & n4351 ) | ( n2989 & n10842 ) | ( n4351 & n10842 ) ;
  assign n11259 = n11257 & n11258 ;
  assign n11260 = n11259 ^ n4723 ^ 1'b0 ;
  assign n11261 = n485 | n8214 ;
  assign n11262 = n11155 ^ n2919 ^ 1'b0 ;
  assign n11263 = n11262 ^ n5216 ^ 1'b0 ;
  assign n11264 = ~n1337 & n11263 ;
  assign n11265 = ( n1548 & ~n2399 ) | ( n1548 & n6379 ) | ( ~n2399 & n6379 ) ;
  assign n11266 = n5445 ^ n3213 ^ n3146 ;
  assign n11267 = n11266 ^ n3654 ^ x87 ;
  assign n11268 = n6672 ^ n1570 ^ 1'b0 ;
  assign n11274 = n2587 ^ x95 ^ 1'b0 ;
  assign n11275 = ~n7018 & n11274 ;
  assign n11269 = n1385 | n5078 ;
  assign n11270 = n302 | n11269 ;
  assign n11271 = n1925 & n3712 ;
  assign n11272 = n1384 & n11271 ;
  assign n11273 = ( ~n8730 & n11270 ) | ( ~n8730 & n11272 ) | ( n11270 & n11272 ) ;
  assign n11276 = n11275 ^ n11273 ^ 1'b0 ;
  assign n11277 = n11276 ^ n5124 ^ n1006 ;
  assign n11278 = n728 & ~n1455 ;
  assign n11282 = ( ~n783 & n4034 ) | ( ~n783 & n6148 ) | ( n4034 & n6148 ) ;
  assign n11279 = ~n405 & n5859 ;
  assign n11280 = n11279 ^ n7145 ^ x74 ;
  assign n11281 = n3748 | n11280 ;
  assign n11283 = n11282 ^ n11281 ^ 1'b0 ;
  assign n11284 = ~n2361 & n8282 ;
  assign n11285 = n10761 ^ n565 ^ 1'b0 ;
  assign n11286 = ~n2503 & n11285 ;
  assign n11287 = n1630 & ~n6456 ;
  assign n11288 = n8865 & n11287 ;
  assign n11289 = ~n2532 & n11288 ;
  assign n11290 = n11286 & ~n11289 ;
  assign n11291 = n11290 ^ x64 ^ 1'b0 ;
  assign n11292 = ( n1392 & n7457 ) | ( n1392 & n9761 ) | ( n7457 & n9761 ) ;
  assign n11293 = n11292 ^ n7857 ^ n1635 ;
  assign n11294 = n5159 & ~n11293 ;
  assign n11295 = n5113 & n11294 ;
  assign n11296 = n837 | n8982 ;
  assign n11297 = n3068 & ~n11296 ;
  assign n11298 = n11297 ^ n6853 ^ 1'b0 ;
  assign n11299 = n2015 & ~n2790 ;
  assign n11300 = n11299 ^ n2438 ^ 1'b0 ;
  assign n11301 = n11300 ^ n10159 ^ n2756 ;
  assign n11302 = n5547 ^ n3120 ^ n1069 ;
  assign n11303 = n2956 ^ n1785 ^ 1'b0 ;
  assign n11304 = n11302 | n11303 ;
  assign n11305 = n8142 | n11304 ;
  assign n11308 = ( n703 & n5676 ) | ( n703 & ~n6239 ) | ( n5676 & ~n6239 ) ;
  assign n11309 = n11308 ^ n4772 ^ 1'b0 ;
  assign n11310 = ~n3365 & n11309 ;
  assign n11306 = n2434 & ~n6116 ;
  assign n11307 = n11306 ^ n4212 ^ 1'b0 ;
  assign n11311 = n11310 ^ n11307 ^ n467 ;
  assign n11312 = n7652 ^ n4853 ^ 1'b0 ;
  assign n11313 = n9723 | n11312 ;
  assign n11314 = n11313 ^ n1923 ^ 1'b0 ;
  assign n11315 = n7940 & n11314 ;
  assign n11316 = ( n5674 & n10903 ) | ( n5674 & n11315 ) | ( n10903 & n11315 ) ;
  assign n11317 = n1188 & n5771 ;
  assign n11318 = n11317 ^ n7152 ^ 1'b0 ;
  assign n11319 = n7033 ^ n2761 ^ 1'b0 ;
  assign n11320 = n11319 ^ n7679 ^ n308 ;
  assign n11321 = n1444 | n11320 ;
  assign n11322 = n11321 ^ n7151 ^ 1'b0 ;
  assign n11323 = ( n1955 & n7580 ) | ( n1955 & n7960 ) | ( n7580 & n7960 ) ;
  assign n11325 = ( n514 & ~n1152 ) | ( n514 & n1456 ) | ( ~n1152 & n1456 ) ;
  assign n11326 = ( n4283 & ~n7941 ) | ( n4283 & n11325 ) | ( ~n7941 & n11325 ) ;
  assign n11324 = n7241 | n7269 ;
  assign n11327 = n11326 ^ n11324 ^ 1'b0 ;
  assign n11328 = n961 & ~n8053 ;
  assign n11329 = ~x21 & n11328 ;
  assign n11330 = n10334 ^ n8622 ^ n8426 ;
  assign n11331 = n5812 ^ n5789 ^ 1'b0 ;
  assign n11332 = n6562 & ~n10346 ;
  assign n11333 = n11331 | n11332 ;
  assign n11334 = n11333 ^ n6527 ^ 1'b0 ;
  assign n11335 = n10469 ^ n6794 ^ 1'b0 ;
  assign n11336 = n3112 & ~n11335 ;
  assign n11337 = n11334 & n11336 ;
  assign n11343 = n2960 & ~n8706 ;
  assign n11338 = n7353 ^ n664 ^ 1'b0 ;
  assign n11339 = ~n804 & n11338 ;
  assign n11340 = n6728 | n11339 ;
  assign n11341 = ( n4592 & n6485 ) | ( n4592 & n11340 ) | ( n6485 & n11340 ) ;
  assign n11342 = n169 & n11341 ;
  assign n11344 = n11343 ^ n11342 ^ n2939 ;
  assign n11345 = n477 ^ n348 ^ 1'b0 ;
  assign n11346 = ~n256 & n11345 ;
  assign n11347 = n11346 ^ n11283 ^ n5984 ;
  assign n11348 = n8301 ^ n5440 ^ 1'b0 ;
  assign n11349 = n3045 & n11348 ;
  assign n11350 = ( n8508 & n10610 ) | ( n8508 & ~n11349 ) | ( n10610 & ~n11349 ) ;
  assign n11351 = n6726 ^ n3613 ^ n3124 ;
  assign n11352 = ( n8422 & ~n8823 ) | ( n8422 & n11351 ) | ( ~n8823 & n11351 ) ;
  assign n11355 = n196 | n4286 ;
  assign n11356 = n1054 | n11355 ;
  assign n11357 = n11356 ^ n6331 ^ n3775 ;
  assign n11353 = ~n3653 & n5958 ;
  assign n11354 = n11353 ^ n6303 ^ 1'b0 ;
  assign n11358 = n11357 ^ n11354 ^ n7039 ;
  assign n11363 = n5428 ^ n2096 ^ 1'b0 ;
  assign n11364 = n877 & ~n11363 ;
  assign n11361 = ( ~n687 & n3473 ) | ( ~n687 & n5054 ) | ( n3473 & n5054 ) ;
  assign n11359 = n2375 ^ n743 ^ 1'b0 ;
  assign n11360 = n972 & ~n11359 ;
  assign n11362 = n11361 ^ n11360 ^ n7521 ;
  assign n11365 = n11364 ^ n11362 ^ n1580 ;
  assign n11366 = n11351 & ~n11365 ;
  assign n11373 = n6910 ^ n5596 ^ 1'b0 ;
  assign n11374 = n11373 ^ n11234 ^ 1'b0 ;
  assign n11367 = n1232 ^ x7 ^ 1'b0 ;
  assign n11368 = n469 & n11367 ;
  assign n11369 = ( n3222 & n5216 ) | ( n3222 & ~n6971 ) | ( n5216 & ~n6971 ) ;
  assign n11370 = n11369 ^ n5887 ^ 1'b0 ;
  assign n11371 = n11368 & ~n11370 ;
  assign n11372 = ~n10807 & n11371 ;
  assign n11375 = n11374 ^ n11372 ^ 1'b0 ;
  assign n11376 = n1529 | n3380 ;
  assign n11377 = n6304 | n11376 ;
  assign n11378 = ~n5050 & n11377 ;
  assign n11379 = ~n3027 & n11378 ;
  assign n11380 = ~n2220 & n5384 ;
  assign n11381 = ~n4615 & n11380 ;
  assign n11382 = n994 | n4434 ;
  assign n11383 = n5411 | n6685 ;
  assign n11384 = n11382 & ~n11383 ;
  assign n11385 = ~n639 & n3311 ;
  assign n11386 = n11385 ^ n2366 ^ 1'b0 ;
  assign n11387 = ~n8019 & n11386 ;
  assign n11388 = ( ~n11381 & n11384 ) | ( ~n11381 & n11387 ) | ( n11384 & n11387 ) ;
  assign n11389 = n10411 | n11388 ;
  assign n11390 = n733 | n6879 ;
  assign n11391 = n1204 & ~n11390 ;
  assign n11392 = n3235 & n11391 ;
  assign n11393 = ( n3043 & ~n3953 ) | ( n3043 & n11200 ) | ( ~n3953 & n11200 ) ;
  assign n11394 = n5941 | n11393 ;
  assign n11395 = n11392 | n11394 ;
  assign n11399 = n4033 & ~n9719 ;
  assign n11400 = n2047 & n2168 ;
  assign n11401 = n11399 & n11400 ;
  assign n11396 = n5230 & ~n6401 ;
  assign n11397 = n11396 ^ n7654 ^ 1'b0 ;
  assign n11398 = n4250 | n11397 ;
  assign n11402 = n11401 ^ n11398 ^ 1'b0 ;
  assign n11403 = n4265 ^ n629 ^ 1'b0 ;
  assign n11404 = ~n346 & n11403 ;
  assign n11405 = n4181 ^ n2884 ^ 1'b0 ;
  assign n11406 = n11404 & ~n11405 ;
  assign n11407 = ~n1298 & n11406 ;
  assign n11408 = n2832 & n11407 ;
  assign n11409 = n3349 ^ n1431 ^ 1'b0 ;
  assign n11410 = ~n11408 & n11409 ;
  assign n11411 = ~n1272 & n8407 ;
  assign n11412 = ~n11410 & n11411 ;
  assign n11413 = n10355 ^ n9722 ^ n4885 ;
  assign n11418 = n1754 ^ n1635 ^ n1032 ;
  assign n11419 = n11418 ^ n5811 ^ n4966 ;
  assign n11420 = n1345 | n8069 ;
  assign n11421 = n11420 ^ n3045 ^ 1'b0 ;
  assign n11422 = ( ~n9876 & n11419 ) | ( ~n9876 & n11421 ) | ( n11419 & n11421 ) ;
  assign n11414 = n1153 & ~n2605 ;
  assign n11415 = n2627 & n11414 ;
  assign n11416 = n10874 | n11415 ;
  assign n11417 = n10225 & ~n11416 ;
  assign n11423 = n11422 ^ n11417 ^ n3413 ;
  assign n11424 = n7582 | n11319 ;
  assign n11425 = n2252 | n11424 ;
  assign n11426 = n1661 | n4423 ;
  assign n11427 = n987 | n11426 ;
  assign n11430 = n5650 ^ n1569 ^ 1'b0 ;
  assign n11431 = n2141 & ~n2702 ;
  assign n11432 = ( n1605 & n11430 ) | ( n1605 & ~n11431 ) | ( n11430 & ~n11431 ) ;
  assign n11428 = n4263 ^ n624 ^ 1'b0 ;
  assign n11429 = n744 & ~n11428 ;
  assign n11433 = n11432 ^ n11429 ^ 1'b0 ;
  assign n11434 = n5890 ^ n5213 ^ n2805 ;
  assign n11435 = ( n2897 & n11433 ) | ( n2897 & n11434 ) | ( n11433 & n11434 ) ;
  assign n11436 = n6475 ^ n419 ^ 1'b0 ;
  assign n11437 = n689 & n11436 ;
  assign n11438 = n227 & n11437 ;
  assign n11439 = n8112 ^ n6110 ^ n2794 ;
  assign n11440 = n2480 & ~n11439 ;
  assign n11441 = n11440 ^ n7806 ^ 1'b0 ;
  assign n11442 = ~n852 & n1724 ;
  assign n11443 = n11441 & n11442 ;
  assign n11444 = n11443 ^ n7698 ^ n5140 ;
  assign n11445 = n11444 ^ n2982 ^ 1'b0 ;
  assign n11446 = x52 & n1585 ;
  assign n11447 = n11446 ^ n8571 ^ 1'b0 ;
  assign n11448 = n9545 & ~n11447 ;
  assign n11449 = n8047 & ~n10003 ;
  assign n11450 = ( ~n1628 & n3991 ) | ( ~n1628 & n11449 ) | ( n3991 & n11449 ) ;
  assign n11451 = n2593 & ~n6261 ;
  assign n11452 = n11451 ^ n5397 ^ n2025 ;
  assign n11453 = n11452 ^ n6186 ^ n1187 ;
  assign n11454 = n11453 ^ n5774 ^ 1'b0 ;
  assign n11455 = ~n3829 & n11454 ;
  assign n11456 = n9243 & ~n11455 ;
  assign n11457 = n11456 ^ n2845 ^ 1'b0 ;
  assign n11458 = ~n4140 & n10058 ;
  assign n11459 = n2876 & ~n11458 ;
  assign n11460 = n1774 & n11459 ;
  assign n11461 = n9123 ^ n349 ^ 1'b0 ;
  assign n11462 = n2868 & ~n11461 ;
  assign n11463 = n11462 ^ n11434 ^ 1'b0 ;
  assign n11464 = ( n386 & ~n610 ) | ( n386 & n5904 ) | ( ~n610 & n5904 ) ;
  assign n11465 = ( n6420 & n7943 ) | ( n6420 & n11464 ) | ( n7943 & n11464 ) ;
  assign n11468 = n6668 ^ n3242 ^ 1'b0 ;
  assign n11469 = n2835 & ~n11468 ;
  assign n11470 = ( ~n3964 & n7251 ) | ( ~n3964 & n11469 ) | ( n7251 & n11469 ) ;
  assign n11466 = n951 & n1724 ;
  assign n11467 = n2027 & ~n11466 ;
  assign n11471 = n11470 ^ n11467 ^ n10172 ;
  assign n11472 = n7317 ^ n4530 ^ 1'b0 ;
  assign n11473 = n6045 & ~n11472 ;
  assign n11474 = ~n10209 & n11473 ;
  assign n11475 = n11474 ^ n687 ^ 1'b0 ;
  assign n11478 = n8061 | n10687 ;
  assign n11479 = n4172 ^ n749 ^ 1'b0 ;
  assign n11480 = n2773 & n11479 ;
  assign n11481 = ( x126 & n1774 ) | ( x126 & n2560 ) | ( n1774 & n2560 ) ;
  assign n11482 = n2361 & ~n11481 ;
  assign n11483 = n5723 & n11482 ;
  assign n11484 = n11480 & ~n11483 ;
  assign n11485 = ~n11478 & n11484 ;
  assign n11476 = n2558 ^ n1650 ^ 1'b0 ;
  assign n11477 = n11476 ^ n5674 ^ n2621 ;
  assign n11486 = n11485 ^ n11477 ^ n865 ;
  assign n11495 = n6122 ^ n5428 ^ 1'b0 ;
  assign n11496 = n164 | n11495 ;
  assign n11490 = ~n437 & n2683 ;
  assign n11491 = n11490 ^ n3044 ^ 1'b0 ;
  assign n11492 = n8054 ^ n5360 ^ n4415 ;
  assign n11493 = n11491 & ~n11492 ;
  assign n11494 = n11493 ^ n3854 ^ 1'b0 ;
  assign n11487 = n540 | n3363 ;
  assign n11488 = ~n2354 & n11487 ;
  assign n11489 = n11488 ^ n1289 ^ 1'b0 ;
  assign n11497 = n11496 ^ n11494 ^ n11489 ;
  assign n11498 = n7227 ^ n5118 ^ n3459 ;
  assign n11499 = ~n10250 & n11498 ;
  assign n11500 = n11499 ^ n1717 ^ 1'b0 ;
  assign n11501 = n6018 ^ n4605 ^ 1'b0 ;
  assign n11502 = n11500 & ~n11501 ;
  assign n11503 = n5831 ^ n2515 ^ 1'b0 ;
  assign n11504 = ( n1121 & ~n5969 ) | ( n1121 & n11503 ) | ( ~n5969 & n11503 ) ;
  assign n11505 = n4933 & n10120 ;
  assign n11506 = n10839 ^ n10619 ^ n6312 ;
  assign n11507 = n7303 ^ n6099 ^ 1'b0 ;
  assign n11508 = n6604 & ~n6723 ;
  assign n11509 = n11508 ^ n10812 ^ 1'b0 ;
  assign n11510 = n10258 ^ n6319 ^ n6100 ;
  assign n11511 = n11510 ^ n6777 ^ 1'b0 ;
  assign n11512 = n10154 | n11511 ;
  assign n11513 = n11512 ^ n6107 ^ n3579 ;
  assign n11514 = ( n4956 & ~n8622 ) | ( n4956 & n11102 ) | ( ~n8622 & n11102 ) ;
  assign n11515 = n5235 & n5655 ;
  assign n11516 = n11515 ^ n7325 ^ 1'b0 ;
  assign n11521 = ( x37 & ~n372 ) | ( x37 & n1664 ) | ( ~n372 & n1664 ) ;
  assign n11522 = n1845 | n11521 ;
  assign n11517 = n3446 ^ n472 ^ 1'b0 ;
  assign n11518 = n4823 | n11517 ;
  assign n11519 = ( n4777 & ~n9226 ) | ( n4777 & n11518 ) | ( ~n9226 & n11518 ) ;
  assign n11520 = n3468 | n11519 ;
  assign n11523 = n11522 ^ n11520 ^ 1'b0 ;
  assign n11524 = ( n266 & n1283 ) | ( n266 & n3060 ) | ( n1283 & n3060 ) ;
  assign n11525 = n11524 ^ n4822 ^ n4637 ;
  assign n11526 = n11525 ^ n8364 ^ n6497 ;
  assign n11527 = ~n7086 & n11526 ;
  assign n11528 = n2165 & n2886 ;
  assign n11529 = ~n7251 & n11528 ;
  assign n11530 = n11529 ^ n9954 ^ n4121 ;
  assign n11531 = n11530 ^ n7748 ^ 1'b0 ;
  assign n11532 = ~n5035 & n7207 ;
  assign n11533 = ~n2175 & n11532 ;
  assign n11534 = n11533 ^ n4179 ^ n2401 ;
  assign n11535 = ( n7412 & ~n8502 ) | ( n7412 & n11534 ) | ( ~n8502 & n11534 ) ;
  assign n11536 = n5928 & ~n11535 ;
  assign n11537 = n5023 & n11536 ;
  assign n11538 = ( n3135 & ~n5230 ) | ( n3135 & n7940 ) | ( ~n5230 & n7940 ) ;
  assign n11539 = n11538 ^ n5521 ^ n2627 ;
  assign n11540 = n11539 ^ n9639 ^ 1'b0 ;
  assign n11541 = n6131 | n11540 ;
  assign n11542 = ( ~n787 & n2962 ) | ( ~n787 & n11541 ) | ( n2962 & n11541 ) ;
  assign n11543 = n5118 & ~n6327 ;
  assign n11544 = n11543 ^ n227 ^ 1'b0 ;
  assign n11545 = ( n1585 & n11292 ) | ( n1585 & ~n11544 ) | ( n11292 & ~n11544 ) ;
  assign n11546 = ( n1287 & n4792 ) | ( n1287 & ~n4873 ) | ( n4792 & ~n4873 ) ;
  assign n11547 = ~n7508 & n11546 ;
  assign n11548 = ~n2794 & n11547 ;
  assign n11549 = n11548 ^ n6191 ^ 1'b0 ;
  assign n11557 = ( n1002 & ~n9736 ) | ( n1002 & n10881 ) | ( ~n9736 & n10881 ) ;
  assign n11555 = n2732 & ~n3282 ;
  assign n11556 = n7705 & n11555 ;
  assign n11550 = n4881 ^ n291 ^ 1'b0 ;
  assign n11551 = n3027 & n11550 ;
  assign n11552 = n7812 ^ n3272 ^ n474 ;
  assign n11553 = n8081 & n11552 ;
  assign n11554 = ~n11551 & n11553 ;
  assign n11558 = n11557 ^ n11556 ^ n11554 ;
  assign n11559 = n8830 ^ n1100 ^ 1'b0 ;
  assign n11560 = ~n5791 & n11559 ;
  assign n11561 = n4391 ^ n2041 ^ 1'b0 ;
  assign n11562 = ( n2199 & n6886 ) | ( n2199 & ~n9239 ) | ( n6886 & ~n9239 ) ;
  assign n11563 = n11562 ^ n8644 ^ 1'b0 ;
  assign n11564 = ~n11561 & n11563 ;
  assign n11565 = n7406 ^ n6800 ^ 1'b0 ;
  assign n11566 = n8067 ^ n7174 ^ 1'b0 ;
  assign n11567 = n1288 ^ n1004 ^ 1'b0 ;
  assign n11568 = n3904 | n11567 ;
  assign n11569 = n898 & n8765 ;
  assign n11570 = n11569 ^ n9390 ^ 1'b0 ;
  assign n11571 = n11570 ^ n10708 ^ 1'b0 ;
  assign n11572 = ( n1203 & ~n7278 ) | ( n1203 & n7759 ) | ( ~n7278 & n7759 ) ;
  assign n11573 = n11572 ^ n1791 ^ 1'b0 ;
  assign n11574 = n6055 | n6333 ;
  assign n11575 = ~n4566 & n5016 ;
  assign n11576 = n9811 ^ n7149 ^ 1'b0 ;
  assign n11577 = n8547 & ~n8664 ;
  assign n11578 = n5414 | n11577 ;
  assign n11579 = n11118 & n11578 ;
  assign n11580 = n3689 | n9901 ;
  assign n11581 = n2558 & n7462 ;
  assign n11582 = n11581 ^ n3285 ^ 1'b0 ;
  assign n11583 = n7928 | n11582 ;
  assign n11590 = n6170 ^ n3124 ^ n977 ;
  assign n11591 = n1475 & n11590 ;
  assign n11592 = ~n8510 & n11591 ;
  assign n11587 = n1390 | n3388 ;
  assign n11588 = n3919 & ~n11587 ;
  assign n11584 = n1095 & ~n1110 ;
  assign n11585 = n8975 & n11584 ;
  assign n11586 = n7624 & ~n11585 ;
  assign n11589 = n11588 ^ n11586 ^ 1'b0 ;
  assign n11593 = n11592 ^ n11589 ^ n5212 ;
  assign n11594 = ~n1318 & n3299 ;
  assign n11595 = n5208 & n11594 ;
  assign n11596 = n9418 & ~n11595 ;
  assign n11597 = n2535 & n11596 ;
  assign n11598 = n11387 | n11597 ;
  assign n11599 = n7806 ^ n2929 ^ n676 ;
  assign n11600 = n11599 ^ n7513 ^ n4257 ;
  assign n11601 = ( ~n2060 & n7192 ) | ( ~n2060 & n11600 ) | ( n7192 & n11600 ) ;
  assign n11602 = n11601 ^ n4236 ^ 1'b0 ;
  assign n11603 = n5076 & ~n11131 ;
  assign n11604 = x24 & n339 ;
  assign n11605 = n11604 ^ n7313 ^ 1'b0 ;
  assign n11606 = n4978 ^ n1054 ^ 1'b0 ;
  assign n11607 = ( n6450 & n8002 ) | ( n6450 & n11606 ) | ( n8002 & n11606 ) ;
  assign n11608 = n11605 & ~n11607 ;
  assign n11609 = n11608 ^ n2331 ^ 1'b0 ;
  assign n11610 = n2345 & ~n3109 ;
  assign n11611 = n11610 ^ n2860 ^ 1'b0 ;
  assign n11612 = ( n6114 & n10371 ) | ( n6114 & ~n11611 ) | ( n10371 & ~n11611 ) ;
  assign n11613 = n5497 & ~n11612 ;
  assign n11614 = n2934 & n11613 ;
  assign n11615 = n3504 ^ n1630 ^ n703 ;
  assign n11616 = ( n9374 & n11093 ) | ( n9374 & ~n11615 ) | ( n11093 & ~n11615 ) ;
  assign n11617 = n11616 ^ n5655 ^ n4123 ;
  assign n11618 = n5915 & ~n10373 ;
  assign n11619 = n11618 ^ n8156 ^ 1'b0 ;
  assign n11620 = n204 & ~n11619 ;
  assign n11622 = n6051 ^ n4278 ^ 1'b0 ;
  assign n11621 = n4154 & n10206 ;
  assign n11623 = n11622 ^ n11621 ^ 1'b0 ;
  assign n11624 = n5457 ^ n495 ^ 1'b0 ;
  assign n11625 = ~n9528 & n11624 ;
  assign n11626 = n901 | n4878 ;
  assign n11627 = ( n4433 & n11625 ) | ( n4433 & n11626 ) | ( n11625 & n11626 ) ;
  assign n11628 = n4821 | n5678 ;
  assign n11629 = n1309 & n11628 ;
  assign n11630 = ( ~n2062 & n3045 ) | ( ~n2062 & n10529 ) | ( n3045 & n10529 ) ;
  assign n11631 = n8957 & ~n11630 ;
  assign n11633 = n3486 ^ n2659 ^ x40 ;
  assign n11632 = n465 | n1223 ;
  assign n11634 = n11633 ^ n11632 ^ 1'b0 ;
  assign n11635 = ( n2462 & n7578 ) | ( n2462 & n11464 ) | ( n7578 & n11464 ) ;
  assign n11636 = n3423 & n5353 ;
  assign n11638 = n230 | n9288 ;
  assign n11639 = n11638 ^ n3309 ^ 1'b0 ;
  assign n11637 = n7338 ^ n6477 ^ 1'b0 ;
  assign n11640 = n11639 ^ n11637 ^ n2884 ;
  assign n11641 = n1285 & n5776 ;
  assign n11642 = n11641 ^ n10767 ^ 1'b0 ;
  assign n11651 = n8763 ^ n1187 ^ 1'b0 ;
  assign n11647 = n4757 ^ n2811 ^ x11 ;
  assign n11648 = n11647 ^ n5453 ^ n2718 ;
  assign n11649 = n11648 ^ n10989 ^ n6226 ;
  assign n11643 = n9799 ^ n1881 ^ 1'b0 ;
  assign n11644 = n5764 & n11643 ;
  assign n11645 = ~n669 & n11644 ;
  assign n11646 = n11645 ^ n4370 ^ 1'b0 ;
  assign n11650 = n11649 ^ n11646 ^ n7691 ;
  assign n11652 = n11651 ^ n11650 ^ n4050 ;
  assign n11653 = n6258 & n6953 ;
  assign n11654 = n7429 | n11653 ;
  assign n11655 = n11654 ^ n5832 ^ 1'b0 ;
  assign n11659 = ( n1068 & n1632 ) | ( n1068 & n10439 ) | ( n1632 & n10439 ) ;
  assign n11660 = n4313 | n11659 ;
  assign n11656 = n4280 ^ n875 ^ 1'b0 ;
  assign n11657 = n3165 & n11656 ;
  assign n11658 = n3606 | n11657 ;
  assign n11661 = n11660 ^ n11658 ^ n4917 ;
  assign n11662 = ~n9607 & n11661 ;
  assign n11663 = n4299 ^ n3861 ^ 1'b0 ;
  assign n11664 = n6223 ^ n6202 ^ 1'b0 ;
  assign n11665 = n6580 | n11664 ;
  assign n11666 = n11665 ^ n5500 ^ 1'b0 ;
  assign n11667 = n5133 ^ n4121 ^ 1'b0 ;
  assign n11668 = n9660 & ~n9945 ;
  assign n11669 = n7483 ^ n7301 ^ 1'b0 ;
  assign n11670 = n5821 & ~n5905 ;
  assign n11671 = ~n2085 & n4928 ;
  assign n11672 = n7483 | n11671 ;
  assign n11673 = n11672 ^ n3682 ^ 1'b0 ;
  assign n11674 = n4172 & n4877 ;
  assign n11675 = n11674 ^ n2981 ^ n1035 ;
  assign n11676 = n9173 ^ n8454 ^ 1'b0 ;
  assign n11679 = ( ~x25 & n4693 ) | ( ~x25 & n11151 ) | ( n4693 & n11151 ) ;
  assign n11677 = ( ~n743 & n3645 ) | ( ~n743 & n8621 ) | ( n3645 & n8621 ) ;
  assign n11678 = n11677 ^ n1609 ^ 1'b0 ;
  assign n11680 = n11679 ^ n11678 ^ 1'b0 ;
  assign n11681 = n11680 ^ n8216 ^ 1'b0 ;
  assign n11682 = ~n5254 & n11681 ;
  assign n11683 = n4959 & n10426 ;
  assign n11684 = n1396 & n11683 ;
  assign n11685 = n447 & ~n2390 ;
  assign n11686 = ~n1298 & n5788 ;
  assign n11687 = n11686 ^ n1877 ^ 1'b0 ;
  assign n11688 = ~n11685 & n11687 ;
  assign n11689 = n5478 & ~n5762 ;
  assign n11690 = n8227 ^ n8035 ^ 1'b0 ;
  assign n11691 = n5704 & ~n11690 ;
  assign n11692 = n3640 ^ n178 ^ 1'b0 ;
  assign n11693 = n11692 ^ n712 ^ 1'b0 ;
  assign n11694 = n11691 & ~n11693 ;
  assign n11695 = n5655 & n11694 ;
  assign n11696 = n11689 & n11695 ;
  assign n11697 = n11696 ^ n3384 ^ 1'b0 ;
  assign n11698 = n4458 ^ n213 ^ 1'b0 ;
  assign n11699 = ( n1185 & n8803 ) | ( n1185 & ~n11698 ) | ( n8803 & ~n11698 ) ;
  assign n11700 = n537 & n2360 ;
  assign n11701 = n10917 & n11700 ;
  assign n11702 = n11701 ^ n3285 ^ n439 ;
  assign n11703 = n8530 ^ n7064 ^ 1'b0 ;
  assign n11705 = ~n5832 & n7496 ;
  assign n11706 = n5832 & n11705 ;
  assign n11704 = n5017 & ~n6137 ;
  assign n11707 = n11706 ^ n11704 ^ 1'b0 ;
  assign n11709 = n6332 ^ n5482 ^ n2660 ;
  assign n11708 = n2111 & n10000 ;
  assign n11710 = n11709 ^ n11708 ^ n3903 ;
  assign n11711 = n6673 & ~n8138 ;
  assign n11712 = n1642 | n4028 ;
  assign n11713 = n11712 ^ n3700 ^ 1'b0 ;
  assign n11714 = n4681 & n11713 ;
  assign n11715 = n11714 ^ n4605 ^ 1'b0 ;
  assign n11716 = n8401 ^ n3581 ^ 1'b0 ;
  assign n11717 = ( n1690 & n3881 ) | ( n1690 & n8387 ) | ( n3881 & n8387 ) ;
  assign n11718 = n1976 | n11717 ;
  assign n11719 = n1476 & n11718 ;
  assign n11720 = n5542 & ~n6159 ;
  assign n11721 = ( n3656 & n5505 ) | ( n3656 & n11720 ) | ( n5505 & n11720 ) ;
  assign n11722 = n519 | n3276 ;
  assign n11723 = n3179 | n11722 ;
  assign n11724 = n11721 | n11723 ;
  assign n11725 = n2752 ^ n1310 ^ 1'b0 ;
  assign n11726 = n538 & n11725 ;
  assign n11727 = ( n1121 & n3309 ) | ( n1121 & n11726 ) | ( n3309 & n11726 ) ;
  assign n11728 = n2262 | n11727 ;
  assign n11729 = n11728 ^ n9254 ^ 1'b0 ;
  assign n11730 = n4865 ^ n1547 ^ 1'b0 ;
  assign n11731 = n11730 ^ n7521 ^ n6170 ;
  assign n11732 = ( n2824 & ~n6873 ) | ( n2824 & n11731 ) | ( ~n6873 & n11731 ) ;
  assign n11733 = n6835 ^ n2972 ^ 1'b0 ;
  assign n11734 = n890 & n11733 ;
  assign n11735 = n11083 & n11734 ;
  assign n11736 = n4754 ^ n1236 ^ 1'b0 ;
  assign n11737 = n3507 ^ n680 ^ 1'b0 ;
  assign n11738 = n2736 ^ n1930 ^ 1'b0 ;
  assign n11739 = ( n2275 & n9672 ) | ( n2275 & n11738 ) | ( n9672 & n11738 ) ;
  assign n11740 = n11375 & n11739 ;
  assign n11741 = ~n11737 & n11740 ;
  assign n11742 = n11736 | n11741 ;
  assign n11743 = n11742 ^ n10149 ^ 1'b0 ;
  assign n11744 = n5889 & ~n7018 ;
  assign n11745 = n8919 ^ n4457 ^ 1'b0 ;
  assign n11746 = ( n5475 & ~n9552 ) | ( n5475 & n11745 ) | ( ~n9552 & n11745 ) ;
  assign n11751 = ~n4327 & n9115 ;
  assign n11752 = ~n8117 & n11751 ;
  assign n11747 = n4262 ^ n654 ^ 1'b0 ;
  assign n11748 = n11747 ^ n7806 ^ n2307 ;
  assign n11749 = n7285 | n11748 ;
  assign n11750 = n11749 ^ n2290 ^ 1'b0 ;
  assign n11753 = n11752 ^ n11750 ^ n2272 ;
  assign n11755 = n1134 | n2793 ;
  assign n11756 = n5575 & ~n11755 ;
  assign n11757 = n10860 ^ n3498 ^ 1'b0 ;
  assign n11758 = n318 & n11757 ;
  assign n11759 = ( n869 & n4921 ) | ( n869 & n7299 ) | ( n4921 & n7299 ) ;
  assign n11760 = n11758 & ~n11759 ;
  assign n11761 = n11756 & n11760 ;
  assign n11762 = n11761 ^ n2715 ^ 1'b0 ;
  assign n11763 = n3605 & n11762 ;
  assign n11754 = n1731 & ~n4550 ;
  assign n11764 = n11763 ^ n11754 ^ 1'b0 ;
  assign n11765 = n1298 | n5032 ;
  assign n11766 = n11765 ^ n5071 ^ 1'b0 ;
  assign n11767 = n8967 ^ n8272 ^ n1611 ;
  assign n11768 = ( n1062 & n5332 ) | ( n1062 & ~n6010 ) | ( n5332 & ~n6010 ) ;
  assign n11769 = n11768 ^ n7788 ^ 1'b0 ;
  assign n11770 = ~n11767 & n11769 ;
  assign n11771 = ( n6034 & n11766 ) | ( n6034 & n11770 ) | ( n11766 & n11770 ) ;
  assign n11772 = n11771 ^ n5364 ^ 1'b0 ;
  assign n11773 = n10459 ^ n3749 ^ n1952 ;
  assign n11774 = n3829 | n4710 ;
  assign n11775 = x112 | n11774 ;
  assign n11776 = n5492 ^ n2713 ^ 1'b0 ;
  assign n11777 = n11776 ^ n10856 ^ 1'b0 ;
  assign n11778 = ( n1223 & n5593 ) | ( n1223 & ~n11777 ) | ( n5593 & ~n11777 ) ;
  assign n11779 = n1588 ^ n1079 ^ 1'b0 ;
  assign n11782 = ( n388 & n469 ) | ( n388 & n1143 ) | ( n469 & n1143 ) ;
  assign n11783 = ( n1886 & n3554 ) | ( n1886 & n11782 ) | ( n3554 & n11782 ) ;
  assign n11780 = n2413 & ~n5547 ;
  assign n11781 = n11780 ^ n5786 ^ 1'b0 ;
  assign n11784 = n11783 ^ n11781 ^ n6455 ;
  assign n11785 = ( n1897 & ~n11779 ) | ( n1897 & n11784 ) | ( ~n11779 & n11784 ) ;
  assign n11786 = ( n4567 & n6388 ) | ( n4567 & ~n8759 ) | ( n6388 & ~n8759 ) ;
  assign n11787 = n11786 ^ n11570 ^ n5723 ;
  assign n11788 = ( n8643 & n9881 ) | ( n8643 & n11787 ) | ( n9881 & n11787 ) ;
  assign n11789 = n2168 ^ n457 ^ n233 ;
  assign n11790 = n11789 ^ n11432 ^ 1'b0 ;
  assign n11791 = x6 & ~n11790 ;
  assign n11792 = n11791 ^ n10435 ^ n9145 ;
  assign n11794 = n227 & n11192 ;
  assign n11795 = n11794 ^ n4848 ^ 1'b0 ;
  assign n11793 = n607 & n3251 ;
  assign n11796 = n11795 ^ n11793 ^ 1'b0 ;
  assign n11797 = ~n4847 & n6841 ;
  assign n11798 = n11797 ^ n7129 ^ 1'b0 ;
  assign n11799 = n7883 ^ n2701 ^ n1000 ;
  assign n11800 = n7136 | n11799 ;
  assign n11801 = n4952 | n11800 ;
  assign n11802 = n187 & n11801 ;
  assign n11803 = n2170 & n11802 ;
  assign n11804 = n487 | n3602 ;
  assign n11805 = ( ~n1548 & n4626 ) | ( ~n1548 & n11804 ) | ( n4626 & n11804 ) ;
  assign n11806 = ( ~n3367 & n5474 ) | ( ~n3367 & n6617 ) | ( n5474 & n6617 ) ;
  assign n11807 = n1611 & ~n3756 ;
  assign n11808 = ~n7738 & n11807 ;
  assign n11809 = n11808 ^ n5711 ^ n4843 ;
  assign n11810 = n11809 ^ n8929 ^ 1'b0 ;
  assign n11811 = n2433 | n11810 ;
  assign n11812 = n7379 & ~n9167 ;
  assign n11813 = ( ~n8074 & n9855 ) | ( ~n8074 & n11812 ) | ( n9855 & n11812 ) ;
  assign n11814 = n7193 ^ n5979 ^ n2553 ;
  assign n11815 = ~n8634 & n11814 ;
  assign n11816 = n11815 ^ n9805 ^ n3709 ;
  assign n11817 = n11816 ^ n5588 ^ 1'b0 ;
  assign n11818 = n6103 ^ n4605 ^ 1'b0 ;
  assign n11819 = n3040 & ~n11818 ;
  assign n11820 = n11819 ^ n3780 ^ 1'b0 ;
  assign n11821 = n11820 ^ n3378 ^ 1'b0 ;
  assign n11822 = ( n1690 & n2934 ) | ( n1690 & ~n3402 ) | ( n2934 & ~n3402 ) ;
  assign n11823 = n11822 ^ n2413 ^ 1'b0 ;
  assign n11824 = n4632 & n11823 ;
  assign n11825 = n2600 & ~n8702 ;
  assign n11826 = n10811 ^ n8825 ^ n4007 ;
  assign n11827 = ~n3602 & n8008 ;
  assign n11828 = ~n11826 & n11827 ;
  assign n11830 = n2247 & ~n2423 ;
  assign n11831 = n11830 ^ n1602 ^ 1'b0 ;
  assign n11829 = n7575 ^ n903 ^ 1'b0 ;
  assign n11832 = n11831 ^ n11829 ^ n2186 ;
  assign n11833 = n2381 ^ n1625 ^ 1'b0 ;
  assign n11834 = n11833 ^ n4914 ^ x74 ;
  assign n11835 = ( ~n738 & n2418 ) | ( ~n738 & n2499 ) | ( n2418 & n2499 ) ;
  assign n11836 = n11835 ^ n6697 ^ 1'b0 ;
  assign n11837 = ~n752 & n11836 ;
  assign n11838 = n10891 & n11837 ;
  assign n11839 = n11838 ^ n3168 ^ 1'b0 ;
  assign n11840 = n10497 ^ n1523 ^ 1'b0 ;
  assign n11844 = n318 | n1789 ;
  assign n11845 = ~n7171 & n11844 ;
  assign n11846 = n11845 ^ n6586 ^ 1'b0 ;
  assign n11847 = n11846 ^ n7449 ^ n4286 ;
  assign n11841 = ( ~n487 & n4155 ) | ( ~n487 & n9626 ) | ( n4155 & n9626 ) ;
  assign n11842 = ( n6623 & n8896 ) | ( n6623 & n11841 ) | ( n8896 & n11841 ) ;
  assign n11843 = n3272 & n11842 ;
  assign n11848 = n11847 ^ n11843 ^ 1'b0 ;
  assign n11849 = ~n2209 & n5596 ;
  assign n11850 = ( n7634 & n8152 ) | ( n7634 & ~n11849 ) | ( n8152 & ~n11849 ) ;
  assign n11851 = ( n1827 & ~n8439 ) | ( n1827 & n11850 ) | ( ~n8439 & n11850 ) ;
  assign n11853 = n6824 & ~n8803 ;
  assign n11854 = n11091 ^ n5247 ^ 1'b0 ;
  assign n11855 = n11853 | n11854 ;
  assign n11852 = n9103 & ~n9734 ;
  assign n11856 = n11855 ^ n11852 ^ 1'b0 ;
  assign n11857 = n7332 ^ n1923 ^ 1'b0 ;
  assign n11861 = ( n1243 & n5154 ) | ( n1243 & ~n5360 ) | ( n5154 & ~n5360 ) ;
  assign n11858 = n6345 | n11469 ;
  assign n11859 = n11858 ^ n4013 ^ 1'b0 ;
  assign n11860 = n409 & ~n11859 ;
  assign n11862 = n11861 ^ n11860 ^ 1'b0 ;
  assign n11863 = n11621 ^ n1751 ^ 1'b0 ;
  assign n11864 = n10979 & n11863 ;
  assign n11865 = n1392 ^ n1032 ^ 1'b0 ;
  assign n11866 = ~n411 & n1411 ;
  assign n11867 = n849 & n11866 ;
  assign n11868 = n5168 ^ n2704 ^ 1'b0 ;
  assign n11869 = n11868 ^ n2438 ^ 1'b0 ;
  assign n11870 = n11869 ^ n6169 ^ n3860 ;
  assign n11871 = ( n11300 & ~n11853 ) | ( n11300 & n11870 ) | ( ~n11853 & n11870 ) ;
  assign n11872 = ( n3654 & n11867 ) | ( n3654 & n11871 ) | ( n11867 & n11871 ) ;
  assign n11873 = n1777 & n10372 ;
  assign n11874 = n2746 & ~n7174 ;
  assign n11875 = n11874 ^ n2132 ^ 1'b0 ;
  assign n11876 = n6641 & n7070 ;
  assign n11877 = n11876 ^ n3259 ^ 1'b0 ;
  assign n11878 = x66 & n2618 ;
  assign n11879 = n11878 ^ n7507 ^ 1'b0 ;
  assign n11880 = n10197 ^ n2668 ^ 1'b0 ;
  assign n11881 = ( ~n401 & n11879 ) | ( ~n401 & n11880 ) | ( n11879 & n11880 ) ;
  assign n11882 = n11881 ^ n11437 ^ 1'b0 ;
  assign n11883 = n11877 & n11882 ;
  assign n11893 = n10443 ^ n468 ^ 1'b0 ;
  assign n11888 = n3003 ^ n357 ^ 1'b0 ;
  assign n11886 = ~n1503 & n2417 ;
  assign n11887 = n131 & n11886 ;
  assign n11889 = n11888 ^ n11887 ^ 1'b0 ;
  assign n11884 = ~n5340 & n8517 ;
  assign n11885 = n11884 ^ n11120 ^ 1'b0 ;
  assign n11890 = n11889 ^ n11885 ^ n2840 ;
  assign n11891 = n11890 ^ n8238 ^ n873 ;
  assign n11892 = n3031 & n11891 ;
  assign n11894 = n11893 ^ n11892 ^ 1'b0 ;
  assign n11895 = ~n7525 & n11894 ;
  assign n11896 = n11895 ^ x23 ^ 1'b0 ;
  assign n11897 = n2521 | n4811 ;
  assign n11898 = n6363 & n10040 ;
  assign n11899 = n11898 ^ n9615 ^ 1'b0 ;
  assign n11900 = n10068 ^ n4754 ^ 1'b0 ;
  assign n11901 = ~n390 & n11900 ;
  assign n11902 = ~n2020 & n6791 ;
  assign n11903 = n11902 ^ n7580 ^ 1'b0 ;
  assign n11904 = ~n6477 & n11369 ;
  assign n11905 = n5294 ^ n3994 ^ 1'b0 ;
  assign n11906 = n11905 ^ n2346 ^ 1'b0 ;
  assign n11907 = n11906 ^ n10084 ^ n5272 ;
  assign n11908 = n3602 & ~n7186 ;
  assign n11909 = n4583 | n11908 ;
  assign n11910 = n11909 ^ x67 ^ 1'b0 ;
  assign n11911 = n2608 & n4066 ;
  assign n11912 = ~n8441 & n11911 ;
  assign n11914 = n1909 ^ n977 ^ 1'b0 ;
  assign n11915 = n306 & n11914 ;
  assign n11913 = ~n3847 & n4174 ;
  assign n11916 = n11915 ^ n11913 ^ 1'b0 ;
  assign n11917 = ~n1154 & n8713 ;
  assign n11918 = ~n6455 & n11917 ;
  assign n11919 = n11918 ^ n3237 ^ n2887 ;
  assign n11920 = n11919 ^ n7269 ^ 1'b0 ;
  assign n11921 = ( n2136 & ~n10210 ) | ( n2136 & n11691 ) | ( ~n10210 & n11691 ) ;
  assign n11922 = n11921 ^ n618 ^ 1'b0 ;
  assign n11923 = n194 & n11922 ;
  assign n11927 = n1034 & n6126 ;
  assign n11924 = n1264 | n5052 ;
  assign n11925 = n11924 ^ n2140 ^ 1'b0 ;
  assign n11926 = ~n2810 & n11925 ;
  assign n11928 = n11927 ^ n11926 ^ 1'b0 ;
  assign n11929 = n2334 & ~n5203 ;
  assign n11930 = n11929 ^ n4370 ^ 1'b0 ;
  assign n11931 = n9573 ^ n8910 ^ 1'b0 ;
  assign n11932 = ( n5476 & n6351 ) | ( n5476 & ~n11931 ) | ( n6351 & ~n11931 ) ;
  assign n11933 = n3418 ^ n2025 ^ 1'b0 ;
  assign n11934 = n1586 | n7956 ;
  assign n11935 = n8859 | n11934 ;
  assign n11936 = ( n7077 & n11933 ) | ( n7077 & n11935 ) | ( n11933 & n11935 ) ;
  assign n11937 = ~n1253 & n11936 ;
  assign n11938 = n4396 ^ n307 ^ 1'b0 ;
  assign n11939 = n11937 | n11938 ;
  assign n11940 = n11612 | n11939 ;
  assign n11943 = n3475 ^ n3007 ^ x97 ;
  assign n11941 = n399 & n2350 ;
  assign n11942 = n5281 & n11941 ;
  assign n11944 = n11943 ^ n11942 ^ x9 ;
  assign n11945 = n4097 ^ n1596 ^ 1'b0 ;
  assign n11946 = n11054 ^ n1319 ^ n1110 ;
  assign n11947 = ~n3857 & n8316 ;
  assign n11948 = n915 & n11947 ;
  assign n11949 = n10640 ^ n1110 ^ 1'b0 ;
  assign n11950 = n7510 ^ n4300 ^ 1'b0 ;
  assign n11951 = n11949 & n11950 ;
  assign n11952 = n7278 ^ n908 ^ 1'b0 ;
  assign n11953 = n565 & ~n5151 ;
  assign n11954 = n794 & ~n10084 ;
  assign n11955 = n5835 & n11954 ;
  assign n11956 = n11955 ^ n3713 ^ 1'b0 ;
  assign n11957 = n1754 & ~n11956 ;
  assign n11958 = ( ~n5714 & n11300 ) | ( ~n5714 & n11957 ) | ( n11300 & n11957 ) ;
  assign n11959 = n655 & n6442 ;
  assign n11960 = ~n2733 & n11959 ;
  assign n11961 = n11960 ^ n1930 ^ 1'b0 ;
  assign n11962 = ( n11953 & n11958 ) | ( n11953 & ~n11961 ) | ( n11958 & ~n11961 ) ;
  assign n11963 = n8555 ^ n3762 ^ n3380 ;
  assign n11964 = n5386 | n11963 ;
  assign n11965 = ( n3684 & n9515 ) | ( n3684 & n11964 ) | ( n9515 & n11964 ) ;
  assign n11966 = ( n2184 & ~n6116 ) | ( n2184 & n11965 ) | ( ~n6116 & n11965 ) ;
  assign n11967 = n5302 | n11086 ;
  assign n11968 = n4323 | n11967 ;
  assign n11969 = n11966 & ~n11968 ;
  assign n11970 = n11962 & n11969 ;
  assign n11971 = n8141 ^ n4070 ^ 1'b0 ;
  assign n11972 = n1329 | n11971 ;
  assign n11973 = x82 & ~n458 ;
  assign n11974 = n11973 ^ n292 ^ 1'b0 ;
  assign n11975 = n11972 | n11974 ;
  assign n11976 = n11758 | n11975 ;
  assign n11977 = n380 & n3076 ;
  assign n11978 = ~x58 & n11977 ;
  assign n11979 = n2145 | n11978 ;
  assign n11983 = ~n319 & n2786 ;
  assign n11984 = n11983 ^ n2455 ^ 1'b0 ;
  assign n11985 = ( ~n2623 & n7000 ) | ( ~n2623 & n11984 ) | ( n7000 & n11984 ) ;
  assign n11980 = n8824 ^ n1860 ^ 1'b0 ;
  assign n11981 = n5576 | n11980 ;
  assign n11982 = ( n1018 & ~n7765 ) | ( n1018 & n11981 ) | ( ~n7765 & n11981 ) ;
  assign n11986 = n11985 ^ n11982 ^ 1'b0 ;
  assign n11987 = ~n9263 & n11986 ;
  assign n11988 = ~n5148 & n6635 ;
  assign n11989 = n6926 | n11988 ;
  assign n11990 = n1664 | n11989 ;
  assign n11991 = n11653 ^ n6109 ^ 1'b0 ;
  assign n11992 = n11990 & n11991 ;
  assign n11993 = n2466 ^ n2343 ^ n2096 ;
  assign n11994 = n11933 | n11993 ;
  assign n11995 = n8067 ^ n3727 ^ 1'b0 ;
  assign n11996 = n5948 ^ n2030 ^ 1'b0 ;
  assign n11997 = n8457 & n11996 ;
  assign n11998 = n5952 ^ n3070 ^ 1'b0 ;
  assign n11999 = n11997 | n11998 ;
  assign n12000 = n6649 ^ n3749 ^ 1'b0 ;
  assign n12001 = n4696 ^ n669 ^ 1'b0 ;
  assign n12002 = n1576 & ~n11539 ;
  assign n12003 = ( n6947 & ~n12001 ) | ( n6947 & n12002 ) | ( ~n12001 & n12002 ) ;
  assign n12004 = n2363 ^ n1971 ^ n307 ;
  assign n12005 = n12004 ^ n6446 ^ n4365 ;
  assign n12006 = n4482 & ~n12005 ;
  assign n12007 = n12006 ^ n7857 ^ 1'b0 ;
  assign n12008 = n5104 ^ n2970 ^ 1'b0 ;
  assign n12009 = n12008 ^ n8113 ^ 1'b0 ;
  assign n12010 = n12009 ^ n8331 ^ 1'b0 ;
  assign n12011 = n10674 | n12010 ;
  assign n12012 = n1885 ^ n826 ^ 1'b0 ;
  assign n12013 = n2970 & n12012 ;
  assign n12014 = n12013 ^ n5505 ^ 1'b0 ;
  assign n12015 = ~n5812 & n7216 ;
  assign n12016 = n12015 ^ n7050 ^ 1'b0 ;
  assign n12017 = n3296 & n5336 ;
  assign n12018 = n12017 ^ n2294 ^ 1'b0 ;
  assign n12019 = n12018 ^ n5024 ^ n1656 ;
  assign n12020 = n12019 ^ n9514 ^ n1923 ;
  assign n12021 = ( n666 & ~n7156 ) | ( n666 & n7730 ) | ( ~n7156 & n7730 ) ;
  assign n12022 = n12021 ^ n8571 ^ n5942 ;
  assign n12023 = n3753 & ~n12022 ;
  assign n12024 = ~n296 & n1499 ;
  assign n12025 = ~n8229 & n12024 ;
  assign n12026 = n4441 & ~n10597 ;
  assign n12027 = n10997 & ~n12026 ;
  assign n12028 = n538 & n11894 ;
  assign n12029 = n12028 ^ n11529 ^ 1'b0 ;
  assign n12030 = ~n207 & n2787 ;
  assign n12031 = ~n7775 & n12030 ;
  assign n12032 = ~n5379 & n6744 ;
  assign n12033 = n12032 ^ x27 ^ 1'b0 ;
  assign n12034 = n715 | n4127 ;
  assign n12035 = n12034 ^ n637 ^ 1'b0 ;
  assign n12036 = n6579 ^ n5137 ^ 1'b0 ;
  assign n12037 = ( ~n12033 & n12035 ) | ( ~n12033 & n12036 ) | ( n12035 & n12036 ) ;
  assign n12038 = n2863 ^ x119 ^ 1'b0 ;
  assign n12039 = n12037 & ~n12038 ;
  assign n12040 = n8264 | n11331 ;
  assign n12041 = n12039 | n12040 ;
  assign n12042 = n4335 & n6248 ;
  assign n12043 = n12042 ^ n8076 ^ 1'b0 ;
  assign n12044 = n3351 ^ n1274 ^ 1'b0 ;
  assign n12045 = n9761 | n12044 ;
  assign n12046 = n5938 | n12045 ;
  assign n12047 = ( n3595 & ~n12043 ) | ( n3595 & n12046 ) | ( ~n12043 & n12046 ) ;
  assign n12048 = n12047 ^ n9719 ^ 1'b0 ;
  assign n12049 = n12041 & ~n12048 ;
  assign n12050 = n9065 ^ n3552 ^ 1'b0 ;
  assign n12051 = n6641 & n12050 ;
  assign n12052 = n2699 & ~n10508 ;
  assign n12053 = n12052 ^ n7136 ^ 1'b0 ;
  assign n12054 = n6503 ^ n1990 ^ n803 ;
  assign n12055 = n227 & ~n12054 ;
  assign n12056 = n12055 ^ n9315 ^ 1'b0 ;
  assign n12058 = n10272 ^ n4545 ^ n1348 ;
  assign n12057 = n724 | n3564 ;
  assign n12059 = n12058 ^ n12057 ^ n3909 ;
  assign n12060 = n12059 ^ n1473 ^ 1'b0 ;
  assign n12061 = n12056 & n12060 ;
  assign n12063 = n6965 ^ n5423 ^ n1761 ;
  assign n12062 = n5920 ^ n2639 ^ n2072 ;
  assign n12064 = n12063 ^ n12062 ^ 1'b0 ;
  assign n12065 = n8429 & n12064 ;
  assign n12066 = n7484 ^ n5454 ^ n4799 ;
  assign n12067 = n207 & n12066 ;
  assign n12068 = ( n2929 & n9384 ) | ( n2929 & ~n9955 ) | ( n9384 & ~n9955 ) ;
  assign n12069 = ( n1193 & n4154 ) | ( n1193 & n12068 ) | ( n4154 & n12068 ) ;
  assign n12070 = n9327 ^ n6168 ^ 1'b0 ;
  assign n12071 = n4856 | n12070 ;
  assign n12072 = n3322 & ~n12071 ;
  assign n12073 = n2251 & n3892 ;
  assign n12074 = n9607 ^ n4341 ^ 1'b0 ;
  assign n12075 = n12073 & ~n12074 ;
  assign n12076 = n8938 ^ n6027 ^ n1628 ;
  assign n12077 = n6786 | n11469 ;
  assign n12078 = ( n6413 & n7380 ) | ( n6413 & ~n12077 ) | ( n7380 & ~n12077 ) ;
  assign n12079 = n1120 & n3542 ;
  assign n12080 = n6494 & n12079 ;
  assign n12081 = n4469 ^ n3055 ^ n2463 ;
  assign n12082 = n12081 ^ n10528 ^ 1'b0 ;
  assign n12083 = ~n12080 & n12082 ;
  assign n12084 = n6030 & ~n12083 ;
  assign n12085 = n10850 ^ n7622 ^ 1'b0 ;
  assign n12086 = n2332 & ~n12085 ;
  assign n12087 = n1445 & ~n10080 ;
  assign n12088 = n8126 ^ n6418 ^ n6256 ;
  assign n12089 = n12088 ^ n7951 ^ n3853 ;
  assign n12090 = n2727 | n7796 ;
  assign n12091 = n12089 | n12090 ;
  assign n12092 = n174 & ~n2541 ;
  assign n12093 = n7279 | n12092 ;
  assign n12094 = n12093 ^ n1503 ^ 1'b0 ;
  assign n12095 = ~n1533 & n6005 ;
  assign n12096 = n1002 & ~n12095 ;
  assign n12097 = n6438 & ~n6518 ;
  assign n12098 = n6751 ^ n1785 ^ 1'b0 ;
  assign n12099 = ~n2662 & n12098 ;
  assign n12100 = ( ~n8155 & n12097 ) | ( ~n8155 & n12099 ) | ( n12097 & n12099 ) ;
  assign n12101 = n5131 & n7513 ;
  assign n12102 = n4029 & n12101 ;
  assign n12103 = n4270 | n6655 ;
  assign n12104 = n2910 ^ x49 ^ 1'b0 ;
  assign n12105 = ~n7832 & n12104 ;
  assign n12106 = n12105 ^ n6835 ^ n6091 ;
  assign n12112 = n3972 & n4121 ;
  assign n12108 = n541 | n5631 ;
  assign n12107 = n8067 & n8765 ;
  assign n12109 = n12108 ^ n12107 ^ 1'b0 ;
  assign n12110 = x62 & ~n3207 ;
  assign n12111 = n12109 & n12110 ;
  assign n12113 = n12112 ^ n12111 ^ 1'b0 ;
  assign n12114 = ( n1803 & ~n8198 ) | ( n1803 & n11915 ) | ( ~n8198 & n11915 ) ;
  assign n12116 = n6503 ^ n4020 ^ 1'b0 ;
  assign n12115 = ~n3074 & n9295 ;
  assign n12117 = n12116 ^ n12115 ^ 1'b0 ;
  assign n12118 = ~n1274 & n7088 ;
  assign n12119 = n12118 ^ n1717 ^ 1'b0 ;
  assign n12120 = n12119 ^ n5230 ^ 1'b0 ;
  assign n12121 = n4827 & ~n12120 ;
  assign n12122 = ( n12114 & n12117 ) | ( n12114 & n12121 ) | ( n12117 & n12121 ) ;
  assign n12123 = n2069 ^ n1204 ^ n599 ;
  assign n12124 = n12123 ^ x108 ^ 1'b0 ;
  assign n12125 = n3219 & n12124 ;
  assign n12126 = n12125 ^ n1283 ^ 1'b0 ;
  assign n12127 = n2017 | n12126 ;
  assign n12128 = n4961 & n9269 ;
  assign n12129 = n11469 | n12128 ;
  assign n12130 = n12129 ^ n7216 ^ 1'b0 ;
  assign n12131 = n1670 & ~n3416 ;
  assign n12132 = n12131 ^ n2848 ^ 1'b0 ;
  assign n12133 = ( n845 & ~n9552 ) | ( n845 & n12132 ) | ( ~n9552 & n12132 ) ;
  assign n12134 = n12133 ^ n574 ^ 1'b0 ;
  assign n12135 = ~n5270 & n12134 ;
  assign n12136 = n1032 & n7845 ;
  assign n12137 = n12136 ^ n9756 ^ 1'b0 ;
  assign n12138 = ( n9622 & n12135 ) | ( n9622 & ~n12137 ) | ( n12135 & ~n12137 ) ;
  assign n12139 = n11441 ^ n3212 ^ 1'b0 ;
  assign n12140 = ~n3992 & n6754 ;
  assign n12141 = n12140 ^ n10926 ^ n2499 ;
  assign n12142 = ~n3500 & n5395 ;
  assign n12143 = n12142 ^ n912 ^ 1'b0 ;
  assign n12144 = n12143 ^ n830 ^ x32 ;
  assign n12145 = n9784 ^ n3235 ^ 1'b0 ;
  assign n12146 = ~n12144 & n12145 ;
  assign n12147 = ( n1296 & n6877 ) | ( n1296 & n12146 ) | ( n6877 & n12146 ) ;
  assign n12148 = n12147 ^ n6961 ^ 1'b0 ;
  assign n12149 = ~n12036 & n12148 ;
  assign n12150 = n12149 ^ n555 ^ 1'b0 ;
  assign n12151 = n10007 ^ n6472 ^ n1914 ;
  assign n12152 = n12151 ^ n5227 ^ n4594 ;
  assign n12153 = n12152 ^ n11816 ^ n5065 ;
  assign n12154 = ( n916 & n923 ) | ( n916 & n1575 ) | ( n923 & n1575 ) ;
  assign n12155 = n4699 & ~n12154 ;
  assign n12156 = n1749 & n12155 ;
  assign n12157 = n12156 ^ n4770 ^ n155 ;
  assign n12158 = n6275 & n12157 ;
  assign n12159 = n12158 ^ n4964 ^ n3003 ;
  assign n12160 = ( ~n131 & n973 ) | ( ~n131 & n12159 ) | ( n973 & n12159 ) ;
  assign n12161 = n12160 ^ n7190 ^ n6145 ;
  assign n12162 = n9211 ^ n7214 ^ 1'b0 ;
  assign n12163 = ~n2319 & n12162 ;
  assign n12164 = n11327 ^ n4837 ^ 1'b0 ;
  assign n12165 = n1514 & n11231 ;
  assign n12166 = n3423 | n6953 ;
  assign n12167 = n12166 ^ n8422 ^ 1'b0 ;
  assign n12168 = ~x108 & n12167 ;
  assign n12169 = n1466 & n3357 ;
  assign n12170 = n12169 ^ n2627 ^ 1'b0 ;
  assign n12171 = n12170 ^ n3424 ^ 1'b0 ;
  assign n12172 = n12168 | n12171 ;
  assign n12173 = n8008 & ~n12076 ;
  assign n12174 = n12173 ^ n10374 ^ 1'b0 ;
  assign n12176 = x119 & ~n3738 ;
  assign n12175 = n719 & ~n1870 ;
  assign n12177 = n12176 ^ n12175 ^ 1'b0 ;
  assign n12178 = n9485 ^ n9226 ^ 1'b0 ;
  assign n12179 = ~n10004 & n12178 ;
  assign n12182 = n1561 & ~n6093 ;
  assign n12183 = ~x28 & n12182 ;
  assign n12181 = ~n3744 & n4891 ;
  assign n12184 = n12183 ^ n12181 ^ 1'b0 ;
  assign n12180 = ~n1542 & n4577 ;
  assign n12185 = n12184 ^ n12180 ^ 1'b0 ;
  assign n12186 = n1870 & ~n3402 ;
  assign n12187 = ( x51 & ~n2923 ) | ( x51 & n4230 ) | ( ~n2923 & n4230 ) ;
  assign n12188 = n12187 ^ n5704 ^ n5449 ;
  assign n12189 = n10370 ^ n4527 ^ 1'b0 ;
  assign n12190 = n6330 & n12189 ;
  assign n12191 = n3188 | n7159 ;
  assign n12192 = n5771 | n12191 ;
  assign n12195 = n9163 ^ n5124 ^ 1'b0 ;
  assign n12193 = n2420 & n5596 ;
  assign n12194 = n12193 ^ n7724 ^ 1'b0 ;
  assign n12196 = n12195 ^ n12194 ^ n1966 ;
  assign n12197 = n9384 & n10020 ;
  assign n12198 = n12197 ^ n620 ^ 1'b0 ;
  assign n12199 = ( n4717 & n8634 ) | ( n4717 & n12198 ) | ( n8634 & n12198 ) ;
  assign n12200 = n1432 & ~n9677 ;
  assign n12201 = n12200 ^ n2582 ^ 1'b0 ;
  assign n12202 = n5212 & n12201 ;
  assign n12203 = ~n12199 & n12202 ;
  assign n12204 = n11086 ^ n2394 ^ 1'b0 ;
  assign n12205 = n12204 ^ n1527 ^ 1'b0 ;
  assign n12206 = n12203 | n12205 ;
  assign n12209 = n10372 ^ n3295 ^ n1601 ;
  assign n12207 = n4729 ^ n631 ^ 1'b0 ;
  assign n12208 = n1673 & ~n12207 ;
  assign n12210 = n12209 ^ n12208 ^ 1'b0 ;
  assign n12211 = n270 | n5936 ;
  assign n12212 = n12211 ^ n1792 ^ 1'b0 ;
  assign n12213 = n11406 ^ n3547 ^ n2377 ;
  assign n12214 = ~n6344 & n12213 ;
  assign n12215 = n12212 & n12214 ;
  assign n12217 = x117 & ~n9594 ;
  assign n12218 = n139 & n12217 ;
  assign n12219 = n8191 & ~n12218 ;
  assign n12216 = n667 | n4175 ;
  assign n12220 = n12219 ^ n12216 ^ 1'b0 ;
  assign n12221 = n5323 ^ n1599 ^ 1'b0 ;
  assign n12222 = n2798 ^ n2072 ^ n1516 ;
  assign n12223 = n8297 ^ n5909 ^ n1859 ;
  assign n12224 = ( n2859 & n12222 ) | ( n2859 & n12223 ) | ( n12222 & n12223 ) ;
  assign n12225 = ( ~n2366 & n8475 ) | ( ~n2366 & n11967 ) | ( n8475 & n11967 ) ;
  assign n12226 = n12225 ^ n7574 ^ 1'b0 ;
  assign n12227 = n4458 | n12226 ;
  assign n12228 = n12227 ^ n7864 ^ 1'b0 ;
  assign n12229 = n1649 & n4010 ;
  assign n12230 = n2093 ^ n723 ^ 1'b0 ;
  assign n12231 = n2968 & n12230 ;
  assign n12232 = n4493 ^ n3354 ^ 1'b0 ;
  assign n12233 = n5036 & ~n12232 ;
  assign n12234 = n3835 ^ n2515 ^ 1'b0 ;
  assign n12235 = n10049 & n12234 ;
  assign n12236 = n5563 & n6261 ;
  assign n12237 = ~n12235 & n12236 ;
  assign n12238 = ~n12233 & n12237 ;
  assign n12239 = n3988 ^ x114 ^ 1'b0 ;
  assign n12240 = ~n5701 & n12239 ;
  assign n12241 = n12240 ^ n4715 ^ 1'b0 ;
  assign n12244 = n3283 | n6378 ;
  assign n12245 = n3677 & ~n12244 ;
  assign n12242 = n2722 | n9365 ;
  assign n12243 = n8287 | n12242 ;
  assign n12246 = n12245 ^ n12243 ^ 1'b0 ;
  assign n12255 = n1083 & ~n9600 ;
  assign n12256 = n5840 & n12255 ;
  assign n12251 = n3215 ^ n214 ^ 1'b0 ;
  assign n12252 = n241 | n12251 ;
  assign n12250 = n2545 ^ n2092 ^ 1'b0 ;
  assign n12253 = n12252 ^ n12250 ^ n10733 ;
  assign n12247 = ~n531 & n2212 ;
  assign n12248 = n12247 ^ n5106 ^ 1'b0 ;
  assign n12249 = n1645 & n12248 ;
  assign n12254 = n12253 ^ n12249 ^ 1'b0 ;
  assign n12257 = n12256 ^ n12254 ^ n2194 ;
  assign n12259 = ~n948 & n9522 ;
  assign n12258 = ~n749 & n3351 ;
  assign n12260 = n12259 ^ n12258 ^ n4689 ;
  assign n12261 = n5045 ^ n4770 ^ n1223 ;
  assign n12262 = ~n10004 & n12261 ;
  assign n12263 = n12260 & n12262 ;
  assign n12264 = n5686 | n10850 ;
  assign n12265 = n9670 & ~n12264 ;
  assign n12266 = ( n924 & ~n3649 ) | ( n924 & n5148 ) | ( ~n3649 & n5148 ) ;
  assign n12267 = n12266 ^ n10315 ^ n2296 ;
  assign n12274 = n4287 ^ n2215 ^ 1'b0 ;
  assign n12275 = n4252 & n12274 ;
  assign n12276 = ( n498 & n1004 ) | ( n498 & ~n12275 ) | ( n1004 & ~n12275 ) ;
  assign n12277 = n12276 ^ n3778 ^ 1'b0 ;
  assign n12278 = n9308 & ~n12277 ;
  assign n12271 = n2498 & ~n4541 ;
  assign n12272 = ~n1591 & n12271 ;
  assign n12270 = n8858 ^ n7096 ^ 1'b0 ;
  assign n12268 = n7802 & n10497 ;
  assign n12269 = n1374 & n12268 ;
  assign n12273 = n12272 ^ n12270 ^ n12269 ;
  assign n12279 = n12278 ^ n12273 ^ n7067 ;
  assign n12280 = n4141 & n10764 ;
  assign n12281 = n6207 | n8254 ;
  assign n12282 = n12281 ^ n746 ^ 1'b0 ;
  assign n12283 = ~n543 & n5026 ;
  assign n12284 = n12283 ^ n3595 ^ x19 ;
  assign n12285 = n12284 ^ n5878 ^ 1'b0 ;
  assign n12286 = n1236 ^ n908 ^ 1'b0 ;
  assign n12287 = n1547 | n12286 ;
  assign n12288 = n1438 | n12287 ;
  assign n12289 = n149 | n12288 ;
  assign n12290 = ( n11748 & ~n12285 ) | ( n11748 & n12289 ) | ( ~n12285 & n12289 ) ;
  assign n12291 = n12290 ^ n4841 ^ n4671 ;
  assign n12292 = ~n11109 & n12291 ;
  assign n12293 = ~n3281 & n12292 ;
  assign n12294 = n11766 ^ n3265 ^ n522 ;
  assign n12295 = ( n2151 & ~n3748 ) | ( n2151 & n4150 ) | ( ~n3748 & n4150 ) ;
  assign n12296 = ~n3249 & n8571 ;
  assign n12297 = ~n5753 & n12296 ;
  assign n12298 = n12297 ^ n5057 ^ n2950 ;
  assign n12299 = ( x108 & n12295 ) | ( x108 & ~n12298 ) | ( n12295 & ~n12298 ) ;
  assign n12300 = ( n1121 & n7628 ) | ( n1121 & n8899 ) | ( n7628 & n8899 ) ;
  assign n12301 = ( n3010 & ~n3163 ) | ( n3010 & n3677 ) | ( ~n3163 & n3677 ) ;
  assign n12302 = n12301 ^ n5391 ^ n797 ;
  assign n12310 = ( ~n2508 & n4060 ) | ( ~n2508 & n8620 ) | ( n4060 & n8620 ) ;
  assign n12308 = n6761 ^ n5800 ^ n3739 ;
  assign n12309 = ~n6705 & n12308 ;
  assign n12311 = n12310 ^ n12309 ^ n7148 ;
  assign n12303 = ~n2423 & n8722 ;
  assign n12304 = n12303 ^ n11030 ^ 1'b0 ;
  assign n12305 = n6511 | n9477 ;
  assign n12306 = n6048 | n12305 ;
  assign n12307 = ~n12304 & n12306 ;
  assign n12312 = n12311 ^ n12307 ^ 1'b0 ;
  assign n12315 = n4327 ^ n3192 ^ 1'b0 ;
  assign n12316 = n7959 | n12315 ;
  assign n12313 = ( n692 & n2036 ) | ( n692 & ~n7820 ) | ( n2036 & ~n7820 ) ;
  assign n12314 = n9357 & ~n12313 ;
  assign n12317 = n12316 ^ n12314 ^ 1'b0 ;
  assign n12318 = n3924 ^ n679 ^ 1'b0 ;
  assign n12319 = ~n4182 & n12318 ;
  assign n12320 = n12319 ^ n10650 ^ n8785 ;
  assign n12321 = ( n4761 & n5301 ) | ( n4761 & ~n11561 ) | ( n5301 & ~n11561 ) ;
  assign n12322 = n8733 & ~n12321 ;
  assign n12323 = ~n10381 & n12147 ;
  assign n12324 = n4242 & n5735 ;
  assign n12325 = ( n7743 & n12323 ) | ( n7743 & n12324 ) | ( n12323 & n12324 ) ;
  assign n12326 = n3461 & ~n6083 ;
  assign n12327 = n8992 & n12326 ;
  assign n12328 = n3982 ^ n618 ^ 1'b0 ;
  assign n12329 = n4502 ^ n2254 ^ n1717 ;
  assign n12330 = n4269 ^ n3033 ^ 1'b0 ;
  assign n12331 = ( n12328 & ~n12329 ) | ( n12328 & n12330 ) | ( ~n12329 & n12330 ) ;
  assign n12332 = n12331 ^ n7816 ^ n1936 ;
  assign n12333 = n7682 & n12332 ;
  assign n12334 = n3437 | n12333 ;
  assign n12335 = n12334 ^ n2346 ^ 1'b0 ;
  assign n12336 = n12335 ^ n3173 ^ 1'b0 ;
  assign n12337 = ( ~n1354 & n5213 ) | ( ~n1354 & n5913 ) | ( n5213 & n5913 ) ;
  assign n12338 = n12336 & ~n12337 ;
  assign n12339 = ( ~n409 & n1291 ) | ( ~n409 & n5897 ) | ( n1291 & n5897 ) ;
  assign n12340 = n12339 ^ n5099 ^ 1'b0 ;
  assign n12341 = ~n6306 & n12340 ;
  assign n12342 = n9986 ^ n1796 ^ 1'b0 ;
  assign n12343 = n4897 & n8049 ;
  assign n12344 = ~n5102 & n12343 ;
  assign n12345 = n10426 | n12344 ;
  assign n12346 = ~n1973 & n12345 ;
  assign n12347 = n9523 | n12346 ;
  assign n12348 = n12347 ^ n8681 ^ n6289 ;
  assign n12349 = ~n11778 & n12348 ;
  assign n12350 = n12349 ^ n1829 ^ 1'b0 ;
  assign n12351 = ( ~n6495 & n9645 ) | ( ~n6495 & n12350 ) | ( n9645 & n12350 ) ;
  assign n12352 = n2229 | n8816 ;
  assign n12353 = n12352 ^ n1445 ^ 1'b0 ;
  assign n12354 = n4181 & ~n4784 ;
  assign n12355 = n12354 ^ n1515 ^ 1'b0 ;
  assign n12356 = ( n3837 & ~n8245 ) | ( n3837 & n12355 ) | ( ~n8245 & n12355 ) ;
  assign n12364 = n6658 ^ n260 ^ n218 ;
  assign n12361 = ( n784 & n1920 ) | ( n784 & ~n8262 ) | ( n1920 & ~n8262 ) ;
  assign n12362 = n12361 ^ n4255 ^ 1'b0 ;
  assign n12357 = n5013 ^ n2118 ^ n1590 ;
  assign n12358 = n1023 & n12357 ;
  assign n12359 = n6469 & n12358 ;
  assign n12360 = n281 & ~n12359 ;
  assign n12363 = n12362 ^ n12360 ^ 1'b0 ;
  assign n12365 = n12364 ^ n12363 ^ n8535 ;
  assign n12366 = ( n1581 & n2113 ) | ( n1581 & n4677 ) | ( n2113 & n4677 ) ;
  assign n12367 = n3544 & ~n12366 ;
  assign n12368 = ~n8113 & n12367 ;
  assign n12369 = ( n8801 & n10708 ) | ( n8801 & n12368 ) | ( n10708 & n12368 ) ;
  assign n12370 = n2467 & ~n2682 ;
  assign n12371 = n12370 ^ n993 ^ 1'b0 ;
  assign n12372 = n12371 ^ n2634 ^ 1'b0 ;
  assign n12373 = n12372 ^ n9098 ^ n2194 ;
  assign n12374 = n12373 ^ n4175 ^ 1'b0 ;
  assign n12375 = n6306 | n12374 ;
  assign n12376 = n6947 ^ n3365 ^ 1'b0 ;
  assign n12377 = ~n8964 & n12376 ;
  assign n12378 = n12375 & n12377 ;
  assign n12383 = n3331 ^ n1073 ^ 1'b0 ;
  assign n12379 = n4713 & ~n7629 ;
  assign n12380 = ~n380 & n12379 ;
  assign n12381 = ~n5249 & n12380 ;
  assign n12382 = n12381 ^ n12290 ^ n10698 ;
  assign n12384 = n12383 ^ n12382 ^ n3488 ;
  assign n12385 = n3260 & ~n10212 ;
  assign n12386 = ~n2616 & n12385 ;
  assign n12387 = ( ~n1515 & n6164 ) | ( ~n1515 & n12386 ) | ( n6164 & n12386 ) ;
  assign n12388 = n512 ^ x55 ^ 1'b0 ;
  assign n12389 = ~n9331 & n12388 ;
  assign n12390 = ~n7285 & n12389 ;
  assign n12391 = n4416 ^ n3349 ^ n218 ;
  assign n12392 = ~n2499 & n7735 ;
  assign n12393 = n12392 ^ n9026 ^ n5476 ;
  assign n12394 = n265 | n1423 ;
  assign n12395 = n12394 ^ n328 ^ 1'b0 ;
  assign n12396 = n8158 | n12395 ;
  assign n12397 = n12396 ^ n4290 ^ 1'b0 ;
  assign n12398 = n1038 & ~n3554 ;
  assign n12399 = ~n12397 & n12398 ;
  assign n12400 = n3896 ^ n2149 ^ n213 ;
  assign n12401 = n8957 & ~n9312 ;
  assign n12402 = ~n3831 & n5234 ;
  assign n12403 = n10895 & n12402 ;
  assign n12404 = ( ~n1683 & n2240 ) | ( ~n1683 & n11392 ) | ( n2240 & n11392 ) ;
  assign n12405 = ( ~n4869 & n12403 ) | ( ~n4869 & n12404 ) | ( n12403 & n12404 ) ;
  assign n12406 = n12405 ^ n1427 ^ 1'b0 ;
  assign n12407 = ( n5128 & ~n6178 ) | ( n5128 & n12406 ) | ( ~n6178 & n12406 ) ;
  assign n12408 = n9427 | n10209 ;
  assign n12409 = n8434 | n12408 ;
  assign n12410 = n12409 ^ x59 ^ 1'b0 ;
  assign n12411 = ~n10092 & n12410 ;
  assign n12412 = n574 & ~n9326 ;
  assign n12413 = n5915 | n8839 ;
  assign n12414 = n12413 ^ n5235 ^ 1'b0 ;
  assign n12415 = ~n9341 & n12414 ;
  assign n12416 = n12415 ^ n9324 ^ 1'b0 ;
  assign n12417 = ( ~x85 & n6469 ) | ( ~x85 & n12416 ) | ( n6469 & n12416 ) ;
  assign n12418 = n1845 | n5287 ;
  assign n12419 = n5421 ^ n1057 ^ 1'b0 ;
  assign n12420 = n3385 & ~n12419 ;
  assign n12421 = ( n4387 & ~n12418 ) | ( n4387 & n12420 ) | ( ~n12418 & n12420 ) ;
  assign n12422 = n4448 & ~n11150 ;
  assign n12423 = ~n11856 & n12422 ;
  assign n12424 = ( ~n1548 & n8973 ) | ( ~n1548 & n10881 ) | ( n8973 & n10881 ) ;
  assign n12426 = n2143 & n5421 ;
  assign n12427 = ( n588 & ~n1541 ) | ( n588 & n12426 ) | ( ~n1541 & n12426 ) ;
  assign n12425 = ( n370 & n4307 ) | ( n370 & n4313 ) | ( n4307 & n4313 ) ;
  assign n12428 = n12427 ^ n12425 ^ 1'b0 ;
  assign n12429 = n5948 | n12428 ;
  assign n12430 = n12429 ^ n1781 ^ 1'b0 ;
  assign n12431 = n7693 & n7948 ;
  assign n12432 = ( n5743 & ~n7380 ) | ( n5743 & n8243 ) | ( ~n7380 & n8243 ) ;
  assign n12433 = n12431 & ~n12432 ;
  assign n12434 = n8999 ^ n1626 ^ 1'b0 ;
  assign n12435 = ~n12433 & n12434 ;
  assign n12436 = n994 | n1915 ;
  assign n12437 = n12436 ^ n8065 ^ 1'b0 ;
  assign n12438 = ~n2897 & n4014 ;
  assign n12439 = n5873 & n6186 ;
  assign n12440 = ~n9551 & n12439 ;
  assign n12441 = n5910 | n12440 ;
  assign n12442 = n5286 & n11507 ;
  assign n12443 = n12441 & n12442 ;
  assign n12444 = ( n3602 & n4129 ) | ( n3602 & n11209 ) | ( n4129 & n11209 ) ;
  assign n12448 = n2455 & ~n3035 ;
  assign n12449 = ~n4747 & n12448 ;
  assign n12450 = ( n1214 & ~n5718 ) | ( n1214 & n12449 ) | ( ~n5718 & n12449 ) ;
  assign n12446 = n9096 ^ n3128 ^ 1'b0 ;
  assign n12445 = n3297 & n12258 ;
  assign n12447 = n12446 ^ n12445 ^ 1'b0 ;
  assign n12451 = n12450 ^ n12447 ^ n9558 ;
  assign n12452 = n7521 | n12451 ;
  assign n12453 = n7721 & ~n12452 ;
  assign n12454 = ~x67 & n5370 ;
  assign n12455 = ~n953 & n6779 ;
  assign n12456 = n12455 ^ n8535 ^ 1'b0 ;
  assign n12457 = ( ~n3071 & n12454 ) | ( ~n3071 & n12456 ) | ( n12454 & n12456 ) ;
  assign n12458 = n12453 & ~n12457 ;
  assign n12459 = n476 | n1905 ;
  assign n12460 = n5889 & ~n12459 ;
  assign n12461 = n7913 | n12460 ;
  assign n12462 = n506 & ~n12461 ;
  assign n12463 = ( n230 & ~n2744 ) | ( n230 & n8308 ) | ( ~n2744 & n8308 ) ;
  assign n12464 = n3463 & ~n12463 ;
  assign n12465 = n12464 ^ x114 ^ 1'b0 ;
  assign n12466 = n12465 ^ n6032 ^ 1'b0 ;
  assign n12467 = n4869 | n12466 ;
  assign n12468 = ( ~n5442 & n6555 ) | ( ~n5442 & n10494 ) | ( n6555 & n10494 ) ;
  assign n12469 = n12468 ^ n6359 ^ 1'b0 ;
  assign n12470 = n8570 | n12469 ;
  assign n12471 = ( n550 & n3633 ) | ( n550 & n12470 ) | ( n3633 & n12470 ) ;
  assign n12472 = n696 | n6221 ;
  assign n12473 = n2697 & n8736 ;
  assign n12474 = n9372 ^ n5554 ^ 1'b0 ;
  assign n12475 = ~n1624 & n12474 ;
  assign n12476 = n12475 ^ n1454 ^ 1'b0 ;
  assign n12477 = n12476 ^ n12184 ^ 1'b0 ;
  assign n12478 = ( ~n12472 & n12473 ) | ( ~n12472 & n12477 ) | ( n12473 & n12477 ) ;
  assign n12479 = n10762 ^ n8359 ^ 1'b0 ;
  assign n12480 = n10351 ^ n8512 ^ 1'b0 ;
  assign n12481 = n9041 & n12480 ;
  assign n12482 = n4394 | n12481 ;
  assign n12483 = n11548 ^ n3909 ^ 1'b0 ;
  assign n12484 = n1198 | n9984 ;
  assign n12485 = n12484 ^ n3580 ^ n2650 ;
  assign n12486 = n262 | n9475 ;
  assign n12487 = n862 | n12486 ;
  assign n12488 = ~n2013 & n12487 ;
  assign n12499 = n6711 ^ n6331 ^ n3439 ;
  assign n12500 = ( ~n349 & n1783 ) | ( ~n349 & n6811 ) | ( n1783 & n6811 ) ;
  assign n12501 = n12499 & ~n12500 ;
  assign n12494 = n1288 & n6316 ;
  assign n12495 = n12494 ^ x126 ^ 1'b0 ;
  assign n12496 = n10272 | n12495 ;
  assign n12489 = n4665 ^ n2500 ^ 1'b0 ;
  assign n12490 = x101 & ~n3001 ;
  assign n12491 = ~n12489 & n12490 ;
  assign n12492 = n7066 ^ n2422 ^ 1'b0 ;
  assign n12493 = n12491 & ~n12492 ;
  assign n12497 = n12496 ^ n12493 ^ 1'b0 ;
  assign n12498 = n4811 | n12497 ;
  assign n12502 = n12501 ^ n12498 ^ 1'b0 ;
  assign n12503 = n4747 ^ n2110 ^ x18 ;
  assign n12504 = ( n1721 & n8043 ) | ( n1721 & n12503 ) | ( n8043 & n12503 ) ;
  assign n12505 = ( n3696 & ~n6371 ) | ( n3696 & n12504 ) | ( ~n6371 & n12504 ) ;
  assign n12506 = n8196 & ~n12505 ;
  assign n12507 = n12033 ^ n8611 ^ 1'b0 ;
  assign n12508 = ( n2421 & n6049 ) | ( n2421 & ~n7763 ) | ( n6049 & ~n7763 ) ;
  assign n12509 = x50 & ~n12508 ;
  assign n12510 = n1402 & n12509 ;
  assign n12511 = n7947 & n12510 ;
  assign n12512 = n7968 ^ n1299 ^ 1'b0 ;
  assign n12513 = n2978 | n12512 ;
  assign n12514 = ( x14 & ~n7380 ) | ( x14 & n12513 ) | ( ~n7380 & n12513 ) ;
  assign n12515 = ( n3831 & ~n5057 ) | ( n3831 & n12514 ) | ( ~n5057 & n12514 ) ;
  assign n12516 = n7930 ^ n5690 ^ 1'b0 ;
  assign n12517 = n12515 | n12516 ;
  assign n12518 = n2011 & n5958 ;
  assign n12519 = n12518 ^ n11726 ^ 1'b0 ;
  assign n12520 = n306 & ~n9324 ;
  assign n12521 = n12520 ^ n575 ^ 1'b0 ;
  assign n12522 = ( ~n1423 & n8695 ) | ( ~n1423 & n12521 ) | ( n8695 & n12521 ) ;
  assign n12523 = n2163 ^ n755 ^ 1'b0 ;
  assign n12524 = ~n12522 & n12523 ;
  assign n12527 = n2988 & ~n11191 ;
  assign n12528 = n2373 & n12527 ;
  assign n12525 = n7786 ^ n7087 ^ n3587 ;
  assign n12526 = ( ~n4990 & n5886 ) | ( ~n4990 & n12525 ) | ( n5886 & n12525 ) ;
  assign n12529 = n12528 ^ n12526 ^ n3362 ;
  assign n12530 = ( n9622 & n12524 ) | ( n9622 & n12529 ) | ( n12524 & n12529 ) ;
  assign n12531 = ( n1900 & n6656 ) | ( n1900 & ~n6726 ) | ( n6656 & ~n6726 ) ;
  assign n12532 = ~n5607 & n12531 ;
  assign n12533 = ( ~n739 & n751 ) | ( ~n739 & n12532 ) | ( n751 & n12532 ) ;
  assign n12537 = n8762 ^ n5175 ^ n360 ;
  assign n12534 = n6442 & n6843 ;
  assign n12535 = n3566 & n12534 ;
  assign n12536 = ( n2019 & n4055 ) | ( n2019 & ~n12535 ) | ( n4055 & ~n12535 ) ;
  assign n12538 = n12537 ^ n12536 ^ n10185 ;
  assign n12540 = n1330 & ~n4744 ;
  assign n12539 = n8092 | n9406 ;
  assign n12541 = n12540 ^ n12539 ^ n675 ;
  assign n12542 = n7016 & ~n12541 ;
  assign n12543 = n12542 ^ n1601 ^ 1'b0 ;
  assign n12544 = n12543 ^ n10512 ^ n1084 ;
  assign n12545 = n3556 & ~n4921 ;
  assign n12546 = n12545 ^ n10730 ^ 1'b0 ;
  assign n12547 = x17 & ~n5067 ;
  assign n12548 = n12547 ^ n1025 ^ 1'b0 ;
  assign n12549 = n1478 | n8836 ;
  assign n12550 = n12549 ^ n1501 ^ n570 ;
  assign n12551 = n12550 ^ n5080 ^ 1'b0 ;
  assign n12552 = n9413 & n12551 ;
  assign n12553 = x122 ^ x111 ^ 1'b0 ;
  assign n12554 = ~n7388 & n12553 ;
  assign n12555 = n3242 & n12554 ;
  assign n12556 = n12555 ^ n7076 ^ 1'b0 ;
  assign n12557 = ~n2077 & n2481 ;
  assign n12558 = n2315 ^ n2006 ^ 1'b0 ;
  assign n12559 = n7419 | n12558 ;
  assign n12560 = n12559 ^ n8638 ^ 1'b0 ;
  assign n12561 = n12560 ^ n10825 ^ n1756 ;
  assign n12562 = ( ~n141 & n5374 ) | ( ~n141 & n8199 ) | ( n5374 & n8199 ) ;
  assign n12565 = n10234 ^ n10093 ^ 1'b0 ;
  assign n12566 = x1 & n12565 ;
  assign n12567 = n12566 ^ n10980 ^ n6279 ;
  assign n12563 = n3098 ^ x53 ^ 1'b0 ;
  assign n12564 = n7913 & ~n12563 ;
  assign n12568 = n12567 ^ n12564 ^ 1'b0 ;
  assign n12569 = ~n3848 & n9781 ;
  assign n12570 = n12121 ^ n9693 ^ 1'b0 ;
  assign n12571 = n9123 & ~n12570 ;
  assign n12572 = n5702 ^ n1182 ^ x93 ;
  assign n12573 = ( ~n3264 & n9713 ) | ( ~n3264 & n12572 ) | ( n9713 & n12572 ) ;
  assign n12574 = ( n7902 & n10469 ) | ( n7902 & n12157 ) | ( n10469 & n12157 ) ;
  assign n12575 = ( n4696 & n11822 ) | ( n4696 & ~n12559 ) | ( n11822 & ~n12559 ) ;
  assign n12576 = n945 | n3352 ;
  assign n12577 = n12576 ^ n7530 ^ 1'b0 ;
  assign n12578 = ~n10825 & n12577 ;
  assign n12579 = n12578 ^ n131 ^ 1'b0 ;
  assign n12580 = ~n6864 & n12579 ;
  assign n12581 = ~n1580 & n6239 ;
  assign n12582 = ~n7064 & n12581 ;
  assign n12585 = n2778 ^ n2545 ^ 1'b0 ;
  assign n12583 = n4093 ^ n3287 ^ n1065 ;
  assign n12584 = ( n3534 & ~n9662 ) | ( n3534 & n12583 ) | ( ~n9662 & n12583 ) ;
  assign n12586 = n12585 ^ n12584 ^ n5369 ;
  assign n12587 = ( n7075 & ~n9216 ) | ( n7075 & n11879 ) | ( ~n9216 & n11879 ) ;
  assign n12588 = n10720 ^ n4261 ^ 1'b0 ;
  assign n12589 = n3943 & n12588 ;
  assign n12590 = n3212 & n12589 ;
  assign n12591 = n4608 & ~n10077 ;
  assign n12592 = n12590 & n12591 ;
  assign n12593 = n6095 ^ n2801 ^ n2770 ;
  assign n12594 = n3892 & n12593 ;
  assign n12595 = ( n327 & n455 ) | ( n327 & n936 ) | ( n455 & n936 ) ;
  assign n12596 = n11599 & n12595 ;
  assign n12597 = n12596 ^ n2811 ^ 1'b0 ;
  assign n12598 = n12597 ^ n9838 ^ n694 ;
  assign n12599 = n5381 & ~n12598 ;
  assign n12600 = n12599 ^ n11012 ^ n2638 ;
  assign n12601 = n12567 ^ n3598 ^ 1'b0 ;
  assign n12602 = n6198 | n12601 ;
  assign n12603 = ~n1217 & n2271 ;
  assign n12604 = n1227 ^ n315 ^ 1'b0 ;
  assign n12605 = n6384 & n12604 ;
  assign n12606 = n5665 & ~n12605 ;
  assign n12607 = n12603 & ~n12606 ;
  assign n12608 = n466 & n12607 ;
  assign n12609 = ( n9205 & n10203 ) | ( n9205 & n12608 ) | ( n10203 & n12608 ) ;
  assign n12610 = n4254 ^ n3575 ^ 1'b0 ;
  assign n12611 = n1615 & ~n12610 ;
  assign n12612 = ( ~n5490 & n8033 ) | ( ~n5490 & n12611 ) | ( n8033 & n12611 ) ;
  assign n12613 = ( n4463 & ~n7724 ) | ( n4463 & n12612 ) | ( ~n7724 & n12612 ) ;
  assign n12614 = n10698 ^ n4539 ^ 1'b0 ;
  assign n12615 = n537 & n12614 ;
  assign n12616 = n12615 ^ n4086 ^ 1'b0 ;
  assign n12617 = n11452 ^ n11125 ^ 1'b0 ;
  assign n12618 = n8390 | n12617 ;
  assign n12619 = n12616 | n12618 ;
  assign n12620 = n12619 ^ n5149 ^ 1'b0 ;
  assign n12621 = ( n1740 & ~n2658 ) | ( n1740 & n4941 ) | ( ~n2658 & n4941 ) ;
  assign n12622 = ( n10029 & ~n12284 ) | ( n10029 & n12621 ) | ( ~n12284 & n12621 ) ;
  assign n12623 = ~n11701 & n12622 ;
  assign n12624 = n1573 & n12623 ;
  assign n12625 = ( ~n2625 & n3176 ) | ( ~n2625 & n7484 ) | ( n3176 & n7484 ) ;
  assign n12626 = n12625 ^ n2396 ^ n1692 ;
  assign n12627 = n10558 ^ n7791 ^ 1'b0 ;
  assign n12628 = n3567 ^ n552 ^ 1'b0 ;
  assign n12629 = ( n1105 & n2807 ) | ( n1105 & ~n12628 ) | ( n2807 & ~n12628 ) ;
  assign n12630 = n448 & n2567 ;
  assign n12631 = n752 ^ n469 ^ 1'b0 ;
  assign n12632 = n6034 | n12631 ;
  assign n12633 = n12630 & ~n12632 ;
  assign n12634 = n8108 | n12633 ;
  assign n12635 = n6759 ^ n523 ^ 1'b0 ;
  assign n12636 = n12635 ^ n5104 ^ 1'b0 ;
  assign n12637 = n211 & ~n4653 ;
  assign n12638 = n3111 & ~n8095 ;
  assign n12639 = n12637 & n12638 ;
  assign n12640 = n12639 ^ n4605 ^ n1468 ;
  assign n12641 = ~n1542 & n5097 ;
  assign n12642 = n7947 & n9429 ;
  assign n12643 = ~n11150 & n12642 ;
  assign n12644 = ( n4932 & n8791 ) | ( n4932 & ~n10404 ) | ( n8791 & ~n10404 ) ;
  assign n12645 = n4166 & n7433 ;
  assign n12649 = ~n800 & n11257 ;
  assign n12650 = n12649 ^ n2503 ^ 1'b0 ;
  assign n12651 = ~n8534 & n12650 ;
  assign n12646 = ( n1824 & n3740 ) | ( n1824 & n6144 ) | ( n3740 & n6144 ) ;
  assign n12647 = ( ~n1054 & n9706 ) | ( ~n1054 & n12646 ) | ( n9706 & n12646 ) ;
  assign n12648 = n12647 ^ n5782 ^ n4933 ;
  assign n12652 = n12651 ^ n12648 ^ n8702 ;
  assign n12653 = n11151 & ~n12057 ;
  assign n12654 = n11870 ^ n9662 ^ 1'b0 ;
  assign n12655 = n10158 ^ n3173 ^ 1'b0 ;
  assign n12656 = n620 ^ n516 ^ n401 ;
  assign n12657 = n5365 | n12656 ;
  assign n12658 = n10860 ^ n8249 ^ n4105 ;
  assign n12659 = n12658 ^ n3475 ^ 1'b0 ;
  assign n12660 = n12657 & n12659 ;
  assign n12661 = n10708 ^ n1713 ^ n1493 ;
  assign n12662 = n2424 ^ n1849 ^ 1'b0 ;
  assign n12663 = ( n197 & n920 ) | ( n197 & n6690 ) | ( n920 & n6690 ) ;
  assign n12664 = n11599 & n12663 ;
  assign n12665 = ~n1798 & n12664 ;
  assign n12666 = n6021 & ~n12665 ;
  assign n12667 = n12666 ^ n3451 ^ 1'b0 ;
  assign n12668 = n12662 & n12667 ;
  assign n12669 = n7448 ^ n7067 ^ 1'b0 ;
  assign n12670 = ~n396 & n12669 ;
  assign n12671 = ~n1555 & n10631 ;
  assign n12672 = n12670 & n12671 ;
  assign n12673 = n739 & n5971 ;
  assign n12674 = n3643 & n9312 ;
  assign n12675 = ( n6466 & n11844 ) | ( n6466 & ~n12674 ) | ( n11844 & ~n12674 ) ;
  assign n12676 = ( ~n589 & n8697 ) | ( ~n589 & n12675 ) | ( n8697 & n12675 ) ;
  assign n12677 = ( n964 & ~n1540 ) | ( n964 & n2020 ) | ( ~n1540 & n2020 ) ;
  assign n12678 = n12677 ^ n12674 ^ n8478 ;
  assign n12679 = n7163 & n9467 ;
  assign n12680 = n9473 ^ n5699 ^ 1'b0 ;
  assign n12681 = ( n3511 & n12679 ) | ( n3511 & n12680 ) | ( n12679 & n12680 ) ;
  assign n12682 = n378 & ~n3352 ;
  assign n12683 = n12682 ^ n5023 ^ 1'b0 ;
  assign n12684 = ( n5535 & n11098 ) | ( n5535 & ~n12683 ) | ( n11098 & ~n12683 ) ;
  assign n12685 = n8662 & n12684 ;
  assign n12686 = n1484 & n12685 ;
  assign n12687 = ~n3077 & n12686 ;
  assign n12688 = n12687 ^ n8351 ^ 1'b0 ;
  assign n12689 = n3925 & ~n7022 ;
  assign n12690 = x72 & ~n1814 ;
  assign n12691 = ( n800 & n11957 ) | ( n800 & n12690 ) | ( n11957 & n12690 ) ;
  assign n12692 = n12691 ^ n4834 ^ 1'b0 ;
  assign n12693 = n3723 & ~n12692 ;
  assign n12694 = n12693 ^ n5566 ^ 1'b0 ;
  assign n12695 = n7216 & ~n11034 ;
  assign n12697 = n4728 ^ n3778 ^ 1'b0 ;
  assign n12698 = n10642 | n12697 ;
  assign n12699 = n12698 ^ n9053 ^ n2738 ;
  assign n12700 = n1471 & ~n12699 ;
  assign n12696 = n2901 & n10060 ;
  assign n12701 = n12700 ^ n12696 ^ 1'b0 ;
  assign n12702 = n12701 ^ n5437 ^ n1697 ;
  assign n12703 = n6421 ^ n3099 ^ 1'b0 ;
  assign n12704 = n3573 & n12703 ;
  assign n12705 = n12704 ^ n6815 ^ 1'b0 ;
  assign n12706 = ~n6860 & n10180 ;
  assign n12707 = ( n1420 & ~n5051 ) | ( n1420 & n9958 ) | ( ~n5051 & n9958 ) ;
  assign n12708 = n12707 ^ n12075 ^ 1'b0 ;
  assign n12709 = n9429 | n12708 ;
  assign n12710 = ( ~n3255 & n5254 ) | ( ~n3255 & n9001 ) | ( n5254 & n9001 ) ;
  assign n12711 = n809 & ~n12710 ;
  assign n12712 = n1542 & ~n3671 ;
  assign n12713 = ( n2119 & n4169 ) | ( n2119 & ~n9136 ) | ( n4169 & ~n9136 ) ;
  assign n12714 = n12713 ^ n6144 ^ 1'b0 ;
  assign n12715 = n3587 | n12714 ;
  assign n12716 = ( n3732 & n6769 ) | ( n3732 & n9859 ) | ( n6769 & n9859 ) ;
  assign n12717 = n12716 ^ n5520 ^ n1505 ;
  assign n12718 = ~n12715 & n12717 ;
  assign n12719 = n980 ^ n147 ^ 1'b0 ;
  assign n12720 = n12719 ^ n4705 ^ 1'b0 ;
  assign n12721 = ~n5616 & n12720 ;
  assign n12722 = ( ~n1711 & n4062 ) | ( ~n1711 & n12721 ) | ( n4062 & n12721 ) ;
  assign n12723 = n12722 ^ n12384 ^ 1'b0 ;
  assign n12724 = n5614 ^ n2269 ^ 1'b0 ;
  assign n12725 = n779 & ~n5699 ;
  assign n12726 = n12725 ^ n7822 ^ 1'b0 ;
  assign n12727 = ( n5058 & ~n12500 ) | ( n5058 & n12726 ) | ( ~n12500 & n12726 ) ;
  assign n12728 = ~n1499 & n12727 ;
  assign n12729 = ~n1071 & n6294 ;
  assign n12730 = ~n6555 & n12729 ;
  assign n12731 = n12730 ^ n8253 ^ 1'b0 ;
  assign n12732 = n8073 ^ n3440 ^ 1'b0 ;
  assign n12733 = n12731 & ~n12732 ;
  assign n12734 = n2443 & ~n9845 ;
  assign n12735 = ( n4334 & n10619 ) | ( n4334 & n10887 ) | ( n10619 & n10887 ) ;
  assign n12736 = n12734 & ~n12735 ;
  assign n12737 = n12736 ^ x29 ^ 1'b0 ;
  assign n12738 = x67 & n12737 ;
  assign n12739 = n5208 | n12037 ;
  assign n12740 = n12363 ^ n5050 ^ 1'b0 ;
  assign n12741 = n12739 & ~n12740 ;
  assign n12742 = n2896 | n10915 ;
  assign n12743 = n4505 ^ n1107 ^ 1'b0 ;
  assign n12744 = ~n9670 & n12743 ;
  assign n12747 = n8554 ^ n599 ^ 1'b0 ;
  assign n12745 = ( n2565 & ~n2724 ) | ( n2565 & n7157 ) | ( ~n2724 & n7157 ) ;
  assign n12746 = n2115 | n12745 ;
  assign n12748 = n12747 ^ n12746 ^ n468 ;
  assign n12749 = n796 | n1685 ;
  assign n12750 = n12749 ^ n8919 ^ 1'b0 ;
  assign n12751 = n5940 ^ n4666 ^ 1'b0 ;
  assign n12752 = ~n10103 & n12751 ;
  assign n12753 = n12752 ^ n6824 ^ n529 ;
  assign n12754 = n4139 | n9562 ;
  assign n12755 = n4699 | n12754 ;
  assign n12756 = n6189 ^ n3030 ^ 1'b0 ;
  assign n12758 = n9226 ^ n5888 ^ n4535 ;
  assign n12757 = n3347 & n5300 ;
  assign n12759 = n12758 ^ n12757 ^ 1'b0 ;
  assign n12760 = ( n10398 & ~n12756 ) | ( n10398 & n12759 ) | ( ~n12756 & n12759 ) ;
  assign n12761 = n11053 ^ n1810 ^ 1'b0 ;
  assign n12762 = n11736 ^ n5634 ^ n846 ;
  assign n12763 = ( ~n10481 & n12761 ) | ( ~n10481 & n12762 ) | ( n12761 & n12762 ) ;
  assign n12764 = ( ~n2083 & n8100 ) | ( ~n2083 & n12763 ) | ( n8100 & n12763 ) ;
  assign n12765 = n12764 ^ n4408 ^ n1758 ;
  assign n12766 = n5249 & n11054 ;
  assign n12767 = n12766 ^ n5257 ^ 1'b0 ;
  assign n12768 = ( ~n3406 & n5597 ) | ( ~n3406 & n11789 ) | ( n5597 & n11789 ) ;
  assign n12769 = ~n5663 & n12768 ;
  assign n12770 = n7968 & n12769 ;
  assign n12771 = n5030 ^ n1617 ^ 1'b0 ;
  assign n12772 = n11392 & ~n12771 ;
  assign n12773 = n10609 ^ n3074 ^ 1'b0 ;
  assign n12774 = n3340 | n12773 ;
  assign n12775 = n4700 ^ n4408 ^ 1'b0 ;
  assign n12776 = ~n12774 & n12775 ;
  assign n12778 = n9634 ^ n4240 ^ n755 ;
  assign n12777 = ~n2869 & n9151 ;
  assign n12779 = n12778 ^ n12777 ^ 1'b0 ;
  assign n12780 = n12779 ^ n11213 ^ n1035 ;
  assign n12781 = ~n4464 & n7054 ;
  assign n12782 = n12781 ^ n1437 ^ 1'b0 ;
  assign n12783 = n1034 & ~n12782 ;
  assign n12784 = n3335 & n12783 ;
  assign n12785 = n12784 ^ n1075 ^ 1'b0 ;
  assign n12786 = ~n5127 & n12785 ;
  assign n12787 = n7785 ^ n7122 ^ 1'b0 ;
  assign n12788 = n6529 & ~n12787 ;
  assign n12793 = n9698 ^ n7963 ^ 1'b0 ;
  assign n12792 = n5351 ^ n2938 ^ 1'b0 ;
  assign n12794 = n12793 ^ n12792 ^ 1'b0 ;
  assign n12795 = n375 & n12794 ;
  assign n12789 = n5281 ^ n2974 ^ 1'b0 ;
  assign n12790 = ~n3513 & n12789 ;
  assign n12791 = ~n3806 & n12790 ;
  assign n12796 = n12795 ^ n12791 ^ 1'b0 ;
  assign n12797 = n8121 ^ n2413 ^ 1'b0 ;
  assign n12798 = n7293 & n12797 ;
  assign n12799 = ~n612 & n12798 ;
  assign n12800 = n3840 & ~n8685 ;
  assign n12801 = n12800 ^ n6823 ^ n4641 ;
  assign n12802 = n11730 ^ n5397 ^ x74 ;
  assign n12803 = ~n4166 & n12802 ;
  assign n12804 = n12803 ^ n10506 ^ n8058 ;
  assign n12805 = ~n5176 & n7108 ;
  assign n12806 = n12805 ^ n4389 ^ 1'b0 ;
  assign n12807 = n12806 ^ n5075 ^ 1'b0 ;
  assign n12808 = ~n12147 & n12807 ;
  assign n12809 = n12808 ^ n5768 ^ 1'b0 ;
  assign n12810 = ( n158 & n7496 ) | ( n158 & ~n12809 ) | ( n7496 & ~n12809 ) ;
  assign n12811 = ~n6781 & n8350 ;
  assign n12812 = n12811 ^ n9174 ^ n5248 ;
  assign n12813 = n5687 | n12812 ;
  assign n12814 = n9675 ^ n8615 ^ 1'b0 ;
  assign n12815 = ~n8220 & n12814 ;
  assign n12816 = n5679 ^ n2197 ^ 1'b0 ;
  assign n12817 = n6773 | n9097 ;
  assign n12824 = n5311 | n8163 ;
  assign n12825 = n5440 | n12824 ;
  assign n12820 = ( ~n537 & n952 ) | ( ~n537 & n5437 ) | ( n952 & n5437 ) ;
  assign n12821 = n12820 ^ n8464 ^ x112 ;
  assign n12822 = ( n4946 & n6393 ) | ( n4946 & n12821 ) | ( n6393 & n12821 ) ;
  assign n12818 = n3999 ^ n3965 ^ n329 ;
  assign n12819 = n2077 & n12818 ;
  assign n12823 = n12822 ^ n12819 ^ 1'b0 ;
  assign n12826 = n12825 ^ n12823 ^ n5014 ;
  assign n12828 = ( ~n1172 & n3602 ) | ( ~n1172 & n4584 ) | ( n3602 & n4584 ) ;
  assign n12829 = n12828 ^ n6772 ^ n6089 ;
  assign n12827 = n12083 ^ n6219 ^ n5385 ;
  assign n12830 = n12829 ^ n12827 ^ n9887 ;
  assign n12831 = n1986 & ~n4823 ;
  assign n12832 = n5946 | n12831 ;
  assign n12833 = n6475 & n10234 ;
  assign n12834 = ~n12832 & n12833 ;
  assign n12835 = n3410 ^ n786 ^ 1'b0 ;
  assign n12836 = ~n565 & n12835 ;
  assign n12837 = ( n4380 & n9508 ) | ( n4380 & n12836 ) | ( n9508 & n12836 ) ;
  assign n12838 = n8461 & ~n11783 ;
  assign n12839 = n12838 ^ n4936 ^ 1'b0 ;
  assign n12840 = ( n1205 & n1609 ) | ( n1205 & ~n2442 ) | ( n1609 & ~n2442 ) ;
  assign n12841 = n6262 ^ n3974 ^ 1'b0 ;
  assign n12842 = n1048 | n12841 ;
  assign n12843 = n3670 | n12842 ;
  assign n12844 = n4479 | n12843 ;
  assign n12845 = n12844 ^ n2616 ^ n525 ;
  assign n12846 = n12628 ^ n2938 ^ n2883 ;
  assign n12847 = n4221 ^ n3999 ^ n304 ;
  assign n12848 = ~n338 & n1108 ;
  assign n12849 = n2811 & n4144 ;
  assign n12850 = n4982 | n6357 ;
  assign n12851 = n12849 | n12850 ;
  assign n12852 = ~n8753 & n12851 ;
  assign n12853 = n12722 ^ n4132 ^ n321 ;
  assign n12854 = n12853 ^ n12641 ^ 1'b0 ;
  assign n12855 = n9867 ^ n3218 ^ n1138 ;
  assign n12856 = n11955 ^ n3964 ^ 1'b0 ;
  assign n12857 = n12855 | n12856 ;
  assign n12858 = n2949 ^ n2168 ^ n1559 ;
  assign n12859 = ( n3204 & ~n12857 ) | ( n3204 & n12858 ) | ( ~n12857 & n12858 ) ;
  assign n12861 = ~n6479 & n6672 ;
  assign n12860 = ~n4996 & n8536 ;
  assign n12862 = n12861 ^ n12860 ^ n11649 ;
  assign n12863 = n7980 ^ n2936 ^ 1'b0 ;
  assign n12864 = n1571 & ~n3703 ;
  assign n12865 = n10581 & ~n12864 ;
  assign n12866 = ( n7432 & ~n10764 ) | ( n7432 & n11872 ) | ( ~n10764 & n11872 ) ;
  assign n12867 = n5468 ^ n3533 ^ n1686 ;
  assign n12868 = n4165 & n12867 ;
  assign n12869 = ~n8170 & n12868 ;
  assign n12870 = n3244 | n12869 ;
  assign n12871 = n12870 ^ n3507 ^ 1'b0 ;
  assign n12872 = n4449 & n6760 ;
  assign n12873 = ~n2712 & n12872 ;
  assign n12877 = n1673 & n4491 ;
  assign n12878 = ~n1647 & n12877 ;
  assign n12874 = ( n1199 & ~n3682 ) | ( n1199 & n3984 ) | ( ~n3682 & n3984 ) ;
  assign n12875 = n12426 ^ n5588 ^ 1'b0 ;
  assign n12876 = n12874 & n12875 ;
  assign n12879 = n12878 ^ n12876 ^ 1'b0 ;
  assign n12880 = n8832 & n12879 ;
  assign n12881 = n9158 ^ n6434 ^ 1'b0 ;
  assign n12882 = n831 & ~n12881 ;
  assign n12883 = n7746 ^ n6586 ^ n1354 ;
  assign n12884 = n12883 ^ n8575 ^ n637 ;
  assign n12885 = ( n7853 & n12841 ) | ( n7853 & n12884 ) | ( n12841 & n12884 ) ;
  assign n12890 = ( n693 & n8555 ) | ( n693 & ~n9817 ) | ( n8555 & ~n9817 ) ;
  assign n12888 = n3209 ^ n2401 ^ 1'b0 ;
  assign n12889 = ~n5564 & n12888 ;
  assign n12886 = n3804 & ~n8256 ;
  assign n12887 = n12886 ^ n2856 ^ 1'b0 ;
  assign n12891 = n12890 ^ n12889 ^ n12887 ;
  assign n12892 = ( n982 & n1683 ) | ( n982 & ~n7697 ) | ( n1683 & ~n7697 ) ;
  assign n12893 = n12892 ^ n10329 ^ 1'b0 ;
  assign n12894 = ~n10272 & n12893 ;
  assign n12895 = n2093 & ~n2244 ;
  assign n12896 = n12895 ^ n9100 ^ n740 ;
  assign n12898 = ~n4097 & n6202 ;
  assign n12899 = n7404 & n12898 ;
  assign n12897 = n4858 & n12081 ;
  assign n12900 = n12899 ^ n12897 ^ 1'b0 ;
  assign n12901 = ~n12896 & n12900 ;
  assign n12902 = n11393 ^ n10716 ^ n4651 ;
  assign n12903 = ( n214 & n320 ) | ( n214 & ~n516 ) | ( n320 & ~n516 ) ;
  assign n12904 = n3812 | n12903 ;
  assign n12905 = n5903 | n12904 ;
  assign n12906 = ~n732 & n12905 ;
  assign n12907 = n6891 & n12906 ;
  assign n12908 = ( n5067 & n8916 ) | ( n5067 & ~n12907 ) | ( n8916 & ~n12907 ) ;
  assign n12909 = n2388 & ~n3990 ;
  assign n12910 = ~n4260 & n12909 ;
  assign n12911 = ( n5453 & n7612 ) | ( n5453 & n12910 ) | ( n7612 & n12910 ) ;
  assign n12912 = ~n8590 & n12911 ;
  assign n12913 = n1271 & n6413 ;
  assign n12914 = n5913 | n12913 ;
  assign n12915 = n12912 | n12914 ;
  assign n12916 = n11671 ^ n8471 ^ n6851 ;
  assign n12917 = n6371 | n11308 ;
  assign n12918 = n12916 | n12917 ;
  assign n12919 = n7318 ^ n5319 ^ n3475 ;
  assign n12920 = n4133 | n12919 ;
  assign n12921 = ~n2072 & n10401 ;
  assign n12922 = n3376 & ~n3447 ;
  assign n12923 = ~n11028 & n12922 ;
  assign n12924 = ( ~n1955 & n5176 ) | ( ~n1955 & n12923 ) | ( n5176 & n12923 ) ;
  assign n12925 = n4087 | n12924 ;
  assign n12926 = n4822 & ~n12925 ;
  assign n12927 = n12926 ^ n4351 ^ n998 ;
  assign n12929 = n7682 ^ n6125 ^ n991 ;
  assign n12928 = n3235 ^ n306 ^ 1'b0 ;
  assign n12930 = n12929 ^ n12928 ^ n9470 ;
  assign n12935 = n2343 & n5308 ;
  assign n12936 = n331 & n12935 ;
  assign n12931 = ~n2642 & n9350 ;
  assign n12932 = n12931 ^ n1547 ^ 1'b0 ;
  assign n12933 = ~n8137 & n12932 ;
  assign n12934 = ~n1437 & n12933 ;
  assign n12937 = n12936 ^ n12934 ^ n9170 ;
  assign n12938 = n2547 & ~n7865 ;
  assign n12939 = n12938 ^ n1218 ^ 1'b0 ;
  assign n12940 = n12939 ^ n1745 ^ 1'b0 ;
  assign n12941 = n4233 & n4296 ;
  assign n12942 = n12941 ^ x55 ^ 1'b0 ;
  assign n12943 = n3572 | n9113 ;
  assign n12944 = x38 & n3597 ;
  assign n12945 = n12944 ^ n894 ^ 1'b0 ;
  assign n12946 = ~n409 & n4595 ;
  assign n12947 = n12195 ^ n307 ^ 1'b0 ;
  assign n12948 = n12946 | n12947 ;
  assign n12949 = ( n11541 & ~n12945 ) | ( n11541 & n12948 ) | ( ~n12945 & n12948 ) ;
  assign n12950 = n12949 ^ n7955 ^ 1'b0 ;
  assign n12951 = n858 | n11044 ;
  assign n12952 = ( ~n535 & n10057 ) | ( ~n535 & n11215 ) | ( n10057 & n11215 ) ;
  assign n12953 = ~n2615 & n6972 ;
  assign n12954 = n12953 ^ n11869 ^ 1'b0 ;
  assign n12955 = n12954 ^ n1894 ^ 1'b0 ;
  assign n12956 = n12952 & n12955 ;
  assign n12957 = ( ~n2219 & n2294 ) | ( ~n2219 & n7597 ) | ( n2294 & n7597 ) ;
  assign n12958 = n7742 ^ n6705 ^ 1'b0 ;
  assign n12959 = n12958 ^ n164 ^ 1'b0 ;
  assign n12960 = n4262 | n6273 ;
  assign n12961 = n5395 & ~n12960 ;
  assign n12962 = n12961 ^ n2767 ^ 1'b0 ;
  assign n12963 = ( n1811 & ~n2720 ) | ( n1811 & n3194 ) | ( ~n2720 & n3194 ) ;
  assign n12964 = n7951 & n12963 ;
  assign n12965 = n12964 ^ n774 ^ 1'b0 ;
  assign n12966 = ( n1562 & ~n10830 ) | ( n1562 & n12965 ) | ( ~n10830 & n12965 ) ;
  assign n12967 = n5864 & n12966 ;
  assign n12968 = ~n707 & n12967 ;
  assign n12969 = n1467 | n7314 ;
  assign n12970 = n12969 ^ n522 ^ 1'b0 ;
  assign n12971 = ( n8417 & n12968 ) | ( n8417 & ~n12970 ) | ( n12968 & ~n12970 ) ;
  assign n12972 = n12971 ^ n10489 ^ 1'b0 ;
  assign n12973 = n4106 & n4459 ;
  assign n12974 = n12973 ^ n11215 ^ n3167 ;
  assign n12975 = n12812 ^ n2386 ^ n275 ;
  assign n12976 = ~n1076 & n12975 ;
  assign n12977 = ~n12974 & n12976 ;
  assign n12978 = ( n1384 & n1864 ) | ( n1384 & n3658 ) | ( n1864 & n3658 ) ;
  assign n12979 = n12978 ^ n5395 ^ n4936 ;
  assign n12980 = n12979 ^ n6989 ^ n3505 ;
  assign n12981 = ~n1419 & n12721 ;
  assign n12982 = ~n1189 & n12981 ;
  assign n12983 = n5570 ^ n5159 ^ 1'b0 ;
  assign n12984 = n12983 ^ n4363 ^ 1'b0 ;
  assign n12985 = n8600 & n12984 ;
  assign n12986 = ( n6409 & n12982 ) | ( n6409 & ~n12985 ) | ( n12982 & ~n12985 ) ;
  assign n12987 = n1811 & ~n3613 ;
  assign n12988 = n5021 & n12987 ;
  assign n12989 = n2901 & ~n3054 ;
  assign n12992 = ( n1182 & n3870 ) | ( n1182 & ~n6889 ) | ( n3870 & ~n6889 ) ;
  assign n12990 = ( n758 & n1918 ) | ( n758 & n7673 ) | ( n1918 & n7673 ) ;
  assign n12991 = ( n1385 & n3432 ) | ( n1385 & n12990 ) | ( n3432 & n12990 ) ;
  assign n12993 = n12992 ^ n12991 ^ n11714 ;
  assign n12994 = n3054 & ~n3137 ;
  assign n12996 = ( n5407 & n7062 ) | ( n5407 & n10637 ) | ( n7062 & n10637 ) ;
  assign n12995 = n6216 ^ n5962 ^ n5390 ;
  assign n12997 = n12996 ^ n12995 ^ 1'b0 ;
  assign n12998 = ( n6147 & n8619 ) | ( n6147 & n11812 ) | ( n8619 & n11812 ) ;
  assign n12999 = n11936 ^ n10020 ^ n4259 ;
  assign n13004 = n10137 ^ n7346 ^ 1'b0 ;
  assign n13005 = n3084 & ~n13004 ;
  assign n13000 = ~n3500 & n3925 ;
  assign n13001 = n3247 & n13000 ;
  assign n13002 = n13001 ^ n11747 ^ n8528 ;
  assign n13003 = n13002 ^ n12572 ^ n6422 ;
  assign n13006 = n13005 ^ n13003 ^ 1'b0 ;
  assign n13007 = n10817 & n13006 ;
  assign n13008 = n9309 ^ n7064 ^ x111 ;
  assign n13009 = n5281 ^ n2561 ^ n1124 ;
  assign n13010 = n7952 ^ n1925 ^ 1'b0 ;
  assign n13011 = n6700 & ~n13010 ;
  assign n13012 = n7905 ^ n4681 ^ 1'b0 ;
  assign n13013 = ( n6016 & n8603 ) | ( n6016 & n13012 ) | ( n8603 & n13012 ) ;
  assign n13014 = n10980 ^ n9100 ^ n6547 ;
  assign n13015 = n12853 ^ n6403 ^ n2578 ;
  assign n13016 = ~n1682 & n4441 ;
  assign n13017 = n2077 ^ n1679 ^ n1366 ;
  assign n13018 = n13017 ^ n7954 ^ n3360 ;
  assign n13019 = n1171 & ~n4558 ;
  assign n13020 = n13019 ^ n10093 ^ 1'b0 ;
  assign n13021 = n968 | n13020 ;
  assign n13022 = n9303 ^ n2480 ^ n658 ;
  assign n13023 = ( ~n3390 & n13021 ) | ( ~n3390 & n13022 ) | ( n13021 & n13022 ) ;
  assign n13024 = n194 & n1592 ;
  assign n13025 = n13024 ^ n1709 ^ 1'b0 ;
  assign n13026 = n13025 ^ n4705 ^ n949 ;
  assign n13027 = n7378 | n9567 ;
  assign n13028 = n6930 | n13027 ;
  assign n13029 = ( n954 & n1484 ) | ( n954 & ~n4278 ) | ( n1484 & ~n4278 ) ;
  assign n13030 = n13029 ^ n9252 ^ 1'b0 ;
  assign n13031 = ( n2277 & n8913 ) | ( n2277 & n10218 ) | ( n8913 & n10218 ) ;
  assign n13032 = n11738 ^ n9928 ^ 1'b0 ;
  assign n13033 = n2181 | n10019 ;
  assign n13034 = n13033 ^ n8191 ^ x113 ;
  assign n13035 = ( ~n3774 & n10322 ) | ( ~n3774 & n13034 ) | ( n10322 & n13034 ) ;
  assign n13036 = n2820 & n9161 ;
  assign n13037 = n6892 & ~n10030 ;
  assign n13038 = n13037 ^ n1961 ^ 1'b0 ;
  assign n13039 = n5267 | n13038 ;
  assign n13040 = n8129 & ~n13039 ;
  assign n13041 = ~n3554 & n6378 ;
  assign n13042 = n3287 & n13041 ;
  assign n13043 = ( n1425 & n3321 ) | ( n1425 & n11178 ) | ( n3321 & n11178 ) ;
  assign n13044 = n13043 ^ n8952 ^ 1'b0 ;
  assign n13045 = ~n9984 & n13044 ;
  assign n13046 = n13045 ^ n9603 ^ n2296 ;
  assign n13050 = n9053 ^ n431 ^ 1'b0 ;
  assign n13051 = n2830 | n13050 ;
  assign n13047 = n4344 ^ n3986 ^ 1'b0 ;
  assign n13048 = n13047 ^ n5749 ^ 1'b0 ;
  assign n13049 = n222 & n13048 ;
  assign n13052 = n13051 ^ n13049 ^ n6908 ;
  assign n13053 = ( n3706 & n4290 ) | ( n3706 & n8018 ) | ( n4290 & n8018 ) ;
  assign n13054 = ~n1073 & n7712 ;
  assign n13055 = n13053 & n13054 ;
  assign n13056 = n3161 | n13055 ;
  assign n13057 = n13056 ^ n8023 ^ 1'b0 ;
  assign n13064 = n2541 & ~n12140 ;
  assign n13065 = n4561 & n13064 ;
  assign n13061 = n2763 ^ n968 ^ 1'b0 ;
  assign n13059 = n1646 ^ n1484 ^ 1'b0 ;
  assign n13060 = n12572 & ~n13059 ;
  assign n13058 = n5024 & n8572 ;
  assign n13062 = n13061 ^ n13060 ^ n13058 ;
  assign n13063 = n1929 & ~n13062 ;
  assign n13066 = n13065 ^ n13063 ^ n10000 ;
  assign n13069 = n11215 ^ n3114 ^ 1'b0 ;
  assign n13067 = n8872 ^ n1586 ^ 1'b0 ;
  assign n13068 = n2878 & n13067 ;
  assign n13070 = n13069 ^ n13068 ^ 1'b0 ;
  assign n13071 = n13070 ^ n7864 ^ 1'b0 ;
  assign n13072 = n1036 | n9038 ;
  assign n13073 = n13072 ^ n838 ^ 1'b0 ;
  assign n13074 = ( n1113 & n2980 ) | ( n1113 & ~n13073 ) | ( n2980 & ~n13073 ) ;
  assign n13075 = n6656 ^ n1389 ^ 1'b0 ;
  assign n13076 = ~n13074 & n13075 ;
  assign n13077 = n6057 ^ n987 ^ 1'b0 ;
  assign n13078 = ~n3249 & n13077 ;
  assign n13079 = n2095 ^ n889 ^ 1'b0 ;
  assign n13080 = n5687 & ~n13079 ;
  assign n13081 = n13080 ^ n2053 ^ 1'b0 ;
  assign n13082 = n13081 ^ n6510 ^ 1'b0 ;
  assign n13083 = ( n2502 & n5632 ) | ( n2502 & ~n7339 ) | ( n5632 & ~n7339 ) ;
  assign n13084 = n13083 ^ n6398 ^ n4481 ;
  assign n13085 = n5729 & n11448 ;
  assign n13086 = n13085 ^ n11918 ^ 1'b0 ;
  assign n13088 = n10803 ^ n3815 ^ n527 ;
  assign n13089 = n13088 ^ n4878 ^ 1'b0 ;
  assign n13090 = n6877 | n13089 ;
  assign n13087 = n4335 & n7890 ;
  assign n13091 = n13090 ^ n13087 ^ 1'b0 ;
  assign n13095 = n7913 & n9000 ;
  assign n13092 = n2187 | n9660 ;
  assign n13093 = n1399 & ~n13092 ;
  assign n13094 = n2167 | n13093 ;
  assign n13096 = n13095 ^ n13094 ^ 1'b0 ;
  assign n13097 = ( ~n4660 & n13091 ) | ( ~n4660 & n13096 ) | ( n13091 & n13096 ) ;
  assign n13098 = n7998 | n10258 ;
  assign n13099 = n2371 & ~n13098 ;
  assign n13100 = ( n2071 & n10527 ) | ( n2071 & ~n12572 ) | ( n10527 & ~n12572 ) ;
  assign n13101 = n13100 ^ n8563 ^ n5410 ;
  assign n13102 = ~n13099 & n13101 ;
  assign n13103 = ~n5314 & n6768 ;
  assign n13104 = ~n7459 & n13103 ;
  assign n13105 = n13104 ^ n3583 ^ 1'b0 ;
  assign n13106 = ~n4459 & n11605 ;
  assign n13107 = n8796 ^ n5133 ^ 1'b0 ;
  assign n13108 = n13106 & ~n13107 ;
  assign n13109 = ( n5122 & ~n5891 ) | ( n5122 & n6402 ) | ( ~n5891 & n6402 ) ;
  assign n13110 = n6701 ^ n5062 ^ n4521 ;
  assign n13111 = ~n1272 & n12595 ;
  assign n13112 = ~n5844 & n13111 ;
  assign n13113 = n13112 ^ n1381 ^ 1'b0 ;
  assign n13114 = n10300 & ~n13113 ;
  assign n13115 = ( n13109 & n13110 ) | ( n13109 & n13114 ) | ( n13110 & n13114 ) ;
  assign n13116 = ~n369 & n1382 ;
  assign n13117 = n13116 ^ n9860 ^ 1'b0 ;
  assign n13119 = n2429 ^ n673 ^ 1'b0 ;
  assign n13118 = n8058 ^ n363 ^ n132 ;
  assign n13120 = n13119 ^ n13118 ^ n10982 ;
  assign n13121 = ( n5186 & ~n13117 ) | ( n5186 & n13120 ) | ( ~n13117 & n13120 ) ;
  assign n13122 = n7108 & n10730 ;
  assign n13125 = n3365 ^ n2170 ^ 1'b0 ;
  assign n13123 = n5979 ^ n1013 ^ 1'b0 ;
  assign n13124 = n13123 ^ n10593 ^ 1'b0 ;
  assign n13126 = n13125 ^ n13124 ^ 1'b0 ;
  assign n13127 = n2009 ^ n1308 ^ 1'b0 ;
  assign n13128 = n13127 ^ x113 ^ 1'b0 ;
  assign n13129 = ~n13126 & n13128 ;
  assign n13130 = ( n612 & n1221 ) | ( n612 & ~n3994 ) | ( n1221 & ~n3994 ) ;
  assign n13131 = ~n2048 & n7974 ;
  assign n13132 = n13130 & n13131 ;
  assign n13148 = ~n4772 & n5678 ;
  assign n13149 = n8141 & n13148 ;
  assign n13150 = n6830 & ~n13149 ;
  assign n13133 = n5304 | n7022 ;
  assign n13134 = ( n834 & n1246 ) | ( n834 & n13133 ) | ( n1246 & n13133 ) ;
  assign n13139 = n5263 & n6263 ;
  assign n13140 = n13139 ^ n6178 ^ 1'b0 ;
  assign n13141 = n13140 ^ n2738 ^ 1'b0 ;
  assign n13142 = n6222 | n13141 ;
  assign n13143 = n4455 & n13142 ;
  assign n13144 = n13143 ^ n4521 ^ 1'b0 ;
  assign n13138 = ~n3416 & n9664 ;
  assign n13137 = n3188 & ~n3858 ;
  assign n13145 = n13144 ^ n13138 ^ n13137 ;
  assign n13135 = n8837 ^ n2106 ^ 1'b0 ;
  assign n13136 = ~n977 & n13135 ;
  assign n13146 = n13145 ^ n13136 ^ 1'b0 ;
  assign n13147 = ( n12499 & n13134 ) | ( n12499 & ~n13146 ) | ( n13134 & ~n13146 ) ;
  assign n13151 = n13150 ^ n13147 ^ 1'b0 ;
  assign n13152 = n6586 ^ n1100 ^ 1'b0 ;
  assign n13153 = n10993 & n13152 ;
  assign n13154 = ~n9804 & n13153 ;
  assign n13155 = n9524 ^ n2561 ^ 1'b0 ;
  assign n13156 = ~n13154 & n13155 ;
  assign n13157 = n6022 ^ n4974 ^ 1'b0 ;
  assign n13159 = n6366 ^ n1458 ^ n255 ;
  assign n13158 = n4925 ^ n2831 ^ 1'b0 ;
  assign n13160 = n13159 ^ n13158 ^ n5641 ;
  assign n13161 = n6260 & ~n10056 ;
  assign n13162 = ~n13160 & n13161 ;
  assign n13163 = n617 & ~n13162 ;
  assign n13164 = n13163 ^ n5984 ^ 1'b0 ;
  assign n13165 = n5821 & n13100 ;
  assign n13166 = n13165 ^ n8306 ^ n3953 ;
  assign n13167 = n4269 & ~n13166 ;
  assign n13168 = n1007 | n1481 ;
  assign n13169 = ~n1578 & n12524 ;
  assign n13170 = ~n13168 & n13169 ;
  assign n13171 = n4765 ^ n3629 ^ 1'b0 ;
  assign n13172 = ~n4195 & n13171 ;
  assign n13173 = ( ~n3754 & n13170 ) | ( ~n3754 & n13172 ) | ( n13170 & n13172 ) ;
  assign n13174 = ( ~n1714 & n2963 ) | ( ~n1714 & n9093 ) | ( n2963 & n9093 ) ;
  assign n13175 = n3628 & ~n6704 ;
  assign n13176 = n13175 ^ n994 ^ 1'b0 ;
  assign n13177 = ( n572 & n6217 ) | ( n572 & n13176 ) | ( n6217 & n13176 ) ;
  assign n13178 = n13177 ^ n4236 ^ n734 ;
  assign n13179 = n9901 ^ n7845 ^ 1'b0 ;
  assign n13180 = n13178 & ~n13179 ;
  assign n13181 = ~n5206 & n6364 ;
  assign n13182 = n13181 ^ n10863 ^ 1'b0 ;
  assign n13183 = n9948 | n13182 ;
  assign n13184 = n13183 ^ n10993 ^ 1'b0 ;
  assign n13185 = n8364 | n13184 ;
  assign n13186 = n10212 ^ n3964 ^ 1'b0 ;
  assign n13187 = n9687 ^ n1288 ^ 1'b0 ;
  assign n13188 = n13187 ^ n11616 ^ n2220 ;
  assign n13189 = n13186 | n13188 ;
  assign n13190 = ( x51 & ~n176 ) | ( x51 & n8490 ) | ( ~n176 & n8490 ) ;
  assign n13191 = n12889 ^ n5367 ^ n4290 ;
  assign n13192 = n13190 & n13191 ;
  assign n13193 = ~n4167 & n13192 ;
  assign n13194 = n13193 ^ n2951 ^ n1209 ;
  assign n13195 = ~n4990 & n13194 ;
  assign n13196 = n4563 & n13195 ;
  assign n13197 = n13196 ^ n8457 ^ 1'b0 ;
  assign n13198 = n12184 & ~n13197 ;
  assign n13199 = ( ~x100 & n4150 ) | ( ~x100 & n13198 ) | ( n4150 & n13198 ) ;
  assign n13200 = n3271 ^ n370 ^ 1'b0 ;
  assign n13201 = n2944 | n13200 ;
  assign n13202 = n13201 ^ n5630 ^ n1451 ;
  assign n13203 = n4512 ^ n2202 ^ 1'b0 ;
  assign n13204 = n12650 & n13203 ;
  assign n13205 = n13204 ^ n574 ^ 1'b0 ;
  assign n13206 = ~n13202 & n13205 ;
  assign n13207 = n13206 ^ n11642 ^ 1'b0 ;
  assign n13208 = ( ~n5403 & n5899 ) | ( ~n5403 & n10831 ) | ( n5899 & n10831 ) ;
  assign n13209 = n4955 | n10238 ;
  assign n13210 = n13209 ^ n2360 ^ 1'b0 ;
  assign n13211 = x57 & n13210 ;
  assign n13212 = ( ~n8653 & n13208 ) | ( ~n8653 & n13211 ) | ( n13208 & n13211 ) ;
  assign n13213 = n13212 ^ n2095 ^ 1'b0 ;
  assign n13215 = n454 | n940 ;
  assign n13216 = n4222 | n13215 ;
  assign n13214 = n7034 | n12372 ;
  assign n13217 = n13216 ^ n13214 ^ n5376 ;
  assign n13218 = n13217 ^ n7512 ^ n356 ;
  assign n13219 = ( n1605 & n3415 ) | ( n1605 & ~n12499 ) | ( n3415 & ~n12499 ) ;
  assign n13220 = n13219 ^ n4718 ^ 1'b0 ;
  assign n13221 = n4465 ^ n833 ^ 1'b0 ;
  assign n13222 = ~n4081 & n13221 ;
  assign n13223 = n13222 ^ n10084 ^ n2222 ;
  assign n13224 = n7639 & ~n13223 ;
  assign n13225 = ~n13220 & n13224 ;
  assign n13226 = n8910 ^ n3689 ^ 1'b0 ;
  assign n13227 = ~n11115 & n13226 ;
  assign n13228 = ( ~n2436 & n8786 ) | ( ~n2436 & n13227 ) | ( n8786 & n13227 ) ;
  assign n13229 = n1449 & n4118 ;
  assign n13230 = n11019 & n13229 ;
  assign n13231 = n466 ^ n170 ^ 1'b0 ;
  assign n13232 = n2389 & ~n13231 ;
  assign n13233 = ( n2762 & n3991 ) | ( n2762 & ~n13232 ) | ( n3991 & ~n13232 ) ;
  assign n13234 = n13233 ^ n8782 ^ n2205 ;
  assign n13235 = ( n7239 & ~n12135 ) | ( n7239 & n13234 ) | ( ~n12135 & n13234 ) ;
  assign n13236 = n9914 & ~n13235 ;
  assign n13237 = n6785 & ~n10339 ;
  assign n13238 = n13237 ^ n7203 ^ 1'b0 ;
  assign n13239 = ( n4828 & ~n8637 ) | ( n4828 & n9065 ) | ( ~n8637 & n9065 ) ;
  assign n13240 = n13239 ^ n6725 ^ 1'b0 ;
  assign n13241 = n4878 ^ n1508 ^ 1'b0 ;
  assign n13242 = n8049 & ~n13241 ;
  assign n13244 = ( n307 & ~n5153 ) | ( n307 & n8133 ) | ( ~n5153 & n8133 ) ;
  assign n13243 = ( n679 & n5229 ) | ( n679 & ~n9391 ) | ( n5229 & ~n9391 ) ;
  assign n13245 = n13244 ^ n13243 ^ n7469 ;
  assign n13246 = n5724 ^ n4064 ^ 1'b0 ;
  assign n13247 = ( ~n3996 & n6497 ) | ( ~n3996 & n13246 ) | ( n6497 & n13246 ) ;
  assign n13248 = ( n13242 & ~n13245 ) | ( n13242 & n13247 ) | ( ~n13245 & n13247 ) ;
  assign n13249 = n3799 ^ n861 ^ 1'b0 ;
  assign n13250 = n3204 ^ n689 ^ 1'b0 ;
  assign n13251 = n571 & ~n13250 ;
  assign n13252 = ~n597 & n6082 ;
  assign n13253 = n13252 ^ n12059 ^ 1'b0 ;
  assign n13254 = n3980 | n6654 ;
  assign n13255 = n13254 ^ n10488 ^ 1'b0 ;
  assign n13256 = n13255 ^ n4365 ^ 1'b0 ;
  assign n13257 = n3887 | n4800 ;
  assign n13258 = n13257 ^ n6971 ^ 1'b0 ;
  assign n13259 = n5453 & n6649 ;
  assign n13260 = n8776 ^ n670 ^ 1'b0 ;
  assign n13265 = n5108 ^ n296 ^ 1'b0 ;
  assign n13266 = n12683 & n13265 ;
  assign n13267 = n13266 ^ n6672 ^ n5670 ;
  assign n13263 = n2682 ^ n2222 ^ 1'b0 ;
  assign n13261 = n6659 ^ n3321 ^ n791 ;
  assign n13262 = n13261 ^ n6475 ^ 1'b0 ;
  assign n13264 = n13263 ^ n13262 ^ 1'b0 ;
  assign n13268 = n13267 ^ n13264 ^ 1'b0 ;
  assign n13269 = n5342 & ~n10830 ;
  assign n13270 = n10961 ^ n5604 ^ 1'b0 ;
  assign n13271 = n4888 ^ n4036 ^ n3698 ;
  assign n13272 = n4297 ^ n3003 ^ n2614 ;
  assign n13273 = n4804 & n13272 ;
  assign n13274 = n13273 ^ n6492 ^ 1'b0 ;
  assign n13275 = n6014 & ~n8055 ;
  assign n13276 = n11931 ^ n5867 ^ n3060 ;
  assign n13277 = n8978 ^ n2174 ^ 1'b0 ;
  assign n13278 = n3455 & ~n13277 ;
  assign n13279 = n452 & n13278 ;
  assign n13280 = n10196 ^ n8632 ^ 1'b0 ;
  assign n13281 = n5843 & n13280 ;
  assign n13282 = n13281 ^ n11668 ^ n8648 ;
  assign n13283 = n4853 & n12890 ;
  assign n13284 = n13283 ^ n10373 ^ 1'b0 ;
  assign n13285 = ( n1518 & n2400 ) | ( n1518 & n4784 ) | ( n2400 & n4784 ) ;
  assign n13286 = n13285 ^ n7381 ^ 1'b0 ;
  assign n13287 = n9588 | n13286 ;
  assign n13288 = n12550 ^ n6193 ^ n3968 ;
  assign n13289 = ( n1689 & n10634 ) | ( n1689 & ~n13288 ) | ( n10634 & ~n13288 ) ;
  assign n13290 = n144 | n13289 ;
  assign n13291 = n2674 | n13290 ;
  assign n13292 = n11391 ^ n6577 ^ n341 ;
  assign n13293 = n7507 & n13141 ;
  assign n13294 = n3605 ^ n339 ^ n304 ;
  assign n13295 = n3104 ^ x108 ^ 1'b0 ;
  assign n13296 = n13295 ^ n10218 ^ 1'b0 ;
  assign n13297 = n13296 ^ n2102 ^ 1'b0 ;
  assign n13298 = ( n173 & n7626 ) | ( n173 & n8472 ) | ( n7626 & n8472 ) ;
  assign n13299 = n13298 ^ n2702 ^ 1'b0 ;
  assign n13300 = n5721 & n13299 ;
  assign n13301 = n13300 ^ n1861 ^ 1'b0 ;
  assign n13302 = ~n1542 & n9250 ;
  assign n13303 = ~n3974 & n4957 ;
  assign n13304 = n12860 & n13303 ;
  assign n13305 = ( n2951 & ~n9113 ) | ( n2951 & n11626 ) | ( ~n9113 & n11626 ) ;
  assign n13306 = ( ~n2623 & n6079 ) | ( ~n2623 & n13305 ) | ( n6079 & n13305 ) ;
  assign n13307 = n1682 | n4397 ;
  assign n13308 = n4397 & ~n13307 ;
  assign n13309 = n13308 ^ n13011 ^ n6529 ;
  assign n13310 = n6924 & ~n7180 ;
  assign n13311 = ~n2547 & n13310 ;
  assign n13312 = n4925 & n8444 ;
  assign n13313 = n13312 ^ n12423 ^ 1'b0 ;
  assign n13315 = ( n1082 & n3029 ) | ( n1082 & n4267 ) | ( n3029 & n4267 ) ;
  assign n13314 = ( n1213 & ~n2497 ) | ( n1213 & n4655 ) | ( ~n2497 & n4655 ) ;
  assign n13316 = n13315 ^ n13314 ^ n714 ;
  assign n13317 = n11325 ^ n8895 ^ 1'b0 ;
  assign n13318 = n1894 & ~n9170 ;
  assign n13319 = n13318 ^ n1223 ^ 1'b0 ;
  assign n13320 = ( ~x75 & n7174 ) | ( ~x75 & n13319 ) | ( n7174 & n13319 ) ;
  assign n13321 = ~n4259 & n7644 ;
  assign n13322 = n13321 ^ n4743 ^ 1'b0 ;
  assign n13324 = ( n1419 & n2499 ) | ( n1419 & n6785 ) | ( n2499 & n6785 ) ;
  assign n13325 = ( n3630 & ~n3824 ) | ( n3630 & n13324 ) | ( ~n3824 & n13324 ) ;
  assign n13323 = ~n511 & n12164 ;
  assign n13326 = n13325 ^ n13323 ^ 1'b0 ;
  assign n13327 = n12505 ^ n9327 ^ n1798 ;
  assign n13328 = ( n6142 & ~n6233 ) | ( n6142 & n12779 ) | ( ~n6233 & n12779 ) ;
  assign n13329 = ~n1547 & n2114 ;
  assign n13330 = ~n11637 & n13329 ;
  assign n13334 = n4044 ^ n3225 ^ n1568 ;
  assign n13331 = n2996 | n7134 ;
  assign n13332 = n4446 & ~n13331 ;
  assign n13333 = n13332 ^ n13285 ^ n9007 ;
  assign n13335 = n13334 ^ n13333 ^ 1'b0 ;
  assign n13336 = n13330 | n13335 ;
  assign n13337 = ~n3067 & n4938 ;
  assign n13338 = n517 & ~n13337 ;
  assign n13339 = ~n4567 & n10193 ;
  assign n13340 = n2947 ^ n2138 ^ n1810 ;
  assign n13341 = ( ~n13338 & n13339 ) | ( ~n13338 & n13340 ) | ( n13339 & n13340 ) ;
  assign n13342 = n2767 | n4403 ;
  assign n13343 = n13342 ^ n12663 ^ 1'b0 ;
  assign n13344 = n5311 & ~n5345 ;
  assign n13345 = ~n9273 & n13344 ;
  assign n13346 = ~n13343 & n13345 ;
  assign n13347 = n7112 ^ n2242 ^ 1'b0 ;
  assign n13348 = n1212 | n13347 ;
  assign n13349 = ( n6644 & n7025 ) | ( n6644 & ~n9041 ) | ( n7025 & ~n9041 ) ;
  assign n13350 = n3010 | n12166 ;
  assign n13351 = n4633 | n13350 ;
  assign n13352 = n10411 & ~n13351 ;
  assign n13353 = n6494 & ~n7824 ;
  assign n13354 = n13353 ^ n10742 ^ n9343 ;
  assign n13355 = n13354 ^ n9683 ^ 1'b0 ;
  assign n13356 = n6368 | n13355 ;
  assign n13357 = n13034 ^ n2718 ^ 1'b0 ;
  assign n13358 = n3276 & ~n3558 ;
  assign n13359 = ~n5675 & n6815 ;
  assign n13360 = ~x61 & n13359 ;
  assign n13361 = n5821 & ~n13360 ;
  assign n13362 = n1355 | n3503 ;
  assign n13363 = n13362 ^ n2100 ^ 1'b0 ;
  assign n13364 = n264 | n13363 ;
  assign n13365 = n10139 & ~n13364 ;
  assign n13366 = n9258 ^ n8104 ^ 1'b0 ;
  assign n13367 = n305 & n13366 ;
  assign n13368 = n13367 ^ x64 ^ 1'b0 ;
  assign n13369 = n13368 ^ n4183 ^ n375 ;
  assign n13370 = n4254 ^ n781 ^ 1'b0 ;
  assign n13371 = ( n758 & n3131 ) | ( n758 & n5519 ) | ( n3131 & n5519 ) ;
  assign n13372 = n13371 ^ n9217 ^ 1'b0 ;
  assign n13373 = n13370 & ~n13372 ;
  assign n13374 = n7320 ^ n4566 ^ 1'b0 ;
  assign n13375 = n7721 | n13374 ;
  assign n13376 = n1149 | n5367 ;
  assign n13377 = n13376 ^ n2896 ^ 1'b0 ;
  assign n13378 = ~n10370 & n13377 ;
  assign n13379 = n5782 ^ n5660 ^ 1'b0 ;
  assign n13380 = ~n8558 & n13379 ;
  assign n13381 = n10382 ^ n668 ^ 1'b0 ;
  assign n13382 = n13381 ^ n1979 ^ 1'b0 ;
  assign n13383 = n983 & ~n13382 ;
  assign n13384 = n9857 ^ n6180 ^ 1'b0 ;
  assign n13385 = n5952 | n13384 ;
  assign n13386 = n12662 ^ n5101 ^ 1'b0 ;
  assign n13387 = n8672 ^ n3611 ^ 1'b0 ;
  assign n13388 = ( n2564 & n3366 ) | ( n2564 & ~n4609 ) | ( n3366 & ~n4609 ) ;
  assign n13389 = ( n7959 & n12690 ) | ( n7959 & ~n13388 ) | ( n12690 & ~n13388 ) ;
  assign n13390 = n13389 ^ n9233 ^ 1'b0 ;
  assign n13391 = ~n2870 & n13390 ;
  assign n13392 = n227 & n7729 ;
  assign n13393 = n4819 & n13392 ;
  assign n13394 = n11105 & ~n13393 ;
  assign n13395 = n13394 ^ n3876 ^ 1'b0 ;
  assign n13396 = ( x3 & ~n500 ) | ( x3 & n4877 ) | ( ~n500 & n4877 ) ;
  assign n13397 = n5118 & n13396 ;
  assign n13398 = n11420 & n13397 ;
  assign n13399 = ( ~x75 & n5792 ) | ( ~x75 & n13398 ) | ( n5792 & n13398 ) ;
  assign n13400 = n13399 ^ n4666 ^ n1542 ;
  assign n13401 = ~n8046 & n13400 ;
  assign n13402 = ~n6768 & n13401 ;
  assign n13403 = ( n675 & n3218 ) | ( n675 & ~n7417 ) | ( n3218 & ~n7417 ) ;
  assign n13404 = n4726 | n10194 ;
  assign n13405 = n1379 | n13404 ;
  assign n13406 = n157 & ~n2585 ;
  assign n13407 = ( n1172 & ~n11730 ) | ( n1172 & n13406 ) | ( ~n11730 & n13406 ) ;
  assign n13408 = n13407 ^ n1978 ^ 1'b0 ;
  assign n13409 = x56 & n3682 ;
  assign n13410 = ( n3027 & n8869 ) | ( n3027 & n8912 ) | ( n8869 & n8912 ) ;
  assign n13411 = n1278 & n13410 ;
  assign n13416 = ( n390 & n2905 ) | ( n390 & n5539 ) | ( n2905 & n5539 ) ;
  assign n13417 = n13416 ^ n10467 ^ n8191 ;
  assign n13418 = n10918 ^ n6848 ^ 1'b0 ;
  assign n13419 = n13417 & n13418 ;
  assign n13412 = n272 | n2337 ;
  assign n13413 = n13412 ^ n905 ^ 1'b0 ;
  assign n13414 = ~n2811 & n13413 ;
  assign n13415 = n7671 & ~n13414 ;
  assign n13420 = n13419 ^ n13415 ^ 1'b0 ;
  assign n13421 = ( n2136 & n4625 ) | ( n2136 & ~n6704 ) | ( n4625 & ~n6704 ) ;
  assign n13422 = ( n2994 & n5398 ) | ( n2994 & ~n8323 ) | ( n5398 & ~n8323 ) ;
  assign n13423 = n13422 ^ n1132 ^ 1'b0 ;
  assign n13424 = n10815 & ~n13423 ;
  assign n13425 = ( n384 & n3183 ) | ( n384 & ~n8844 ) | ( n3183 & ~n8844 ) ;
  assign n13426 = n13425 ^ n10562 ^ n7599 ;
  assign n13427 = ( ~n7644 & n13424 ) | ( ~n7644 & n13426 ) | ( n13424 & n13426 ) ;
  assign n13428 = n13427 ^ n5215 ^ 1'b0 ;
  assign n13429 = ~n13421 & n13428 ;
  assign n13430 = n3229 ^ n650 ^ n318 ;
  assign n13431 = ( n180 & ~n10321 ) | ( n180 & n12218 ) | ( ~n10321 & n12218 ) ;
  assign n13432 = n13431 ^ n10388 ^ n1962 ;
  assign n13433 = ( n4177 & n6085 ) | ( n4177 & ~n10480 ) | ( n6085 & ~n10480 ) ;
  assign n13434 = n13433 ^ n13413 ^ n531 ;
  assign n13435 = n13434 ^ n4918 ^ 1'b0 ;
  assign n13436 = n871 & ~n13435 ;
  assign n13437 = n13199 ^ n9347 ^ 1'b0 ;
  assign n13438 = n3301 & ~n13437 ;
  assign n13439 = n3239 & n10991 ;
  assign n13441 = ( ~n567 & n2132 ) | ( ~n567 & n7639 ) | ( n2132 & n7639 ) ;
  assign n13442 = n6607 | n13441 ;
  assign n13443 = n13442 ^ n2344 ^ 1'b0 ;
  assign n13440 = n11949 ^ n10926 ^ n2402 ;
  assign n13444 = n13443 ^ n13440 ^ 1'b0 ;
  assign n13445 = n12635 & ~n13444 ;
  assign n13446 = n11525 & ~n13445 ;
  assign n13448 = n664 & ~n6566 ;
  assign n13447 = n878 & ~n13152 ;
  assign n13449 = n13448 ^ n13447 ^ 1'b0 ;
  assign n13450 = n1902 | n13449 ;
  assign n13451 = n11250 | n13450 ;
  assign n13452 = n13451 ^ n6590 ^ n5561 ;
  assign n13458 = ( ~x52 & n3439 ) | ( ~x52 & n11632 ) | ( n3439 & n11632 ) ;
  assign n13453 = n6256 ^ n3084 ^ 1'b0 ;
  assign n13454 = n6187 | n13453 ;
  assign n13455 = n13454 ^ n3325 ^ 1'b0 ;
  assign n13456 = n13204 ^ n12245 ^ 1'b0 ;
  assign n13457 = n13455 & ~n13456 ;
  assign n13459 = n13458 ^ n13457 ^ n5661 ;
  assign n13460 = ( n2334 & n3555 ) | ( n2334 & ~n6271 ) | ( n3555 & ~n6271 ) ;
  assign n13461 = n7168 ^ x42 ^ 1'b0 ;
  assign n13462 = ( ~n2718 & n9423 ) | ( ~n2718 & n13461 ) | ( n9423 & n13461 ) ;
  assign n13463 = ( n422 & ~n13460 ) | ( n422 & n13462 ) | ( ~n13460 & n13462 ) ;
  assign n13464 = n2712 | n3572 ;
  assign n13465 = n10790 ^ n4758 ^ n2027 ;
  assign n13466 = n8467 ^ n2897 ^ 1'b0 ;
  assign n13467 = n6755 | n13466 ;
  assign n13468 = n4509 & ~n5727 ;
  assign n13469 = n3035 | n13468 ;
  assign n13470 = n8065 & ~n13469 ;
  assign n13471 = n13470 ^ n3879 ^ 1'b0 ;
  assign n13472 = n5381 | n6592 ;
  assign n13473 = ( n2050 & ~n9144 ) | ( n2050 & n13472 ) | ( ~n9144 & n13472 ) ;
  assign n13474 = n1490 & ~n2515 ;
  assign n13475 = ~n4962 & n13474 ;
  assign n13476 = n3003 & ~n3020 ;
  assign n13477 = n13476 ^ n5942 ^ 1'b0 ;
  assign n13478 = n4653 ^ n1431 ^ n352 ;
  assign n13479 = n13478 ^ n2787 ^ 1'b0 ;
  assign n13480 = n13479 ^ n10374 ^ 1'b0 ;
  assign n13481 = ( n6947 & n13477 ) | ( n6947 & ~n13480 ) | ( n13477 & ~n13480 ) ;
  assign n13482 = ( n6835 & n12453 ) | ( n6835 & ~n13481 ) | ( n12453 & ~n13481 ) ;
  assign n13483 = n9065 ^ n1406 ^ 1'b0 ;
  assign n13484 = ( n1509 & n2638 ) | ( n1509 & n3817 ) | ( n2638 & n3817 ) ;
  assign n13490 = n11342 ^ n7839 ^ n2674 ;
  assign n13485 = n6551 ^ n3746 ^ n3137 ;
  assign n13486 = ~n4401 & n12484 ;
  assign n13487 = n10175 & n13486 ;
  assign n13488 = n13485 & ~n13487 ;
  assign n13489 = n13488 ^ n1387 ^ 1'b0 ;
  assign n13491 = n13490 ^ n13489 ^ n9829 ;
  assign n13492 = n8454 ^ n1050 ^ 1'b0 ;
  assign n13493 = n9042 ^ n8225 ^ n1267 ;
  assign n13499 = ( ~n454 & n1704 ) | ( ~n454 & n3672 ) | ( n1704 & n3672 ) ;
  assign n13494 = n986 ^ n779 ^ 1'b0 ;
  assign n13495 = n5034 & n6829 ;
  assign n13496 = n13495 ^ n432 ^ 1'b0 ;
  assign n13497 = n13496 ^ n3698 ^ 1'b0 ;
  assign n13498 = ( n5131 & ~n13494 ) | ( n5131 & n13497 ) | ( ~n13494 & n13497 ) ;
  assign n13500 = n13499 ^ n13498 ^ 1'b0 ;
  assign n13501 = ~n13493 & n13500 ;
  assign n13502 = n12301 ^ n269 ^ 1'b0 ;
  assign n13503 = n6532 ^ n1935 ^ n310 ;
  assign n13504 = n13503 ^ n7951 ^ 1'b0 ;
  assign n13505 = ~n5905 & n13504 ;
  assign n13506 = ~n3476 & n5474 ;
  assign n13507 = ~n13505 & n13506 ;
  assign n13508 = n13507 ^ n4725 ^ n4085 ;
  assign n13509 = n13238 ^ n6003 ^ 1'b0 ;
  assign n13510 = n12222 ^ n9607 ^ 1'b0 ;
  assign n13511 = ~n10850 & n13510 ;
  assign n13512 = ~n5600 & n13511 ;
  assign n13513 = ~n2072 & n13512 ;
  assign n13514 = ~n3648 & n3707 ;
  assign n13515 = n13514 ^ n462 ^ 1'b0 ;
  assign n13516 = n13467 ^ n9571 ^ 1'b0 ;
  assign n13517 = n13515 & n13516 ;
  assign n13518 = n4725 ^ n4371 ^ 1'b0 ;
  assign n13519 = n1901 & n13518 ;
  assign n13520 = n13177 & ~n13519 ;
  assign n13524 = ~n458 & n2882 ;
  assign n13525 = n13524 ^ n328 ^ 1'b0 ;
  assign n13526 = ~n256 & n13525 ;
  assign n13521 = n9857 & n10843 ;
  assign n13522 = n5040 & n13521 ;
  assign n13523 = n373 | n13522 ;
  assign n13527 = n13526 ^ n13523 ^ 1'b0 ;
  assign n13528 = n12450 ^ n3597 ^ 1'b0 ;
  assign n13529 = n3264 & ~n13528 ;
  assign n13530 = n13529 ^ n11421 ^ n3636 ;
  assign n13531 = n13530 ^ n7721 ^ 1'b0 ;
  assign n13532 = n10432 & ~n13531 ;
  assign n13533 = n5799 ^ n514 ^ 1'b0 ;
  assign n13534 = n6178 & n7450 ;
  assign n13535 = n2975 | n13534 ;
  assign n13536 = n13535 ^ n8264 ^ 1'b0 ;
  assign n13537 = ~n8490 & n9698 ;
  assign n13538 = n1842 ^ n1135 ^ 1'b0 ;
  assign n13539 = n10689 ^ n1717 ^ n1511 ;
  assign n13540 = ~n2679 & n10777 ;
  assign n13541 = n13539 & n13540 ;
  assign n13542 = n13541 ^ n11834 ^ n7178 ;
  assign n13543 = ~n7211 & n13542 ;
  assign n13545 = n6547 ^ n6309 ^ n2416 ;
  assign n13544 = n4942 & n5582 ;
  assign n13546 = n13545 ^ n13544 ^ 1'b0 ;
  assign n13548 = ~n1201 & n3116 ;
  assign n13549 = n13548 ^ n1874 ^ 1'b0 ;
  assign n13547 = n3101 & ~n4693 ;
  assign n13550 = n13549 ^ n13547 ^ 1'b0 ;
  assign n13551 = n13550 ^ n9987 ^ n1101 ;
  assign n13552 = n13551 ^ n9740 ^ 1'b0 ;
  assign n13553 = ~n12104 & n13472 ;
  assign n13554 = n10087 ^ n9876 ^ 1'b0 ;
  assign n13555 = n13553 & n13554 ;
  assign n13556 = n6797 ^ n1553 ^ 1'b0 ;
  assign n13557 = ( n8969 & n13555 ) | ( n8969 & ~n13556 ) | ( n13555 & ~n13556 ) ;
  assign n13558 = ~n6121 & n10827 ;
  assign n13559 = n13558 ^ n12965 ^ 1'b0 ;
  assign n13560 = ( n2352 & n4274 ) | ( n2352 & ~n10767 ) | ( n4274 & ~n10767 ) ;
  assign n13561 = n13559 & ~n13560 ;
  assign n13562 = n13561 ^ n10053 ^ 1'b0 ;
  assign n13564 = n4457 ^ n289 ^ 1'b0 ;
  assign n13563 = n6911 | n11203 ;
  assign n13565 = n13564 ^ n13563 ^ 1'b0 ;
  assign n13566 = n9111 ^ n6570 ^ n2175 ;
  assign n13567 = n13566 ^ n9829 ^ 1'b0 ;
  assign n13568 = n8932 & ~n10576 ;
  assign n13569 = n8046 & n13568 ;
  assign n13570 = ~n5434 & n9434 ;
  assign n13571 = ~n8606 & n13570 ;
  assign n13572 = n13571 ^ n497 ^ 1'b0 ;
  assign n13573 = n1264 & n13572 ;
  assign n13574 = n13573 ^ n6916 ^ 1'b0 ;
  assign n13575 = n1076 & ~n13574 ;
  assign n13580 = n7735 | n8007 ;
  assign n13576 = n584 | n5356 ;
  assign n13577 = n13576 ^ n11038 ^ n4265 ;
  assign n13578 = n3299 & ~n13577 ;
  assign n13579 = n6197 & n13578 ;
  assign n13581 = n13580 ^ n13579 ^ n3018 ;
  assign n13582 = n3171 ^ x106 ^ 1'b0 ;
  assign n13583 = n704 & n2317 ;
  assign n13584 = n12647 | n13583 ;
  assign n13585 = n13584 ^ n1276 ^ 1'b0 ;
  assign n13586 = ~n13582 & n13585 ;
  assign n13587 = n10708 & n11098 ;
  assign n13588 = ~n5099 & n13587 ;
  assign n13589 = n10465 & n13588 ;
  assign n13590 = ( ~n2521 & n5071 ) | ( ~n2521 & n6196 ) | ( n5071 & n6196 ) ;
  assign n13591 = n13590 ^ n2539 ^ x84 ;
  assign n13592 = n2263 & n13591 ;
  assign n13593 = ~n8836 & n13592 ;
  assign n13594 = n11297 ^ n4008 ^ n1998 ;
  assign n13595 = n13594 ^ n7695 ^ n915 ;
  assign n13596 = n10871 & ~n13595 ;
  assign n13597 = ( n188 & n5868 ) | ( n188 & n8296 ) | ( n5868 & n8296 ) ;
  assign n13598 = ~n6600 & n13597 ;
  assign n13599 = ( n8908 & n10445 ) | ( n8908 & ~n12047 ) | ( n10445 & ~n12047 ) ;
  assign n13600 = n8600 ^ n4745 ^ n3409 ;
  assign n13601 = n13600 ^ n2840 ^ n1019 ;
  assign n13602 = ( ~n1232 & n12287 ) | ( ~n1232 & n13601 ) | ( n12287 & n13601 ) ;
  assign n13603 = ~n10017 & n12392 ;
  assign n13604 = n13603 ^ n8966 ^ 1'b0 ;
  assign n13605 = ~n560 & n13604 ;
  assign n13606 = n4242 & n5909 ;
  assign n13607 = ~n908 & n13606 ;
  assign n13608 = n12749 ^ n4158 ^ 1'b0 ;
  assign n13609 = n13607 | n13608 ;
  assign n13610 = n6990 & ~n9014 ;
  assign n13613 = n198 | n1846 ;
  assign n13611 = n6388 ^ n1784 ^ n809 ;
  assign n13612 = n13611 ^ n1961 ^ n1388 ;
  assign n13614 = n13613 ^ n13612 ^ n4691 ;
  assign n13615 = n7776 ^ n4900 ^ n3060 ;
  assign n13616 = n4691 ^ n2450 ^ 1'b0 ;
  assign n13617 = n13615 & n13616 ;
  assign n13618 = ( n154 & ~n13614 ) | ( n154 & n13617 ) | ( ~n13614 & n13617 ) ;
  assign n13619 = n5933 ^ n4190 ^ 1'b0 ;
  assign n13620 = ~n2378 & n13619 ;
  assign n13621 = n421 & n13620 ;
  assign n13622 = n13621 ^ n2458 ^ 1'b0 ;
  assign n13623 = ~n3026 & n9067 ;
  assign n13624 = n13421 ^ n5458 ^ 1'b0 ;
  assign n13625 = n13624 ^ n11886 ^ n11031 ;
  assign n13626 = ~n1671 & n13625 ;
  assign n13629 = n1097 & ~n3565 ;
  assign n13627 = n7053 & n12578 ;
  assign n13628 = n13627 ^ n10343 ^ n316 ;
  assign n13630 = n13629 ^ n13628 ^ n1374 ;
  assign n13631 = n4192 ^ n3515 ^ n144 ;
  assign n13632 = n13631 ^ n4256 ^ n3974 ;
  assign n13633 = n1288 | n13632 ;
  assign n13634 = n13633 ^ n5095 ^ 1'b0 ;
  assign n13635 = n1855 | n13634 ;
  assign n13646 = n8522 ^ n6018 ^ n4176 ;
  assign n13647 = ~n1828 & n13646 ;
  assign n13641 = n8856 ^ n1645 ^ 1'b0 ;
  assign n13642 = n7929 | n13641 ;
  assign n13643 = ( n468 & n1743 ) | ( n468 & ~n2627 ) | ( n1743 & ~n2627 ) ;
  assign n13644 = n13642 & n13643 ;
  assign n13636 = n11712 ^ n2752 ^ 1'b0 ;
  assign n13637 = n9635 | n13636 ;
  assign n13638 = n9860 ^ n1740 ^ 1'b0 ;
  assign n13639 = n13637 | n13638 ;
  assign n13640 = n2738 | n13639 ;
  assign n13645 = n13644 ^ n13640 ^ 1'b0 ;
  assign n13648 = n13647 ^ n13645 ^ n13470 ;
  assign n13649 = n256 | n8580 ;
  assign n13650 = n13649 ^ n6858 ^ 1'b0 ;
  assign n13651 = n5782 ^ n819 ^ 1'b0 ;
  assign n13652 = n8030 & n10763 ;
  assign n13658 = n1550 ^ n551 ^ 1'b0 ;
  assign n13653 = n4175 ^ n2051 ^ 1'b0 ;
  assign n13654 = n1966 & n13653 ;
  assign n13655 = ~n739 & n13654 ;
  assign n13656 = ~n7969 & n13655 ;
  assign n13657 = n849 | n13656 ;
  assign n13659 = n13658 ^ n13657 ^ 1'b0 ;
  assign n13660 = n511 ^ n373 ^ 1'b0 ;
  assign n13661 = n13660 ^ n5229 ^ n2141 ;
  assign n13662 = n13661 ^ n5322 ^ n2372 ;
  assign n13663 = n7627 ^ n6911 ^ n971 ;
  assign n13664 = n4645 & n5275 ;
  assign n13665 = ( n2829 & n13663 ) | ( n2829 & ~n13664 ) | ( n13663 & ~n13664 ) ;
  assign n13666 = n9183 ^ n5079 ^ n878 ;
  assign n13667 = n6103 ^ n615 ^ 1'b0 ;
  assign n13668 = n13667 ^ n10189 ^ 1'b0 ;
  assign n13669 = ~n11302 & n13668 ;
  assign n13670 = n9536 ^ n4592 ^ 1'b0 ;
  assign n13673 = ( ~n2647 & n4176 ) | ( ~n2647 & n5616 ) | ( n4176 & n5616 ) ;
  assign n13674 = n13673 ^ n9281 ^ n1132 ;
  assign n13671 = n2925 | n9315 ;
  assign n13672 = n13671 ^ n2370 ^ 1'b0 ;
  assign n13675 = n13674 ^ n13672 ^ n1720 ;
  assign n13676 = ( n1287 & n11720 ) | ( n1287 & ~n12287 ) | ( n11720 & ~n12287 ) ;
  assign n13677 = n13676 ^ n4832 ^ 1'b0 ;
  assign n13678 = n8431 ^ n7806 ^ 1'b0 ;
  assign n13679 = n5042 & n13678 ;
  assign n13681 = n10355 ^ n5853 ^ n5721 ;
  assign n13680 = ~n1553 & n5956 ;
  assign n13682 = n13681 ^ n13680 ^ n5439 ;
  assign n13683 = n1449 & ~n11607 ;
  assign n13684 = n132 | n3684 ;
  assign n13685 = ( n6093 & n12104 ) | ( n6093 & n13684 ) | ( n12104 & n13684 ) ;
  assign n13686 = n2222 & ~n12418 ;
  assign n13687 = ~n2558 & n13686 ;
  assign n13688 = n13685 | n13687 ;
  assign n13689 = n13021 & ~n13688 ;
  assign n13690 = n9200 & n10395 ;
  assign n13691 = n13413 & n13690 ;
  assign n13692 = n4989 ^ n1426 ^ 1'b0 ;
  assign n13693 = n5463 | n13692 ;
  assign n13694 = n6277 & n8228 ;
  assign n13695 = n2636 & n13694 ;
  assign n13696 = n13693 & ~n13695 ;
  assign n13697 = n13696 ^ n3858 ^ 1'b0 ;
  assign n13698 = n11343 ^ n227 ^ 1'b0 ;
  assign n13699 = n266 & n3738 ;
  assign n13700 = n13699 ^ n1856 ^ 1'b0 ;
  assign n13701 = n13700 ^ n10983 ^ n3750 ;
  assign n13702 = n13701 ^ n8661 ^ 1'b0 ;
  assign n13703 = n2511 & n13591 ;
  assign n13704 = n348 & ~n5014 ;
  assign n13705 = n13704 ^ n2340 ^ 1'b0 ;
  assign n13706 = n13705 ^ n6102 ^ 1'b0 ;
  assign n13707 = n13703 | n13706 ;
  assign n13708 = n13702 | n13707 ;
  assign n13709 = n10713 & ~n13095 ;
  assign n13710 = n13709 ^ n9179 ^ 1'b0 ;
  assign n13711 = ~n3637 & n6034 ;
  assign n13712 = n1094 & ~n5663 ;
  assign n13713 = n5071 & n13712 ;
  assign n13714 = n3169 | n13713 ;
  assign n13715 = n5427 & ~n13714 ;
  assign n13716 = ( ~n2222 & n9553 ) | ( ~n2222 & n12083 ) | ( n9553 & n12083 ) ;
  assign n13717 = n4544 ^ n169 ^ 1'b0 ;
  assign n13718 = n13717 ^ n10881 ^ n3637 ;
  assign n13719 = n5351 & ~n13718 ;
  assign n13720 = ~n9413 & n13719 ;
  assign n13721 = n13720 ^ n9588 ^ n1804 ;
  assign n13722 = ~n13716 & n13721 ;
  assign n13723 = n8807 & n13722 ;
  assign n13724 = ~n4462 & n8342 ;
  assign n13725 = n3312 & ~n12183 ;
  assign n13726 = ~n2152 & n13725 ;
  assign n13727 = ( n2191 & ~n12662 ) | ( n2191 & n13726 ) | ( ~n12662 & n13726 ) ;
  assign n13728 = n8957 ^ n4111 ^ 1'b0 ;
  assign n13729 = n8032 & n13728 ;
  assign n13730 = ( n5928 & ~n13526 ) | ( n5928 & n13729 ) | ( ~n13526 & n13729 ) ;
  assign n13731 = n5322 | n9475 ;
  assign n13732 = ~n5224 & n7061 ;
  assign n13733 = n3212 & n13732 ;
  assign n13734 = n11721 | n13733 ;
  assign n13735 = n5118 | n13734 ;
  assign n13736 = ( n7959 & n9664 ) | ( n7959 & ~n10503 ) | ( n9664 & ~n10503 ) ;
  assign n13737 = n7757 ^ n1385 ^ 1'b0 ;
  assign n13738 = n12146 | n13737 ;
  assign n13739 = ( n3043 & n9690 ) | ( n3043 & n10166 ) | ( n9690 & n10166 ) ;
  assign n13740 = n5441 | n13739 ;
  assign n13741 = n3798 & ~n13740 ;
  assign n13742 = n13741 ^ n1545 ^ 1'b0 ;
  assign n13743 = ~n4986 & n9483 ;
  assign n13744 = ~n3964 & n13743 ;
  assign n13745 = n13742 & n13744 ;
  assign n13746 = ~n1413 & n6330 ;
  assign n13747 = n13746 ^ n1117 ^ 1'b0 ;
  assign n13748 = n1862 | n4185 ;
  assign n13749 = ( ~n3371 & n11421 ) | ( ~n3371 & n13748 ) | ( n11421 & n13748 ) ;
  assign n13750 = n13702 ^ n928 ^ 1'b0 ;
  assign n13753 = ( n1176 & n4642 ) | ( n1176 & ~n6675 ) | ( n4642 & ~n6675 ) ;
  assign n13751 = n2816 & ~n10915 ;
  assign n13752 = n899 & n13751 ;
  assign n13754 = n13753 ^ n13752 ^ n9207 ;
  assign n13755 = n10199 & ~n13754 ;
  assign n13756 = n5336 ^ n1074 ^ 1'b0 ;
  assign n13757 = ( n2458 & n2749 ) | ( n2458 & n11307 ) | ( n2749 & n11307 ) ;
  assign n13758 = ( ~n2481 & n2921 ) | ( ~n2481 & n4433 ) | ( n2921 & n4433 ) ;
  assign n13759 = n13758 ^ n846 ^ 1'b0 ;
  assign n13760 = n5603 | n13759 ;
  assign n13761 = n13760 ^ n4094 ^ 1'b0 ;
  assign n13762 = n13738 & n13761 ;
  assign n13763 = n299 & n2239 ;
  assign n13764 = n6146 & n13763 ;
  assign n13765 = n9450 | n13764 ;
  assign n13766 = n13765 ^ n1883 ^ 1'b0 ;
  assign n13767 = n9678 ^ n5057 ^ 1'b0 ;
  assign n13768 = n378 & n4328 ;
  assign n13769 = n6796 & n13768 ;
  assign n13770 = n2023 & ~n13769 ;
  assign n13771 = ~n3285 & n13770 ;
  assign n13772 = n10134 ^ n1035 ^ 1'b0 ;
  assign n13773 = n6808 & ~n10689 ;
  assign n13774 = n10288 & n13773 ;
  assign n13775 = ( ~n4912 & n12405 ) | ( ~n4912 & n13774 ) | ( n12405 & n13774 ) ;
  assign n13776 = n6598 | n9343 ;
  assign n13777 = ~n1342 & n7568 ;
  assign n13778 = n13777 ^ n1738 ^ 1'b0 ;
  assign n13779 = n1979 | n3645 ;
  assign n13780 = n6884 | n13779 ;
  assign n13781 = ( n1718 & n2273 ) | ( n1718 & n6506 ) | ( n2273 & n6506 ) ;
  assign n13782 = n987 & ~n13781 ;
  assign n13783 = n13782 ^ n577 ^ 1'b0 ;
  assign n13784 = n8828 ^ n7048 ^ 1'b0 ;
  assign n13785 = ( n11126 & ~n13783 ) | ( n11126 & n13784 ) | ( ~n13783 & n13784 ) ;
  assign n13786 = n3274 & n3704 ;
  assign n13787 = n13786 ^ n2205 ^ 1'b0 ;
  assign n13788 = n13654 ^ n11039 ^ n7744 ;
  assign n13789 = ( n1819 & ~n13787 ) | ( n1819 & n13788 ) | ( ~n13787 & n13788 ) ;
  assign n13790 = n12002 & n12065 ;
  assign n13791 = n1745 & n13790 ;
  assign n13792 = n3994 & ~n5048 ;
  assign n13793 = ( n6918 & n12044 ) | ( n6918 & ~n13792 ) | ( n12044 & ~n13792 ) ;
  assign n13794 = n9965 ^ n4854 ^ 1'b0 ;
  assign n13795 = n5519 | n13794 ;
  assign n13796 = n13795 ^ n11775 ^ 1'b0 ;
  assign n13797 = n12685 ^ n11341 ^ 1'b0 ;
  assign n13798 = n10394 ^ n1517 ^ 1'b0 ;
  assign n13799 = n7838 ^ n848 ^ 1'b0 ;
  assign n13800 = ~n8802 & n13799 ;
  assign n13801 = n13798 & n13800 ;
  assign n13803 = ~n2329 & n5234 ;
  assign n13804 = n5713 & n13803 ;
  assign n13802 = n5228 | n11776 ;
  assign n13805 = n13804 ^ n13802 ^ n12053 ;
  assign n13806 = n7257 | n8343 ;
  assign n13807 = ~n390 & n11386 ;
  assign n13808 = n5778 & n13807 ;
  assign n13809 = n13263 ^ n5819 ^ 1'b0 ;
  assign n13810 = n1928 ^ n1525 ^ 1'b0 ;
  assign n13811 = ( n5632 & n7928 ) | ( n5632 & ~n13810 ) | ( n7928 & ~n13810 ) ;
  assign n13812 = n8415 & n11325 ;
  assign n13813 = n3363 & n6370 ;
  assign n13814 = ( ~n3582 & n7268 ) | ( ~n3582 & n11691 ) | ( n7268 & n11691 ) ;
  assign n13815 = ~n12522 & n13814 ;
  assign n13816 = n13815 ^ n6036 ^ n1319 ;
  assign n13817 = ( ~n3681 & n3715 ) | ( ~n3681 & n13255 ) | ( n3715 & n13255 ) ;
  assign n13818 = ( ~n1454 & n13816 ) | ( ~n1454 & n13817 ) | ( n13816 & n13817 ) ;
  assign n13819 = n10132 ^ n9364 ^ n2662 ;
  assign n13820 = n1564 ^ n462 ^ 1'b0 ;
  assign n13821 = n1907 | n13820 ;
  assign n13822 = n9427 & ~n13821 ;
  assign n13823 = n4946 ^ n3217 ^ 1'b0 ;
  assign n13824 = n347 | n13823 ;
  assign n13825 = n13824 ^ n6986 ^ 1'b0 ;
  assign n13826 = n141 | n3959 ;
  assign n13827 = n1764 ^ n985 ^ 1'b0 ;
  assign n13828 = n6596 & ~n7350 ;
  assign n13829 = ~n7022 & n13828 ;
  assign n13830 = ( ~n2929 & n13827 ) | ( ~n2929 & n13829 ) | ( n13827 & n13829 ) ;
  assign n13834 = ( n2805 & n8822 ) | ( n2805 & ~n12144 ) | ( n8822 & ~n12144 ) ;
  assign n13831 = n563 | n6306 ;
  assign n13832 = n4299 & ~n13831 ;
  assign n13833 = n2613 | n13832 ;
  assign n13835 = n13834 ^ n13833 ^ 1'b0 ;
  assign n13836 = ( n4221 & ~n4251 ) | ( n4221 & n10391 ) | ( ~n4251 & n10391 ) ;
  assign n13837 = n13836 ^ n5026 ^ 1'b0 ;
  assign n13838 = n1084 & n4747 ;
  assign n13839 = n13837 & n13838 ;
  assign n13840 = ~n3069 & n10986 ;
  assign n13841 = n1088 & n13840 ;
  assign n13842 = n7853 & ~n13841 ;
  assign n13843 = n7542 ^ n6144 ^ 1'b0 ;
  assign n13844 = n9501 ^ n4583 ^ n3507 ;
  assign n13845 = n11957 ^ x3 ^ 1'b0 ;
  assign n13846 = ~n8563 & n13845 ;
  assign n13847 = n2072 & n12693 ;
  assign n13848 = n5136 ^ n3943 ^ 1'b0 ;
  assign n13849 = n13848 ^ n5900 ^ n2737 ;
  assign n13850 = n833 & ~n8086 ;
  assign n13851 = n13850 ^ n307 ^ 1'b0 ;
  assign n13852 = n3156 ^ n1143 ^ 1'b0 ;
  assign n13853 = ( n5064 & ~n9039 ) | ( n5064 & n13852 ) | ( ~n9039 & n13852 ) ;
  assign n13854 = n13853 ^ n10218 ^ n1877 ;
  assign n13855 = n1714 | n6668 ;
  assign n13856 = n13855 ^ n1681 ^ 1'b0 ;
  assign n13857 = n641 ^ n274 ^ 1'b0 ;
  assign n13858 = ( n1781 & n13856 ) | ( n1781 & n13857 ) | ( n13856 & n13857 ) ;
  assign n13859 = n4636 ^ n1558 ^ 1'b0 ;
  assign n13860 = n2328 | n13859 ;
  assign n13861 = n522 & n2788 ;
  assign n13862 = ~n2091 & n13861 ;
  assign n13863 = n13862 ^ n11128 ^ 1'b0 ;
  assign n13864 = n10216 ^ n7482 ^ n2364 ;
  assign n13865 = n13864 ^ n11562 ^ n11487 ;
  assign n13866 = ( n4154 & ~n7528 ) | ( n4154 & n13865 ) | ( ~n7528 & n13865 ) ;
  assign n13867 = n11696 ^ n10911 ^ 1'b0 ;
  assign n13868 = n13823 ^ n5532 ^ 1'b0 ;
  assign n13869 = n2205 & ~n13868 ;
  assign n13870 = n13869 ^ n12465 ^ 1'b0 ;
  assign n13871 = n8546 & ~n13870 ;
  assign n13872 = n12549 ^ n10472 ^ 1'b0 ;
  assign n13873 = n13871 & ~n13872 ;
  assign n13874 = n7827 ^ n7411 ^ n4675 ;
  assign n13875 = ~n2470 & n7958 ;
  assign n13876 = ~n3991 & n13875 ;
  assign n13877 = ( n4716 & n13874 ) | ( n4716 & ~n13876 ) | ( n13874 & ~n13876 ) ;
  assign n13878 = n13877 ^ n5282 ^ 1'b0 ;
  assign n13879 = ~n8719 & n13878 ;
  assign n13880 = ~n13873 & n13879 ;
  assign n13881 = n589 | n3437 ;
  assign n13882 = n9167 | n13881 ;
  assign n13883 = n1754 | n13882 ;
  assign n13884 = n12752 | n13883 ;
  assign n13885 = n1032 | n3803 ;
  assign n13886 = n13885 ^ n5431 ^ 1'b0 ;
  assign n13887 = n4338 & ~n13582 ;
  assign n13888 = ( n2831 & n8502 ) | ( n2831 & n13739 ) | ( n8502 & n13739 ) ;
  assign n13889 = ~n4545 & n13888 ;
  assign n13890 = n3812 & n13889 ;
  assign n13891 = ( n3173 & n6750 ) | ( n3173 & ~n11622 ) | ( n6750 & ~n11622 ) ;
  assign n13893 = n5760 ^ n141 ^ 1'b0 ;
  assign n13892 = n8076 ^ n6967 ^ n538 ;
  assign n13894 = n13893 ^ n13892 ^ n6922 ;
  assign n13895 = ( n9354 & n10637 ) | ( n9354 & ~n13894 ) | ( n10637 & ~n13894 ) ;
  assign n13896 = ( n4272 & ~n9615 ) | ( n4272 & n13895 ) | ( ~n9615 & n13895 ) ;
  assign n13897 = ( n13666 & ~n13891 ) | ( n13666 & n13896 ) | ( ~n13891 & n13896 ) ;
  assign n13899 = n367 | n7532 ;
  assign n13900 = n13899 ^ n234 ^ 1'b0 ;
  assign n13898 = ( n840 & n3646 ) | ( n840 & ~n8733 ) | ( n3646 & ~n8733 ) ;
  assign n13901 = n13900 ^ n13898 ^ n3926 ;
  assign n13904 = n5564 | n7719 ;
  assign n13902 = n921 & n2530 ;
  assign n13903 = n3264 & n13902 ;
  assign n13905 = n13904 ^ n13903 ^ 1'b0 ;
  assign n13906 = n6947 | n10790 ;
  assign n13907 = n4526 | n13906 ;
  assign n13908 = n786 ^ x48 ^ 1'b0 ;
  assign n13909 = ( n3774 & n10792 ) | ( n3774 & n13908 ) | ( n10792 & n13908 ) ;
  assign n13910 = n7848 | n13909 ;
  assign n13911 = n13910 ^ n1068 ^ 1'b0 ;
  assign n13912 = n13911 ^ n13672 ^ 1'b0 ;
  assign n13913 = n4539 | n13912 ;
  assign n13914 = ~n154 & n3616 ;
  assign n13915 = ~n11927 & n13914 ;
  assign n13916 = n13915 ^ n5012 ^ n3027 ;
  assign n13917 = n6103 ^ n626 ^ 1'b0 ;
  assign n13918 = n13916 & ~n13917 ;
  assign n13919 = n8361 ^ n1364 ^ 1'b0 ;
  assign n13920 = n6218 ^ n4063 ^ 1'b0 ;
  assign n13921 = n2200 & n7794 ;
  assign n13922 = n13921 ^ n9529 ^ 1'b0 ;
  assign n13923 = n8058 & n13922 ;
  assign n13924 = n257 | n5002 ;
  assign n13925 = n13924 ^ n2822 ^ 1'b0 ;
  assign n13926 = n13208 ^ n6503 ^ n3679 ;
  assign n13929 = n2657 | n13051 ;
  assign n13927 = n10295 ^ n4114 ^ n1225 ;
  assign n13928 = n3979 & ~n13927 ;
  assign n13930 = n13929 ^ n13928 ^ 1'b0 ;
  assign n13931 = ~n348 & n13930 ;
  assign n13932 = ( ~n11781 & n11936 ) | ( ~n11781 & n13931 ) | ( n11936 & n13931 ) ;
  assign n13933 = ( n834 & n1773 ) | ( n834 & ~n2168 ) | ( n1773 & ~n2168 ) ;
  assign n13934 = n12895 & ~n13933 ;
  assign n13937 = n7153 ^ n6750 ^ x18 ;
  assign n13938 = ( ~n2975 & n6399 ) | ( ~n2975 & n13937 ) | ( n6399 & n13937 ) ;
  assign n13935 = n694 & n2508 ;
  assign n13936 = ~n250 & n13935 ;
  assign n13939 = n13938 ^ n13936 ^ n180 ;
  assign n13940 = ~n3163 & n13939 ;
  assign n13942 = n3449 ^ n1207 ^ 1'b0 ;
  assign n13941 = n259 | n6024 ;
  assign n13943 = n13942 ^ n13941 ^ n1938 ;
  assign n13944 = n4524 | n13943 ;
  assign n13945 = n13944 ^ n7939 ^ n6204 ;
  assign n13946 = n13945 ^ n3607 ^ 1'b0 ;
  assign n13947 = n13144 ^ n12508 ^ x22 ;
  assign n13948 = n418 | n7085 ;
  assign n13949 = ~n1603 & n11722 ;
  assign n13950 = n2739 & n8528 ;
  assign n13951 = n13950 ^ n2657 ^ 1'b0 ;
  assign n13952 = n5259 ^ n2573 ^ 1'b0 ;
  assign n13953 = n13951 & n13952 ;
  assign n13954 = ~n295 & n11067 ;
  assign n13955 = n13954 ^ n6218 ^ 1'b0 ;
  assign n13956 = n2317 ^ n1168 ^ 1'b0 ;
  assign n13957 = n13955 & n13956 ;
  assign n13958 = n8909 & ~n9406 ;
  assign n13959 = ~n5859 & n13958 ;
  assign n13964 = ~n5157 & n5532 ;
  assign n13965 = n2499 & n13964 ;
  assign n13962 = n1929 & ~n7333 ;
  assign n13963 = n13962 ^ n7467 ^ 1'b0 ;
  assign n13960 = ( n1422 & n3188 ) | ( n1422 & n6628 ) | ( n3188 & n6628 ) ;
  assign n13961 = n13960 ^ n5831 ^ n1759 ;
  assign n13966 = n13965 ^ n13963 ^ n13961 ;
  assign n13967 = n8951 ^ n2681 ^ 1'b0 ;
  assign n13968 = ~n6120 & n13967 ;
  assign n13969 = n9398 ^ n8772 ^ n1089 ;
  assign n13970 = n4518 ^ n3340 ^ 1'b0 ;
  assign n13971 = n6338 & ~n11987 ;
  assign n13972 = n307 | n8432 ;
  assign n13973 = n13972 ^ n3984 ^ 1'b0 ;
  assign n13974 = n13973 ^ n5338 ^ n3158 ;
  assign n13975 = n13441 & ~n13974 ;
  assign n13976 = n12497 & n13975 ;
  assign n13977 = n6193 & ~n12329 ;
  assign n13978 = ( n758 & n1571 ) | ( n758 & ~n13977 ) | ( n1571 & ~n13977 ) ;
  assign n13979 = ( n958 & n3303 ) | ( n958 & ~n6879 ) | ( n3303 & ~n6879 ) ;
  assign n13980 = n6294 & ~n11651 ;
  assign n13981 = n13980 ^ n10459 ^ 1'b0 ;
  assign n13982 = ~n13979 & n13981 ;
  assign n13983 = n2847 | n13815 ;
  assign n13984 = n3267 & ~n13983 ;
  assign n13985 = n4096 ^ n1173 ^ 1'b0 ;
  assign n13986 = n13984 | n13985 ;
  assign n13987 = n13986 ^ n2402 ^ 1'b0 ;
  assign n13988 = n9502 | n13987 ;
  assign n13989 = ( n986 & ~n5900 ) | ( n986 & n13988 ) | ( ~n5900 & n13988 ) ;
  assign n13990 = n3235 & ~n13989 ;
  assign n13991 = n3900 | n12603 ;
  assign n13992 = n13991 ^ n4959 ^ 1'b0 ;
  assign n13993 = ( n1317 & n3857 ) | ( n1317 & n13701 ) | ( n3857 & n13701 ) ;
  assign n13994 = n13993 ^ n2315 ^ 1'b0 ;
  assign n13995 = n9103 & ~n13994 ;
  assign n13996 = n13995 ^ n13991 ^ 1'b0 ;
  assign n13997 = n6273 ^ n2833 ^ 1'b0 ;
  assign n13998 = n13997 ^ n7528 ^ 1'b0 ;
  assign n13999 = n6819 & n13998 ;
  assign n14000 = n349 | n13999 ;
  assign n14001 = x114 & n9216 ;
  assign n14002 = ( n11588 & n11791 ) | ( n11588 & ~n14001 ) | ( n11791 & ~n14001 ) ;
  assign n14003 = n6461 ^ n4946 ^ n3152 ;
  assign n14004 = n14003 ^ n13187 ^ n1554 ;
  assign n14005 = ( n6517 & n6635 ) | ( n6517 & ~n8084 ) | ( n6635 & ~n8084 ) ;
  assign n14006 = n3504 & ~n4774 ;
  assign n14007 = n14006 ^ n3354 ^ 1'b0 ;
  assign n14008 = n14007 ^ n6359 ^ 1'b0 ;
  assign n14010 = n9552 ^ n2948 ^ n584 ;
  assign n14011 = n14010 ^ n3428 ^ 1'b0 ;
  assign n14009 = n4717 ^ n738 ^ 1'b0 ;
  assign n14012 = n14011 ^ n14009 ^ n7661 ;
  assign n14013 = n5433 | n8051 ;
  assign n14014 = n3438 & ~n8918 ;
  assign n14015 = ( n5893 & n14013 ) | ( n5893 & ~n14014 ) | ( n14013 & ~n14014 ) ;
  assign n14016 = n8113 ^ n6148 ^ 1'b0 ;
  assign n14017 = ( n2475 & n4339 ) | ( n2475 & n7186 ) | ( n4339 & n7186 ) ;
  assign n14018 = n619 & n2476 ;
  assign n14019 = n7357 & n14018 ;
  assign n14020 = x37 & ~n14019 ;
  assign n14021 = n14020 ^ n10049 ^ 1'b0 ;
  assign n14022 = n7116 ^ n2478 ^ n807 ;
  assign n14023 = n14022 ^ n10382 ^ n6121 ;
  assign n14024 = n14023 ^ n10475 ^ 1'b0 ;
  assign n14025 = n5083 | n14024 ;
  assign n14026 = n11150 ^ n6264 ^ n2785 ;
  assign n14027 = n5332 & ~n11421 ;
  assign n14028 = ~n390 & n14027 ;
  assign n14029 = n708 | n9307 ;
  assign n14030 = ( n14026 & ~n14028 ) | ( n14026 & n14029 ) | ( ~n14028 & n14029 ) ;
  assign n14031 = ( ~n3291 & n7198 ) | ( ~n3291 & n9723 ) | ( n7198 & n9723 ) ;
  assign n14033 = ( n242 & n3748 ) | ( n242 & ~n3798 ) | ( n3748 & ~n3798 ) ;
  assign n14034 = n14033 ^ n7404 ^ n2822 ;
  assign n14035 = n14034 ^ n9798 ^ 1'b0 ;
  assign n14032 = n2671 & ~n10599 ;
  assign n14036 = n14035 ^ n14032 ^ 1'b0 ;
  assign n14037 = n3853 ^ n721 ^ n207 ;
  assign n14038 = n9047 | n14037 ;
  assign n14039 = n8170 | n14038 ;
  assign n14040 = n7732 ^ n6797 ^ 1'b0 ;
  assign n14041 = n7484 | n14040 ;
  assign n14042 = n14041 ^ n5956 ^ n2283 ;
  assign n14043 = ( n1527 & ~n2130 ) | ( n1527 & n3160 ) | ( ~n2130 & n3160 ) ;
  assign n14044 = n14043 ^ n12297 ^ 1'b0 ;
  assign n14045 = n4367 ^ n2153 ^ 1'b0 ;
  assign n14046 = ( ~n2390 & n4251 ) | ( ~n2390 & n14045 ) | ( n4251 & n14045 ) ;
  assign n14047 = n6193 | n9237 ;
  assign n14048 = n6475 ^ n4982 ^ n178 ;
  assign n14049 = n5679 & n8208 ;
  assign n14050 = ~n14048 & n14049 ;
  assign n14051 = n9053 ^ n5736 ^ x83 ;
  assign n14052 = n5995 ^ n4894 ^ 1'b0 ;
  assign n14053 = ~n2894 & n14052 ;
  assign n14054 = n14053 ^ n1116 ^ 1'b0 ;
  assign n14055 = n1966 & n14054 ;
  assign n14056 = ~n2373 & n14055 ;
  assign n14057 = n14056 ^ n8545 ^ 1'b0 ;
  assign n14058 = n9569 ^ n6877 ^ n2896 ;
  assign n14059 = ~n6140 & n14058 ;
  assign n14060 = n14059 ^ n394 ^ 1'b0 ;
  assign n14061 = ( n14051 & n14057 ) | ( n14051 & n14060 ) | ( n14057 & n14060 ) ;
  assign n14062 = n10316 ^ n6422 ^ 1'b0 ;
  assign n14063 = n14062 ^ n12970 ^ n9838 ;
  assign n14069 = ( ~n5396 & n5714 ) | ( ~n5396 & n11814 ) | ( n5714 & n11814 ) ;
  assign n14064 = ~n1696 & n6075 ;
  assign n14065 = n14064 ^ n7936 ^ n6541 ;
  assign n14066 = n2160 & ~n2509 ;
  assign n14067 = n14066 ^ n3332 ^ 1'b0 ;
  assign n14068 = n14065 | n14067 ;
  assign n14070 = n14069 ^ n14068 ^ n9284 ;
  assign n14071 = ( n863 & ~n6018 ) | ( n863 & n6770 ) | ( ~n6018 & n6770 ) ;
  assign n14072 = n14071 ^ n5332 ^ n4023 ;
  assign n14073 = n3314 & ~n13433 ;
  assign n14074 = n4497 & n14073 ;
  assign n14076 = n7792 ^ n2293 ^ 1'b0 ;
  assign n14077 = n14076 ^ n13594 ^ n270 ;
  assign n14078 = n7819 & n14077 ;
  assign n14079 = n3321 & n14078 ;
  assign n14075 = n1749 | n7691 ;
  assign n14080 = n14079 ^ n14075 ^ 1'b0 ;
  assign n14081 = n2077 | n2561 ;
  assign n14082 = n1334 | n4427 ;
  assign n14083 = n14082 ^ n7049 ^ n5381 ;
  assign n14084 = n12621 | n14083 ;
  assign n14085 = n14081 | n14084 ;
  assign n14086 = n4237 | n14085 ;
  assign n14087 = n11480 ^ n3645 ^ n3323 ;
  assign n14088 = n1605 ^ n341 ^ 1'b0 ;
  assign n14089 = n6578 ^ n5128 ^ n1451 ;
  assign n14090 = n14089 ^ n10590 ^ n9672 ;
  assign n14091 = n14088 & ~n14090 ;
  assign n14094 = n4049 | n10439 ;
  assign n14093 = n1469 & n5282 ;
  assign n14095 = n14094 ^ n14093 ^ 1'b0 ;
  assign n14092 = ( ~n1182 & n5564 ) | ( ~n1182 & n12704 ) | ( n5564 & n12704 ) ;
  assign n14096 = n14095 ^ n14092 ^ n12494 ;
  assign n14098 = ( ~x93 & n1285 ) | ( ~x93 & n3242 ) | ( n1285 & n3242 ) ;
  assign n14097 = n632 | n4387 ;
  assign n14099 = n14098 ^ n14097 ^ 1'b0 ;
  assign n14100 = n4692 ^ n2563 ^ 1'b0 ;
  assign n14101 = n4908 ^ n2762 ^ n1704 ;
  assign n14102 = n14101 ^ n2440 ^ 1'b0 ;
  assign n14103 = n14100 & n14102 ;
  assign n14104 = n11680 ^ n8812 ^ 1'b0 ;
  assign n14105 = n5706 ^ n1870 ^ 1'b0 ;
  assign n14106 = n4564 ^ n2272 ^ 1'b0 ;
  assign n14107 = n14106 ^ n13899 ^ n523 ;
  assign n14108 = n6746 & ~n7726 ;
  assign n14109 = n13625 ^ n5161 ^ n4194 ;
  assign n14110 = n7636 ^ n6966 ^ 1'b0 ;
  assign n14111 = ( n14108 & ~n14109 ) | ( n14108 & n14110 ) | ( ~n14109 & n14110 ) ;
  assign n14112 = n2213 | n3780 ;
  assign n14113 = n7091 & ~n14112 ;
  assign n14114 = n14113 ^ n7863 ^ 1'b0 ;
  assign n14115 = n11344 ^ n5793 ^ 1'b0 ;
  assign n14116 = ~n5259 & n10060 ;
  assign n14117 = ( x103 & n3900 ) | ( x103 & ~n11694 ) | ( n3900 & ~n11694 ) ;
  assign n14118 = n14117 ^ n9756 ^ n6953 ;
  assign n14119 = ~n338 & n2232 ;
  assign n14120 = n14119 ^ n6733 ^ 1'b0 ;
  assign n14121 = n11346 ^ n7415 ^ n4859 ;
  assign n14122 = n6649 & ~n9789 ;
  assign n14123 = n14122 ^ n8844 ^ 1'b0 ;
  assign n14124 = n14121 | n14123 ;
  assign n14125 = n12022 ^ n6176 ^ n5867 ;
  assign n14126 = x15 & n10715 ;
  assign n14127 = n14126 ^ n5240 ^ 1'b0 ;
  assign n14128 = n14127 ^ n11369 ^ n5095 ;
  assign n14129 = n14128 ^ n12853 ^ n4712 ;
  assign n14130 = n13239 ^ n12159 ^ n12154 ;
  assign n14131 = n734 & ~n2891 ;
  assign n14132 = n14131 ^ n1554 ^ 1'b0 ;
  assign n14133 = n3637 | n12593 ;
  assign n14134 = n14132 & ~n14133 ;
  assign n14135 = n241 | n8573 ;
  assign n14136 = ~n2999 & n4472 ;
  assign n14137 = n6330 ^ x77 ^ 1'b0 ;
  assign n14138 = ( n1626 & n14136 ) | ( n1626 & n14137 ) | ( n14136 & n14137 ) ;
  assign n14139 = n3542 ^ n3224 ^ n1396 ;
  assign n14140 = n1770 & ~n11687 ;
  assign n14141 = n2947 & n9231 ;
  assign n14142 = n14140 & ~n14141 ;
  assign n14143 = ( n5609 & n5714 ) | ( n5609 & n14142 ) | ( n5714 & n14142 ) ;
  assign n14144 = n6271 | n10156 ;
  assign n14145 = ~n12311 & n14144 ;
  assign n14146 = ~n12285 & n14145 ;
  assign n14147 = n14146 ^ n6495 ^ 1'b0 ;
  assign n14148 = n3984 & n7421 ;
  assign n14149 = n14148 ^ n7641 ^ 1'b0 ;
  assign n14150 = n14149 ^ n10962 ^ n6294 ;
  assign n14151 = ( ~n3546 & n5004 ) | ( ~n3546 & n14150 ) | ( n5004 & n14150 ) ;
  assign n14152 = n14147 & ~n14151 ;
  assign n14153 = n14152 ^ n826 ^ 1'b0 ;
  assign n14154 = n6503 ^ n3971 ^ 1'b0 ;
  assign n14155 = ( n1212 & n2396 ) | ( n1212 & ~n3625 ) | ( n2396 & ~n3625 ) ;
  assign n14156 = ( n295 & n11537 ) | ( n295 & ~n14155 ) | ( n11537 & ~n14155 ) ;
  assign n14157 = n14149 ^ n6317 ^ n153 ;
  assign n14158 = n14157 ^ n8439 ^ n3738 ;
  assign n14159 = n14158 ^ n8611 ^ n4491 ;
  assign n14160 = n3664 | n14159 ;
  assign n14161 = n8314 ^ n1201 ^ 1'b0 ;
  assign n14162 = n10785 & n14161 ;
  assign n14163 = n9881 ^ n2429 ^ 1'b0 ;
  assign n14164 = n14162 & ~n14163 ;
  assign n14165 = ( n4182 & ~n10675 ) | ( n4182 & n14164 ) | ( ~n10675 & n14164 ) ;
  assign n14166 = n6198 ^ n274 ^ 1'b0 ;
  assign n14167 = n7157 & ~n14166 ;
  assign n14168 = n11181 ^ n2572 ^ 1'b0 ;
  assign n14169 = n1883 & ~n14168 ;
  assign n14170 = ( n754 & ~n5122 ) | ( n754 & n12910 ) | ( ~n5122 & n12910 ) ;
  assign n14171 = n14170 ^ n9963 ^ n1947 ;
  assign n14172 = n3040 ^ n2688 ^ 1'b0 ;
  assign n14173 = n14172 ^ n10875 ^ 1'b0 ;
  assign n14176 = ~n4006 & n9957 ;
  assign n14177 = n3166 & ~n14176 ;
  assign n14178 = ~n2662 & n10408 ;
  assign n14179 = ~n14177 & n14178 ;
  assign n14174 = n8929 | n9627 ;
  assign n14175 = n14174 ^ n5532 ^ 1'b0 ;
  assign n14180 = n14179 ^ n14175 ^ n6706 ;
  assign n14183 = ~n2197 & n9902 ;
  assign n14181 = ~n5088 & n13214 ;
  assign n14182 = n14181 ^ n11984 ^ 1'b0 ;
  assign n14184 = n14183 ^ n14182 ^ 1'b0 ;
  assign n14185 = ( ~n356 & n7848 ) | ( ~n356 & n10327 ) | ( n7848 & n10327 ) ;
  assign n14189 = n332 & n3152 ;
  assign n14190 = ~n6559 & n14189 ;
  assign n14186 = ~n2188 & n9471 ;
  assign n14187 = n1848 & n14186 ;
  assign n14188 = n14187 ^ n14122 ^ n9465 ;
  assign n14191 = n14190 ^ n14188 ^ 1'b0 ;
  assign n14192 = ~n14185 & n14191 ;
  assign n14193 = n2539 & n4839 ;
  assign n14194 = ~n7717 & n14193 ;
  assign n14195 = ( n1407 & n2071 ) | ( n1407 & ~n12755 ) | ( n2071 & ~n12755 ) ;
  assign n14196 = n8478 & ~n9827 ;
  assign n14197 = n9951 ^ n3142 ^ 1'b0 ;
  assign n14198 = n3325 | n13001 ;
  assign n14199 = n11816 | n14198 ;
  assign n14200 = n11585 & ~n14199 ;
  assign n14201 = n184 | n6510 ;
  assign n14202 = n3768 & ~n10886 ;
  assign n14203 = n4049 | n7555 ;
  assign n14204 = n10911 & ~n14203 ;
  assign n14205 = n14204 ^ n1317 ^ n328 ;
  assign n14206 = n4457 & ~n11747 ;
  assign n14207 = ( ~n4705 & n8239 ) | ( ~n4705 & n14206 ) | ( n8239 & n14206 ) ;
  assign n14208 = ( ~n942 & n5326 ) | ( ~n942 & n11896 ) | ( n5326 & n11896 ) ;
  assign n14210 = x20 & ~n5230 ;
  assign n14211 = n6086 ^ x76 ^ 1'b0 ;
  assign n14212 = n7395 & ~n14211 ;
  assign n14213 = ~n14210 & n14212 ;
  assign n14209 = n3738 & n4506 ;
  assign n14214 = n14213 ^ n14209 ^ 1'b0 ;
  assign n14215 = n2118 & n2402 ;
  assign n14216 = ~x14 & n14215 ;
  assign n14217 = n14216 ^ n3418 ^ 1'b0 ;
  assign n14218 = n6074 & n7462 ;
  assign n14219 = n14218 ^ n11747 ^ n9097 ;
  assign n14220 = n2790 | n5099 ;
  assign n14221 = n1511 & ~n14220 ;
  assign n14222 = n6439 & ~n14221 ;
  assign n14223 = n12259 & n14222 ;
  assign n14226 = n1936 | n2113 ;
  assign n14227 = n14226 ^ n11320 ^ 1'b0 ;
  assign n14224 = n3246 | n10231 ;
  assign n14225 = n6607 | n14224 ;
  assign n14228 = n14227 ^ n14225 ^ n3230 ;
  assign n14229 = n5766 & n11478 ;
  assign n14230 = n5147 & n14229 ;
  assign n14231 = n5664 | n14230 ;
  assign n14232 = n8908 & ~n14231 ;
  assign n14233 = n13477 ^ n1131 ^ 1'b0 ;
  assign n14234 = n14232 & ~n14233 ;
  assign n14235 = n2536 ^ n2246 ^ n1674 ;
  assign n14236 = n862 & n5108 ;
  assign n14237 = ( n6194 & n8915 ) | ( n6194 & n14236 ) | ( n8915 & n14236 ) ;
  assign n14238 = ( n6780 & n14235 ) | ( n6780 & n14237 ) | ( n14235 & n14237 ) ;
  assign n14239 = n14238 ^ n10051 ^ 1'b0 ;
  assign n14240 = n2149 | n10022 ;
  assign n14241 = n14240 ^ n13445 ^ 1'b0 ;
  assign n14242 = n11480 ^ n1310 ^ 1'b0 ;
  assign n14243 = ~n2805 & n14242 ;
  assign n14244 = n6858 & n14243 ;
  assign n14245 = n14244 ^ n7306 ^ n3636 ;
  assign n14246 = ( n2463 & ~n3666 ) | ( n2463 & n6249 ) | ( ~n3666 & n6249 ) ;
  assign n14247 = n2632 ^ n1889 ^ 1'b0 ;
  assign n14248 = n14247 ^ n9048 ^ 1'b0 ;
  assign n14249 = n2903 ^ n2239 ^ n2182 ;
  assign n14250 = ~n2025 & n14249 ;
  assign n14251 = n5275 ^ n5218 ^ n289 ;
  assign n14252 = ( n2178 & n10216 ) | ( n2178 & ~n10308 ) | ( n10216 & ~n10308 ) ;
  assign n14253 = ( n852 & n14251 ) | ( n852 & n14252 ) | ( n14251 & n14252 ) ;
  assign n14254 = n14253 ^ n8975 ^ 1'b0 ;
  assign n14255 = n520 & ~n14254 ;
  assign n14256 = ~n7132 & n14255 ;
  assign n14257 = ~n1798 & n14256 ;
  assign n14258 = n650 & ~n14257 ;
  assign n14259 = n12258 ^ n7251 ^ n485 ;
  assign n14260 = n14259 ^ n9220 ^ n604 ;
  assign n14261 = ( n6040 & ~n13643 ) | ( n6040 & n14260 ) | ( ~n13643 & n14260 ) ;
  assign n14262 = n14261 ^ n3176 ^ 1'b0 ;
  assign n14263 = x79 & n14262 ;
  assign n14264 = n4529 | n12309 ;
  assign n14265 = ~n2072 & n4976 ;
  assign n14266 = n14265 ^ n3569 ^ 1'b0 ;
  assign n14267 = ( n3004 & ~n11871 ) | ( n3004 & n14266 ) | ( ~n11871 & n14266 ) ;
  assign n14268 = n3181 ^ n1165 ^ 1'b0 ;
  assign n14269 = n2463 & n14268 ;
  assign n14270 = n131 & n3864 ;
  assign n14271 = ~n12044 & n14270 ;
  assign n14272 = n14271 ^ n9331 ^ 1'b0 ;
  assign n14273 = n1372 | n14272 ;
  assign n14274 = n2329 | n14273 ;
  assign n14275 = n3232 | n14274 ;
  assign n14276 = n1139 & n9850 ;
  assign n14277 = n13539 ^ n1438 ^ 1'b0 ;
  assign n14279 = n4887 ^ n2023 ^ 1'b0 ;
  assign n14278 = n2776 & ~n3724 ;
  assign n14280 = n14279 ^ n14278 ^ 1'b0 ;
  assign n14281 = n381 | n3200 ;
  assign n14282 = n595 | n12501 ;
  assign n14283 = n2609 ^ n1566 ^ 1'b0 ;
  assign n14284 = n10036 ^ n7795 ^ 1'b0 ;
  assign n14285 = n2851 ^ n474 ^ n174 ;
  assign n14286 = n14285 ^ n11031 ^ 1'b0 ;
  assign n14287 = n14284 & ~n14286 ;
  assign n14288 = ( n420 & n1797 ) | ( n420 & n14287 ) | ( n1797 & n14287 ) ;
  assign n14289 = n4508 ^ n1201 ^ 1'b0 ;
  assign n14290 = n14289 ^ n6322 ^ n1553 ;
  assign n14291 = n14290 ^ n13370 ^ 1'b0 ;
  assign n14292 = n2222 ^ n1385 ^ n1332 ;
  assign n14293 = n14292 ^ n3620 ^ 1'b0 ;
  assign n14294 = n3343 | n14293 ;
  assign n14295 = n2681 & n12350 ;
  assign n14300 = n6759 ^ n6455 ^ 1'b0 ;
  assign n14301 = n5714 | n14300 ;
  assign n14296 = n6012 & n8730 ;
  assign n14297 = n14296 ^ n2242 ^ 1'b0 ;
  assign n14298 = n14297 ^ n11649 ^ 1'b0 ;
  assign n14299 = n8411 & ~n14298 ;
  assign n14302 = n14301 ^ n14299 ^ 1'b0 ;
  assign n14303 = n9955 ^ n5448 ^ n3148 ;
  assign n14304 = n1636 & n11748 ;
  assign n14305 = n13747 | n13825 ;
  assign n14306 = n889 | n14305 ;
  assign n14307 = n5133 ^ n3946 ^ 1'b0 ;
  assign n14308 = n4201 ^ n3046 ^ n218 ;
  assign n14309 = ~n1573 & n14308 ;
  assign n14310 = n14309 ^ n12752 ^ 1'b0 ;
  assign n14311 = n14310 ^ n1137 ^ 1'b0 ;
  assign n14312 = n6619 ^ n1939 ^ 1'b0 ;
  assign n14313 = ~n6309 & n14312 ;
  assign n14314 = ( n3438 & ~n3630 ) | ( n3438 & n14313 ) | ( ~n3630 & n14313 ) ;
  assign n14315 = n14314 ^ n4591 ^ 1'b0 ;
  assign n14316 = ( n2884 & n11328 ) | ( n2884 & n13233 ) | ( n11328 & n13233 ) ;
  assign n14317 = n3330 | n4397 ;
  assign n14324 = n10812 ^ n3599 ^ n2127 ;
  assign n14318 = n9081 ^ n2688 ^ n1666 ;
  assign n14319 = n6657 | n7233 ;
  assign n14320 = n14318 & ~n14319 ;
  assign n14321 = n2638 & n4234 ;
  assign n14322 = n14320 & n14321 ;
  assign n14323 = n11886 | n14322 ;
  assign n14325 = n14324 ^ n14323 ^ 1'b0 ;
  assign n14326 = n3951 ^ n3341 ^ n1054 ;
  assign n14327 = n2451 & ~n14326 ;
  assign n14328 = ~n14325 & n14327 ;
  assign n14329 = n14328 ^ n12836 ^ 1'b0 ;
  assign n14330 = n4371 ^ n2438 ^ n658 ;
  assign n14331 = x57 | n8198 ;
  assign n14332 = n6882 ^ n6625 ^ 1'b0 ;
  assign n14333 = n14331 & n14332 ;
  assign n14334 = ( n12001 & ~n14330 ) | ( n12001 & n14333 ) | ( ~n14330 & n14333 ) ;
  assign n14335 = n6267 ^ n1789 ^ 1'b0 ;
  assign n14336 = n4041 | n14335 ;
  assign n14337 = n10103 ^ n9105 ^ 1'b0 ;
  assign n14338 = n11212 & ~n14337 ;
  assign n14339 = n14338 ^ n4694 ^ 1'b0 ;
  assign n14340 = ~n9037 & n14339 ;
  assign n14348 = n2969 ^ n870 ^ 1'b0 ;
  assign n14341 = ( n5402 & n8158 ) | ( n5402 & n11270 ) | ( n8158 & n11270 ) ;
  assign n14343 = n545 ^ n492 ^ 1'b0 ;
  assign n14344 = ~n1252 & n14343 ;
  assign n14345 = n4304 & n14344 ;
  assign n14342 = n9901 ^ n4636 ^ 1'b0 ;
  assign n14346 = n14345 ^ n14342 ^ 1'b0 ;
  assign n14347 = ( n392 & n14341 ) | ( n392 & ~n14346 ) | ( n14341 & ~n14346 ) ;
  assign n14349 = n14348 ^ n14347 ^ n11072 ;
  assign n14350 = n2797 & n6248 ;
  assign n14351 = n9526 & ~n14350 ;
  assign n14352 = n2365 & n12176 ;
  assign n14353 = n7591 & ~n13849 ;
  assign n14354 = n984 & n1445 ;
  assign n14355 = n14354 ^ n4782 ^ 1'b0 ;
  assign n14356 = n5492 ^ n3473 ^ n2996 ;
  assign n14357 = n981 & ~n14356 ;
  assign n14358 = n6053 & n14357 ;
  assign n14360 = n12490 ^ n9183 ^ n6449 ;
  assign n14359 = x50 & ~n5485 ;
  assign n14361 = n14360 ^ n14359 ^ 1'b0 ;
  assign n14362 = ~n708 & n3186 ;
  assign n14363 = n14362 ^ n7094 ^ 1'b0 ;
  assign n14364 = ~n14361 & n14363 ;
  assign n14365 = n5347 ^ n4123 ^ 1'b0 ;
  assign n14366 = n12928 & n14365 ;
  assign n14369 = n10271 ^ n6596 ^ 1'b0 ;
  assign n14367 = n6699 ^ n4106 ^ 1'b0 ;
  assign n14368 = n7189 | n14367 ;
  assign n14370 = n14369 ^ n14368 ^ 1'b0 ;
  assign n14378 = n8630 ^ n2017 ^ 1'b0 ;
  assign n14379 = n10979 & n14378 ;
  assign n14376 = ~n5647 & n6439 ;
  assign n14374 = ( ~n2331 & n6159 ) | ( ~n2331 & n12001 ) | ( n6159 & n12001 ) ;
  assign n14371 = n6473 | n7162 ;
  assign n14372 = n940 & ~n14371 ;
  assign n14373 = n5049 | n14372 ;
  assign n14375 = n14374 ^ n14373 ^ 1'b0 ;
  assign n14377 = n14376 ^ n14375 ^ n9111 ;
  assign n14380 = n14379 ^ n14377 ^ 1'b0 ;
  assign n14381 = n6642 & ~n7116 ;
  assign n14382 = n7040 & ~n14381 ;
  assign n14383 = n14382 ^ n9161 ^ n7657 ;
  assign n14384 = ( n5257 & ~n5458 ) | ( n5257 & n13165 ) | ( ~n5458 & n13165 ) ;
  assign n14385 = n3826 ^ n1126 ^ 1'b0 ;
  assign n14386 = ~n13698 & n14385 ;
  assign n14391 = n7038 ^ n2768 ^ n1601 ;
  assign n14392 = ~n12943 & n14391 ;
  assign n14387 = n760 | n8839 ;
  assign n14388 = n14387 ^ n2292 ^ 1'b0 ;
  assign n14389 = n14388 ^ n7913 ^ n3265 ;
  assign n14390 = n11689 | n14389 ;
  assign n14393 = n14392 ^ n14390 ^ 1'b0 ;
  assign n14394 = n3811 & ~n13262 ;
  assign n14395 = n12252 ^ n7914 ^ 1'b0 ;
  assign n14396 = n9307 ^ n1514 ^ 1'b0 ;
  assign n14397 = n1111 | n14396 ;
  assign n14398 = n8772 & ~n9528 ;
  assign n14399 = n6590 & n14398 ;
  assign n14400 = n14399 ^ n3731 ^ 1'b0 ;
  assign n14401 = n6482 & n14400 ;
  assign n14402 = n14401 ^ n4775 ^ 1'b0 ;
  assign n14403 = n14402 ^ n8478 ^ 1'b0 ;
  assign n14404 = n13232 & ~n14403 ;
  assign n14405 = ~n10784 & n14404 ;
  assign n14406 = n9101 ^ n7620 ^ n1434 ;
  assign n14407 = ( ~n8108 & n9588 ) | ( ~n8108 & n14406 ) | ( n9588 & n14406 ) ;
  assign n14408 = n3788 | n6878 ;
  assign n14409 = n14408 ^ n5238 ^ 1'b0 ;
  assign n14410 = n5533 & n5597 ;
  assign n14411 = ( n12918 & n14409 ) | ( n12918 & ~n14410 ) | ( n14409 & ~n14410 ) ;
  assign n14412 = n3097 ^ n1519 ^ n129 ;
  assign n14413 = ( n635 & n7012 ) | ( n635 & ~n14412 ) | ( n7012 & ~n14412 ) ;
  assign n14414 = n14413 ^ n1135 ^ 1'b0 ;
  assign n14415 = n11549 & ~n13243 ;
  assign n14416 = ~n14414 & n14415 ;
  assign n14417 = ~n2296 & n14416 ;
  assign n14418 = n4653 ^ n798 ^ 1'b0 ;
  assign n14419 = n2459 | n14418 ;
  assign n14420 = n12572 | n14419 ;
  assign n14421 = n12919 | n14420 ;
  assign n14422 = n6705 ^ n388 ^ 1'b0 ;
  assign n14423 = n4579 & n14422 ;
  assign n14424 = ~n4226 & n14423 ;
  assign n14425 = n8949 ^ n717 ^ n495 ;
  assign n14426 = n14425 ^ n1691 ^ 1'b0 ;
  assign n14427 = n2093 | n14426 ;
  assign n14428 = n5868 ^ n5764 ^ n2989 ;
  assign n14429 = n14428 ^ n930 ^ 1'b0 ;
  assign n14430 = n12874 & ~n14429 ;
  assign n14431 = n13528 ^ n1162 ^ 1'b0 ;
  assign n14432 = ~n895 & n14431 ;
  assign n14433 = n14432 ^ n1666 ^ 1'b0 ;
  assign n14434 = ~n14137 & n14433 ;
  assign n14435 = n8660 & ~n11005 ;
  assign n14436 = n14435 ^ n10521 ^ 1'b0 ;
  assign n14437 = n2894 | n13011 ;
  assign n14438 = n774 & ~n5173 ;
  assign n14439 = n11933 ^ n5824 ^ 1'b0 ;
  assign n14440 = n7252 & ~n14439 ;
  assign n14448 = ~n1420 & n7760 ;
  assign n14449 = n14448 ^ n9338 ^ 1'b0 ;
  assign n14450 = ~n9675 & n14449 ;
  assign n14445 = ~n4784 & n9778 ;
  assign n14446 = n14445 ^ n874 ^ 1'b0 ;
  assign n14444 = n12063 ^ n4121 ^ 1'b0 ;
  assign n14447 = n14446 ^ n14444 ^ n8029 ;
  assign n14441 = n3935 & n6931 ;
  assign n14442 = n5545 & n14441 ;
  assign n14443 = n14442 ^ n6182 ^ 1'b0 ;
  assign n14451 = n14450 ^ n14447 ^ n14443 ;
  assign n14452 = n9564 ^ n8413 ^ n2818 ;
  assign n14453 = n9129 ^ n8657 ^ n5631 ;
  assign n14454 = n14453 ^ n6986 ^ n2212 ;
  assign n14455 = ( ~n3161 & n6888 ) | ( ~n3161 & n8039 ) | ( n6888 & n8039 ) ;
  assign n14456 = n2780 & ~n4086 ;
  assign n14457 = n2896 | n5438 ;
  assign n14458 = n1428 & ~n14457 ;
  assign n14459 = n12187 ^ n11889 ^ n451 ;
  assign n14461 = ~n456 & n3063 ;
  assign n14462 = n14461 ^ n1438 ^ 1'b0 ;
  assign n14463 = ~n3506 & n14462 ;
  assign n14460 = n8919 ^ n4052 ^ n3033 ;
  assign n14464 = n14463 ^ n14460 ^ 1'b0 ;
  assign n14465 = n641 & n3824 ;
  assign n14466 = n5661 & ~n14465 ;
  assign n14467 = n14466 ^ n14331 ^ n12133 ;
  assign n14468 = ( n4465 & ~n9541 ) | ( n4465 & n14467 ) | ( ~n9541 & n14467 ) ;
  assign n14469 = n8590 ^ n7883 ^ n3611 ;
  assign n14470 = ~n196 & n8970 ;
  assign n14471 = n14469 & n14470 ;
  assign n14472 = n6396 | n13529 ;
  assign n14473 = n12528 & ~n14472 ;
  assign n14474 = ( n888 & ~n2508 ) | ( n888 & n7774 ) | ( ~n2508 & n7774 ) ;
  assign n14475 = n14473 | n14474 ;
  assign n14476 = n14475 ^ n7293 ^ 1'b0 ;
  assign n14477 = ~n380 & n14476 ;
  assign n14478 = n2953 & n4902 ;
  assign n14479 = n14477 & n14478 ;
  assign n14480 = n3177 & ~n11288 ;
  assign n14481 = n1363 & n14480 ;
  assign n14482 = n4127 & n5234 ;
  assign n14483 = n14482 ^ n7197 ^ 1'b0 ;
  assign n14484 = n7110 | n10508 ;
  assign n14485 = n14484 ^ n3763 ^ 1'b0 ;
  assign n14486 = n14485 ^ n13503 ^ 1'b0 ;
  assign n14487 = n4912 ^ n3279 ^ 1'b0 ;
  assign n14488 = n11790 ^ n7780 ^ n2468 ;
  assign n14489 = n14488 ^ n6248 ^ 1'b0 ;
  assign n14490 = ~n7224 & n14489 ;
  assign n14491 = n14490 ^ n2067 ^ 1'b0 ;
  assign n14492 = n6338 ^ n3596 ^ n2756 ;
  assign n14493 = ~n6824 & n12663 ;
  assign n14494 = ~n4214 & n14493 ;
  assign n14495 = n14492 & n14494 ;
  assign n14496 = ( x115 & n2788 ) | ( x115 & ~n3671 ) | ( n2788 & ~n3671 ) ;
  assign n14497 = ( n4628 & n4666 ) | ( n4628 & ~n14496 ) | ( n4666 & ~n14496 ) ;
  assign n14498 = ( n4714 & n4838 ) | ( n4714 & ~n14497 ) | ( n4838 & ~n14497 ) ;
  assign n14499 = ( n2542 & n4106 ) | ( n2542 & n9406 ) | ( n4106 & n9406 ) ;
  assign n14500 = ~n7360 & n7593 ;
  assign n14501 = n9324 | n14500 ;
  assign n14502 = n11605 | n14501 ;
  assign n14503 = ~n798 & n7497 ;
  assign n14504 = ~n9729 & n14503 ;
  assign n14505 = ( n2955 & n14502 ) | ( n2955 & n14504 ) | ( n14502 & n14504 ) ;
  assign n14506 = n2271 ^ n1352 ^ n1139 ;
  assign n14507 = n14506 ^ n2108 ^ n1252 ;
  assign n14512 = n14345 ^ n13396 ^ n856 ;
  assign n14513 = ~n1425 & n14512 ;
  assign n14514 = n14513 ^ n10118 ^ 1'b0 ;
  assign n14515 = ~n4094 & n7623 ;
  assign n14516 = ~n14514 & n14515 ;
  assign n14508 = n11747 ^ n3497 ^ n2378 ;
  assign n14509 = n14508 ^ n7152 ^ 1'b0 ;
  assign n14510 = ~n5248 & n7051 ;
  assign n14511 = n14509 & n14510 ;
  assign n14517 = n14516 ^ n14511 ^ 1'b0 ;
  assign n14523 = n6822 ^ n1913 ^ 1'b0 ;
  assign n14524 = ( n208 & ~n3797 ) | ( n208 & n14523 ) | ( ~n3797 & n14523 ) ;
  assign n14525 = n8202 ^ n4033 ^ 1'b0 ;
  assign n14526 = ~n14524 & n14525 ;
  assign n14520 = n2673 ^ n315 ^ 1'b0 ;
  assign n14521 = n9230 & n14520 ;
  assign n14518 = n596 & n7985 ;
  assign n14519 = n10300 & ~n14518 ;
  assign n14522 = n14521 ^ n14519 ^ 1'b0 ;
  assign n14527 = n14526 ^ n14522 ^ n3750 ;
  assign n14528 = n5844 | n7192 ;
  assign n14529 = n14527 | n14528 ;
  assign n14530 = ~n4464 & n6031 ;
  assign n14531 = ~n7578 & n14530 ;
  assign n14532 = n14531 ^ n8970 ^ 1'b0 ;
  assign n14533 = n7668 ^ n1167 ^ 1'b0 ;
  assign n14534 = n5008 & n6559 ;
  assign n14535 = n14533 & n14534 ;
  assign n14536 = n14532 | n14535 ;
  assign n14537 = n10205 ^ n2704 ^ 1'b0 ;
  assign n14538 = n9488 | n14537 ;
  assign n14539 = ( ~n10218 & n11648 ) | ( ~n10218 & n13352 ) | ( n11648 & n13352 ) ;
  assign n14541 = n5241 ^ n1772 ^ 1'b0 ;
  assign n14542 = n14541 ^ n9880 ^ 1'b0 ;
  assign n14543 = ~n4839 & n14542 ;
  assign n14544 = n14543 ^ n11927 ^ 1'b0 ;
  assign n14545 = ~n662 & n14544 ;
  assign n14540 = n9569 & ~n11050 ;
  assign n14546 = n14545 ^ n14540 ^ 1'b0 ;
  assign n14547 = n10776 ^ n5674 ^ 1'b0 ;
  assign n14549 = ~n644 & n3052 ;
  assign n14550 = n14549 ^ n2859 ^ 1'b0 ;
  assign n14548 = n6299 ^ n3044 ^ 1'b0 ;
  assign n14551 = n14550 ^ n14548 ^ 1'b0 ;
  assign n14552 = n12456 | n14551 ;
  assign n14554 = n8796 ^ n3489 ^ 1'b0 ;
  assign n14553 = ~n628 & n14289 ;
  assign n14555 = n14554 ^ n14553 ^ 1'b0 ;
  assign n14556 = n3321 ^ n1797 ^ 1'b0 ;
  assign n14557 = x115 & n14556 ;
  assign n14558 = n3645 | n14557 ;
  assign n14559 = n2543 | n5855 ;
  assign n14560 = n14559 ^ n6256 ^ 1'b0 ;
  assign n14561 = n9811 ^ n2438 ^ n406 ;
  assign n14562 = n11453 | n14561 ;
  assign n14563 = n14562 ^ n469 ^ 1'b0 ;
  assign n14564 = n1391 | n2345 ;
  assign n14565 = ( ~n14560 & n14563 ) | ( ~n14560 & n14564 ) | ( n14563 & n14564 ) ;
  assign n14566 = n10708 ^ n8867 ^ 1'b0 ;
  assign n14567 = n13232 ^ n4555 ^ n4338 ;
  assign n14568 = n2571 & ~n13123 ;
  assign n14569 = n14567 & n14568 ;
  assign n14570 = ~n1046 & n14569 ;
  assign n14571 = ~n1818 & n2539 ;
  assign n14572 = n350 & n3629 ;
  assign n14573 = ~n2521 & n14572 ;
  assign n14574 = n3515 & ~n5897 ;
  assign n14575 = n14574 ^ n13700 ^ n3904 ;
  assign n14576 = n6122 ^ n1603 ^ 1'b0 ;
  assign n14577 = ~n4386 & n14576 ;
  assign n14578 = ( ~n5131 & n14575 ) | ( ~n5131 & n14577 ) | ( n14575 & n14577 ) ;
  assign n14579 = n14578 ^ n13564 ^ n3202 ;
  assign n14580 = n14579 ^ n9936 ^ n1922 ;
  assign n14581 = ~n1876 & n14580 ;
  assign n14582 = n14581 ^ n8032 ^ 1'b0 ;
  assign n14583 = n13334 | n14582 ;
  assign n14584 = n7376 | n14583 ;
  assign n14585 = n1898 & ~n9414 ;
  assign n14586 = ~n204 & n14585 ;
  assign n14587 = n12150 ^ n7513 ^ n2858 ;
  assign n14588 = n5713 ^ n3806 ^ 1'b0 ;
  assign n14589 = ~n12978 & n14588 ;
  assign n14590 = n7855 ^ n275 ^ 1'b0 ;
  assign n14591 = n2433 | n14590 ;
  assign n14592 = n6249 & ~n14591 ;
  assign n14593 = ~n7269 & n12879 ;
  assign n14594 = n14593 ^ n194 ^ 1'b0 ;
  assign n14595 = ( n14589 & n14592 ) | ( n14589 & n14594 ) | ( n14592 & n14594 ) ;
  assign n14596 = ( x21 & n10230 ) | ( x21 & n14522 ) | ( n10230 & n14522 ) ;
  assign n14597 = n1280 & n1670 ;
  assign n14598 = n7966 ^ n3990 ^ 1'b0 ;
  assign n14599 = n2835 & ~n14598 ;
  assign n14600 = ( n12828 & ~n14597 ) | ( n12828 & n14599 ) | ( ~n14597 & n14599 ) ;
  assign n14601 = n7347 ^ n1304 ^ 1'b0 ;
  assign n14602 = n291 | n14601 ;
  assign n14603 = n14602 ^ x114 ^ 1'b0 ;
  assign n14604 = ~n14600 & n14603 ;
  assign n14605 = ~n2472 & n9848 ;
  assign n14606 = n1004 & ~n14605 ;
  assign n14607 = n3646 ^ n1215 ^ 1'b0 ;
  assign n14608 = n9001 ^ n7006 ^ 1'b0 ;
  assign n14609 = ( n329 & n7580 ) | ( n329 & ~n7959 ) | ( n7580 & ~n7959 ) ;
  assign n14610 = n14608 & n14609 ;
  assign n14611 = n6010 & n14610 ;
  assign n14612 = n6048 ^ n5533 ^ 1'b0 ;
  assign n14613 = ( ~n10584 & n12453 ) | ( ~n10584 & n14612 ) | ( n12453 & n14612 ) ;
  assign n14614 = n13145 ^ n11928 ^ n10320 ;
  assign n14615 = n11061 ^ n5550 ^ 1'b0 ;
  assign n14616 = n7381 & ~n14615 ;
  assign n14617 = n2660 ^ n1791 ^ 1'b0 ;
  assign n14618 = n4526 & ~n14617 ;
  assign n14619 = n4956 ^ n1712 ^ 1'b0 ;
  assign n14620 = n14618 | n14619 ;
  assign n14621 = n1223 | n14620 ;
  assign n14622 = n6463 & ~n12185 ;
  assign n14623 = n173 & ~n10915 ;
  assign n14624 = n14623 ^ n1426 ^ 1'b0 ;
  assign n14625 = ~n2259 & n7213 ;
  assign n14626 = n14625 ^ n5303 ^ 1'b0 ;
  assign n14627 = ( ~n3796 & n4689 ) | ( ~n3796 & n6333 ) | ( n4689 & n6333 ) ;
  assign n14628 = n3980 | n14627 ;
  assign n14629 = n4029 & ~n14628 ;
  assign n14630 = n5353 ^ n5106 ^ n1925 ;
  assign n14631 = n4762 ^ n436 ^ 1'b0 ;
  assign n14632 = n2443 & ~n2757 ;
  assign n14633 = n14631 & n14632 ;
  assign n14634 = n14633 ^ x25 ^ 1'b0 ;
  assign n14635 = n14630 & ~n14634 ;
  assign n14636 = ( n2896 & ~n14629 ) | ( n2896 & n14635 ) | ( ~n14629 & n14635 ) ;
  assign n14637 = ~n11542 & n14636 ;
  assign n14638 = n8780 & n14637 ;
  assign n14639 = ( n3840 & n7251 ) | ( n3840 & ~n11027 ) | ( n7251 & ~n11027 ) ;
  assign n14640 = n6330 & n8538 ;
  assign n14641 = n4279 | n7702 ;
  assign n14642 = ( ~n14639 & n14640 ) | ( ~n14639 & n14641 ) | ( n14640 & n14641 ) ;
  assign n14646 = n12208 ^ n11605 ^ 1'b0 ;
  assign n14643 = n3222 ^ n1757 ^ n1612 ;
  assign n14644 = n3833 & n14643 ;
  assign n14645 = n14644 ^ n945 ^ 1'b0 ;
  assign n14647 = n14646 ^ n14645 ^ n8151 ;
  assign n14648 = n13973 ^ n13114 ^ n4342 ;
  assign n14649 = n13185 ^ n7358 ^ n858 ;
  assign n14650 = ( n808 & n1602 ) | ( n808 & n5484 ) | ( n1602 & n5484 ) ;
  assign n14651 = n2010 | n14650 ;
  assign n14652 = ( n8212 & n9665 ) | ( n8212 & n14651 ) | ( n9665 & n14651 ) ;
  assign n14653 = n3704 & n6503 ;
  assign n14654 = n960 & n14653 ;
  assign n14655 = n14654 ^ n8424 ^ n5993 ;
  assign n14657 = ( x120 & n171 ) | ( x120 & n4400 ) | ( n171 & n4400 ) ;
  assign n14658 = n11996 ^ n6272 ^ 1'b0 ;
  assign n14659 = n14657 & n14658 ;
  assign n14656 = ~n584 & n10079 ;
  assign n14660 = n14659 ^ n14656 ^ 1'b0 ;
  assign n14661 = ( n6301 & ~n12723 ) | ( n6301 & n14660 ) | ( ~n12723 & n14660 ) ;
  assign n14663 = n9762 ^ n1929 ^ 1'b0 ;
  assign n14664 = n1527 & ~n14663 ;
  assign n14662 = n13194 ^ n12088 ^ 1'b0 ;
  assign n14665 = n14664 ^ n14662 ^ n8211 ;
  assign n14666 = n8865 ^ n8318 ^ n4390 ;
  assign n14667 = n14666 ^ n13936 ^ 1'b0 ;
  assign n14668 = x1 & n14667 ;
  assign n14671 = n9037 ^ n5266 ^ 1'b0 ;
  assign n14672 = ~n4591 & n14671 ;
  assign n14669 = n5122 ^ n3426 ^ 1'b0 ;
  assign n14670 = n5960 | n14669 ;
  assign n14673 = n14672 ^ n14670 ^ n11544 ;
  assign n14674 = ( n3741 & ~n14668 ) | ( n3741 & n14673 ) | ( ~n14668 & n14673 ) ;
  assign n14675 = ~n1337 & n12787 ;
  assign n14676 = n14675 ^ n7701 ^ 1'b0 ;
  assign n14677 = ( n1600 & n3230 ) | ( n1600 & ~n14331 ) | ( n3230 & ~n14331 ) ;
  assign n14678 = n14677 ^ n1253 ^ 1'b0 ;
  assign n14679 = n12767 & ~n14678 ;
  assign n14680 = n14679 ^ n9744 ^ 1'b0 ;
  assign n14681 = n7599 ^ n3065 ^ 1'b0 ;
  assign n14682 = n9243 & ~n14681 ;
  assign n14683 = n14682 ^ n8086 ^ n5929 ;
  assign n14684 = n9594 | n14683 ;
  assign n14685 = n6415 ^ n3689 ^ 1'b0 ;
  assign n14686 = n3135 | n14685 ;
  assign n14687 = n11678 ^ n10622 ^ 1'b0 ;
  assign n14688 = n2884 | n4705 ;
  assign n14689 = n14688 ^ n6256 ^ 1'b0 ;
  assign n14690 = n14689 ^ n8007 ^ n5507 ;
  assign n14691 = n7813 ^ n3124 ^ 1'b0 ;
  assign n14692 = n2752 & n14691 ;
  assign n14693 = n3625 & n14692 ;
  assign n14694 = ( n6583 & n6652 ) | ( n6583 & ~n7119 ) | ( n6652 & ~n7119 ) ;
  assign n14695 = n3114 & ~n13147 ;
  assign n14696 = n14361 ^ n5868 ^ 1'b0 ;
  assign n14697 = ( n4727 & n6570 ) | ( n4727 & ~n9249 ) | ( n6570 & ~n9249 ) ;
  assign n14698 = n13354 | n14697 ;
  assign n14699 = n14698 ^ n4684 ^ 1'b0 ;
  assign n14700 = n10398 ^ n3502 ^ 1'b0 ;
  assign n14701 = n4557 | n14700 ;
  assign n14702 = n8655 & ~n14701 ;
  assign n14703 = n14702 ^ n13813 ^ 1'b0 ;
  assign n14704 = n635 & ~n14703 ;
  assign n14705 = ( n5017 & n5177 ) | ( n5017 & ~n11626 ) | ( n5177 & ~n11626 ) ;
  assign n14706 = n14705 ^ n3037 ^ n2242 ;
  assign n14707 = n11117 ^ n10004 ^ n5495 ;
  assign n14708 = ~n6145 & n11837 ;
  assign n14709 = n1385 & n14708 ;
  assign n14710 = n14709 ^ n11319 ^ 1'b0 ;
  assign n14711 = ~n2211 & n14710 ;
  assign n14712 = ~n7427 & n9964 ;
  assign n14713 = n14712 ^ n4177 ^ 1'b0 ;
  assign n14714 = n6754 ^ n812 ^ 1'b0 ;
  assign n14715 = n1035 & n14714 ;
  assign n14716 = n14715 ^ n11349 ^ n10263 ;
  assign n14718 = n846 ^ x78 ^ 1'b0 ;
  assign n14719 = ~n1252 & n14718 ;
  assign n14717 = n5956 & ~n10593 ;
  assign n14720 = n14719 ^ n14717 ^ 1'b0 ;
  assign n14723 = n10371 ^ n4739 ^ n2102 ;
  assign n14724 = ( n8582 & n10271 ) | ( n8582 & n14723 ) | ( n10271 & n14723 ) ;
  assign n14721 = ~n2378 & n11651 ;
  assign n14722 = ~n1267 & n14721 ;
  assign n14725 = n14724 ^ n14722 ^ n3410 ;
  assign n14726 = n3598 ^ n1154 ^ n869 ;
  assign n14727 = n9757 ^ n2500 ^ 1'b0 ;
  assign n14728 = n14726 | n14727 ;
  assign n14729 = n6100 ^ n3307 ^ 1'b0 ;
  assign n14730 = ~n14728 & n14729 ;
  assign n14731 = n8460 ^ n5866 ^ 1'b0 ;
  assign n14732 = n14366 & ~n14731 ;
  assign n14733 = n6093 & n14732 ;
  assign n14735 = n8113 & ~n9789 ;
  assign n14736 = n14735 ^ n10788 ^ n2557 ;
  assign n14734 = n3718 ^ n2112 ^ n872 ;
  assign n14737 = n14736 ^ n14734 ^ 1'b0 ;
  assign n14738 = n5969 ^ n5122 ^ n2499 ;
  assign n14739 = ( n1357 & n13073 ) | ( n1357 & n14738 ) | ( n13073 & n14738 ) ;
  assign n14740 = n6853 ^ n5748 ^ n3994 ;
  assign n14741 = n4187 & n14740 ;
  assign n14742 = n6415 & n14741 ;
  assign n14745 = n6886 & ~n8842 ;
  assign n14743 = ( ~n2063 & n7151 ) | ( ~n2063 & n8196 ) | ( n7151 & n8196 ) ;
  assign n14744 = n5723 | n14743 ;
  assign n14746 = n14745 ^ n14744 ^ 1'b0 ;
  assign n14747 = n14746 ^ n2447 ^ 1'b0 ;
  assign n14748 = n14747 ^ n9033 ^ n835 ;
  assign n14757 = ~n3393 & n5325 ;
  assign n14754 = n7459 & ~n13882 ;
  assign n14755 = n3396 & n14754 ;
  assign n14753 = ~n3799 & n9251 ;
  assign n14756 = n14755 ^ n14753 ^ 1'b0 ;
  assign n14749 = ( x75 & n815 ) | ( x75 & ~n1761 ) | ( n815 & ~n1761 ) ;
  assign n14750 = n14749 ^ n4804 ^ n4727 ;
  assign n14751 = ~n10219 & n14750 ;
  assign n14752 = ( x56 & n3065 ) | ( x56 & ~n14751 ) | ( n3065 & ~n14751 ) ;
  assign n14758 = n14757 ^ n14756 ^ n14752 ;
  assign n14759 = n12916 ^ n5157 ^ 1'b0 ;
  assign n14760 = n2273 & ~n14759 ;
  assign n14761 = n11464 ^ n4086 ^ 1'b0 ;
  assign n14762 = n1184 | n4961 ;
  assign n14763 = n14762 ^ n993 ^ 1'b0 ;
  assign n14764 = n10364 ^ n5566 ^ 1'b0 ;
  assign n14765 = n2527 & n3964 ;
  assign n14766 = n10586 ^ n8597 ^ 1'b0 ;
  assign n14767 = n10785 & ~n14766 ;
  assign n14768 = ( n8099 & n12948 ) | ( n8099 & n14767 ) | ( n12948 & n14767 ) ;
  assign n14769 = n3701 | n4598 ;
  assign n14770 = ( ~n1448 & n9501 ) | ( ~n1448 & n14769 ) | ( n9501 & n14769 ) ;
  assign n14771 = x31 & ~n3938 ;
  assign n14772 = n416 & n14771 ;
  assign n14773 = ~n5313 & n14772 ;
  assign n14774 = n6447 & ~n14773 ;
  assign n14778 = ( n2496 & n3806 ) | ( n2496 & ~n8084 ) | ( n3806 & ~n8084 ) ;
  assign n14775 = n2041 ^ n255 ^ x11 ;
  assign n14776 = n14775 ^ n2629 ^ 1'b0 ;
  assign n14777 = ( ~n7795 & n12505 ) | ( ~n7795 & n14776 ) | ( n12505 & n14776 ) ;
  assign n14779 = n14778 ^ n14777 ^ n9775 ;
  assign n14780 = n12073 & ~n13427 ;
  assign n14781 = n14780 ^ n6296 ^ 1'b0 ;
  assign n14782 = ~n7998 & n11009 ;
  assign n14783 = n14782 ^ n2342 ^ 1'b0 ;
  assign n14784 = n1076 | n4658 ;
  assign n14785 = n14784 ^ n5615 ^ n3194 ;
  assign n14786 = n12454 | n14785 ;
  assign n14787 = n14786 ^ n256 ^ 1'b0 ;
  assign n14788 = n14787 ^ n9741 ^ 1'b0 ;
  assign n14789 = n14320 | n14788 ;
  assign n14790 = n13781 ^ n8661 ^ 1'b0 ;
  assign n14791 = ( ~n1278 & n11868 ) | ( ~n1278 & n14790 ) | ( n11868 & n14790 ) ;
  assign n14796 = n7832 ^ n6231 ^ 1'b0 ;
  assign n14794 = n226 & ~n7770 ;
  assign n14795 = n14794 ^ n6861 ^ n3238 ;
  assign n14792 = ~n3051 & n7361 ;
  assign n14793 = n14792 ^ n5686 ^ 1'b0 ;
  assign n14797 = n14796 ^ n14795 ^ n14793 ;
  assign n14798 = x7 & ~n4705 ;
  assign n14799 = n14798 ^ n12043 ^ 1'b0 ;
  assign n14800 = n3668 | n14799 ;
  assign n14801 = n2748 ^ n1581 ^ 1'b0 ;
  assign n14802 = ~n1286 & n11481 ;
  assign n14803 = n10679 | n14425 ;
  assign n14804 = n1057 & ~n14803 ;
  assign n14805 = n8626 ^ n8342 ^ 1'b0 ;
  assign n14806 = n5421 & n14805 ;
  assign n14807 = n14806 ^ n1019 ^ 1'b0 ;
  assign n14808 = ( n4661 & n4784 ) | ( n4661 & n14807 ) | ( n4784 & n14807 ) ;
  assign n14809 = x83 & n14808 ;
  assign n14810 = ~n1932 & n8669 ;
  assign n14811 = n14810 ^ n9157 ^ 1'b0 ;
  assign n14812 = n4508 ^ n4127 ^ n2154 ;
  assign n14813 = n14812 ^ n6632 ^ 1'b0 ;
  assign n14814 = ( n8039 & n13674 ) | ( n8039 & n14813 ) | ( n13674 & n14813 ) ;
  assign n14815 = n14814 ^ n8441 ^ 1'b0 ;
  assign n14816 = ( ~n586 & n3321 ) | ( ~n586 & n14815 ) | ( n3321 & n14815 ) ;
  assign n14819 = n7990 & n13133 ;
  assign n14817 = n4830 & n7903 ;
  assign n14818 = n14817 ^ n9147 ^ 1'b0 ;
  assign n14820 = n14819 ^ n14818 ^ 1'b0 ;
  assign n14821 = n1543 & n5461 ;
  assign n14822 = n3703 & n14821 ;
  assign n14823 = n10601 ^ n1927 ^ 1'b0 ;
  assign n14824 = n14822 | n14823 ;
  assign n14825 = n7762 ^ n1286 ^ 1'b0 ;
  assign n14826 = n869 & n14825 ;
  assign n14827 = n8008 ^ n1439 ^ n998 ;
  assign n14828 = n11262 & ~n14827 ;
  assign n14829 = n2113 ^ n872 ^ 1'b0 ;
  assign n14830 = ( n2039 & ~n13971 ) | ( n2039 & n14829 ) | ( ~n13971 & n14829 ) ;
  assign n14831 = n6068 & n10240 ;
  assign n14832 = n4359 & ~n6385 ;
  assign n14833 = n14831 & n14832 ;
  assign n14834 = n13477 ^ n12936 ^ n2813 ;
  assign n14835 = ~n367 & n14834 ;
  assign n14836 = n14833 & ~n14835 ;
  assign n14837 = n8763 ^ n7591 ^ n5857 ;
  assign n14838 = n14837 ^ n11101 ^ 1'b0 ;
  assign n14839 = n10779 ^ n4592 ^ n2624 ;
  assign n14840 = ( n2927 & ~n3971 ) | ( n2927 & n14839 ) | ( ~n3971 & n14839 ) ;
  assign n14841 = n13381 ^ x14 ^ 1'b0 ;
  assign n14842 = ~n8112 & n14841 ;
  assign n14843 = n14842 ^ n8308 ^ 1'b0 ;
  assign n14844 = ~n2156 & n8507 ;
  assign n14845 = n14844 ^ n6702 ^ 1'b0 ;
  assign n14846 = ( x99 & ~n4578 ) | ( x99 & n11905 ) | ( ~n4578 & n11905 ) ;
  assign n14847 = ~n11572 & n14846 ;
  assign n14848 = n14847 ^ n14749 ^ 1'b0 ;
  assign n14849 = n5361 ^ n4441 ^ 1'b0 ;
  assign n14850 = ( ~n533 & n1885 ) | ( ~n533 & n4107 ) | ( n1885 & n4107 ) ;
  assign n14851 = ( ~n2487 & n5858 ) | ( ~n2487 & n14850 ) | ( n5858 & n14850 ) ;
  assign n14852 = ( n232 & n13367 ) | ( n232 & n14851 ) | ( n13367 & n14851 ) ;
  assign n14853 = ( n12656 & n14849 ) | ( n12656 & n14852 ) | ( n14849 & n14852 ) ;
  assign n14854 = ( n851 & ~n1079 ) | ( n851 & n10260 ) | ( ~n1079 & n10260 ) ;
  assign n14855 = n681 | n7284 ;
  assign n14856 = ~n1716 & n14855 ;
  assign n14857 = n14856 ^ n7299 ^ 1'b0 ;
  assign n14858 = n14835 ^ n5915 ^ 1'b0 ;
  assign n14859 = n270 & n14858 ;
  assign n14860 = n6828 ^ n319 ^ 1'b0 ;
  assign n14861 = n7614 ^ n5655 ^ 1'b0 ;
  assign n14862 = ~n8995 & n11835 ;
  assign n14863 = n14862 ^ n5054 ^ 1'b0 ;
  assign n14864 = ( n2381 & n14861 ) | ( n2381 & ~n14863 ) | ( n14861 & ~n14863 ) ;
  assign n14865 = ~x60 & n6909 ;
  assign n14866 = n14865 ^ n2826 ^ 1'b0 ;
  assign n14867 = ~n10976 & n14866 ;
  assign n14868 = n14867 ^ n6621 ^ n5182 ;
  assign n14869 = ( n5168 & ~n7524 ) | ( n5168 & n14868 ) | ( ~n7524 & n14868 ) ;
  assign n14870 = n11241 ^ n7022 ^ 1'b0 ;
  assign n14872 = n983 & ~n2496 ;
  assign n14871 = n803 | n3540 ;
  assign n14873 = n14872 ^ n14871 ^ 1'b0 ;
  assign n14874 = n1870 & ~n8437 ;
  assign n14875 = ( n322 & n719 ) | ( n322 & ~n6362 ) | ( n719 & ~n6362 ) ;
  assign n14876 = n14875 ^ n13421 ^ n2057 ;
  assign n14877 = n4552 | n5723 ;
  assign n14878 = n5331 ^ n4116 ^ n2742 ;
  assign n14879 = n12297 & ~n14878 ;
  assign n14880 = ~n531 & n14879 ;
  assign n14881 = n11609 & n14880 ;
  assign n14882 = n5796 & n14144 ;
  assign n14883 = n11622 & n14882 ;
  assign n14884 = n2969 | n14883 ;
  assign n14885 = ~n259 & n2091 ;
  assign n14886 = ~n2074 & n14885 ;
  assign n14887 = n7072 ^ n1824 ^ 1'b0 ;
  assign n14888 = n9448 | n12823 ;
  assign n14889 = ( n14886 & ~n14887 ) | ( n14886 & n14888 ) | ( ~n14887 & n14888 ) ;
  assign n14890 = ~n3337 & n4583 ;
  assign n14891 = n14890 ^ n912 ^ 1'b0 ;
  assign n14892 = ~n1036 & n14891 ;
  assign n14894 = n8785 ^ n7963 ^ 1'b0 ;
  assign n14895 = ~n8365 & n14894 ;
  assign n14893 = n227 | n8821 ;
  assign n14896 = n14895 ^ n14893 ^ 1'b0 ;
  assign n14897 = n366 | n2209 ;
  assign n14898 = ~n2323 & n14897 ;
  assign n14899 = ( n6183 & ~n14117 ) | ( n6183 & n14898 ) | ( ~n14117 & n14898 ) ;
  assign n14900 = n11588 ^ n4686 ^ n1574 ;
  assign n14901 = n14900 ^ n9008 ^ n5166 ;
  assign n14902 = ( n808 & n7902 ) | ( n808 & n14901 ) | ( n7902 & n14901 ) ;
  assign n14903 = ( n12489 & ~n14899 ) | ( n12489 & n14902 ) | ( ~n14899 & n14902 ) ;
  assign n14905 = ( n7942 & n9536 ) | ( n7942 & ~n9608 ) | ( n9536 & ~n9608 ) ;
  assign n14904 = n13172 ^ n9913 ^ n346 ;
  assign n14906 = n14905 ^ n14904 ^ n2745 ;
  assign n14908 = n8336 ^ n3681 ^ 1'b0 ;
  assign n14907 = n7982 ^ n129 ^ 1'b0 ;
  assign n14909 = n14908 ^ n14907 ^ n4290 ;
  assign n14910 = n14909 ^ n10681 ^ n5116 ;
  assign n14911 = n4576 ^ n747 ^ 1'b0 ;
  assign n14912 = n14911 ^ n1360 ^ 1'b0 ;
  assign n14913 = n8370 ^ n3055 ^ n1574 ;
  assign n14914 = n1332 & n14913 ;
  assign n14915 = ( ~n849 & n1780 ) | ( ~n849 & n14914 ) | ( n1780 & n14914 ) ;
  assign n14916 = n3976 ^ n514 ^ 1'b0 ;
  assign n14917 = n14915 & ~n14916 ;
  assign n14918 = n9925 ^ n4602 ^ 1'b0 ;
  assign n14919 = n4199 | n14918 ;
  assign n14920 = n14919 ^ n2398 ^ n2051 ;
  assign n14921 = ( ~n4413 & n4795 ) | ( ~n4413 & n5928 ) | ( n4795 & n5928 ) ;
  assign n14922 = n14921 ^ n14007 ^ n8577 ;
  assign n14923 = ( ~n2003 & n7376 ) | ( ~n2003 & n12707 ) | ( n7376 & n12707 ) ;
  assign n14924 = n14923 ^ n10060 ^ 1'b0 ;
  assign n14925 = n2972 | n4253 ;
  assign n14926 = ( n11377 & n14183 ) | ( n11377 & n14925 ) | ( n14183 & n14925 ) ;
  assign n14927 = n9757 ^ n655 ^ 1'b0 ;
  assign n14928 = ( n4413 & n11061 ) | ( n4413 & n14601 ) | ( n11061 & n14601 ) ;
  assign n14929 = ( ~n5689 & n14927 ) | ( ~n5689 & n14928 ) | ( n14927 & n14928 ) ;
  assign n14930 = n2082 | n2644 ;
  assign n14931 = n14930 ^ n13413 ^ 1'b0 ;
  assign n14932 = n14931 ^ n6252 ^ n2882 ;
  assign n14933 = ~n6436 & n14932 ;
  assign n14934 = n8523 & n14933 ;
  assign n14935 = n13991 & n14934 ;
  assign n14936 = n2076 & n11231 ;
  assign n14937 = n14936 ^ n12427 ^ 1'b0 ;
  assign n14938 = ~n1762 & n7812 ;
  assign n14939 = n14938 ^ n3664 ^ 1'b0 ;
  assign n14940 = n14273 ^ n11953 ^ 1'b0 ;
  assign n14941 = ~n6673 & n14940 ;
  assign n14942 = n1454 & ~n6938 ;
  assign n14943 = n7100 ^ n6396 ^ 1'b0 ;
  assign n14944 = ( n13613 & n14942 ) | ( n13613 & n14943 ) | ( n14942 & n14943 ) ;
  assign n14945 = n14944 ^ n9553 ^ n7430 ;
  assign n14946 = n14945 ^ n14919 ^ 1'b0 ;
  assign n14947 = n2870 | n5054 ;
  assign n14948 = n14947 ^ n3888 ^ 1'b0 ;
  assign n14949 = n2626 & ~n14948 ;
  assign n14950 = n8990 | n14949 ;
  assign n14951 = n14950 ^ n3820 ^ 1'b0 ;
  assign n14952 = n2797 ^ n2782 ^ 1'b0 ;
  assign n14953 = n3338 & n14952 ;
  assign n14954 = ~n14951 & n14953 ;
  assign n14955 = ~n6941 & n10346 ;
  assign n14956 = ( n2645 & ~n14954 ) | ( n2645 & n14955 ) | ( ~n14954 & n14955 ) ;
  assign n14957 = ~n11190 & n14956 ;
  assign n14958 = n12861 ^ n9125 ^ 1'b0 ;
  assign n14959 = ( n454 & n7913 ) | ( n454 & n14958 ) | ( n7913 & n14958 ) ;
  assign n14960 = n1699 ^ n977 ^ 1'b0 ;
  assign n14961 = n4931 & ~n14960 ;
  assign n14962 = ( ~n5283 & n13145 ) | ( ~n5283 & n14961 ) | ( n13145 & n14961 ) ;
  assign n14963 = n12094 & ~n14962 ;
  assign n14964 = n4087 & n7326 ;
  assign n14965 = n11557 ^ n7854 ^ 1'b0 ;
  assign n14966 = n7180 ^ n2654 ^ 1'b0 ;
  assign n14967 = n14966 ^ n6344 ^ n758 ;
  assign n14968 = n14967 ^ n5059 ^ n1138 ;
  assign n14969 = ( n11053 & n14965 ) | ( n11053 & n14968 ) | ( n14965 & n14968 ) ;
  assign n14970 = n8393 ^ n6493 ^ 1'b0 ;
  assign n14971 = n2063 & n14970 ;
  assign n14972 = n14971 ^ n1319 ^ 1'b0 ;
  assign n14973 = n14972 ^ n11868 ^ n11698 ;
  assign n14974 = ( n3036 & ~n3256 ) | ( n3036 & n4942 ) | ( ~n3256 & n4942 ) ;
  assign n14975 = ( ~n11202 & n14407 ) | ( ~n11202 & n14974 ) | ( n14407 & n14974 ) ;
  assign n14976 = n14509 ^ n12503 ^ n3290 ;
  assign n14977 = n14976 ^ n9137 ^ 1'b0 ;
  assign n14979 = n1449 & ~n4614 ;
  assign n14980 = n14979 ^ n620 ^ 1'b0 ;
  assign n14978 = n6458 & n12736 ;
  assign n14981 = n14980 ^ n14978 ^ 1'b0 ;
  assign n14982 = ( n6026 & n7624 ) | ( n6026 & ~n14981 ) | ( n7624 & ~n14981 ) ;
  assign n14983 = ( ~n6099 & n6226 ) | ( ~n6099 & n6623 ) | ( n6226 & n6623 ) ;
  assign n14984 = n1732 ^ n1513 ^ 1'b0 ;
  assign n14985 = n14983 & n14984 ;
  assign n14986 = n9948 | n14374 ;
  assign n14987 = n14985 | n14986 ;
  assign n14988 = ( n2453 & n8833 ) | ( n2453 & n14001 ) | ( n8833 & n14001 ) ;
  assign n14989 = n9151 ^ n2319 ^ 1'b0 ;
  assign n14990 = n1036 & n12095 ;
  assign n14991 = n14990 ^ n8552 ^ n1355 ;
  assign n14992 = n2387 ^ n1626 ^ 1'b0 ;
  assign n14993 = ~n4678 & n7108 ;
  assign n14994 = n14993 ^ x80 ^ 1'b0 ;
  assign n14995 = n14994 ^ n2272 ^ 1'b0 ;
  assign n14999 = n12563 ^ n888 ^ 1'b0 ;
  assign n15000 = n6434 | n8412 ;
  assign n15001 = n14999 & ~n15000 ;
  assign n14996 = n7080 ^ n3441 ^ 1'b0 ;
  assign n14997 = n9911 & n14996 ;
  assign n14998 = ~n3566 & n14997 ;
  assign n15002 = n15001 ^ n14998 ^ 1'b0 ;
  assign n15003 = n7865 ^ n337 ^ 1'b0 ;
  assign n15004 = ( n11379 & n13141 ) | ( n11379 & ~n15003 ) | ( n13141 & ~n15003 ) ;
  assign n15005 = n15004 ^ n9521 ^ 1'b0 ;
  assign n15006 = n3168 & ~n3870 ;
  assign n15007 = n12473 ^ n701 ^ 1'b0 ;
  assign n15008 = n4554 & ~n15007 ;
  assign n15009 = n1968 & n8066 ;
  assign n15010 = n1240 & n15009 ;
  assign n15011 = n2170 | n8038 ;
  assign n15012 = n3532 ^ n2559 ^ 1'b0 ;
  assign n15013 = n5824 & ~n8076 ;
  assign n15014 = ~n3062 & n15013 ;
  assign n15015 = n9082 | n15014 ;
  assign n15016 = n15015 ^ n8399 ^ 1'b0 ;
  assign n15017 = n15016 ^ n12726 ^ n2417 ;
  assign n15018 = ( ~n2475 & n2949 ) | ( ~n2475 & n7968 ) | ( n2949 & n7968 ) ;
  assign n15019 = n15018 ^ n5596 ^ n3602 ;
  assign n15020 = n4217 ^ n2000 ^ n1056 ;
  assign n15021 = n3399 & ~n4650 ;
  assign n15022 = n15021 ^ n6572 ^ 1'b0 ;
  assign n15023 = n15022 ^ n14846 ^ n14460 ;
  assign n15024 = ( n15019 & n15020 ) | ( n15019 & ~n15023 ) | ( n15020 & ~n15023 ) ;
  assign n15025 = ~n1639 & n5729 ;
  assign n15026 = n13832 & n15025 ;
  assign n15029 = n6058 ^ n589 ^ 1'b0 ;
  assign n15030 = ~n14318 & n15029 ;
  assign n15027 = n1944 | n5660 ;
  assign n15028 = n15027 ^ n2555 ^ 1'b0 ;
  assign n15031 = n15030 ^ n15028 ^ 1'b0 ;
  assign n15032 = n15031 ^ n10132 ^ n1903 ;
  assign n15033 = n15026 & n15032 ;
  assign n15034 = ( n3314 & n4167 ) | ( n3314 & n9670 ) | ( n4167 & n9670 ) ;
  assign n15035 = ( n3218 & ~n3691 ) | ( n3218 & n5381 ) | ( ~n3691 & n5381 ) ;
  assign n15036 = ( n3947 & ~n9827 ) | ( n3947 & n15035 ) | ( ~n9827 & n15035 ) ;
  assign n15037 = n15036 ^ n9007 ^ 1'b0 ;
  assign n15038 = n567 | n8130 ;
  assign n15039 = n10767 | n15038 ;
  assign n15040 = n15039 ^ n9465 ^ n3641 ;
  assign n15041 = ~n7659 & n15040 ;
  assign n15042 = n2865 & n15041 ;
  assign n15043 = n6120 | n15042 ;
  assign n15044 = n7646 & ~n15043 ;
  assign n15045 = n4083 & n8651 ;
  assign n15046 = n15045 ^ n12543 ^ n3990 ;
  assign n15047 = n6856 ^ n3959 ^ 1'b0 ;
  assign n15048 = n15047 ^ n3694 ^ n207 ;
  assign n15049 = n7009 ^ n2923 ^ 1'b0 ;
  assign n15050 = n3351 | n15049 ;
  assign n15052 = n3106 | n5932 ;
  assign n15053 = n15052 ^ n5523 ^ 1'b0 ;
  assign n15054 = ~n14561 & n15053 ;
  assign n15051 = n3860 & ~n7801 ;
  assign n15055 = n15054 ^ n15051 ^ 1'b0 ;
  assign n15056 = n12923 ^ n3424 ^ 1'b0 ;
  assign n15057 = n6488 & n15056 ;
  assign n15058 = n4934 | n5284 ;
  assign n15059 = n4100 | n15058 ;
  assign n15060 = ( ~n2900 & n3980 ) | ( ~n2900 & n15059 ) | ( n3980 & n15059 ) ;
  assign n15061 = x51 & ~n6085 ;
  assign n15062 = n13244 & n15061 ;
  assign n15063 = n4334 & ~n6197 ;
  assign n15064 = ~n9819 & n15063 ;
  assign n15065 = n3734 | n15064 ;
  assign n15066 = n15065 ^ n987 ^ 1'b0 ;
  assign n15069 = n5313 & n6060 ;
  assign n15070 = n15069 ^ n11717 ^ 1'b0 ;
  assign n15067 = n830 | n13701 ;
  assign n15068 = n7855 | n15067 ;
  assign n15071 = n15070 ^ n15068 ^ 1'b0 ;
  assign n15072 = ~n2718 & n15071 ;
  assign n15073 = ( n1311 & n1673 ) | ( n1311 & n15072 ) | ( n1673 & n15072 ) ;
  assign n15074 = ~n897 & n3597 ;
  assign n15075 = ( n10453 & n13017 ) | ( n10453 & n15074 ) | ( n13017 & n15074 ) ;
  assign n15076 = ( n5356 & n6652 ) | ( n5356 & n15075 ) | ( n6652 & n15075 ) ;
  assign n15077 = n14934 ^ n4961 ^ 1'b0 ;
  assign n15078 = n8255 ^ n2453 ^ 1'b0 ;
  assign n15079 = ~n13902 & n15078 ;
  assign n15080 = n15079 ^ n15024 ^ 1'b0 ;
  assign n15081 = ~n1264 & n4207 ;
  assign n15082 = n797 ^ n307 ^ 1'b0 ;
  assign n15083 = n15081 & n15082 ;
  assign n15084 = n11779 ^ n3323 ^ 1'b0 ;
  assign n15087 = n10192 ^ n3567 ^ n3448 ;
  assign n15086 = n666 & ~n3031 ;
  assign n15085 = ( n1947 & ~n4640 ) | ( n1947 & n13396 ) | ( ~n4640 & n13396 ) ;
  assign n15088 = n15087 ^ n15086 ^ n15085 ;
  assign n15089 = n7417 & ~n8786 ;
  assign n15090 = ~n5836 & n15089 ;
  assign n15091 = n1838 | n7490 ;
  assign n15092 = n11546 | n15091 ;
  assign n15093 = n7929 ^ n5672 ^ n1188 ;
  assign n15094 = n15093 ^ n13705 ^ n159 ;
  assign n15099 = n1629 & ~n7501 ;
  assign n15100 = n15099 ^ n522 ^ 1'b0 ;
  assign n15095 = n9933 ^ n2881 ^ n2181 ;
  assign n15096 = n10584 & n15095 ;
  assign n15097 = n1034 & n15096 ;
  assign n15098 = n15097 ^ n11464 ^ 1'b0 ;
  assign n15101 = n15100 ^ n15098 ^ n4210 ;
  assign n15102 = ( n5349 & n5377 ) | ( n5349 & n5714 ) | ( n5377 & n5714 ) ;
  assign n15103 = n7410 ^ n2872 ^ n1638 ;
  assign n15104 = ( n7465 & ~n11198 ) | ( n7465 & n15103 ) | ( ~n11198 & n15103 ) ;
  assign n15105 = n15102 & ~n15104 ;
  assign n15106 = n3872 & n9597 ;
  assign n15107 = ~n10180 & n15106 ;
  assign n15108 = ~n7419 & n9582 ;
  assign n15109 = n15107 & n15108 ;
  assign n15111 = n3573 ^ n1590 ^ 1'b0 ;
  assign n15112 = ~n4727 & n15111 ;
  assign n15110 = n11847 ^ n1792 ^ 1'b0 ;
  assign n15113 = n15112 ^ n15110 ^ n1092 ;
  assign n15114 = n9193 ^ n8240 ^ n7205 ;
  assign n15115 = ( ~n2166 & n8860 ) | ( ~n2166 & n15114 ) | ( n8860 & n15114 ) ;
  assign n15116 = n10978 | n15115 ;
  assign n15117 = n13818 & ~n15116 ;
  assign n15118 = ( n9999 & n10224 ) | ( n9999 & ~n12157 ) | ( n10224 & ~n12157 ) ;
  assign n15119 = n6678 ^ n4270 ^ n2608 ;
  assign n15120 = n15119 ^ n4402 ^ 1'b0 ;
  assign n15121 = ~n15118 & n15120 ;
  assign n15122 = n3848 & ~n4414 ;
  assign n15123 = n15122 ^ n8210 ^ 1'b0 ;
  assign n15124 = n5705 & ~n15123 ;
  assign n15125 = n15124 ^ n14409 ^ 1'b0 ;
  assign n15126 = ( ~n3500 & n3528 ) | ( ~n3500 & n13564 ) | ( n3528 & n13564 ) ;
  assign n15127 = n2167 ^ n2114 ^ 1'b0 ;
  assign n15128 = ~n1578 & n15127 ;
  assign n15129 = ( n717 & n11419 ) | ( n717 & ~n15128 ) | ( n11419 & ~n15128 ) ;
  assign n15130 = ( n1338 & n5832 ) | ( n1338 & n15129 ) | ( n5832 & n15129 ) ;
  assign n15131 = n5392 | n13130 ;
  assign n15132 = n611 & ~n5633 ;
  assign n15133 = n15131 & n15132 ;
  assign n15134 = ( n15126 & ~n15130 ) | ( n15126 & n15133 ) | ( ~n15130 & n15133 ) ;
  assign n15135 = n5519 ^ n2846 ^ n318 ;
  assign n15136 = n15135 ^ n6166 ^ n3752 ;
  assign n15137 = n1929 & ~n10554 ;
  assign n15138 = ~n2845 & n15137 ;
  assign n15139 = n12441 | n15138 ;
  assign n15140 = n15136 & ~n15139 ;
  assign n15141 = n13438 ^ n5189 ^ 1'b0 ;
  assign n15142 = ( n155 & n7618 ) | ( n155 & n10084 ) | ( n7618 & n10084 ) ;
  assign n15145 = ( n1273 & ~n4859 ) | ( n1273 & n5699 ) | ( ~n4859 & n5699 ) ;
  assign n15143 = n2520 | n4461 ;
  assign n15144 = n4978 | n15143 ;
  assign n15146 = n15145 ^ n15144 ^ n6878 ;
  assign n15147 = ( x18 & n5596 ) | ( x18 & n12812 ) | ( n5596 & n12812 ) ;
  assign n15148 = n2122 | n11931 ;
  assign n15149 = n3285 | n15148 ;
  assign n15150 = n6568 ^ n1678 ^ n429 ;
  assign n15151 = n2713 & n15150 ;
  assign n15152 = n15151 ^ n7024 ^ 1'b0 ;
  assign n15153 = n11126 ^ n4982 ^ 1'b0 ;
  assign n15154 = ( n11883 & n13834 ) | ( n11883 & ~n15153 ) | ( n13834 & ~n15153 ) ;
  assign n15155 = n8805 ^ n8735 ^ n4413 ;
  assign n15156 = n9766 & ~n14778 ;
  assign n15157 = n14778 & n15156 ;
  assign n15158 = n12260 ^ n4036 ^ n1214 ;
  assign n15159 = n4756 ^ n3913 ^ 1'b0 ;
  assign n15160 = n9647 ^ n3486 ^ 1'b0 ;
  assign n15161 = n8310 & ~n15160 ;
  assign n15162 = ~n4267 & n8451 ;
  assign n15163 = ( n14177 & n15161 ) | ( n14177 & n15162 ) | ( n15161 & n15162 ) ;
  assign n15167 = n9207 ^ n9203 ^ 1'b0 ;
  assign n15168 = n6384 & ~n15167 ;
  assign n15169 = n15168 ^ n5120 ^ 1'b0 ;
  assign n15164 = n8301 ^ n4306 ^ 1'b0 ;
  assign n15165 = n943 & n15164 ;
  assign n15166 = n15165 ^ n13432 ^ 1'b0 ;
  assign n15170 = n15169 ^ n15166 ^ n6092 ;
  assign n15171 = n8567 ^ n3098 ^ 1'b0 ;
  assign n15172 = n13100 ^ n1488 ^ 1'b0 ;
  assign n15173 = n5542 & n15172 ;
  assign n15174 = n1760 & n15173 ;
  assign n15176 = n3080 ^ n1073 ^ 1'b0 ;
  assign n15177 = n376 & ~n15176 ;
  assign n15178 = n15177 ^ n13701 ^ n10701 ;
  assign n15175 = n9242 & ~n13223 ;
  assign n15179 = n15178 ^ n15175 ^ 1'b0 ;
  assign n15180 = n9463 & n10442 ;
  assign n15181 = n11072 ^ n4704 ^ n3636 ;
  assign n15182 = n9851 ^ n9773 ^ n7099 ;
  assign n15183 = ~n1975 & n15182 ;
  assign n15184 = n15183 ^ n487 ^ 1'b0 ;
  assign n15185 = n5345 | n15184 ;
  assign n15186 = n3299 ^ n514 ^ 1'b0 ;
  assign n15187 = n5086 | n15186 ;
  assign n15188 = ~n1993 & n5704 ;
  assign n15189 = n15188 ^ n6316 ^ 1'b0 ;
  assign n15190 = ~n2917 & n15189 ;
  assign n15191 = ( n3858 & ~n9926 ) | ( n3858 & n15190 ) | ( ~n9926 & n15190 ) ;
  assign n15192 = n2141 & ~n15191 ;
  assign n15193 = n15187 & n15192 ;
  assign n15194 = n8904 | n14413 ;
  assign n15195 = ( n5389 & ~n7883 ) | ( n5389 & n15194 ) | ( ~n7883 & n15194 ) ;
  assign n15196 = n6385 ^ n4789 ^ n1254 ;
  assign n15197 = n14150 ^ n1464 ^ 1'b0 ;
  assign n15198 = ~n15196 & n15197 ;
  assign n15199 = n3109 | n10127 ;
  assign n15200 = n6340 & ~n15199 ;
  assign n15201 = ( n1568 & n13419 ) | ( n1568 & n14678 ) | ( n13419 & n14678 ) ;
  assign n15202 = ( ~n649 & n15200 ) | ( ~n649 & n15201 ) | ( n15200 & n15201 ) ;
  assign n15203 = n285 & n3713 ;
  assign n15204 = n15202 & n15203 ;
  assign n15205 = ( ~n2369 & n2863 ) | ( ~n2369 & n6554 ) | ( n2863 & n6554 ) ;
  assign n15206 = n11341 | n13017 ;
  assign n15207 = n9958 | n15206 ;
  assign n15208 = n15205 & ~n15207 ;
  assign n15209 = ~n7998 & n12371 ;
  assign n15210 = n926 & ~n1235 ;
  assign n15211 = ~n2172 & n15210 ;
  assign n15212 = n15211 ^ n8370 ^ 1'b0 ;
  assign n15213 = ( n6261 & ~n15209 ) | ( n6261 & n15212 ) | ( ~n15209 & n15212 ) ;
  assign n15214 = n14333 & ~n15213 ;
  assign n15215 = n10467 ^ n10154 ^ 1'b0 ;
  assign n15216 = n7988 ^ n4629 ^ n3610 ;
  assign n15221 = n12112 ^ n7852 ^ 1'b0 ;
  assign n15222 = n15221 ^ n8987 ^ n8527 ;
  assign n15220 = n4723 ^ n3722 ^ 1'b0 ;
  assign n15217 = n8466 & ~n12499 ;
  assign n15218 = n5416 & ~n15217 ;
  assign n15219 = n9948 & n15218 ;
  assign n15223 = n15222 ^ n15220 ^ n15219 ;
  assign n15224 = n11602 ^ n8038 ^ 1'b0 ;
  assign n15225 = n15216 | n15224 ;
  assign n15226 = n1030 | n3423 ;
  assign n15227 = n10650 & ~n15226 ;
  assign n15228 = ( n1208 & n5436 ) | ( n1208 & n15227 ) | ( n5436 & n15227 ) ;
  assign n15229 = n3281 ^ n1117 ^ 1'b0 ;
  assign n15230 = ~n15228 & n15229 ;
  assign n15233 = ( ~n1889 & n3449 ) | ( ~n1889 & n10373 ) | ( n3449 & n10373 ) ;
  assign n15231 = n11286 ^ n1416 ^ 1'b0 ;
  assign n15232 = n3357 & ~n15231 ;
  assign n15234 = n15233 ^ n15232 ^ 1'b0 ;
  assign n15235 = n13305 ^ n10288 ^ n4426 ;
  assign n15236 = n7827 ^ n4558 ^ 1'b0 ;
  assign n15237 = n7774 ^ n5482 ^ n2978 ;
  assign n15238 = n890 ^ n194 ^ 1'b0 ;
  assign n15239 = n15237 & n15238 ;
  assign n15240 = n15236 & n15239 ;
  assign n15241 = ~n7855 & n15240 ;
  assign n15242 = n1405 | n11687 ;
  assign n15243 = n15242 ^ n1647 ^ 1'b0 ;
  assign n15244 = n9857 ^ n5704 ^ n583 ;
  assign n15245 = ~n7347 & n7626 ;
  assign n15246 = n12575 ^ n3879 ^ 1'b0 ;
  assign n15247 = n15245 & ~n15246 ;
  assign n15248 = n4185 | n13787 ;
  assign n15249 = x113 | n15248 ;
  assign n15250 = n541 & ~n5769 ;
  assign n15251 = n15250 ^ n4640 ^ 1'b0 ;
  assign n15252 = n15249 & n15251 ;
  assign n15253 = n4930 ^ n3219 ^ 1'b0 ;
  assign n15254 = n15253 ^ n574 ^ 1'b0 ;
  assign n15255 = n4584 & ~n15254 ;
  assign n15257 = ~n1196 & n8946 ;
  assign n15258 = n15257 ^ n3738 ^ n693 ;
  assign n15256 = ( ~n8280 & n8888 ) | ( ~n8280 & n12879 ) | ( n8888 & n12879 ) ;
  assign n15259 = n15258 ^ n15256 ^ n3759 ;
  assign n15260 = n6027 ^ n6024 ^ 1'b0 ;
  assign n15261 = n5765 ^ n5760 ^ n333 ;
  assign n15262 = ( ~n13674 & n15260 ) | ( ~n13674 & n15261 ) | ( n15260 & n15261 ) ;
  assign n15263 = ~n1349 & n6607 ;
  assign n15265 = ( n5062 & n9741 ) | ( n5062 & ~n11597 ) | ( n9741 & ~n11597 ) ;
  assign n15266 = ( n357 & n5652 ) | ( n357 & ~n15265 ) | ( n5652 & ~n15265 ) ;
  assign n15264 = ~n9105 & n9241 ;
  assign n15267 = n15266 ^ n15264 ^ n9828 ;
  assign n15268 = n4015 & n4374 ;
  assign n15269 = ~n10676 & n15268 ;
  assign n15270 = n1872 | n4033 ;
  assign n15271 = ~n1508 & n8088 ;
  assign n15272 = n15271 ^ n6644 ^ 1'b0 ;
  assign n15273 = n2898 & n8287 ;
  assign n15274 = n15273 ^ n8749 ^ 1'b0 ;
  assign n15275 = ( n6562 & n13426 ) | ( n6562 & n15274 ) | ( n13426 & n15274 ) ;
  assign n15276 = ( n3485 & n15272 ) | ( n3485 & n15275 ) | ( n15272 & n15275 ) ;
  assign n15277 = ( n9770 & n10604 ) | ( n9770 & n15138 ) | ( n10604 & n15138 ) ;
  assign n15278 = ( n10687 & n14048 ) | ( n10687 & n14218 ) | ( n14048 & n14218 ) ;
  assign n15279 = n11722 ^ n848 ^ 1'b0 ;
  assign n15280 = ~n844 & n11322 ;
  assign n15281 = ~n5917 & n15280 ;
  assign n15282 = n7471 & n11879 ;
  assign n15283 = ( n661 & n5667 ) | ( n661 & ~n9277 ) | ( n5667 & ~n9277 ) ;
  assign n15284 = ~n2727 & n10918 ;
  assign n15285 = ~x60 & n15284 ;
  assign n15286 = n15285 ^ n6580 ^ n2290 ;
  assign n15287 = ~n12177 & n13538 ;
  assign n15288 = n951 | n4357 ;
  assign n15289 = n1649 | n15288 ;
  assign n15290 = n10799 ^ n2956 ^ 1'b0 ;
  assign n15291 = n1205 | n9298 ;
  assign n15292 = n15290 | n15291 ;
  assign n15293 = n6385 ^ n3507 ^ 1'b0 ;
  assign n15294 = n5231 & ~n15293 ;
  assign n15295 = n4270 & ~n6966 ;
  assign n15296 = n15294 | n15295 ;
  assign n15297 = n9098 ^ n6967 ^ 1'b0 ;
  assign n15298 = ( n3365 & n8298 ) | ( n3365 & ~n15297 ) | ( n8298 & ~n15297 ) ;
  assign n15299 = n2433 ^ n461 ^ 1'b0 ;
  assign n15300 = n15299 ^ n10875 ^ n10645 ;
  assign n15301 = n3052 & n4224 ;
  assign n15302 = ~n15300 & n15301 ;
  assign n15303 = ~n3032 & n13620 ;
  assign n15304 = n8052 ^ n3438 ^ 1'b0 ;
  assign n15305 = n5533 ^ n1839 ^ n739 ;
  assign n15306 = n15305 ^ n2737 ^ 1'b0 ;
  assign n15307 = n15306 ^ n1360 ^ 1'b0 ;
  assign n15308 = n15307 ^ n13864 ^ n4120 ;
  assign n15309 = n3282 ^ n1492 ^ 1'b0 ;
  assign n15310 = n15309 ^ n14621 ^ n11302 ;
  assign n15311 = n13354 ^ n1515 ^ 1'b0 ;
  assign n15312 = n2593 & n10711 ;
  assign n15313 = n8215 ^ n154 ^ 1'b0 ;
  assign n15314 = n7622 & n15313 ;
  assign n15315 = n11087 ^ n1199 ^ 1'b0 ;
  assign n15316 = n15170 & n15315 ;
  assign n15319 = n13632 ^ x45 ^ 1'b0 ;
  assign n15317 = ~n4424 & n8800 ;
  assign n15318 = n8337 & ~n15317 ;
  assign n15320 = n15319 ^ n15318 ^ 1'b0 ;
  assign n15321 = n11246 ^ n10900 ^ n7417 ;
  assign n15322 = ( ~n2304 & n4008 ) | ( ~n2304 & n11921 ) | ( n4008 & n11921 ) ;
  assign n15323 = ( n283 & n1838 ) | ( n283 & ~n2856 ) | ( n1838 & ~n2856 ) ;
  assign n15324 = n8492 & ~n11601 ;
  assign n15325 = n5369 & n15324 ;
  assign n15326 = ( n1867 & ~n5762 ) | ( n1867 & n7876 ) | ( ~n5762 & n7876 ) ;
  assign n15327 = n15325 | n15326 ;
  assign n15328 = ( n1581 & ~n14424 ) | ( n1581 & n15222 ) | ( ~n14424 & n15222 ) ;
  assign n15329 = ( n1902 & ~n2353 ) | ( n1902 & n15328 ) | ( ~n2353 & n15328 ) ;
  assign n15330 = n6413 ^ n1542 ^ 1'b0 ;
  assign n15331 = n9136 ^ n4155 ^ n486 ;
  assign n15332 = n15331 ^ n13744 ^ 1'b0 ;
  assign n15333 = n15330 & ~n15332 ;
  assign n15334 = ( ~n11809 & n14330 ) | ( ~n11809 & n15333 ) | ( n14330 & n15333 ) ;
  assign n15335 = n11025 ^ n10572 ^ n9679 ;
  assign n15336 = n6662 & ~n15335 ;
  assign n15337 = ~n11609 & n15336 ;
  assign n15338 = ~n6198 & n15337 ;
  assign n15339 = ( n3831 & ~n6780 ) | ( n3831 & n9041 ) | ( ~n6780 & n9041 ) ;
  assign n15341 = n6733 ^ n4668 ^ 1'b0 ;
  assign n15340 = n7992 | n11136 ;
  assign n15342 = n15341 ^ n15340 ^ 1'b0 ;
  assign n15343 = n15342 ^ n12256 ^ n8475 ;
  assign n15344 = n5220 ^ n4618 ^ n3657 ;
  assign n15345 = n1425 & n6382 ;
  assign n15346 = ( n773 & ~n9223 ) | ( n773 & n15345 ) | ( ~n9223 & n15345 ) ;
  assign n15347 = n3140 | n15346 ;
  assign n15348 = n15344 & ~n15347 ;
  assign n15349 = ~n6315 & n15348 ;
  assign n15350 = n1374 ^ n184 ^ 1'b0 ;
  assign n15351 = ( n10713 & n13061 ) | ( n10713 & ~n15350 ) | ( n13061 & ~n15350 ) ;
  assign n15352 = ( x121 & ~n13885 ) | ( x121 & n15351 ) | ( ~n13885 & n15351 ) ;
  assign n15353 = n6958 ^ n4157 ^ 1'b0 ;
  assign n15354 = n2748 | n15353 ;
  assign n15355 = ( n3678 & n11777 ) | ( n3678 & n15354 ) | ( n11777 & n15354 ) ;
  assign n15356 = n3065 ^ n1688 ^ 1'b0 ;
  assign n15357 = n6636 & ~n15356 ;
  assign n15358 = n2982 & ~n6133 ;
  assign n15359 = n12942 & n15358 ;
  assign n15360 = n9199 ^ n6196 ^ n3192 ;
  assign n15361 = n4157 ^ n3946 ^ n1966 ;
  assign n15362 = ( ~n10154 & n12275 ) | ( ~n10154 & n15361 ) | ( n12275 & n15361 ) ;
  assign n15363 = n15362 ^ n9722 ^ n1796 ;
  assign n15364 = n1580 & n15363 ;
  assign n15366 = n3525 ^ n2500 ^ 1'b0 ;
  assign n15365 = n6276 & ~n11606 ;
  assign n15367 = n15366 ^ n15365 ^ 1'b0 ;
  assign n15371 = n416 & ~n5674 ;
  assign n15368 = ( n5231 & ~n12309 ) | ( n5231 & n12563 ) | ( ~n12309 & n12563 ) ;
  assign n15369 = ~n5122 & n15368 ;
  assign n15370 = n3385 & n15369 ;
  assign n15372 = n15371 ^ n15370 ^ 1'b0 ;
  assign n15375 = x113 & n1124 ;
  assign n15376 = n15375 ^ n2360 ^ 1'b0 ;
  assign n15373 = n1442 & ~n9220 ;
  assign n15374 = n11477 & ~n15373 ;
  assign n15377 = n15376 ^ n15374 ^ 1'b0 ;
  assign n15378 = n15377 ^ n14836 ^ 1'b0 ;
  assign n15379 = n7216 & n15378 ;
  assign n15380 = n5792 & ~n11799 ;
  assign n15381 = n15380 ^ n6187 ^ 1'b0 ;
  assign n15382 = n15381 ^ n13876 ^ n2045 ;
  assign n15383 = ( n908 & n6700 ) | ( n908 & ~n14053 ) | ( n6700 & ~n14053 ) ;
  assign n15384 = ( n2136 & ~n6374 ) | ( n2136 & n7325 ) | ( ~n6374 & n7325 ) ;
  assign n15385 = n11423 ^ n9406 ^ n8006 ;
  assign n15386 = n15385 ^ n8291 ^ 1'b0 ;
  assign n15387 = ~n447 & n15386 ;
  assign n15388 = ( n15383 & n15384 ) | ( n15383 & n15387 ) | ( n15384 & n15387 ) ;
  assign n15389 = n4668 & ~n6649 ;
  assign n15392 = n5396 ^ n3664 ^ n1291 ;
  assign n15390 = n5584 ^ n2931 ^ 1'b0 ;
  assign n15391 = n998 & n15390 ;
  assign n15393 = n15392 ^ n15391 ^ n6100 ;
  assign n15394 = n13337 | n15393 ;
  assign n15395 = ( n7494 & n8928 ) | ( n7494 & n9116 ) | ( n8928 & n9116 ) ;
  assign n15396 = n15395 ^ n13344 ^ n3648 ;
  assign n15400 = n618 | n8134 ;
  assign n15397 = n3707 & ~n8362 ;
  assign n15398 = n15397 ^ n9039 ^ 1'b0 ;
  assign n15399 = ~n7790 & n15398 ;
  assign n15401 = n15400 ^ n15399 ^ n8796 ;
  assign n15402 = n5051 & n11906 ;
  assign n15403 = n15402 ^ n5821 ^ 1'b0 ;
  assign n15404 = n9186 ^ n6058 ^ 1'b0 ;
  assign n15405 = n15404 ^ n7333 ^ n5021 ;
  assign n15406 = n2977 & n15405 ;
  assign n15407 = n15406 ^ n4959 ^ 1'b0 ;
  assign n15408 = n9041 & ~n13752 ;
  assign n15409 = n11188 ^ n9197 ^ n2257 ;
  assign n15410 = n8460 ^ n5819 ^ n5282 ;
  assign n15411 = ( n7617 & n11759 ) | ( n7617 & n15410 ) | ( n11759 & n15410 ) ;
  assign n15412 = n4851 ^ n2441 ^ 1'b0 ;
  assign n15413 = n10431 | n15412 ;
  assign n15414 = n15413 ^ n9403 ^ n6332 ;
  assign n15415 = ~n971 & n6908 ;
  assign n15416 = n1306 & n15415 ;
  assign n15417 = n15416 ^ n11877 ^ 1'b0 ;
  assign n15418 = n5129 | n15417 ;
  assign n15419 = n15414 & n15418 ;
  assign n15420 = n1688 & ~n1920 ;
  assign n15421 = n3221 & n15420 ;
  assign n15422 = n11879 & ~n15421 ;
  assign n15423 = n11150 & n15422 ;
  assign n15424 = ( n701 & n1385 ) | ( n701 & n15423 ) | ( n1385 & n15423 ) ;
  assign n15425 = n13129 ^ n6304 ^ 1'b0 ;
  assign n15426 = n6500 & n15425 ;
  assign n15427 = n5156 ^ n533 ^ 1'b0 ;
  assign n15428 = ~n11423 & n15427 ;
  assign n15429 = n3734 | n15428 ;
  assign n15430 = ( n821 & n7379 ) | ( n821 & n13433 ) | ( n7379 & n13433 ) ;
  assign n15431 = n15430 ^ n6919 ^ n3413 ;
  assign n15432 = n15431 ^ n13893 ^ n452 ;
  assign n15433 = n11981 ^ n6483 ^ 1'b0 ;
  assign n15434 = n2820 & n15433 ;
  assign n15435 = n8033 & n15434 ;
  assign n15436 = ~n447 & n6275 ;
  assign n15437 = n12109 & n15436 ;
  assign n15438 = n2178 & n8682 ;
  assign n15439 = n15437 & n15438 ;
  assign n15440 = ~n2048 & n6697 ;
  assign n15441 = n15440 ^ n10693 ^ 1'b0 ;
  assign n15443 = ( n7129 & n10105 ) | ( n7129 & ~n13478 ) | ( n10105 & ~n13478 ) ;
  assign n15442 = ( ~n4043 & n4554 ) | ( ~n4043 & n7768 ) | ( n4554 & n7768 ) ;
  assign n15444 = n15443 ^ n15442 ^ n754 ;
  assign n15445 = ~n1176 & n9921 ;
  assign n15446 = ~n6290 & n13485 ;
  assign n15447 = n14232 ^ n10831 ^ 1'b0 ;
  assign n15448 = n238 | n15447 ;
  assign n15449 = ( n299 & ~n2674 ) | ( n299 & n5169 ) | ( ~n2674 & n5169 ) ;
  assign n15450 = ~n7974 & n15449 ;
  assign n15451 = x118 & ~n2172 ;
  assign n15452 = n14713 ^ n10000 ^ 1'b0 ;
  assign n15453 = n13472 | n14787 ;
  assign n15454 = n11004 | n15453 ;
  assign n15455 = n7346 & n15454 ;
  assign n15456 = n12099 & n12570 ;
  assign n15457 = n15456 ^ n10068 ^ 1'b0 ;
  assign n15461 = n11184 ^ n7622 ^ n5907 ;
  assign n15462 = n15461 ^ n5028 ^ n462 ;
  assign n15463 = n4090 | n15462 ;
  assign n15464 = n6206 ^ n4211 ^ n1715 ;
  assign n15465 = n15464 ^ n8946 ^ n4101 ;
  assign n15466 = ~n15463 & n15465 ;
  assign n15458 = n10693 ^ n7287 ^ n5351 ;
  assign n15459 = n12787 ^ n1786 ^ 1'b0 ;
  assign n15460 = ( n11533 & n15458 ) | ( n11533 & n15459 ) | ( n15458 & n15459 ) ;
  assign n15467 = n15466 ^ n15460 ^ n12441 ;
  assign n15468 = n3850 ^ x92 ^ 1'b0 ;
  assign n15469 = n15468 ^ n3590 ^ n2855 ;
  assign n15470 = ( n1160 & n3584 ) | ( n1160 & ~n14171 ) | ( n3584 & ~n14171 ) ;
  assign n15471 = n10199 & ~n10265 ;
  assign n15472 = n9127 ^ n2160 ^ n321 ;
  assign n15473 = n4691 ^ n4529 ^ n663 ;
  assign n15482 = n2038 ^ n1924 ^ 1'b0 ;
  assign n15483 = n15482 ^ n15053 ^ n5418 ;
  assign n15478 = n3697 ^ n2761 ^ n293 ;
  assign n15474 = ~n155 & n4357 ;
  assign n15475 = n15474 ^ n14643 ^ 1'b0 ;
  assign n15476 = n4446 ^ n4069 ^ 1'b0 ;
  assign n15477 = ~n15475 & n15476 ;
  assign n15479 = n15478 ^ n15477 ^ n11455 ;
  assign n15480 = n15479 ^ n13219 ^ 1'b0 ;
  assign n15481 = n15480 ^ n9867 ^ n1530 ;
  assign n15484 = n15483 ^ n15481 ^ 1'b0 ;
  assign n15485 = n3604 | n4256 ;
  assign n15486 = ( n5742 & n14406 ) | ( n5742 & ~n15485 ) | ( n14406 & ~n15485 ) ;
  assign n15487 = n7924 & n15486 ;
  assign n15488 = ~n188 & n15487 ;
  assign n15495 = ( n1580 & ~n2197 ) | ( n1580 & n5909 ) | ( ~n2197 & n5909 ) ;
  assign n15496 = n15495 ^ n13814 ^ 1'b0 ;
  assign n15497 = ( n8312 & ~n9033 ) | ( n8312 & n15496 ) | ( ~n9033 & n15496 ) ;
  assign n15492 = ( n6512 & ~n9804 ) | ( n6512 & n11100 ) | ( ~n9804 & n11100 ) ;
  assign n15489 = n270 & ~n5739 ;
  assign n15490 = n6148 & n15489 ;
  assign n15491 = n8322 | n15490 ;
  assign n15493 = n15492 ^ n15491 ^ 1'b0 ;
  assign n15494 = ~n11420 & n15493 ;
  assign n15498 = n15497 ^ n15494 ^ n15319 ;
  assign n15499 = n5131 & ~n10205 ;
  assign n15500 = ( n4978 & n5041 ) | ( n4978 & ~n15499 ) | ( n5041 & ~n15499 ) ;
  assign n15501 = n6955 ^ n2549 ^ 1'b0 ;
  assign n15502 = n12963 & ~n15501 ;
  assign n15503 = n8253 | n9762 ;
  assign n15504 = n15502 | n15503 ;
  assign n15505 = n4141 & ~n8164 ;
  assign n15506 = ~n14747 & n15505 ;
  assign n15509 = n10822 ^ n1733 ^ 1'b0 ;
  assign n15507 = n2376 & ~n4433 ;
  assign n15508 = ~n3739 & n15507 ;
  assign n15510 = n15509 ^ n15508 ^ n1276 ;
  assign n15511 = n10092 ^ n1292 ^ 1'b0 ;
  assign n15512 = ( n1879 & ~n7943 ) | ( n1879 & n11183 ) | ( ~n7943 & n11183 ) ;
  assign n15513 = ~n5460 & n15512 ;
  assign n15514 = n3736 & n4078 ;
  assign n15515 = n3360 & ~n4370 ;
  assign n15516 = n768 & ~n6546 ;
  assign n15517 = n15516 ^ n2715 ^ 1'b0 ;
  assign n15518 = n12229 & ~n15517 ;
  assign n15519 = n8199 | n15518 ;
  assign n15520 = n15519 ^ n3268 ^ 1'b0 ;
  assign n15521 = n9291 ^ n401 ^ 1'b0 ;
  assign n15522 = ~n4120 & n15521 ;
  assign n15523 = n5024 & n10780 ;
  assign n15524 = n4483 ^ n4123 ^ 1'b0 ;
  assign n15525 = n14175 ^ n8812 ^ n3561 ;
  assign n15526 = n1585 & n8695 ;
  assign n15527 = ~n4135 & n12484 ;
  assign n15528 = n12654 ^ n983 ^ 1'b0 ;
  assign n15529 = ~n15527 & n15528 ;
  assign n15530 = n15529 ^ n1485 ^ 1'b0 ;
  assign n15533 = n4545 & n5960 ;
  assign n15531 = ~n4661 & n11966 ;
  assign n15532 = n15531 ^ n3189 ^ n3047 ;
  assign n15534 = n15533 ^ n15532 ^ 1'b0 ;
  assign n15535 = n1564 & n15534 ;
  assign n15536 = ( ~n3045 & n9457 ) | ( ~n3045 & n15535 ) | ( n9457 & n15535 ) ;
  assign n15537 = n12446 ^ n4605 ^ 1'b0 ;
  assign n15538 = n12308 ^ n5024 ^ n403 ;
  assign n15539 = n13936 ^ n2578 ^ 1'b0 ;
  assign n15540 = n15538 & ~n15539 ;
  assign n15541 = n8966 ^ n6566 ^ 1'b0 ;
  assign n15542 = n12650 & ~n15541 ;
  assign n15543 = n6961 | n13439 ;
  assign n15544 = n15543 ^ n4392 ^ 1'b0 ;
  assign n15548 = ( n3560 & ~n6146 ) | ( n3560 & n9661 ) | ( ~n6146 & n9661 ) ;
  assign n15549 = n3229 ^ n1223 ^ n197 ;
  assign n15550 = n2416 ^ n1212 ^ 1'b0 ;
  assign n15551 = n15549 & n15550 ;
  assign n15552 = n15548 & n15551 ;
  assign n15553 = n15552 ^ n7402 ^ 1'b0 ;
  assign n15554 = n15553 ^ n9236 ^ n4215 ;
  assign n15545 = n404 & ~n5160 ;
  assign n15546 = n15545 ^ n1467 ^ 1'b0 ;
  assign n15547 = n12425 & ~n15546 ;
  assign n15555 = n15554 ^ n15547 ^ 1'b0 ;
  assign n15556 = n8437 ^ n6399 ^ 1'b0 ;
  assign n15557 = ~n539 & n15556 ;
  assign n15558 = n8468 | n12403 ;
  assign n15559 = n15558 ^ n3955 ^ 1'b0 ;
  assign n15560 = n15559 ^ n11996 ^ n10884 ;
  assign n15561 = n633 & n1025 ;
  assign n15562 = ~x116 & n15561 ;
  assign n15563 = n4138 | n15562 ;
  assign n15564 = ( n349 & ~n1832 ) | ( n349 & n3179 ) | ( ~n1832 & n3179 ) ;
  assign n15565 = n15564 ^ n6683 ^ n1146 ;
  assign n15566 = n10020 ^ n1423 ^ 1'b0 ;
  assign n15567 = n15566 ^ n270 ^ 1'b0 ;
  assign n15568 = n15565 & ~n15567 ;
  assign n15569 = n8966 & ~n11612 ;
  assign n15570 = n15569 ^ n7252 ^ 1'b0 ;
  assign n15571 = ( n15563 & n15568 ) | ( n15563 & n15570 ) | ( n15568 & n15570 ) ;
  assign n15572 = ( ~n2363 & n4422 ) | ( ~n2363 & n14757 ) | ( n4422 & n14757 ) ;
  assign n15573 = n6230 ^ n3621 ^ 1'b0 ;
  assign n15574 = n5457 & ~n15573 ;
  assign n15575 = ~n10127 & n13172 ;
  assign n15576 = ~n11733 & n15575 ;
  assign n15577 = n8624 | n15576 ;
  assign n15578 = n15574 | n15577 ;
  assign n15579 = n5476 & ~n11612 ;
  assign n15580 = n15579 ^ n15397 ^ n7913 ;
  assign n15581 = n3719 ^ n901 ^ 1'b0 ;
  assign n15582 = n7024 ^ n2872 ^ 1'b0 ;
  assign n15583 = n11005 | n15582 ;
  assign n15584 = n15581 & ~n15583 ;
  assign n15585 = ~n495 & n15584 ;
  assign n15586 = ( n1423 & n15580 ) | ( n1423 & ~n15585 ) | ( n15580 & ~n15585 ) ;
  assign n15587 = n8323 ^ n914 ^ 1'b0 ;
  assign n15588 = n5390 ^ n2682 ^ 1'b0 ;
  assign n15589 = n1080 | n15588 ;
  assign n15590 = n2836 & ~n8942 ;
  assign n15591 = n15590 ^ n7965 ^ 1'b0 ;
  assign n15592 = n7992 | n12618 ;
  assign n15593 = n15592 ^ n11119 ^ 1'b0 ;
  assign n15595 = n14379 ^ n9627 ^ 1'b0 ;
  assign n15594 = ~n439 & n9336 ;
  assign n15596 = n15595 ^ n15594 ^ 1'b0 ;
  assign n15597 = n13830 | n15596 ;
  assign n15598 = n15593 | n15597 ;
  assign n15599 = ~n2085 & n12990 ;
  assign n15600 = n14249 & n15599 ;
  assign n15601 = n9194 & ~n15600 ;
  assign n15602 = n13279 ^ n9146 ^ n1789 ;
  assign n15603 = n15602 ^ n13105 ^ 1'b0 ;
  assign n15604 = n522 | n10343 ;
  assign n15605 = n15604 ^ n7542 ^ 1'b0 ;
  assign n15606 = ( n3340 & n10481 ) | ( n3340 & ~n13924 ) | ( n10481 & ~n13924 ) ;
  assign n15607 = n15449 ^ n5102 ^ 1'b0 ;
  assign n15608 = n15606 & n15607 ;
  assign n15609 = n15608 ^ n6799 ^ 1'b0 ;
  assign n15612 = n2442 ^ n2022 ^ n436 ;
  assign n15613 = n760 | n15612 ;
  assign n15614 = n15613 ^ n8385 ^ n7669 ;
  assign n15610 = n7007 ^ n4605 ^ n4247 ;
  assign n15611 = n5713 | n15610 ;
  assign n15615 = n15614 ^ n15611 ^ 1'b0 ;
  assign n15616 = n15615 ^ n9105 ^ n2331 ;
  assign n15617 = n7725 & n8310 ;
  assign n15618 = n349 & n15617 ;
  assign n15619 = n2386 & n15618 ;
  assign n15620 = n6555 & n10891 ;
  assign n15621 = n15619 & n15620 ;
  assign n15622 = n10116 ^ n2224 ^ 1'b0 ;
  assign n15623 = n2124 & ~n15622 ;
  assign n15624 = n830 | n1485 ;
  assign n15625 = n5661 | n15624 ;
  assign n15626 = n5796 ^ n315 ^ 1'b0 ;
  assign n15627 = n15625 & ~n15626 ;
  assign n15628 = n5086 & n15627 ;
  assign n15629 = n14511 ^ n8557 ^ n7241 ;
  assign n15630 = n8033 ^ x45 ^ 1'b0 ;
  assign n15631 = n2186 & ~n10045 ;
  assign n15632 = ~n3475 & n15631 ;
  assign n15633 = n15632 ^ n11231 ^ 1'b0 ;
  assign n15634 = n5052 ^ n2813 ^ 1'b0 ;
  assign n15635 = ( ~n306 & n9933 ) | ( ~n306 & n10127 ) | ( n9933 & n10127 ) ;
  assign n15636 = n5231 & ~n8073 ;
  assign n15637 = n7875 ^ n7388 ^ n996 ;
  assign n15638 = n4228 ^ n1925 ^ 1'b0 ;
  assign n15639 = n4658 ^ n2354 ^ 1'b0 ;
  assign n15640 = n15639 ^ n11010 ^ 1'b0 ;
  assign n15641 = ~n2518 & n15640 ;
  assign n15642 = n5314 & n15641 ;
  assign n15643 = n7444 ^ n1044 ^ 1'b0 ;
  assign n15644 = ~n680 & n15643 ;
  assign n15645 = n3303 ^ n2141 ^ n360 ;
  assign n15646 = n7693 ^ n5606 ^ 1'b0 ;
  assign n15647 = n6893 | n15646 ;
  assign n15648 = ~n15645 & n15647 ;
  assign n15650 = ( n1405 & n8467 ) | ( n1405 & n9785 ) | ( n8467 & n9785 ) ;
  assign n15651 = ( n264 & n1205 ) | ( n264 & ~n1663 ) | ( n1205 & ~n1663 ) ;
  assign n15652 = n4424 | n15651 ;
  assign n15653 = n15650 | n15652 ;
  assign n15649 = n2189 & n3740 ;
  assign n15654 = n15653 ^ n15649 ^ 1'b0 ;
  assign n15655 = n15654 ^ n11467 ^ 1'b0 ;
  assign n15656 = n15648 & n15655 ;
  assign n15657 = n14767 ^ n13864 ^ n2848 ;
  assign n15658 = n1898 & n1978 ;
  assign n15659 = ~n5771 & n15658 ;
  assign n15660 = n15659 ^ n7520 ^ n1471 ;
  assign n15661 = n4329 ^ n3311 ^ 1'b0 ;
  assign n15662 = n1243 | n9132 ;
  assign n15663 = n15662 ^ n6303 ^ 1'b0 ;
  assign n15664 = n2172 & n15663 ;
  assign n15665 = ( n12766 & n15661 ) | ( n12766 & n15664 ) | ( n15661 & n15664 ) ;
  assign n15666 = n6575 ^ n1882 ^ n646 ;
  assign n15667 = n7913 | n15666 ;
  assign n15668 = n1949 | n10564 ;
  assign n15669 = ~n1260 & n3722 ;
  assign n15670 = n15669 ^ n2569 ^ 1'b0 ;
  assign n15671 = n3239 | n15670 ;
  assign n15672 = ~n13571 & n15671 ;
  assign n15673 = n12473 ^ n4008 ^ 1'b0 ;
  assign n15674 = n15673 ^ n15212 ^ n5304 ;
  assign n15675 = n4279 ^ n3972 ^ 1'b0 ;
  assign n15676 = n15675 ^ n5428 ^ 1'b0 ;
  assign n15677 = ( ~n5563 & n11680 ) | ( ~n5563 & n15676 ) | ( n11680 & n15676 ) ;
  assign n15678 = ( n1295 & n3091 ) | ( n1295 & ~n15677 ) | ( n3091 & ~n15677 ) ;
  assign n15679 = n9063 ^ n7455 ^ 1'b0 ;
  assign n15680 = n4972 ^ n654 ^ 1'b0 ;
  assign n15681 = n15680 ^ n14066 ^ 1'b0 ;
  assign n15682 = n5746 | n15681 ;
  assign n15683 = n15679 & ~n15682 ;
  assign n15685 = n15538 ^ n9388 ^ n2475 ;
  assign n15684 = n6088 | n7512 ;
  assign n15686 = n15685 ^ n15684 ^ 1'b0 ;
  assign n15687 = n2462 & ~n6469 ;
  assign n15688 = ( n1246 & ~n1936 ) | ( n1246 & n3311 ) | ( ~n1936 & n3311 ) ;
  assign n15689 = n14346 ^ n10002 ^ 1'b0 ;
  assign n15690 = n8665 & n14149 ;
  assign n15691 = ( n6624 & ~n9108 ) | ( n6624 & n11622 ) | ( ~n9108 & n11622 ) ;
  assign n15692 = n15691 ^ n11867 ^ n2178 ;
  assign n15693 = n2031 ^ n999 ^ 1'b0 ;
  assign n15694 = ~n3070 & n15693 ;
  assign n15695 = n15692 | n15694 ;
  assign n15696 = n921 & ~n10088 ;
  assign n15697 = n15696 ^ n9024 ^ 1'b0 ;
  assign n15698 = ( n781 & n2204 ) | ( n781 & n11231 ) | ( n2204 & n11231 ) ;
  assign n15699 = ~n1294 & n14432 ;
  assign n15700 = ~n4198 & n15699 ;
  assign n15701 = n10114 & ~n15700 ;
  assign n15702 = ~n15698 & n15701 ;
  assign n15703 = n12073 & ~n15669 ;
  assign n15704 = n15703 ^ n3349 ^ 1'b0 ;
  assign n15705 = n335 & ~n5502 ;
  assign n15706 = n15705 ^ n6164 ^ 1'b0 ;
  assign n15707 = ( n8482 & n11646 ) | ( n8482 & n15706 ) | ( n11646 & n15706 ) ;
  assign n15708 = n15707 ^ n5133 ^ 1'b0 ;
  assign n15709 = ~n15704 & n15708 ;
  assign n15710 = n1390 | n15709 ;
  assign n15711 = n12927 ^ n3421 ^ 1'b0 ;
  assign n15712 = n11614 ^ n9250 ^ 1'b0 ;
  assign n15713 = n12184 & ~n15712 ;
  assign n15714 = n1580 | n4884 ;
  assign n15715 = n14282 | n15714 ;
  assign n15716 = ~n1992 & n7671 ;
  assign n15717 = n13900 & n15716 ;
  assign n15718 = n15717 ^ n4018 ^ 1'b0 ;
  assign n15719 = n15718 ^ n14376 ^ n1921 ;
  assign n15720 = ( n6082 & n10056 ) | ( n6082 & n15719 ) | ( n10056 & n15719 ) ;
  assign n15721 = n11993 ^ n7646 ^ n7165 ;
  assign n15722 = n6805 ^ n2807 ^ 1'b0 ;
  assign n15723 = n15722 ^ n12427 ^ 1'b0 ;
  assign n15724 = n8440 & ~n8954 ;
  assign n15725 = ( n6252 & n15723 ) | ( n6252 & ~n15724 ) | ( n15723 & ~n15724 ) ;
  assign n15726 = n11326 ^ n5109 ^ 1'b0 ;
  assign n15727 = n3004 | n15726 ;
  assign n15728 = n7307 | n15727 ;
  assign n15729 = n15728 ^ n9402 ^ 1'b0 ;
  assign n15730 = n15729 ^ n12368 ^ 1'b0 ;
  assign n15731 = n6210 & ~n14966 ;
  assign n15732 = n15731 ^ n14066 ^ 1'b0 ;
  assign n15733 = n9721 ^ n9462 ^ 1'b0 ;
  assign n15734 = n5984 ^ n4762 ^ 1'b0 ;
  assign n15735 = n15733 | n15734 ;
  assign n15736 = n7562 | n15735 ;
  assign n15737 = n331 | n15736 ;
  assign n15738 = n15732 | n15737 ;
  assign n15743 = n14702 ^ n7643 ^ 1'b0 ;
  assign n15739 = n10647 ^ n559 ^ 1'b0 ;
  assign n15740 = n3766 | n15739 ;
  assign n15741 = n12603 | n15740 ;
  assign n15742 = ~n4628 & n15741 ;
  assign n15744 = n15743 ^ n15742 ^ 1'b0 ;
  assign n15745 = ~n3136 & n13664 ;
  assign n15746 = n5082 ^ n1747 ^ 1'b0 ;
  assign n15747 = n15746 ^ n7739 ^ n4232 ;
  assign n15748 = ~n4754 & n15747 ;
  assign n15749 = n4305 & n12231 ;
  assign n15750 = ~n3553 & n15749 ;
  assign n15759 = n2129 ^ n1000 ^ 1'b0 ;
  assign n15751 = n4952 ^ n2122 ^ 1'b0 ;
  assign n15752 = n9254 ^ n4660 ^ 1'b0 ;
  assign n15753 = ~n7049 & n15752 ;
  assign n15754 = ~n15751 & n15753 ;
  assign n15755 = n1301 | n15754 ;
  assign n15756 = n15755 ^ n293 ^ 1'b0 ;
  assign n15757 = ( n11747 & ~n13892 ) | ( n11747 & n15756 ) | ( ~n13892 & n15756 ) ;
  assign n15758 = n12421 & ~n15757 ;
  assign n15760 = n15759 ^ n15758 ^ 1'b0 ;
  assign n15761 = ( n981 & n7000 ) | ( n981 & n14776 ) | ( n7000 & n14776 ) ;
  assign n15762 = ( n8645 & ~n8808 ) | ( n8645 & n12001 ) | ( ~n8808 & n12001 ) ;
  assign n15763 = n15081 ^ n1704 ^ 1'b0 ;
  assign n15764 = n10462 ^ n7278 ^ 1'b0 ;
  assign n15765 = n9543 & n15764 ;
  assign n15766 = n15765 ^ n2787 ^ 1'b0 ;
  assign n15767 = n15763 & n15766 ;
  assign n15768 = n9657 ^ n6210 ^ 1'b0 ;
  assign n15769 = n4859 | n15768 ;
  assign n15770 = ( n11279 & n12657 ) | ( n11279 & n15769 ) | ( n12657 & n15769 ) ;
  assign n15771 = ( n11848 & n12381 ) | ( n11848 & n15770 ) | ( n12381 & n15770 ) ;
  assign n15772 = n10915 | n15771 ;
  assign n15773 = n3349 & ~n3409 ;
  assign n15774 = n2305 & n15773 ;
  assign n15778 = ( ~n618 & n4597 ) | ( ~n618 & n6402 ) | ( n4597 & n6402 ) ;
  assign n15776 = n6694 ^ n4190 ^ 1'b0 ;
  assign n15777 = ~n1496 & n15776 ;
  assign n15775 = n3010 ^ n2121 ^ 1'b0 ;
  assign n15779 = n15778 ^ n15777 ^ n15775 ;
  assign n15780 = ~n3200 & n6982 ;
  assign n15781 = n15780 ^ n885 ^ 1'b0 ;
  assign n15782 = ~n898 & n15781 ;
  assign n15783 = ( ~n3542 & n4895 ) | ( ~n3542 & n5782 ) | ( n4895 & n5782 ) ;
  assign n15784 = n15782 & ~n15783 ;
  assign n15786 = n2041 & n7000 ;
  assign n15787 = ~n14310 & n15786 ;
  assign n15788 = n15787 ^ n13634 ^ 1'b0 ;
  assign n15785 = n11226 ^ n9021 ^ 1'b0 ;
  assign n15789 = n15788 ^ n15785 ^ n3003 ;
  assign n15790 = n7806 ^ n436 ^ 1'b0 ;
  assign n15791 = n8298 & ~n15790 ;
  assign n15792 = n15791 ^ n8547 ^ 1'b0 ;
  assign n15793 = n6971 ^ n2147 ^ 1'b0 ;
  assign n15794 = ~n8042 & n15793 ;
  assign n15797 = n10531 ^ n9857 ^ n3496 ;
  assign n15798 = n15797 ^ n10627 ^ 1'b0 ;
  assign n15795 = n14831 ^ n9876 ^ n717 ;
  assign n15796 = ~n4156 & n15795 ;
  assign n15799 = n15798 ^ n15796 ^ 1'b0 ;
  assign n15800 = ( n161 & n7384 ) | ( n161 & n12269 ) | ( n7384 & n12269 ) ;
  assign n15801 = ( n3911 & n5788 ) | ( n3911 & ~n14942 ) | ( n5788 & ~n14942 ) ;
  assign n15802 = n3337 ^ n3016 ^ n707 ;
  assign n15803 = n10622 | n15802 ;
  assign n15804 = n15619 & ~n15803 ;
  assign n15805 = n15801 & ~n15804 ;
  assign n15806 = n15433 ^ n11886 ^ n6340 ;
  assign n15807 = n8922 & ~n15806 ;
  assign n15808 = n11004 ^ n9656 ^ n1833 ;
  assign n15809 = n5124 | n14023 ;
  assign n15810 = ( n984 & n2227 ) | ( n984 & ~n5883 ) | ( n2227 & ~n5883 ) ;
  assign n15811 = n15810 ^ n14482 ^ n8312 ;
  assign n15812 = n5114 ^ n3867 ^ 1'b0 ;
  assign n15813 = n10610 & ~n15812 ;
  assign n15814 = n5495 & n15813 ;
  assign n15815 = n352 | n9485 ;
  assign n15816 = n307 & ~n15815 ;
  assign n15817 = ~n2830 & n13332 ;
  assign n15818 = n2523 & ~n15817 ;
  assign n15819 = n15816 & n15818 ;
  assign n15820 = n7613 ^ n908 ^ 1'b0 ;
  assign n15821 = n15820 ^ n12304 ^ n384 ;
  assign n15822 = n6422 ^ n393 ^ n170 ;
  assign n15823 = n871 ^ x89 ^ 1'b0 ;
  assign n15824 = ( n2941 & ~n5748 ) | ( n2941 & n15823 ) | ( ~n5748 & n15823 ) ;
  assign n15825 = n15824 ^ n701 ^ 1'b0 ;
  assign n15826 = n6241 & n15825 ;
  assign n15827 = n5121 | n9528 ;
  assign n15828 = n15826 | n15827 ;
  assign n15829 = ( n11679 & n15822 ) | ( n11679 & n15828 ) | ( n15822 & n15828 ) ;
  assign n15830 = ( n2780 & n4445 ) | ( n2780 & n15829 ) | ( n4445 & n15829 ) ;
  assign n15831 = ( n676 & n2500 ) | ( n676 & ~n10995 ) | ( n2500 & ~n10995 ) ;
  assign n15832 = n15831 ^ n1628 ^ 1'b0 ;
  assign n15833 = ( n1590 & n5222 ) | ( n1590 & n5948 ) | ( n5222 & n5948 ) ;
  assign n15834 = x53 & ~n6557 ;
  assign n15835 = ( n6368 & ~n15833 ) | ( n6368 & n15834 ) | ( ~n15833 & n15834 ) ;
  assign n15836 = n1274 | n3872 ;
  assign n15837 = ~n3277 & n12376 ;
  assign n15838 = n15837 ^ n7430 ^ 1'b0 ;
  assign n15839 = n15836 & ~n15838 ;
  assign n15840 = ( n238 & ~n7040 ) | ( n238 & n7553 ) | ( ~n7040 & n7553 ) ;
  assign n15841 = n15840 ^ n5122 ^ n4187 ;
  assign n15842 = n9501 & n11286 ;
  assign n15843 = n15842 ^ n6858 ^ n570 ;
  assign n15844 = n8286 & ~n15843 ;
  assign n15845 = n10161 ^ n1816 ^ 1'b0 ;
  assign n15846 = ( ~n541 & n3991 ) | ( ~n541 & n10597 ) | ( n3991 & n10597 ) ;
  assign n15847 = n15846 ^ n14974 ^ n2096 ;
  assign n15848 = n15847 ^ n12146 ^ n4768 ;
  assign n15849 = n15848 ^ n11521 ^ n216 ;
  assign n15850 = n9972 ^ n3258 ^ n2599 ;
  assign n15851 = n10251 | n15850 ;
  assign n15852 = n15851 ^ n8396 ^ 1'b0 ;
  assign n15853 = n6003 ^ n5962 ^ 1'b0 ;
  assign n15854 = n8100 | n15853 ;
  assign n15855 = ( n448 & ~n5485 ) | ( n448 & n15854 ) | ( ~n5485 & n15854 ) ;
  assign n15856 = ~n14906 & n15855 ;
  assign n15860 = n2820 & ~n14966 ;
  assign n15857 = ~n289 & n752 ;
  assign n15858 = n15857 ^ n12491 ^ 1'b0 ;
  assign n15859 = n15858 ^ n4396 ^ 1'b0 ;
  assign n15861 = n15860 ^ n15859 ^ n6862 ;
  assign n15862 = n6871 ^ n2817 ^ 1'b0 ;
  assign n15863 = n10401 ^ n8544 ^ n2962 ;
  assign n15864 = n10364 & ~n15863 ;
  assign n15865 = n15864 ^ n12123 ^ 1'b0 ;
  assign n15866 = ( n8808 & n15862 ) | ( n8808 & ~n15865 ) | ( n15862 & ~n15865 ) ;
  assign n15867 = n13082 ^ n2640 ^ n2243 ;
  assign n15868 = n1078 & ~n3237 ;
  assign n15869 = n4792 | n6816 ;
  assign n15870 = n6119 & ~n15869 ;
  assign n15871 = n10278 & ~n15870 ;
  assign n15872 = n15868 & n15871 ;
  assign n15873 = n11272 ^ n1327 ^ 1'b0 ;
  assign n15874 = n15873 ^ n915 ^ 1'b0 ;
  assign n15875 = n2180 | n3130 ;
  assign n15876 = n15805 ^ n5145 ^ 1'b0 ;
  assign n15877 = n15875 | n15876 ;
  assign n15878 = n7252 ^ n6206 ^ n4701 ;
  assign n15879 = n4096 ^ n2304 ^ n1943 ;
  assign n15880 = n4992 & ~n7586 ;
  assign n15881 = ~n15879 & n15880 ;
  assign n15882 = x32 & n14561 ;
  assign n15883 = ( n14682 & ~n15881 ) | ( n14682 & n15882 ) | ( ~n15881 & n15882 ) ;
  assign n15884 = ( n4728 & ~n12585 ) | ( n4728 & n15883 ) | ( ~n12585 & n15883 ) ;
  assign n15885 = n15884 ^ n525 ^ 1'b0 ;
  assign n15886 = n6529 ^ n1397 ^ 1'b0 ;
  assign n15887 = ( ~n9866 & n10316 ) | ( ~n9866 & n15886 ) | ( n10316 & n15886 ) ;
  assign n15888 = n11246 ^ n7878 ^ n7285 ;
  assign n15889 = n15887 & n15888 ;
  assign n15890 = ( n10016 & n15786 ) | ( n10016 & n15868 ) | ( n15786 & n15868 ) ;
  assign n15895 = ~n951 & n7494 ;
  assign n15896 = n15895 ^ n298 ^ 1'b0 ;
  assign n15897 = n11498 & n15896 ;
  assign n15898 = n12260 & n14252 ;
  assign n15899 = ~n15897 & n15898 ;
  assign n15894 = ( x92 & ~n5805 ) | ( x92 & n9269 ) | ( ~n5805 & n9269 ) ;
  assign n15891 = ( ~n2288 & n2687 ) | ( ~n2288 & n10837 ) | ( n2687 & n10837 ) ;
  assign n15892 = n4341 | n15891 ;
  assign n15893 = n15892 ^ n6702 ^ n1469 ;
  assign n15900 = n15899 ^ n15894 ^ n15893 ;
  assign n15901 = n2692 & n6829 ;
  assign n15902 = n15901 ^ n4010 ^ 1'b0 ;
  assign n15903 = ( n2168 & n9830 ) | ( n2168 & n15902 ) | ( n9830 & n15902 ) ;
  assign n15904 = n13373 ^ n4993 ^ 1'b0 ;
  assign n15905 = n6271 & ~n15904 ;
  assign n15906 = n2970 & n7519 ;
  assign n15907 = n15906 ^ n214 ^ 1'b0 ;
  assign n15908 = n15482 ^ n14743 ^ 1'b0 ;
  assign n15909 = n1586 | n1902 ;
  assign n15910 = n15909 ^ n5760 ^ 1'b0 ;
  assign n15911 = n15910 ^ n8555 ^ n3578 ;
  assign n15912 = n13714 ^ n8414 ^ n6861 ;
  assign n15913 = n11599 ^ n980 ^ 1'b0 ;
  assign n15914 = n11865 & n15913 ;
  assign n15915 = ~n2152 & n15914 ;
  assign n15916 = ~x77 & n5159 ;
  assign n15917 = n15916 ^ n11721 ^ 1'b0 ;
  assign n15918 = ( n1038 & n1717 ) | ( n1038 & n5238 ) | ( n1717 & n5238 ) ;
  assign n15919 = n3444 & ~n6443 ;
  assign n15920 = n15918 & n15919 ;
  assign n15921 = ( n8286 & n10689 ) | ( n8286 & n15920 ) | ( n10689 & n15920 ) ;
  assign n15922 = n15921 ^ n9009 ^ 1'b0 ;
  assign n15923 = n13583 ^ n5679 ^ 1'b0 ;
  assign n15924 = n5382 | n15923 ;
  assign n15925 = n11401 ^ n9142 ^ n4231 ;
  assign n15926 = ~n15924 & n15925 ;
  assign n15927 = ~n3033 & n15926 ;
  assign n15928 = ( ~n2168 & n6382 ) | ( ~n2168 & n8942 ) | ( n6382 & n8942 ) ;
  assign n15929 = n15928 ^ n7594 ^ n2165 ;
  assign n15930 = n15929 ^ n2058 ^ x60 ;
  assign n15931 = n10213 | n15930 ;
  assign n15932 = n4881 | n6446 ;
  assign n15933 = n15932 ^ n9756 ^ n8196 ;
  assign n15934 = ( n6731 & n11329 ) | ( n6731 & ~n15614 ) | ( n11329 & ~n15614 ) ;
  assign n15935 = ~n8388 & n15934 ;
  assign n15936 = n393 & n9921 ;
  assign n15937 = n15936 ^ n11408 ^ n10137 ;
  assign n15938 = n5341 & n15937 ;
  assign n15939 = n15938 ^ n12905 ^ 1'b0 ;
  assign n15940 = ( x97 & n3905 ) | ( x97 & ~n7599 ) | ( n3905 & ~n7599 ) ;
  assign n15941 = n15940 ^ n14943 ^ n10465 ;
  assign n15942 = n393 & ~n1876 ;
  assign n15943 = n15942 ^ x85 ^ 1'b0 ;
  assign n15944 = n5030 | n8916 ;
  assign n15945 = n15944 ^ n4768 ^ 1'b0 ;
  assign n15952 = ~n9312 & n9558 ;
  assign n15946 = ~n237 & n2824 ;
  assign n15947 = n15946 ^ n386 ^ 1'b0 ;
  assign n15948 = n6057 ^ n1246 ^ 1'b0 ;
  assign n15949 = n15947 | n15948 ;
  assign n15950 = n15949 ^ n11601 ^ n8249 ;
  assign n15951 = n15950 ^ n9473 ^ 1'b0 ;
  assign n15953 = n15952 ^ n15951 ^ n15477 ;
  assign n15954 = n14284 ^ n7009 ^ 1'b0 ;
  assign n15955 = n8622 & n15954 ;
  assign n15956 = n5104 & ~n15955 ;
  assign n15957 = n4226 ^ n4038 ^ n2713 ;
  assign n15958 = n10000 ^ n7781 ^ n3689 ;
  assign n15959 = n15957 & ~n15958 ;
  assign n15960 = n5408 & n15959 ;
  assign n15961 = n2426 | n15960 ;
  assign n15962 = n6222 & ~n15961 ;
  assign n15963 = ( n6767 & ~n8410 ) | ( n6767 & n12727 ) | ( ~n8410 & n12727 ) ;
  assign n15964 = n8132 & n15963 ;
  assign n15965 = ( n2056 & ~n7326 ) | ( n2056 & n10360 ) | ( ~n7326 & n10360 ) ;
  assign n15966 = ~n1203 & n11808 ;
  assign n15967 = ~x73 & n9239 ;
  assign n15968 = n15967 ^ n14575 ^ x111 ;
  assign n15969 = ( ~n13045 & n15966 ) | ( ~n13045 & n15968 ) | ( n15966 & n15968 ) ;
  assign n15970 = n14883 ^ n12148 ^ n3154 ;
  assign n15971 = n15970 ^ n15115 ^ 1'b0 ;
  assign n15972 = n15971 ^ n6970 ^ 1'b0 ;
  assign n15973 = n12195 | n15972 ;
  assign n15974 = n2955 | n6166 ;
  assign n15975 = n15974 ^ n1388 ^ 1'b0 ;
  assign n15976 = ~n3909 & n15975 ;
  assign n15977 = n8765 | n13109 ;
  assign n15978 = n2354 & ~n15977 ;
  assign n15979 = ~n6553 & n13177 ;
  assign n15980 = n15978 & n15979 ;
  assign n15981 = n3856 ^ n2887 ^ n329 ;
  assign n15986 = n3710 & ~n4774 ;
  assign n15982 = n3332 & n12316 ;
  assign n15983 = n771 & ~n15982 ;
  assign n15984 = n5707 & n15983 ;
  assign n15985 = n4171 | n15984 ;
  assign n15987 = n15986 ^ n15985 ^ n1762 ;
  assign n15988 = ( n12225 & n15981 ) | ( n12225 & n15987 ) | ( n15981 & n15987 ) ;
  assign n15995 = n1456 ^ n1261 ^ 1'b0 ;
  assign n15993 = n8497 ^ n4270 ^ 1'b0 ;
  assign n15994 = ~n8135 & n15993 ;
  assign n15996 = n15995 ^ n15994 ^ 1'b0 ;
  assign n15989 = n5608 ^ n3493 ^ 1'b0 ;
  assign n15990 = n6123 | n15989 ;
  assign n15991 = n11615 ^ n7326 ^ n3721 ;
  assign n15992 = n15990 & n15991 ;
  assign n15997 = n15996 ^ n15992 ^ n10068 ;
  assign n16001 = n7855 ^ n1548 ^ 1'b0 ;
  assign n16002 = ~n4283 & n16001 ;
  assign n15998 = n4208 ^ n2326 ^ n926 ;
  assign n15999 = x46 | n1365 ;
  assign n16000 = ( n2937 & n15998 ) | ( n2937 & n15999 ) | ( n15998 & n15999 ) ;
  assign n16003 = n16002 ^ n16000 ^ n5032 ;
  assign n16004 = n1689 ^ x52 ^ 1'b0 ;
  assign n16006 = ( n1975 & n7874 ) | ( n1975 & n14001 ) | ( n7874 & n14001 ) ;
  assign n16007 = ( n320 & n10341 ) | ( n320 & n16006 ) | ( n10341 & n16006 ) ;
  assign n16005 = n14172 | n15704 ;
  assign n16008 = n16007 ^ n16005 ^ 1'b0 ;
  assign n16009 = n1159 | n9195 ;
  assign n16010 = n6424 & ~n16009 ;
  assign n16011 = ~n12535 & n16010 ;
  assign n16018 = n2296 & n9914 ;
  assign n16019 = n16018 ^ n12073 ^ 1'b0 ;
  assign n16015 = ( n6892 & n9152 ) | ( n6892 & n11566 ) | ( n9152 & n11566 ) ;
  assign n16016 = n16015 ^ n11922 ^ 1'b0 ;
  assign n16017 = ~n7822 & n16016 ;
  assign n16012 = n2313 ^ n157 ^ 1'b0 ;
  assign n16013 = n4614 & n16012 ;
  assign n16014 = n16013 ^ n14914 ^ n13266 ;
  assign n16020 = n16019 ^ n16017 ^ n16014 ;
  assign n16022 = n3378 ^ n714 ^ 1'b0 ;
  assign n16023 = ( n707 & n1381 ) | ( n707 & ~n16022 ) | ( n1381 & ~n16022 ) ;
  assign n16021 = ( ~n470 & n1208 ) | ( ~n470 & n1894 ) | ( n1208 & n1894 ) ;
  assign n16024 = n16023 ^ n16021 ^ n4857 ;
  assign n16025 = ( n3497 & n4449 ) | ( n3497 & ~n11007 ) | ( n4449 & ~n11007 ) ;
  assign n16026 = n5941 ^ n3040 ^ 1'b0 ;
  assign n16027 = x39 & ~n16026 ;
  assign n16028 = ( n16024 & n16025 ) | ( n16024 & n16027 ) | ( n16025 & n16027 ) ;
  assign n16032 = n5313 | n11086 ;
  assign n16029 = n7324 ^ n5899 ^ n1911 ;
  assign n16030 = n16029 ^ n6773 ^ n747 ;
  assign n16031 = ( n1092 & n3654 ) | ( n1092 & n16030 ) | ( n3654 & n16030 ) ;
  assign n16033 = n16032 ^ n16031 ^ n3137 ;
  assign n16034 = n1851 | n9371 ;
  assign n16035 = n16034 ^ n1466 ^ 1'b0 ;
  assign n16036 = n8699 | n16035 ;
  assign n16037 = n16036 ^ n15719 ^ 1'b0 ;
  assign n16038 = n846 & ~n16037 ;
  assign n16039 = ~n1824 & n2394 ;
  assign n16040 = n16039 ^ n7830 ^ 1'b0 ;
  assign n16041 = ~n5492 & n5500 ;
  assign n16042 = ~n12793 & n16041 ;
  assign n16043 = n10623 ^ n3255 ^ x59 ;
  assign n16044 = n11226 & ~n16043 ;
  assign n16045 = n16044 ^ n2372 ^ 1'b0 ;
  assign n16046 = ( n5654 & n16042 ) | ( n5654 & ~n16045 ) | ( n16042 & ~n16045 ) ;
  assign n16047 = n7526 ^ n6637 ^ n527 ;
  assign n16051 = n2161 & n10467 ;
  assign n16052 = n13590 | n16051 ;
  assign n16053 = n2495 | n16052 ;
  assign n16048 = n2568 ^ n188 ^ 1'b0 ;
  assign n16049 = ( n4111 & n15850 ) | ( n4111 & ~n16048 ) | ( n15850 & ~n16048 ) ;
  assign n16050 = n3010 & ~n16049 ;
  assign n16054 = n16053 ^ n16050 ^ 1'b0 ;
  assign n16055 = n854 | n10416 ;
  assign n16056 = n16055 ^ n13214 ^ 1'b0 ;
  assign n16057 = ~n3440 & n5819 ;
  assign n16058 = n12560 & n16057 ;
  assign n16059 = n16058 ^ n15136 ^ n13055 ;
  assign n16060 = n3923 & ~n14505 ;
  assign n16061 = n8542 & n16060 ;
  assign n16062 = n15509 ^ n13150 ^ 1'b0 ;
  assign n16063 = ~n1740 & n16062 ;
  assign n16064 = n16063 ^ n8316 ^ n8100 ;
  assign n16065 = n11150 ^ n8133 ^ 1'b0 ;
  assign n16066 = n10140 & n10249 ;
  assign n16067 = n10822 ^ n2445 ^ 1'b0 ;
  assign n16068 = n14833 | n16067 ;
  assign n16069 = n16068 ^ n4731 ^ 1'b0 ;
  assign n16070 = x19 & ~n9813 ;
  assign n16071 = ~n16069 & n16070 ;
  assign n16072 = n7417 ^ n144 ^ 1'b0 ;
  assign n16073 = ( n5014 & n16071 ) | ( n5014 & ~n16072 ) | ( n16071 & ~n16072 ) ;
  assign n16074 = ( ~n474 & n5139 ) | ( ~n474 & n5801 ) | ( n5139 & n5801 ) ;
  assign n16075 = n3525 | n9312 ;
  assign n16076 = n1952 & n5765 ;
  assign n16077 = n16076 ^ n13639 ^ 1'b0 ;
  assign n16078 = n4022 & n16077 ;
  assign n16079 = n4588 & n16078 ;
  assign n16080 = n5349 ^ n1827 ^ 1'b0 ;
  assign n16081 = n3820 & n9860 ;
  assign n16082 = n2285 & ~n9002 ;
  assign n16083 = ~n11176 & n16082 ;
  assign n16084 = n1620 | n6075 ;
  assign n16085 = n15028 ^ n2355 ^ 1'b0 ;
  assign n16086 = n10987 | n16085 ;
  assign n16087 = n617 & n15813 ;
  assign n16088 = n16086 & n16087 ;
  assign n16089 = n5450 | n7568 ;
  assign n16090 = n16089 ^ n9028 ^ 1'b0 ;
  assign n16091 = n16090 ^ n5024 ^ 1'b0 ;
  assign n16092 = n14028 ^ n13185 ^ n7955 ;
  assign n16097 = n4370 ^ n2567 ^ 1'b0 ;
  assign n16093 = ~n454 & n3985 ;
  assign n16094 = n16093 ^ n198 ^ 1'b0 ;
  assign n16095 = n866 & ~n1530 ;
  assign n16096 = n16094 | n16095 ;
  assign n16098 = n16097 ^ n16096 ^ n6287 ;
  assign n16099 = n12958 & n14308 ;
  assign n16100 = n3162 & n12306 ;
  assign n16101 = n7853 ^ n6194 ^ 1'b0 ;
  assign n16102 = n16101 ^ n4618 ^ n3625 ;
  assign n16103 = n5796 & n16102 ;
  assign n16104 = ( n1707 & ~n8393 ) | ( n1707 & n12750 ) | ( ~n8393 & n12750 ) ;
  assign n16105 = n12121 ^ n9965 ^ 1'b0 ;
  assign n16106 = n2963 & n8833 ;
  assign n16107 = n16106 ^ n3848 ^ n758 ;
  assign n16111 = n4073 ^ n182 ^ 1'b0 ;
  assign n16112 = ~n14310 & n16111 ;
  assign n16108 = n5885 ^ n5576 ^ n1666 ;
  assign n16109 = n16108 ^ n6759 ^ 1'b0 ;
  assign n16110 = n1767 & ~n16109 ;
  assign n16113 = n16112 ^ n16110 ^ 1'b0 ;
  assign n16114 = ( n4392 & n5056 ) | ( n4392 & ~n7661 ) | ( n5056 & ~n7661 ) ;
  assign n16115 = ( n4818 & n5699 ) | ( n4818 & n16114 ) | ( n5699 & n16114 ) ;
  assign n16116 = n9121 & ~n16115 ;
  assign n16117 = n5588 ^ n3895 ^ n1200 ;
  assign n16118 = ( n1135 & n7827 ) | ( n1135 & ~n16117 ) | ( n7827 & ~n16117 ) ;
  assign n16119 = n15165 ^ n7056 ^ 1'b0 ;
  assign n16121 = n5864 ^ n5023 ^ 1'b0 ;
  assign n16122 = ( n5439 & n5522 ) | ( n5439 & ~n16121 ) | ( n5522 & ~n16121 ) ;
  assign n16120 = n10004 | n11388 ;
  assign n16123 = n16122 ^ n16120 ^ 1'b0 ;
  assign n16124 = ( n9007 & ~n16119 ) | ( n9007 & n16123 ) | ( ~n16119 & n16123 ) ;
  assign n16126 = n4567 | n8554 ;
  assign n16127 = n16126 ^ n3595 ^ 1'b0 ;
  assign n16128 = n16127 ^ n10970 ^ n3991 ;
  assign n16125 = ~n1992 & n15795 ;
  assign n16129 = n16128 ^ n16125 ^ 1'b0 ;
  assign n16130 = ~n3527 & n9003 ;
  assign n16131 = ~n2425 & n8336 ;
  assign n16132 = n16131 ^ n7929 ^ 1'b0 ;
  assign n16133 = n16132 ^ n13127 ^ 1'b0 ;
  assign n16134 = ( n6353 & n7779 ) | ( n6353 & n16133 ) | ( n7779 & n16133 ) ;
  assign n16135 = n3639 ^ n2805 ^ n2723 ;
  assign n16140 = n8763 ^ n5139 ^ n2743 ;
  assign n16138 = n3917 ^ n2292 ^ 1'b0 ;
  assign n16139 = n3727 | n16138 ;
  assign n16136 = n7096 ^ n4216 ^ n3848 ;
  assign n16137 = ( n8616 & n11222 ) | ( n8616 & n16136 ) | ( n11222 & n16136 ) ;
  assign n16141 = n16140 ^ n16139 ^ n16137 ;
  assign n16142 = ( ~n307 & n16135 ) | ( ~n307 & n16141 ) | ( n16135 & n16141 ) ;
  assign n16143 = n3393 ^ n2408 ^ 1'b0 ;
  assign n16144 = n1422 | n16143 ;
  assign n16145 = n10249 ^ n6124 ^ n2917 ;
  assign n16146 = n16145 ^ n7085 ^ n2029 ;
  assign n16147 = n16146 ^ n7215 ^ n2363 ;
  assign n16148 = n16147 ^ n7988 ^ 1'b0 ;
  assign n16149 = ( n5449 & n6768 ) | ( n5449 & ~n7144 ) | ( n6768 & ~n7144 ) ;
  assign n16150 = n16149 ^ n1173 ^ n866 ;
  assign n16151 = ( n473 & n627 ) | ( n473 & n9585 ) | ( n627 & n9585 ) ;
  assign n16152 = ( n11239 & n16150 ) | ( n11239 & n16151 ) | ( n16150 & n16151 ) ;
  assign n16153 = n3996 & n6384 ;
  assign n16154 = ( n1726 & n10760 ) | ( n1726 & ~n16153 ) | ( n10760 & ~n16153 ) ;
  assign n16155 = n16154 ^ n5524 ^ 1'b0 ;
  assign n16156 = ( n2344 & n6311 ) | ( n2344 & n12132 ) | ( n6311 & n12132 ) ;
  assign n16157 = n5356 & n16156 ;
  assign n16158 = ~n4789 & n16157 ;
  assign n16159 = ~n4839 & n9194 ;
  assign n16160 = n16158 & n16159 ;
  assign n16161 = n13902 ^ n2240 ^ 1'b0 ;
  assign n16162 = n2794 & n16161 ;
  assign n16163 = ~n2413 & n16162 ;
  assign n16164 = n16163 ^ n3106 ^ 1'b0 ;
  assign n16166 = n7171 ^ n5723 ^ 1'b0 ;
  assign n16167 = n4365 & n16166 ;
  assign n16168 = n16167 ^ n14055 ^ n7339 ;
  assign n16165 = n11250 ^ n903 ^ 1'b0 ;
  assign n16169 = n16168 ^ n16165 ^ 1'b0 ;
  assign n16170 = ~n8767 & n15150 ;
  assign n16171 = n3715 & n16170 ;
  assign n16172 = n16171 ^ n2784 ^ 1'b0 ;
  assign n16173 = x63 & n16172 ;
  assign n16175 = n13058 | n14644 ;
  assign n16174 = n4137 & n11962 ;
  assign n16176 = n16175 ^ n16174 ^ n12112 ;
  assign n16181 = ~n3585 & n9736 ;
  assign n16182 = n16181 ^ n3069 ^ 1'b0 ;
  assign n16183 = ( n3524 & n6338 ) | ( n3524 & ~n16182 ) | ( n6338 & ~n16182 ) ;
  assign n16177 = ~n1607 & n10373 ;
  assign n16178 = n16177 ^ n11731 ^ n6116 ;
  assign n16179 = n2359 & n16178 ;
  assign n16180 = n16179 ^ n11512 ^ 1'b0 ;
  assign n16184 = n16183 ^ n16180 ^ 1'b0 ;
  assign n16191 = ( ~n5900 & n9581 ) | ( ~n5900 & n11439 ) | ( n9581 & n11439 ) ;
  assign n16186 = ~n165 & n2576 ;
  assign n16187 = ~n4858 & n16186 ;
  assign n16185 = n491 & ~n1311 ;
  assign n16188 = n16187 ^ n16185 ^ 1'b0 ;
  assign n16189 = n751 & n2476 ;
  assign n16190 = ~n16188 & n16189 ;
  assign n16192 = n16191 ^ n16190 ^ n12646 ;
  assign n16193 = ~n2299 & n16192 ;
  assign n16194 = n16193 ^ n14672 ^ 1'b0 ;
  assign n16195 = n5257 & ~n15510 ;
  assign n16196 = n16195 ^ n1070 ^ 1'b0 ;
  assign n16197 = n3306 ^ n2432 ^ 1'b0 ;
  assign n16198 = ~n8052 & n16197 ;
  assign n16199 = n6546 ^ n1110 ^ 1'b0 ;
  assign n16200 = n7874 & ~n16199 ;
  assign n16201 = n6450 & n16200 ;
  assign n16202 = n16201 ^ n15261 ^ n1682 ;
  assign n16203 = n5649 & n7899 ;
  assign n16204 = ( n1009 & n7992 ) | ( n1009 & ~n16203 ) | ( n7992 & ~n16203 ) ;
  assign n16205 = ( x13 & ~n2400 ) | ( x13 & n3198 ) | ( ~n2400 & n3198 ) ;
  assign n16206 = n16205 ^ n14298 ^ n2142 ;
  assign n16207 = n6264 & n11462 ;
  assign n16208 = n16207 ^ n968 ^ 1'b0 ;
  assign n16209 = n4862 | n9628 ;
  assign n16210 = n16209 ^ n1296 ^ 1'b0 ;
  assign n16211 = n7229 ^ n5010 ^ 1'b0 ;
  assign n16212 = n10255 | n16211 ;
  assign n16213 = ( n454 & n12004 ) | ( n454 & n16212 ) | ( n12004 & n16212 ) ;
  assign n16214 = n572 & ~n3728 ;
  assign n16215 = ( ~n3607 & n7536 ) | ( ~n3607 & n16214 ) | ( n7536 & n16214 ) ;
  assign n16216 = n12331 ^ n2030 ^ 1'b0 ;
  assign n16217 = n13752 ^ n8606 ^ 1'b0 ;
  assign n16218 = n9923 & ~n15629 ;
  assign n16219 = n16218 ^ n4048 ^ 1'b0 ;
  assign n16220 = n15836 ^ n5173 ^ 1'b0 ;
  assign n16221 = n16000 ^ n15984 ^ 1'b0 ;
  assign n16222 = ~n8368 & n10947 ;
  assign n16223 = n12556 ^ n964 ^ 1'b0 ;
  assign n16224 = n15395 ^ n14485 ^ 1'b0 ;
  assign n16225 = n13079 ^ n7301 ^ n2619 ;
  assign n16226 = n16225 ^ n15836 ^ n15596 ;
  assign n16227 = ~n137 & n9781 ;
  assign n16228 = ( n4521 & ~n15265 ) | ( n4521 & n16227 ) | ( ~n15265 & n16227 ) ;
  assign n16229 = ( ~n3616 & n6008 ) | ( ~n3616 & n9867 ) | ( n6008 & n9867 ) ;
  assign n16230 = n6284 ^ n3861 ^ n911 ;
  assign n16231 = n16229 & ~n16230 ;
  assign n16232 = n11855 ^ n3429 ^ 1'b0 ;
  assign n16233 = n14617 & ~n16232 ;
  assign n16234 = ( ~n2331 & n4085 ) | ( ~n2331 & n16233 ) | ( n4085 & n16233 ) ;
  assign n16235 = n15591 & n16234 ;
  assign n16236 = n14662 ^ n699 ^ 1'b0 ;
  assign n16237 = n4944 | n16236 ;
  assign n16238 = n2518 | n4819 ;
  assign n16239 = n5216 & ~n7729 ;
  assign n16240 = n7099 | n16239 ;
  assign n16241 = n16238 & ~n16240 ;
  assign n16242 = n4779 & ~n6816 ;
  assign n16243 = n16241 & n16242 ;
  assign n16244 = n8611 ^ n4489 ^ n2160 ;
  assign n16245 = n16244 ^ n14178 ^ 1'b0 ;
  assign n16246 = ( n1209 & ~n9594 ) | ( n1209 & n16245 ) | ( ~n9594 & n16245 ) ;
  assign n16247 = n15231 ^ n10414 ^ n8467 ;
  assign n16248 = n16168 ^ n2466 ^ 1'b0 ;
  assign n16249 = ( n7917 & n10858 ) | ( n7917 & ~n16248 ) | ( n10858 & ~n16248 ) ;
  assign n16250 = n3363 ^ n631 ^ 1'b0 ;
  assign n16251 = n2101 & ~n16250 ;
  assign n16252 = n8307 & n16251 ;
  assign n16253 = n9227 & n16252 ;
  assign n16254 = ( ~n9767 & n10549 ) | ( ~n9767 & n16253 ) | ( n10549 & n16253 ) ;
  assign n16255 = n8151 ^ n2932 ^ n983 ;
  assign n16256 = ( n2371 & ~n13647 ) | ( n2371 & n16255 ) | ( ~n13647 & n16255 ) ;
  assign n16257 = n16254 | n16256 ;
  assign n16258 = n1803 | n5272 ;
  assign n16259 = ~n7249 & n16258 ;
  assign n16260 = n16259 ^ n16014 ^ 1'b0 ;
  assign n16261 = n11101 ^ n8087 ^ 1'b0 ;
  assign n16262 = n7558 | n16261 ;
  assign n16263 = n16262 ^ n11889 ^ n1417 ;
  assign n16264 = ~n1230 & n15824 ;
  assign n16265 = n16264 ^ n12890 ^ 1'b0 ;
  assign n16266 = ( n2457 & n5434 ) | ( n2457 & ~n16265 ) | ( n5434 & ~n16265 ) ;
  assign n16267 = n6570 ^ n1572 ^ 1'b0 ;
  assign n16268 = n16266 & ~n16267 ;
  assign n16269 = ( n3357 & n10517 ) | ( n3357 & ~n16268 ) | ( n10517 & ~n16268 ) ;
  assign n16270 = n16269 ^ n6557 ^ n292 ;
  assign n16271 = n16270 ^ n1625 ^ 1'b0 ;
  assign n16272 = ~n388 & n7918 ;
  assign n16273 = n16272 ^ n11722 ^ 1'b0 ;
  assign n16274 = ~n10803 & n16273 ;
  assign n16276 = ~n2573 & n6420 ;
  assign n16277 = n16276 ^ n8572 ^ 1'b0 ;
  assign n16275 = n8140 | n8791 ;
  assign n16278 = n16277 ^ n16275 ^ n434 ;
  assign n16282 = n5108 ^ n442 ^ 1'b0 ;
  assign n16279 = ( n3932 & n4022 ) | ( n3932 & n10108 ) | ( n4022 & n10108 ) ;
  assign n16280 = ( ~x93 & n7455 ) | ( ~x93 & n16279 ) | ( n7455 & n16279 ) ;
  assign n16281 = ~n1966 & n16280 ;
  assign n16283 = n16282 ^ n16281 ^ 1'b0 ;
  assign n16284 = n8359 | n16283 ;
  assign n16285 = n7096 ^ n6495 ^ 1'b0 ;
  assign n16286 = n2884 ^ n2434 ^ 1'b0 ;
  assign n16287 = n4825 | n16286 ;
  assign n16288 = ( n5560 & n7318 ) | ( n5560 & ~n16287 ) | ( n7318 & ~n16287 ) ;
  assign n16289 = n4550 ^ n3657 ^ n559 ;
  assign n16290 = n10368 ^ n1499 ^ 1'b0 ;
  assign n16291 = n16289 & ~n16290 ;
  assign n16292 = ( x107 & n16288 ) | ( x107 & ~n16291 ) | ( n16288 & ~n16291 ) ;
  assign n16293 = n16292 ^ n2572 ^ 1'b0 ;
  assign n16295 = n4045 & n15894 ;
  assign n16294 = ~n3421 & n7216 ;
  assign n16296 = n16295 ^ n16294 ^ 1'b0 ;
  assign n16297 = n8879 ^ n6734 ^ 1'b0 ;
  assign n16298 = n1484 ^ n739 ^ 1'b0 ;
  assign n16299 = n4455 & ~n9256 ;
  assign n16300 = n3197 & n16299 ;
  assign n16303 = n3183 & ~n7706 ;
  assign n16301 = n5963 ^ n1598 ^ 1'b0 ;
  assign n16302 = n16301 ^ n12329 ^ 1'b0 ;
  assign n16304 = n16303 ^ n16302 ^ 1'b0 ;
  assign n16306 = n710 & n5666 ;
  assign n16307 = ( n4869 & n8630 ) | ( n4869 & ~n16306 ) | ( n8630 & ~n16306 ) ;
  assign n16305 = n4285 & n5453 ;
  assign n16308 = n16307 ^ n16305 ^ 1'b0 ;
  assign n16309 = ( n4544 & ~n16304 ) | ( n4544 & n16308 ) | ( ~n16304 & n16308 ) ;
  assign n16310 = n13507 ^ n8789 ^ n5791 ;
  assign n16311 = n16310 ^ n3136 ^ n1092 ;
  assign n16312 = n6388 & n8298 ;
  assign n16313 = n16312 ^ n4142 ^ 1'b0 ;
  assign n16314 = n4862 ^ n376 ^ 1'b0 ;
  assign n16315 = ~n8112 & n16314 ;
  assign n16316 = n16315 ^ n10494 ^ n5591 ;
  assign n16317 = ~n11920 & n16316 ;
  assign n16318 = ~n16313 & n16317 ;
  assign n16319 = n16318 ^ n15557 ^ 1'b0 ;
  assign n16320 = n8868 & ~n16319 ;
  assign n16321 = ( n6875 & ~n16311 ) | ( n6875 & n16320 ) | ( ~n16311 & n16320 ) ;
  assign n16322 = n13135 ^ n3424 ^ 1'b0 ;
  assign n16323 = ( ~n5080 & n5449 ) | ( ~n5080 & n9999 ) | ( n5449 & n9999 ) ;
  assign n16324 = n16323 ^ n14251 ^ n5102 ;
  assign n16325 = n1426 | n10359 ;
  assign n16326 = n5121 & ~n16325 ;
  assign n16327 = ( ~n3161 & n11644 ) | ( ~n3161 & n16326 ) | ( n11644 & n16326 ) ;
  assign n16328 = n9999 | n16327 ;
  assign n16329 = n16324 | n16328 ;
  assign n16330 = n3732 ^ n872 ^ 1'b0 ;
  assign n16331 = n12009 & n16330 ;
  assign n16332 = n16331 ^ n12066 ^ 1'b0 ;
  assign n16333 = n1261 & n4226 ;
  assign n16334 = n16333 ^ n458 ^ 1'b0 ;
  assign n16346 = x96 & ~n1581 ;
  assign n16338 = ( n2768 & ~n12525 ) | ( n2768 & n13204 ) | ( ~n12525 & n13204 ) ;
  assign n16339 = n9105 ^ n1735 ^ 1'b0 ;
  assign n16340 = n3929 & ~n16339 ;
  assign n16341 = n14650 ^ n327 ^ 1'b0 ;
  assign n16342 = n14058 & n16341 ;
  assign n16343 = ( x92 & n16340 ) | ( x92 & ~n16342 ) | ( n16340 & ~n16342 ) ;
  assign n16344 = ( n11614 & n16338 ) | ( n11614 & n16343 ) | ( n16338 & n16343 ) ;
  assign n16345 = n16344 ^ n12426 ^ n7700 ;
  assign n16335 = n1501 & ~n8699 ;
  assign n16336 = n328 & n16335 ;
  assign n16337 = ( n299 & ~n3812 ) | ( n299 & n16336 ) | ( ~n3812 & n16336 ) ;
  assign n16347 = n16346 ^ n16345 ^ n16337 ;
  assign n16348 = n5562 ^ n3032 ^ 1'b0 ;
  assign n16349 = n15376 ^ n3354 ^ 1'b0 ;
  assign n16350 = ~n16348 & n16349 ;
  assign n16351 = n16350 ^ n7617 ^ 1'b0 ;
  assign n16352 = n16351 ^ n5268 ^ n2481 ;
  assign n16353 = n16106 ^ n16022 ^ n9040 ;
  assign n16354 = n16353 ^ n9658 ^ n3802 ;
  assign n16355 = n12580 & ~n12730 ;
  assign n16356 = n16355 ^ n1861 ^ 1'b0 ;
  assign n16357 = n2572 | n16356 ;
  assign n16358 = n4660 & ~n14611 ;
  assign n16359 = n12578 ^ n12431 ^ n3513 ;
  assign n16360 = n2015 ^ n1221 ^ n420 ;
  assign n16361 = n9962 & ~n16360 ;
  assign n16362 = n16361 ^ n1433 ^ 1'b0 ;
  assign n16363 = ( n2122 & n4750 ) | ( n2122 & n16362 ) | ( n4750 & n16362 ) ;
  assign n16364 = n5903 & ~n16363 ;
  assign n16365 = n12147 ^ n11801 ^ n8071 ;
  assign n16366 = n14522 & ~n16365 ;
  assign n16367 = n2590 & ~n16366 ;
  assign n16368 = n16364 & n16367 ;
  assign n16369 = n3670 & n7960 ;
  assign n16370 = n16369 ^ n8765 ^ 1'b0 ;
  assign n16371 = n2740 & n16370 ;
  assign n16372 = n16371 ^ n6642 ^ n1057 ;
  assign n16373 = ( n4597 & ~n15468 ) | ( n4597 & n16372 ) | ( ~n15468 & n16372 ) ;
  assign n16374 = n4616 & n16373 ;
  assign n16375 = n11726 & n16374 ;
  assign n16376 = n4307 ^ n1916 ^ x41 ;
  assign n16377 = ( n3219 & ~n6477 ) | ( n3219 & n16376 ) | ( ~n6477 & n16376 ) ;
  assign n16378 = n4392 | n16377 ;
  assign n16379 = ~n10320 & n16378 ;
  assign n16380 = ~n2509 & n16379 ;
  assign n16381 = n920 & ~n16380 ;
  assign n16382 = ( n2524 & n6036 ) | ( n2524 & n14252 ) | ( n6036 & n14252 ) ;
  assign n16383 = n15281 ^ n5632 ^ n3770 ;
  assign n16384 = n11894 ^ n289 ^ 1'b0 ;
  assign n16385 = n4999 & ~n16384 ;
  assign n16386 = n354 & ~n5627 ;
  assign n16387 = ~n12761 & n16386 ;
  assign n16388 = n6793 | n16387 ;
  assign n16389 = n16385 | n16388 ;
  assign n16390 = n1986 ^ n1417 ^ 1'b0 ;
  assign n16391 = n10599 ^ n1959 ^ 1'b0 ;
  assign n16392 = n14545 & ~n16391 ;
  assign n16393 = ( n9541 & n10291 ) | ( n9541 & ~n11759 ) | ( n10291 & ~n11759 ) ;
  assign n16394 = ( n3896 & n6173 ) | ( n3896 & n8862 ) | ( n6173 & n8862 ) ;
  assign n16395 = n5706 & n16394 ;
  assign n16396 = ( n3493 & n4328 ) | ( n3493 & ~n7806 ) | ( n4328 & ~n7806 ) ;
  assign n16397 = ~n5079 & n16396 ;
  assign n16398 = n2416 ^ n1903 ^ 1'b0 ;
  assign n16399 = n16397 & n16398 ;
  assign n16400 = n16399 ^ n2088 ^ 1'b0 ;
  assign n16401 = n15614 & n16400 ;
  assign n16402 = ( n1129 & ~n1328 ) | ( n1129 & n15056 ) | ( ~n1328 & n15056 ) ;
  assign n16403 = n6802 ^ n851 ^ 1'b0 ;
  assign n16404 = n7494 ^ n5179 ^ n5148 ;
  assign n16405 = ~n1816 & n16404 ;
  assign n16406 = n8510 ^ n4807 ^ n211 ;
  assign n16407 = n6416 & n12295 ;
  assign n16408 = x50 & n15887 ;
  assign n16409 = ( n4152 & n16407 ) | ( n4152 & n16408 ) | ( n16407 & n16408 ) ;
  assign n16411 = n4742 ^ n4367 ^ 1'b0 ;
  assign n16410 = n7009 ^ n2901 ^ 1'b0 ;
  assign n16412 = n16411 ^ n16410 ^ n9056 ;
  assign n16413 = ( n3515 & ~n15832 ) | ( n3515 & n16412 ) | ( ~n15832 & n16412 ) ;
  assign n16414 = n2071 | n14283 ;
  assign n16415 = n16414 ^ n5395 ^ 1'b0 ;
  assign n16416 = n7489 & n16415 ;
  assign n16417 = n5675 & n16416 ;
  assign n16418 = ( n5961 & n6414 ) | ( n5961 & n8911 ) | ( n6414 & n8911 ) ;
  assign n16419 = n13381 & n16315 ;
  assign n16420 = n16419 ^ n5281 ^ 1'b0 ;
  assign n16421 = n13019 ^ n1597 ^ 1'b0 ;
  assign n16422 = n16421 ^ n9835 ^ n4561 ;
  assign n16423 = ~n7998 & n16422 ;
  assign n16424 = n13421 ^ n9230 ^ 1'b0 ;
  assign n16425 = n6466 | n16424 ;
  assign n16426 = n10109 ^ n8738 ^ 1'b0 ;
  assign n16427 = ( n7232 & n16313 ) | ( n7232 & n16426 ) | ( n16313 & n16426 ) ;
  assign n16428 = n11487 ^ x114 ^ 1'b0 ;
  assign n16429 = n12543 & n16428 ;
  assign n16430 = n887 & ~n2754 ;
  assign n16431 = n15461 ^ n1781 ^ n269 ;
  assign n16432 = n8844 ^ n1302 ^ 1'b0 ;
  assign n16433 = ~n6622 & n16432 ;
  assign n16434 = n512 & ~n1705 ;
  assign n16435 = n13522 & n16434 ;
  assign n16436 = ( ~n6229 & n16433 ) | ( ~n6229 & n16435 ) | ( n16433 & n16435 ) ;
  assign n16437 = ( n16430 & n16431 ) | ( n16430 & n16436 ) | ( n16431 & n16436 ) ;
  assign n16438 = n14042 ^ n3365 ^ 1'b0 ;
  assign n16439 = n3032 & ~n16438 ;
  assign n16440 = n13796 ^ n2666 ^ 1'b0 ;
  assign n16441 = ~n16230 & n16440 ;
  assign n16442 = n202 & n10989 ;
  assign n16443 = ~n4959 & n16442 ;
  assign n16444 = n16443 ^ n13220 ^ n7284 ;
  assign n16448 = ( n2936 & n4899 ) | ( n2936 & ~n7733 ) | ( n4899 & ~n7733 ) ;
  assign n16445 = ( x36 & x94 ) | ( x36 & n659 ) | ( x94 & n659 ) ;
  assign n16446 = ( n5280 & ~n5865 ) | ( n5280 & n16445 ) | ( ~n5865 & n16445 ) ;
  assign n16447 = n16446 ^ n12593 ^ n5866 ;
  assign n16449 = n16448 ^ n16447 ^ n13127 ;
  assign n16450 = n6304 & ~n6970 ;
  assign n16451 = ~n5647 & n16450 ;
  assign n16452 = n10232 | n11783 ;
  assign n16453 = n16452 ^ n8765 ^ 1'b0 ;
  assign n16454 = ~n1223 & n9331 ;
  assign n16455 = ~n5026 & n9161 ;
  assign n16456 = n485 & ~n16455 ;
  assign n16457 = n16456 ^ n10839 ^ 1'b0 ;
  assign n16458 = n11808 ^ n8916 ^ 1'b0 ;
  assign n16459 = n227 & ~n3467 ;
  assign n16460 = ~n2862 & n16459 ;
  assign n16461 = ~n2865 & n8578 ;
  assign n16462 = n16461 ^ n6956 ^ 1'b0 ;
  assign n16463 = ( n3515 & n12719 ) | ( n3515 & n16462 ) | ( n12719 & n16462 ) ;
  assign n16470 = ( n926 & n2019 ) | ( n926 & ~n2688 ) | ( n2019 & ~n2688 ) ;
  assign n16469 = ( n5949 & n10765 ) | ( n5949 & n11304 ) | ( n10765 & n11304 ) ;
  assign n16466 = n11420 ^ n2600 ^ 1'b0 ;
  assign n16467 = n6343 & ~n16466 ;
  assign n16464 = n8306 ^ n6590 ^ 1'b0 ;
  assign n16465 = n15103 & ~n16464 ;
  assign n16468 = n16467 ^ n16465 ^ 1'b0 ;
  assign n16471 = n16470 ^ n16469 ^ n16468 ;
  assign n16472 = ( ~n1083 & n3551 ) | ( ~n1083 & n4365 ) | ( n3551 & n4365 ) ;
  assign n16473 = ( ~n1611 & n4783 ) | ( ~n1611 & n6619 ) | ( n4783 & n6619 ) ;
  assign n16474 = n2776 & ~n9945 ;
  assign n16475 = n10417 & n16474 ;
  assign n16476 = n7478 & ~n16475 ;
  assign n16477 = n16473 & n16476 ;
  assign n16478 = n16065 | n16477 ;
  assign n16479 = n12916 | n16478 ;
  assign n16480 = n2400 & ~n11476 ;
  assign n16481 = n4262 & n16480 ;
  assign n16482 = ( ~n852 & n921 ) | ( ~n852 & n1165 ) | ( n921 & n1165 ) ;
  assign n16483 = n16482 ^ n13123 ^ n2031 ;
  assign n16484 = n10713 & n16483 ;
  assign n16485 = n16481 & n16484 ;
  assign n16486 = n16485 ^ n7197 ^ n5290 ;
  assign n16487 = n474 | n9971 ;
  assign n16488 = n16487 ^ n3935 ^ 1'b0 ;
  assign n16489 = ( n5798 & n10514 ) | ( n5798 & ~n16488 ) | ( n10514 & ~n16488 ) ;
  assign n16490 = n7657 & n15426 ;
  assign n16491 = n16490 ^ n15763 ^ 1'b0 ;
  assign n16492 = n298 & n3942 ;
  assign n16493 = ~n3874 & n16492 ;
  assign n16494 = ~n7649 & n9576 ;
  assign n16495 = n16494 ^ n15709 ^ 1'b0 ;
  assign n16496 = n5954 | n10642 ;
  assign n16497 = n11588 | n16496 ;
  assign n16501 = ( ~n5365 & n5418 ) | ( ~n5365 & n5610 ) | ( n5418 & n5610 ) ;
  assign n16502 = n16501 ^ n8522 ^ 1'b0 ;
  assign n16499 = n7318 ^ n6191 ^ 1'b0 ;
  assign n16498 = n12304 ^ n4438 ^ n1011 ;
  assign n16500 = n16499 ^ n16498 ^ 1'b0 ;
  assign n16503 = n16502 ^ n16500 ^ n14349 ;
  assign n16504 = n15639 ^ n1590 ^ n429 ;
  assign n16505 = ~n363 & n6946 ;
  assign n16506 = n5785 & n13467 ;
  assign n16508 = n10831 ^ x10 ^ 1'b0 ;
  assign n16509 = n5966 & n16508 ;
  assign n16507 = n10152 ^ n5742 ^ n4388 ;
  assign n16510 = n16509 ^ n16507 ^ x68 ;
  assign n16511 = n3926 & n8545 ;
  assign n16512 = ~n7094 & n11873 ;
  assign n16513 = n16512 ^ n3004 ^ 1'b0 ;
  assign n16514 = n7635 ^ n7489 ^ 1'b0 ;
  assign n16515 = n16514 ^ n7178 ^ 1'b0 ;
  assign n16516 = n7095 ^ n4805 ^ 1'b0 ;
  assign n16517 = n5900 | n7259 ;
  assign n16518 = n3288 & ~n16517 ;
  assign n16519 = n2511 ^ n1286 ^ n1175 ;
  assign n16520 = n2255 & n11648 ;
  assign n16521 = n16520 ^ n3265 ^ 1'b0 ;
  assign n16522 = n14618 ^ n11606 ^ 1'b0 ;
  assign n16523 = ~n16521 & n16522 ;
  assign n16524 = ( n7370 & ~n16519 ) | ( n7370 & n16523 ) | ( ~n16519 & n16523 ) ;
  assign n16525 = ~n506 & n5797 ;
  assign n16526 = n16525 ^ n7214 ^ 1'b0 ;
  assign n16527 = n9205 & n16526 ;
  assign n16528 = ( n6394 & n12862 ) | ( n6394 & n16527 ) | ( n12862 & n16527 ) ;
  assign n16529 = n2670 ^ x119 ^ 1'b0 ;
  assign n16530 = n4198 & ~n11658 ;
  assign n16531 = ~n298 & n16530 ;
  assign n16532 = n16531 ^ n16164 ^ 1'b0 ;
  assign n16533 = n9944 ^ n1400 ^ 1'b0 ;
  assign n16534 = n1658 & ~n16533 ;
  assign n16535 = n6609 ^ n2772 ^ 1'b0 ;
  assign n16536 = ( ~n2662 & n11848 ) | ( ~n2662 & n12308 ) | ( n11848 & n12308 ) ;
  assign n16537 = n1083 & n2190 ;
  assign n16538 = ~n2190 & n16537 ;
  assign n16539 = ( ~n3555 & n9964 ) | ( ~n3555 & n16538 ) | ( n9964 & n16538 ) ;
  assign n16541 = n5590 ^ n196 ^ 1'b0 ;
  assign n16540 = ~n9157 & n11992 ;
  assign n16542 = n16541 ^ n16540 ^ 1'b0 ;
  assign n16543 = n908 & n8516 ;
  assign n16544 = n10827 & n12872 ;
  assign n16545 = n16543 & n16544 ;
  assign n16546 = ( ~n1252 & n1974 ) | ( ~n1252 & n2389 ) | ( n1974 & n2389 ) ;
  assign n16547 = n2568 & ~n16546 ;
  assign n16548 = n2107 | n5954 ;
  assign n16549 = n10309 | n16548 ;
  assign n16550 = n16549 ^ n12559 ^ 1'b0 ;
  assign n16551 = n16547 | n16550 ;
  assign n16552 = n15465 ^ n11379 ^ n971 ;
  assign n16560 = n8297 | n15126 ;
  assign n16557 = n8616 ^ n2150 ^ 1'b0 ;
  assign n16558 = n16557 ^ n5020 ^ n669 ;
  assign n16553 = n1419 | n15126 ;
  assign n16554 = n16553 ^ n12966 ^ n335 ;
  assign n16555 = n3742 & ~n16554 ;
  assign n16556 = n14235 & n16555 ;
  assign n16559 = n16558 ^ n16556 ^ 1'b0 ;
  assign n16561 = n16560 ^ n16559 ^ n3447 ;
  assign n16562 = ~n7550 & n11777 ;
  assign n16563 = n16562 ^ n8061 ^ 1'b0 ;
  assign n16564 = n16563 ^ n13799 ^ n10415 ;
  assign n16565 = ~n15788 & n16564 ;
  assign n16566 = n16565 ^ x95 ^ 1'b0 ;
  assign n16567 = n6434 ^ n4764 ^ 1'b0 ;
  assign n16568 = n1493 | n16567 ;
  assign n16569 = ( ~n10491 & n15547 ) | ( ~n10491 & n15718 ) | ( n15547 & n15718 ) ;
  assign n16570 = n4653 ^ n248 ^ 1'b0 ;
  assign n16571 = ( n2718 & ~n8431 ) | ( n2718 & n16570 ) | ( ~n8431 & n16570 ) ;
  assign n16572 = n8434 ^ n5562 ^ n5132 ;
  assign n16576 = ( ~n2229 & n4589 ) | ( ~n2229 & n8885 ) | ( n4589 & n8885 ) ;
  assign n16573 = n14641 ^ n5915 ^ 1'b0 ;
  assign n16574 = n2522 & n16573 ;
  assign n16575 = ~n6861 & n16574 ;
  assign n16577 = n16576 ^ n16575 ^ 1'b0 ;
  assign n16578 = n16577 ^ n15547 ^ n5140 ;
  assign n16579 = n16350 | n16578 ;
  assign n16580 = n7300 | n16579 ;
  assign n16581 = ( n3161 & ~n8214 ) | ( n3161 & n16255 ) | ( ~n8214 & n16255 ) ;
  assign n16582 = ( n5116 & ~n8999 ) | ( n5116 & n12320 ) | ( ~n8999 & n12320 ) ;
  assign n16583 = n7722 ^ n7467 ^ 1'b0 ;
  assign n16584 = ~n6890 & n16583 ;
  assign n16585 = n16584 ^ n11162 ^ n596 ;
  assign n16586 = ( n4176 & n11307 ) | ( n4176 & n16585 ) | ( n11307 & n16585 ) ;
  assign n16587 = n8086 ^ n8026 ^ 1'b0 ;
  assign n16588 = n2023 & n7545 ;
  assign n16589 = ~n2539 & n16588 ;
  assign n16590 = ( n1925 & ~n16587 ) | ( n1925 & n16589 ) | ( ~n16587 & n16589 ) ;
  assign n16591 = ~n3645 & n4733 ;
  assign n16592 = ~n1740 & n16591 ;
  assign n16593 = ( ~n1273 & n10445 ) | ( ~n1273 & n16027 ) | ( n10445 & n16027 ) ;
  assign n16594 = n1598 & n2549 ;
  assign n16595 = n16594 ^ n5328 ^ 1'b0 ;
  assign n16596 = n1954 & n6294 ;
  assign n16597 = n2921 & n16596 ;
  assign n16598 = ( n5963 & ~n16595 ) | ( n5963 & n16597 ) | ( ~n16595 & n16597 ) ;
  assign n16599 = ( n9746 & n16593 ) | ( n9746 & n16598 ) | ( n16593 & n16598 ) ;
  assign n16600 = ( n3999 & ~n9464 ) | ( n3999 & n15820 ) | ( ~n9464 & n15820 ) ;
  assign n16601 = n8773 ^ n2145 ^ 1'b0 ;
  assign n16602 = ~n13151 & n16601 ;
  assign n16603 = n5184 & n16602 ;
  assign n16604 = ( x25 & n260 ) | ( x25 & ~n1146 ) | ( n260 & ~n1146 ) ;
  assign n16605 = n14788 & n16604 ;
  assign n16606 = ( n852 & n1444 ) | ( n852 & ~n8114 ) | ( n1444 & ~n8114 ) ;
  assign n16607 = n4960 | n16606 ;
  assign n16608 = n16607 ^ n6896 ^ 1'b0 ;
  assign n16609 = ~n5821 & n16608 ;
  assign n16610 = n8552 & n15129 ;
  assign n16611 = n16610 ^ n4538 ^ 1'b0 ;
  assign n16612 = ~n1063 & n2167 ;
  assign n16613 = ( x59 & n5291 ) | ( x59 & n16612 ) | ( n5291 & n16612 ) ;
  assign n16614 = n16613 ^ n8763 ^ 1'b0 ;
  assign n16615 = ( n16609 & n16611 ) | ( n16609 & ~n16614 ) | ( n16611 & ~n16614 ) ;
  assign n16617 = n3286 ^ n2660 ^ 1'b0 ;
  assign n16616 = n4482 & n5491 ;
  assign n16618 = n16617 ^ n16616 ^ 1'b0 ;
  assign n16619 = n16618 ^ n8277 ^ 1'b0 ;
  assign n16620 = n10557 & ~n16619 ;
  assign n16621 = n16620 ^ n16024 ^ n15570 ;
  assign n16622 = n16621 ^ n5990 ^ 1'b0 ;
  assign n16623 = n838 & ~n16622 ;
  assign n16624 = x32 & ~n13201 ;
  assign n16625 = n16624 ^ n16369 ^ 1'b0 ;
  assign n16626 = n16625 ^ n14961 ^ n14224 ;
  assign n16627 = ( n3919 & n4616 ) | ( n3919 & n5177 ) | ( n4616 & n5177 ) ;
  assign n16628 = n8112 | n16627 ;
  assign n16629 = n1791 ^ x84 ^ 1'b0 ;
  assign n16630 = n16629 ^ n10283 ^ 1'b0 ;
  assign n16631 = n478 | n16630 ;
  assign n16632 = n16631 ^ n11408 ^ 1'b0 ;
  assign n16633 = n4875 ^ n2110 ^ 1'b0 ;
  assign n16634 = n6457 | n16633 ;
  assign n16635 = n16634 ^ n1861 ^ 1'b0 ;
  assign n16636 = n2116 ^ n1837 ^ 1'b0 ;
  assign n16637 = n16215 & ~n16636 ;
  assign n16638 = ~n3028 & n11351 ;
  assign n16639 = n4810 | n13685 ;
  assign n16640 = n16639 ^ n14757 ^ 1'b0 ;
  assign n16641 = n7882 ^ n6457 ^ 1'b0 ;
  assign n16642 = ( n4294 & n10982 ) | ( n4294 & ~n16641 ) | ( n10982 & ~n16641 ) ;
  assign n16643 = ~n3948 & n6734 ;
  assign n16644 = n16643 ^ n12289 ^ n5208 ;
  assign n16645 = n14111 ^ n4492 ^ 1'b0 ;
  assign n16646 = n8597 ^ n6673 ^ n1730 ;
  assign n16647 = ( n2248 & ~n4684 ) | ( n2248 & n6547 ) | ( ~n4684 & n6547 ) ;
  assign n16648 = n7641 & ~n15854 ;
  assign n16649 = ( n16646 & ~n16647 ) | ( n16646 & n16648 ) | ( ~n16647 & n16648 ) ;
  assign n16650 = n10189 ^ n6562 ^ 1'b0 ;
  assign n16651 = n8126 ^ n2377 ^ 1'b0 ;
  assign n16652 = n851 & ~n9511 ;
  assign n16653 = n16651 & n16652 ;
  assign n16654 = ( n7311 & n12790 ) | ( n7311 & ~n13375 ) | ( n12790 & ~n13375 ) ;
  assign n16655 = ( n5390 & n16653 ) | ( n5390 & n16654 ) | ( n16653 & n16654 ) ;
  assign n16656 = n8555 ^ n1015 ^ 1'b0 ;
  assign n16657 = n4344 & n16656 ;
  assign n16658 = n16657 ^ n1837 ^ 1'b0 ;
  assign n16659 = ~n6562 & n15392 ;
  assign n16660 = n16659 ^ n14898 ^ 1'b0 ;
  assign n16661 = ( n10157 & n16614 ) | ( n10157 & ~n16660 ) | ( n16614 & ~n16660 ) ;
  assign n16662 = n2215 & ~n16661 ;
  assign n16663 = ( n9398 & ~n16658 ) | ( n9398 & n16662 ) | ( ~n16658 & n16662 ) ;
  assign n16667 = n12024 | n15509 ;
  assign n16664 = n7048 ^ n5057 ^ 1'b0 ;
  assign n16665 = ~n13328 & n16664 ;
  assign n16666 = ( n1556 & n8297 ) | ( n1556 & n16665 ) | ( n8297 & n16665 ) ;
  assign n16668 = n16667 ^ n16666 ^ n13440 ;
  assign n16669 = n16668 ^ n320 ^ 1'b0 ;
  assign n16670 = n8691 ^ n6309 ^ n1646 ;
  assign n16671 = n16670 ^ n7448 ^ n2801 ;
  assign n16672 = n13795 ^ n5766 ^ n5097 ;
  assign n16673 = n16672 ^ n15022 ^ n10812 ;
  assign n16674 = n16673 ^ n14901 ^ n1709 ;
  assign n16675 = n12590 ^ n7197 ^ 1'b0 ;
  assign n16676 = n1700 & n16675 ;
  assign n16677 = n16676 ^ n5680 ^ 1'b0 ;
  assign n16678 = n9336 & ~n16677 ;
  assign n16679 = ~n5711 & n11249 ;
  assign n16680 = n8812 ^ n7635 ^ n6189 ;
  assign n16681 = n7485 & n16680 ;
  assign n16682 = n11079 ^ n4285 ^ 1'b0 ;
  assign n16683 = n16681 & ~n16682 ;
  assign n16684 = n16683 ^ n3352 ^ 1'b0 ;
  assign n16685 = n11262 & n16684 ;
  assign n16686 = ~n16679 & n16685 ;
  assign n16687 = n12905 ^ n2290 ^ 1'b0 ;
  assign n16688 = n14579 ^ n4872 ^ n2187 ;
  assign n16689 = ~n10022 & n10556 ;
  assign n16690 = n16689 ^ n1635 ^ 1'b0 ;
  assign n16691 = ( ~n3678 & n4521 ) | ( ~n3678 & n5088 ) | ( n4521 & n5088 ) ;
  assign n16692 = n16691 ^ n6230 ^ 1'b0 ;
  assign n16693 = n3375 | n16692 ;
  assign n16694 = n4952 & ~n16693 ;
  assign n16695 = ~n16690 & n16694 ;
  assign n16697 = ~n1422 & n4121 ;
  assign n16696 = n4156 | n11307 ;
  assign n16698 = n16697 ^ n16696 ^ 1'b0 ;
  assign n16699 = x73 & n16698 ;
  assign n16700 = n620 & n16699 ;
  assign n16701 = n6611 | n16700 ;
  assign n16702 = n3388 & n12047 ;
  assign n16704 = n8954 ^ n6749 ^ n1083 ;
  assign n16705 = n8699 | n16704 ;
  assign n16706 = n16705 ^ n10136 ^ 1'b0 ;
  assign n16703 = ~n7504 & n7652 ;
  assign n16707 = n16706 ^ n16703 ^ 1'b0 ;
  assign n16708 = ~n8270 & n14162 ;
  assign n16709 = ~n301 & n16708 ;
  assign n16710 = n16709 ^ x57 ^ 1'b0 ;
  assign n16711 = n3707 & ~n11525 ;
  assign n16712 = n951 & n16711 ;
  assign n16713 = n295 | n10290 ;
  assign n16714 = n1194 & n3688 ;
  assign n16715 = ~n881 & n16714 ;
  assign n16716 = n12072 & ~n16715 ;
  assign n16719 = ( n776 & n9014 ) | ( n776 & n11250 ) | ( n9014 & n11250 ) ;
  assign n16717 = n12853 ^ n1964 ^ 1'b0 ;
  assign n16718 = ~n14037 & n16717 ;
  assign n16720 = n16719 ^ n16718 ^ n15788 ;
  assign n16721 = n607 & ~n3527 ;
  assign n16722 = n3527 & n16721 ;
  assign n16723 = ~n197 & n3864 ;
  assign n16724 = n16722 & n16723 ;
  assign n16725 = ( n4233 & ~n5441 ) | ( n4233 & n10830 ) | ( ~n5441 & n10830 ) ;
  assign n16726 = ~n1914 & n6475 ;
  assign n16727 = ~n16725 & n16726 ;
  assign n16728 = ( n4515 & n5769 ) | ( n4515 & n14064 ) | ( n5769 & n14064 ) ;
  assign n16729 = n8422 ^ n4378 ^ 1'b0 ;
  assign n16730 = n1264 & ~n16729 ;
  assign n16731 = ~n3491 & n16730 ;
  assign n16732 = n6085 & n16731 ;
  assign n16733 = ( n16727 & ~n16728 ) | ( n16727 & n16732 ) | ( ~n16728 & n16732 ) ;
  assign n16734 = n16733 ^ n1176 ^ 1'b0 ;
  assign n16735 = ~n560 & n4269 ;
  assign n16736 = n5216 & ~n16151 ;
  assign n16737 = ~n16735 & n16736 ;
  assign n16738 = n16737 ^ n15950 ^ n13660 ;
  assign n16739 = n16738 ^ n5343 ^ 1'b0 ;
  assign n16740 = ~n14500 & n16739 ;
  assign n16741 = n9845 ^ n9137 ^ n7362 ;
  assign n16742 = n5975 | n16741 ;
  assign n16743 = n16742 ^ n10610 ^ 1'b0 ;
  assign n16744 = n4658 & ~n10027 ;
  assign n16745 = n16744 ^ n1747 ^ 1'b0 ;
  assign n16746 = ( ~n2758 & n7622 ) | ( ~n2758 & n9363 ) | ( n7622 & n9363 ) ;
  assign n16747 = ( n2522 & n16745 ) | ( n2522 & n16746 ) | ( n16745 & n16746 ) ;
  assign n16748 = ( n4844 & ~n5364 ) | ( n4844 & n8632 ) | ( ~n5364 & n8632 ) ;
  assign n16749 = n9826 ^ n8393 ^ 1'b0 ;
  assign n16750 = n13928 | n16749 ;
  assign n16751 = n15788 ^ n6629 ^ n3360 ;
  assign n16752 = ( ~n840 & n16750 ) | ( ~n840 & n16751 ) | ( n16750 & n16751 ) ;
  assign n16753 = ( ~n7830 & n8429 ) | ( ~n7830 & n15035 ) | ( n8429 & n15035 ) ;
  assign n16754 = n990 | n13334 ;
  assign n16755 = n2199 ^ x26 ^ 1'b0 ;
  assign n16756 = n5904 | n16755 ;
  assign n16757 = ( n455 & n2893 ) | ( n455 & n16756 ) | ( n2893 & n16756 ) ;
  assign n16758 = ( n1902 & n14966 ) | ( n1902 & ~n16757 ) | ( n14966 & ~n16757 ) ;
  assign n16759 = n992 & ~n16758 ;
  assign n16760 = ~n16754 & n16759 ;
  assign n16761 = n16753 & n16760 ;
  assign n16762 = ( n1601 & n5944 ) | ( n1601 & n8334 ) | ( n5944 & n8334 ) ;
  assign n16765 = n451 & n4010 ;
  assign n16763 = n693 & ~n10622 ;
  assign n16764 = n16763 ^ n13407 ^ 1'b0 ;
  assign n16766 = n16765 ^ n16764 ^ n6457 ;
  assign n16767 = n1116 & ~n16766 ;
  assign n16768 = n16762 & n16767 ;
  assign n16769 = n2682 ^ n2262 ^ 1'b0 ;
  assign n16770 = ( n7898 & ~n14425 ) | ( n7898 & n16769 ) | ( ~n14425 & n16769 ) ;
  assign n16771 = n10214 ^ n3321 ^ 1'b0 ;
  assign n16772 = ( ~n1034 & n7725 ) | ( ~n1034 & n9443 ) | ( n7725 & n9443 ) ;
  assign n16773 = n16772 ^ n419 ^ x2 ;
  assign n16774 = n11480 ^ n3560 ^ n1065 ;
  assign n16775 = n16774 ^ n1277 ^ 1'b0 ;
  assign n16776 = n16578 ^ n13560 ^ 1'b0 ;
  assign n16777 = ~n325 & n14560 ;
  assign n16778 = n3382 & n16777 ;
  assign n16779 = n11362 ^ n7945 ^ n6564 ;
  assign n16780 = ( n9053 & n16778 ) | ( n9053 & n16779 ) | ( n16778 & n16779 ) ;
  assign n16781 = ~n13649 & n14514 ;
  assign n16782 = n16781 ^ n11280 ^ 1'b0 ;
  assign n16783 = ( n1505 & n9715 ) | ( n1505 & ~n16782 ) | ( n9715 & ~n16782 ) ;
  assign n16784 = n1067 & n4710 ;
  assign n16786 = n2254 & ~n2951 ;
  assign n16787 = n2346 & n16786 ;
  assign n16785 = ~n678 & n9347 ;
  assign n16788 = n16787 ^ n16785 ^ n10370 ;
  assign n16789 = n5800 ^ n4658 ^ 1'b0 ;
  assign n16790 = n5260 ^ n1176 ^ 1'b0 ;
  assign n16791 = n13862 ^ n9309 ^ n6051 ;
  assign n16792 = n13060 & n16441 ;
  assign n16793 = ~n16791 & n16792 ;
  assign n16794 = n4606 & n15330 ;
  assign n16795 = n16794 ^ n3721 ^ 1'b0 ;
  assign n16796 = n16795 ^ n5843 ^ 1'b0 ;
  assign n16797 = n12836 ^ n8126 ^ 1'b0 ;
  assign n16798 = n4819 & ~n16797 ;
  assign n16799 = ~n2207 & n7664 ;
  assign n16800 = n16799 ^ n2239 ^ 1'b0 ;
  assign n16801 = n7050 & ~n16800 ;
  assign n16802 = n5118 & ~n16191 ;
  assign n16803 = n16802 ^ n10123 ^ 1'b0 ;
  assign n16804 = ~n5221 & n16803 ;
  assign n16818 = n4403 | n15423 ;
  assign n16805 = n1785 & ~n7542 ;
  assign n16810 = n2915 | n10306 ;
  assign n16811 = n16810 ^ n8579 ^ n635 ;
  assign n16812 = n8121 & ~n16811 ;
  assign n16813 = ~n10587 & n16812 ;
  assign n16806 = ( n1273 & ~n4904 ) | ( n1273 & n12287 ) | ( ~n4904 & n12287 ) ;
  assign n16807 = n16806 ^ n2647 ^ n299 ;
  assign n16808 = n11881 & n16807 ;
  assign n16809 = ~n9074 & n16808 ;
  assign n16814 = n16813 ^ n16809 ^ 1'b0 ;
  assign n16815 = n16814 ^ n3020 ^ 1'b0 ;
  assign n16816 = n16805 | n16815 ;
  assign n16817 = n3837 | n16816 ;
  assign n16819 = n16818 ^ n16817 ^ 1'b0 ;
  assign n16820 = n16819 ^ n12539 ^ 1'b0 ;
  assign n16821 = ( n6029 & n9824 ) | ( n6029 & n10472 ) | ( n9824 & n10472 ) ;
  assign n16822 = n928 & ~n4920 ;
  assign n16823 = n9798 & n16822 ;
  assign n16824 = n1120 & n3501 ;
  assign n16825 = n16824 ^ n12508 ^ 1'b0 ;
  assign n16826 = n386 & n2658 ;
  assign n16827 = n2992 & n16826 ;
  assign n16828 = n3955 | n8056 ;
  assign n16829 = n16827 & ~n16828 ;
  assign n16832 = n14685 ^ n4615 ^ 1'b0 ;
  assign n16833 = ~n16727 & n16832 ;
  assign n16834 = n16833 ^ n4270 ^ 1'b0 ;
  assign n16830 = n1182 | n14684 ;
  assign n16831 = n16830 ^ n8941 ^ 1'b0 ;
  assign n16835 = n16834 ^ n16831 ^ n1120 ;
  assign n16836 = ( n1443 & n2077 ) | ( n1443 & n10249 ) | ( n2077 & n10249 ) ;
  assign n16840 = n8679 ^ n5106 ^ n984 ;
  assign n16841 = ( n511 & n942 ) | ( n511 & n3114 ) | ( n942 & n3114 ) ;
  assign n16842 = n7478 ^ n1852 ^ n294 ;
  assign n16843 = n16842 ^ n8926 ^ n232 ;
  assign n16844 = n16843 ^ n647 ^ 1'b0 ;
  assign n16845 = ~n16841 & n16844 ;
  assign n16846 = n16845 ^ n14672 ^ 1'b0 ;
  assign n16847 = n16840 & n16846 ;
  assign n16837 = n2794 & n3972 ;
  assign n16838 = n16837 ^ n4481 ^ 1'b0 ;
  assign n16839 = n7878 | n16838 ;
  assign n16848 = n16847 ^ n16839 ^ 1'b0 ;
  assign n16849 = ( ~n1543 & n6867 ) | ( ~n1543 & n16500 ) | ( n6867 & n16500 ) ;
  assign n16850 = n12321 ^ n6326 ^ 1'b0 ;
  assign n16851 = ~n11556 & n16850 ;
  assign n16852 = n8341 & n12310 ;
  assign n16853 = n11716 ^ n968 ^ 1'b0 ;
  assign n16854 = ~n3422 & n5041 ;
  assign n16855 = n16854 ^ n9179 ^ n7838 ;
  assign n16856 = ( n293 & ~n1312 ) | ( n293 & n5751 ) | ( ~n1312 & n5751 ) ;
  assign n16857 = n6046 & n14094 ;
  assign n16858 = ~n10074 & n16857 ;
  assign n16859 = ( ~n12585 & n16856 ) | ( ~n12585 & n16858 ) | ( n16856 & n16858 ) ;
  assign n16860 = ~n8597 & n16433 ;
  assign n16861 = n16860 ^ n15995 ^ 1'b0 ;
  assign n16866 = n7774 | n10172 ;
  assign n16867 = n14575 | n16866 ;
  assign n16862 = n7256 ^ n4334 ^ n2858 ;
  assign n16863 = n1834 & n11630 ;
  assign n16864 = n16862 & n16863 ;
  assign n16865 = n8722 & ~n16864 ;
  assign n16868 = n16867 ^ n16865 ^ 1'b0 ;
  assign n16870 = n3559 ^ n2022 ^ n1007 ;
  assign n16869 = n214 & ~n6091 ;
  assign n16871 = n16870 ^ n16869 ^ 1'b0 ;
  assign n16872 = ~n12298 & n16871 ;
  assign n16873 = n16872 ^ n15685 ^ 1'b0 ;
  assign n16874 = ~n13288 & n15770 ;
  assign n16875 = n5159 & n16787 ;
  assign n16876 = n10158 & ~n14230 ;
  assign n16877 = ( ~n6897 & n8067 ) | ( ~n6897 & n11272 ) | ( n8067 & n11272 ) ;
  assign n16878 = n2033 & ~n8497 ;
  assign n16879 = n3132 & n16878 ;
  assign n16880 = ~n2483 & n14292 ;
  assign n16881 = ( n12250 & ~n16879 ) | ( n12250 & n16880 ) | ( ~n16879 & n16880 ) ;
  assign n16882 = n16881 ^ n2149 ^ n1263 ;
  assign n16883 = ( n6655 & n16877 ) | ( n6655 & ~n16882 ) | ( n16877 & ~n16882 ) ;
  assign n16884 = n13038 ^ n2167 ^ 1'b0 ;
  assign n16885 = ~n243 & n16884 ;
  assign n16886 = ~n11759 & n16885 ;
  assign n16887 = n16886 ^ n16122 ^ 1'b0 ;
  assign n16890 = n5729 & ~n7368 ;
  assign n16888 = n2011 | n5358 ;
  assign n16889 = n7505 & ~n16888 ;
  assign n16891 = n16890 ^ n16889 ^ 1'b0 ;
  assign n16892 = n8314 ^ n3266 ^ 1'b0 ;
  assign n16893 = ~n16891 & n16892 ;
  assign n16894 = n869 ^ n466 ^ 1'b0 ;
  assign n16895 = n4415 & n16894 ;
  assign n16896 = ~n7621 & n16895 ;
  assign n16897 = n7022 & n16896 ;
  assign n16898 = n4010 & n4559 ;
  assign n16899 = ~n8997 & n16898 ;
  assign n16900 = n13755 ^ n10121 ^ 1'b0 ;
  assign n16902 = n11272 ^ n2918 ^ 1'b0 ;
  assign n16903 = ( n6731 & n7313 ) | ( n6731 & n16902 ) | ( n7313 & n16902 ) ;
  assign n16904 = n16903 ^ n9866 ^ n8961 ;
  assign n16901 = n1330 & ~n9996 ;
  assign n16905 = n16904 ^ n16901 ^ 1'b0 ;
  assign n16906 = n11483 ^ n3692 ^ 1'b0 ;
  assign n16907 = n5793 ^ n2399 ^ 1'b0 ;
  assign n16910 = n8017 ^ n3044 ^ n604 ;
  assign n16908 = n1488 & ~n13590 ;
  assign n16909 = n5338 & n16908 ;
  assign n16911 = n16910 ^ n16909 ^ n15566 ;
  assign n16912 = ~n5746 & n16415 ;
  assign n16913 = n16912 ^ n5229 ^ 1'b0 ;
  assign n16914 = n2263 ^ n1697 ^ 1'b0 ;
  assign n16915 = n2900 & ~n16914 ;
  assign n16916 = n16840 & n16915 ;
  assign n16917 = ~n13111 & n16916 ;
  assign n16921 = n12841 ^ n4633 ^ 1'b0 ;
  assign n16922 = n9082 | n16921 ;
  assign n16923 = n573 & ~n16922 ;
  assign n16924 = ~n10494 & n16923 ;
  assign n16918 = n4521 ^ n3096 ^ 1'b0 ;
  assign n16919 = n367 & n16918 ;
  assign n16920 = ( n7328 & n10543 ) | ( n7328 & ~n16919 ) | ( n10543 & ~n16919 ) ;
  assign n16925 = n16924 ^ n16920 ^ n14132 ;
  assign n16926 = ~n5948 & n14077 ;
  assign n16927 = n15757 ^ n2145 ^ 1'b0 ;
  assign n16930 = ( n6685 & ~n10605 ) | ( n6685 & n15993 ) | ( ~n10605 & n15993 ) ;
  assign n16928 = n1602 & ~n3030 ;
  assign n16929 = n16928 ^ n4448 ^ 1'b0 ;
  assign n16931 = n16930 ^ n16929 ^ n3972 ;
  assign n16932 = n4804 & ~n10575 ;
  assign n16933 = n4660 & n16932 ;
  assign n16934 = n16933 ^ n1302 ^ 1'b0 ;
  assign n16935 = ~n16931 & n16934 ;
  assign n16936 = n15884 & n16935 ;
  assign n16937 = n4569 ^ n2901 ^ 1'b0 ;
  assign n16938 = n16937 ^ n13207 ^ 1'b0 ;
  assign n16939 = ~n5796 & n8002 ;
  assign n16940 = n2200 ^ n679 ^ 1'b0 ;
  assign n16941 = ( n5403 & ~n9319 ) | ( n5403 & n9698 ) | ( ~n9319 & n9698 ) ;
  assign n16942 = ( ~n12721 & n16940 ) | ( ~n12721 & n16941 ) | ( n16940 & n16941 ) ;
  assign n16944 = n9679 ^ n3835 ^ n2785 ;
  assign n16945 = n16944 ^ n1469 ^ n599 ;
  assign n16946 = n16945 ^ n8672 ^ 1'b0 ;
  assign n16947 = n4808 & n16946 ;
  assign n16943 = n6932 & ~n11632 ;
  assign n16948 = n16947 ^ n16943 ^ 1'b0 ;
  assign n16949 = n16948 ^ n6859 ^ n6503 ;
  assign n16950 = n9473 | n15317 ;
  assign n16951 = n1902 & ~n16950 ;
  assign n16952 = n905 & ~n1400 ;
  assign n16953 = n16952 ^ n5124 ^ 1'b0 ;
  assign n16954 = n3521 ^ n2676 ^ n1089 ;
  assign n16955 = n7843 ^ n7492 ^ n1534 ;
  assign n16956 = ( n10491 & ~n16954 ) | ( n10491 & n16955 ) | ( ~n16954 & n16955 ) ;
  assign n16957 = n16956 ^ n10615 ^ 1'b0 ;
  assign n16958 = ( n3832 & n7772 ) | ( n3832 & n8407 ) | ( n7772 & n8407 ) ;
  assign n16961 = n2667 & ~n5675 ;
  assign n16962 = n16961 ^ n12589 ^ 1'b0 ;
  assign n16963 = n16962 ^ n15344 ^ 1'b0 ;
  assign n16959 = ( ~n219 & n1545 ) | ( ~n219 & n12832 ) | ( n1545 & n12832 ) ;
  assign n16960 = n11417 | n16959 ;
  assign n16964 = n16963 ^ n16960 ^ 1'b0 ;
  assign n16968 = n6175 ^ n3807 ^ 1'b0 ;
  assign n16965 = ~n5080 & n5436 ;
  assign n16966 = n16965 ^ n7024 ^ 1'b0 ;
  assign n16967 = ~n11157 & n16966 ;
  assign n16969 = n16968 ^ n16967 ^ 1'b0 ;
  assign n16970 = n11886 ^ n4889 ^ 1'b0 ;
  assign n16971 = n2827 & n16970 ;
  assign n16972 = ~n3428 & n7362 ;
  assign n16973 = n16972 ^ n11530 ^ 1'b0 ;
  assign n16974 = n16973 ^ n13997 ^ n1957 ;
  assign n16975 = n3946 & ~n3971 ;
  assign n16976 = n6451 & n16975 ;
  assign n16977 = n16976 ^ n13587 ^ n10156 ;
  assign n16982 = n2857 & ~n8288 ;
  assign n16983 = n16982 ^ n13145 ^ n2522 ;
  assign n16978 = x82 & n6268 ;
  assign n16979 = n15736 & n16978 ;
  assign n16980 = n10327 ^ n308 ^ 1'b0 ;
  assign n16981 = ( n12500 & n16979 ) | ( n12500 & n16980 ) | ( n16979 & n16980 ) ;
  assign n16984 = n16983 ^ n16981 ^ n2607 ;
  assign n16985 = ( ~n3062 & n5905 ) | ( ~n3062 & n6558 ) | ( n5905 & n6558 ) ;
  assign n16986 = n6291 ^ n4429 ^ 1'b0 ;
  assign n16987 = n5054 | n16986 ;
  assign n16988 = ~n3123 & n16987 ;
  assign n16990 = n633 ^ n404 ^ 1'b0 ;
  assign n16991 = ~n1441 & n16990 ;
  assign n16989 = n3278 ^ n2767 ^ n1973 ;
  assign n16992 = n16991 ^ n16989 ^ 1'b0 ;
  assign n16993 = n294 | n16992 ;
  assign n16994 = ~n6434 & n9878 ;
  assign n16995 = n16993 & n16994 ;
  assign n16996 = n9106 ^ n1378 ^ 1'b0 ;
  assign n16997 = ~n16995 & n16996 ;
  assign n16998 = ~n5184 & n15644 ;
  assign n16999 = n16998 ^ n4972 ^ 1'b0 ;
  assign n17000 = n1529 & ~n7490 ;
  assign n17001 = n6816 ^ n3235 ^ 1'b0 ;
  assign n17002 = n17000 | n17001 ;
  assign n17003 = n724 ^ n550 ^ 1'b0 ;
  assign n17004 = ( n8916 & ~n11942 ) | ( n8916 & n17003 ) | ( ~n11942 & n17003 ) ;
  assign n17005 = n7209 & n12966 ;
  assign n17006 = n15345 & n17005 ;
  assign n17007 = n17006 ^ n12936 ^ x120 ;
  assign n17008 = n4772 & ~n7707 ;
  assign n17009 = n11044 | n17008 ;
  assign n17010 = ~n3637 & n10557 ;
  assign n17011 = n2910 | n10915 ;
  assign n17012 = n683 & ~n17011 ;
  assign n17013 = n3177 | n16067 ;
  assign n17014 = ( n5904 & ~n11226 ) | ( n5904 & n17013 ) | ( ~n11226 & n17013 ) ;
  assign n17015 = n6340 | n7039 ;
  assign n17016 = n17015 ^ n2923 ^ 1'b0 ;
  assign n17017 = n2475 & ~n17016 ;
  assign n17018 = n17017 ^ n6489 ^ 1'b0 ;
  assign n17019 = n1292 & ~n17018 ;
  assign n17020 = n17019 ^ x9 ^ 1'b0 ;
  assign n17021 = ( ~n17012 & n17014 ) | ( ~n17012 & n17020 ) | ( n17014 & n17020 ) ;
  assign n17022 = ( ~n449 & n4762 ) | ( ~n449 & n6327 ) | ( n4762 & n6327 ) ;
  assign n17023 = n9284 ^ n6332 ^ n2160 ;
  assign n17024 = n10218 ^ n2805 ^ 1'b0 ;
  assign n17025 = n17024 ^ n3454 ^ 1'b0 ;
  assign n17026 = n16032 & n17025 ;
  assign n17027 = n15408 & ~n16827 ;
  assign n17028 = n17027 ^ n15315 ^ 1'b0 ;
  assign n17029 = n5714 ^ n2387 ^ 1'b0 ;
  assign n17030 = ( ~n14560 & n16704 ) | ( ~n14560 & n17029 ) | ( n16704 & n17029 ) ;
  assign n17031 = n6119 ^ n4522 ^ 1'b0 ;
  assign n17032 = n17031 ^ n15984 ^ n4811 ;
  assign n17033 = n6055 | n15574 ;
  assign n17034 = n16691 & ~n17033 ;
  assign n17035 = n10729 | n17034 ;
  assign n17036 = n13560 & ~n17035 ;
  assign n17037 = n7998 ^ n2639 ^ 1'b0 ;
  assign n17038 = ~n2944 & n5384 ;
  assign n17039 = n3137 | n17038 ;
  assign n17040 = n17039 ^ n8051 ^ 1'b0 ;
  assign n17041 = n15788 | n17040 ;
  assign n17042 = n17041 ^ n416 ^ 1'b0 ;
  assign n17043 = n4980 ^ n846 ^ 1'b0 ;
  assign n17044 = ( ~n7180 & n12590 ) | ( ~n7180 & n17043 ) | ( n12590 & n17043 ) ;
  assign n17045 = n8775 | n16918 ;
  assign n17046 = ( n551 & n1100 ) | ( n551 & ~n4300 ) | ( n1100 & ~n4300 ) ;
  assign n17047 = ~n8041 & n9517 ;
  assign n17048 = n17047 ^ n5302 ^ 1'b0 ;
  assign n17049 = n17048 ^ n8268 ^ 1'b0 ;
  assign n17050 = n3569 | n17049 ;
  assign n17051 = ( ~n7243 & n17046 ) | ( ~n7243 & n17050 ) | ( n17046 & n17050 ) ;
  assign n17052 = n7984 ^ n6071 ^ x92 ;
  assign n17053 = n16611 ^ n8547 ^ n2640 ;
  assign n17054 = n3324 & n9114 ;
  assign n17055 = ( ~n4705 & n8972 ) | ( ~n4705 & n17054 ) | ( n8972 & n17054 ) ;
  assign n17056 = n1201 | n12646 ;
  assign n17057 = n3406 & ~n7344 ;
  assign n17058 = ( n2423 & n13997 ) | ( n2423 & ~n17057 ) | ( n13997 & ~n17057 ) ;
  assign n17059 = n12802 & ~n14342 ;
  assign n17060 = n17058 & n17059 ;
  assign n17061 = n3355 ^ n2398 ^ 1'b0 ;
  assign n17062 = n17060 | n17061 ;
  assign n17063 = n2752 & n9656 ;
  assign n17064 = ( n227 & n3686 ) | ( n227 & n17063 ) | ( n3686 & n17063 ) ;
  assign n17065 = n9480 & n17064 ;
  assign n17066 = ~n6839 & n17065 ;
  assign n17067 = n17066 ^ n12057 ^ 1'b0 ;
  assign n17070 = n12429 ^ n9222 ^ 1'b0 ;
  assign n17071 = n17070 ^ n7820 ^ n7319 ;
  assign n17068 = n4622 | n8568 ;
  assign n17069 = n17068 ^ n11420 ^ n8017 ;
  assign n17072 = n17071 ^ n17069 ^ n16632 ;
  assign n17073 = n15574 ^ n9948 ^ 1'b0 ;
  assign n17074 = n10398 ^ n6777 ^ 1'b0 ;
  assign n17075 = n2543 | n17074 ;
  assign n17076 = n17075 ^ n5440 ^ 1'b0 ;
  assign n17077 = n17076 ^ n7875 ^ n5870 ;
  assign n17078 = n8981 | n14333 ;
  assign n17079 = n9135 & n17078 ;
  assign n17080 = n17079 ^ n3307 ^ 1'b0 ;
  assign n17081 = ~n5547 & n9404 ;
  assign n17082 = ~n2541 & n17081 ;
  assign n17083 = n17082 ^ n12072 ^ 1'b0 ;
  assign n17084 = ~n942 & n17083 ;
  assign n17085 = n15916 ^ n7399 ^ n911 ;
  assign n17087 = n9139 ^ n4283 ^ 1'b0 ;
  assign n17086 = n3047 | n16554 ;
  assign n17088 = n17087 ^ n17086 ^ 1'b0 ;
  assign n17089 = n15486 ^ n2458 ^ n1365 ;
  assign n17090 = n8890 | n17089 ;
  assign n17091 = n2167 ^ n628 ^ n164 ;
  assign n17092 = n10715 & n17091 ;
  assign n17093 = n12874 ^ n11611 ^ 1'b0 ;
  assign n17094 = ( ~n5224 & n13586 ) | ( ~n5224 & n17093 ) | ( n13586 & n17093 ) ;
  assign n17095 = n1172 & n11112 ;
  assign n17096 = ~n5980 & n17095 ;
  assign n17097 = ~n1203 & n4194 ;
  assign n17098 = ~n6870 & n17097 ;
  assign n17099 = n335 & n7593 ;
  assign n17100 = ( n474 & n636 ) | ( n474 & n3985 ) | ( n636 & n3985 ) ;
  assign n17101 = n14399 ^ n4002 ^ 1'b0 ;
  assign n17102 = n17100 & n17101 ;
  assign n17103 = ~n4472 & n17102 ;
  assign n17104 = n3158 & n17103 ;
  assign n17105 = n10191 ^ n164 ^ 1'b0 ;
  assign n17106 = ~n17104 & n17105 ;
  assign n17109 = n5711 ^ n3116 ^ 1'b0 ;
  assign n17107 = n15437 ^ n9349 ^ 1'b0 ;
  assign n17108 = n4689 & ~n17107 ;
  assign n17110 = n17109 ^ n17108 ^ n9811 ;
  assign n17111 = n6103 ^ n3741 ^ 1'b0 ;
  assign n17112 = n1986 ^ x37 ^ 1'b0 ;
  assign n17113 = n6472 & ~n13296 ;
  assign n17114 = n14177 & n17113 ;
  assign n17115 = n16612 ^ n14900 ^ 1'b0 ;
  assign n17116 = n1713 | n3075 ;
  assign n17117 = n535 | n17116 ;
  assign n17118 = n8967 & ~n17117 ;
  assign n17119 = n932 & ~n13944 ;
  assign n17120 = ( n10719 & ~n12869 ) | ( n10719 & n14983 ) | ( ~n12869 & n14983 ) ;
  assign n17121 = n17120 ^ n7311 ^ n1930 ;
  assign n17122 = ( n12147 & n15405 ) | ( n12147 & n15922 ) | ( n15405 & n15922 ) ;
  assign n17123 = n1368 | n4625 ;
  assign n17124 = n17123 ^ n2462 ^ 1'b0 ;
  assign n17125 = n17124 ^ n9036 ^ 1'b0 ;
  assign n17126 = n3816 | n7530 ;
  assign n17127 = n17126 ^ n3223 ^ 1'b0 ;
  assign n17128 = ( n1909 & n8643 ) | ( n1909 & n15336 ) | ( n8643 & n15336 ) ;
  assign n17129 = n4872 | n7620 ;
  assign n17130 = n3351 ^ n3029 ^ 1'b0 ;
  assign n17131 = ( n1455 & n2198 ) | ( n1455 & ~n4749 ) | ( n2198 & ~n4749 ) ;
  assign n17132 = n7737 & n14144 ;
  assign n17133 = n17131 & n17132 ;
  assign n17134 = ~n569 & n2555 ;
  assign n17135 = n17133 & n17134 ;
  assign n17136 = x67 & n13467 ;
  assign n17137 = n17136 ^ n2018 ^ 1'b0 ;
  assign n17141 = ( ~n8305 & n11208 ) | ( ~n8305 & n11781 ) | ( n11208 & n11781 ) ;
  assign n17138 = n3950 ^ n2573 ^ n1914 ;
  assign n17139 = n17138 ^ n10514 ^ 1'b0 ;
  assign n17140 = n17139 ^ n7460 ^ 1'b0 ;
  assign n17142 = n17141 ^ n17140 ^ 1'b0 ;
  assign n17143 = n14064 ^ n12957 ^ 1'b0 ;
  assign n17144 = ~n8716 & n9194 ;
  assign n17145 = n17144 ^ n9441 ^ 1'b0 ;
  assign n17146 = n5471 ^ n2190 ^ 1'b0 ;
  assign n17148 = ~n5837 & n11297 ;
  assign n17149 = ( n5227 & n16049 ) | ( n5227 & ~n17148 ) | ( n16049 & ~n17148 ) ;
  assign n17147 = n8382 & n14493 ;
  assign n17150 = n17149 ^ n17147 ^ 1'b0 ;
  assign n17152 = n12323 ^ n2409 ^ n2301 ;
  assign n17151 = n8450 ^ n3326 ^ n1160 ;
  assign n17153 = n17152 ^ n17151 ^ 1'b0 ;
  assign n17154 = n8084 ^ n3459 ^ 1'b0 ;
  assign n17155 = n6816 | n17154 ;
  assign n17156 = n4108 & n17155 ;
  assign n17157 = n17156 ^ n15574 ^ 1'b0 ;
  assign n17158 = ( n7641 & n17153 ) | ( n7641 & n17157 ) | ( n17153 & n17157 ) ;
  assign n17159 = n4133 ^ n1229 ^ n1013 ;
  assign n17160 = n10710 | n17159 ;
  assign n17161 = n17160 ^ n1814 ^ 1'b0 ;
  assign n17162 = n17161 ^ n7193 ^ 1'b0 ;
  assign n17163 = ~n4457 & n17162 ;
  assign n17164 = n5474 & n6138 ;
  assign n17165 = n3374 ^ x9 ^ 1'b0 ;
  assign n17166 = n17164 & ~n17165 ;
  assign n17167 = n1006 ^ n710 ^ 1'b0 ;
  assign n17168 = ~n15252 & n17167 ;
  assign n17169 = n15612 ^ n3450 ^ 1'b0 ;
  assign n17170 = ( n1443 & n12463 ) | ( n1443 & n17169 ) | ( n12463 & n17169 ) ;
  assign n17171 = n17170 ^ n9357 ^ 1'b0 ;
  assign n17172 = n4853 ^ n4123 ^ 1'b0 ;
  assign n17173 = n10306 & ~n17172 ;
  assign n17174 = ~n4081 & n11712 ;
  assign n17175 = n730 | n17174 ;
  assign n17176 = n17175 ^ n850 ^ 1'b0 ;
  assign n17177 = n17176 ^ n10852 ^ n4344 ;
  assign n17178 = n17177 ^ n8490 ^ 1'b0 ;
  assign n17179 = n10619 ^ n4281 ^ 1'b0 ;
  assign n17180 = n17179 ^ n11451 ^ n5497 ;
  assign n17181 = ~n6796 & n12371 ;
  assign n17182 = n17181 ^ n16634 ^ 1'b0 ;
  assign n17183 = ( n1041 & n7019 ) | ( n1041 & n17182 ) | ( n7019 & n17182 ) ;
  assign n17184 = n17183 ^ n15150 ^ n15129 ;
  assign n17185 = n12225 ^ n8618 ^ n2853 ;
  assign n17186 = n17185 ^ n2897 ^ 1'b0 ;
  assign n17187 = ~n17184 & n17186 ;
  assign n17188 = n17187 ^ n6229 ^ 1'b0 ;
  assign n17189 = ( n556 & n9403 ) | ( n556 & ~n12946 ) | ( n9403 & ~n12946 ) ;
  assign n17190 = n17189 ^ n13445 ^ 1'b0 ;
  assign n17191 = n1781 ^ n298 ^ 1'b0 ;
  assign n17192 = n3054 & n17191 ;
  assign n17193 = ( n4015 & n10030 ) | ( n4015 & n11074 ) | ( n10030 & n11074 ) ;
  assign n17194 = n4394 ^ n2528 ^ 1'b0 ;
  assign n17195 = ~n1357 & n8447 ;
  assign n17196 = n17195 ^ n4260 ^ n752 ;
  assign n17197 = n15564 ^ n538 ^ 1'b0 ;
  assign n17198 = ~n5128 & n17197 ;
  assign n17199 = n5716 & n17198 ;
  assign n17200 = ( n13498 & n13997 ) | ( n13498 & n16014 ) | ( n13997 & n16014 ) ;
  assign n17201 = n16208 | n16464 ;
  assign n17202 = ( ~n831 & n9597 ) | ( ~n831 & n15334 ) | ( n9597 & n15334 ) ;
  assign n17203 = ( n2231 & ~n3994 ) | ( n2231 & n9880 ) | ( ~n3994 & n9880 ) ;
  assign n17204 = n5678 ^ n655 ^ 1'b0 ;
  assign n17205 = ~n1756 & n17204 ;
  assign n17206 = ( ~n1907 & n4546 ) | ( ~n1907 & n17205 ) | ( n4546 & n17205 ) ;
  assign n17207 = n1643 & n17206 ;
  assign n17208 = n511 & n17207 ;
  assign n17209 = n13232 ^ n2998 ^ 1'b0 ;
  assign n17211 = ( ~n5751 & n8099 ) | ( ~n5751 & n8683 ) | ( n8099 & n8683 ) ;
  assign n17210 = ~n4518 & n7614 ;
  assign n17212 = n17211 ^ n17210 ^ 1'b0 ;
  assign n17213 = n17212 ^ n3677 ^ 1'b0 ;
  assign n17214 = n9904 | n17213 ;
  assign n17215 = n4050 ^ n641 ^ 1'b0 ;
  assign n17216 = n919 & n2862 ;
  assign n17217 = n3173 & n17216 ;
  assign n17218 = n1381 ^ n917 ^ 1'b0 ;
  assign n17219 = n17217 | n17218 ;
  assign n17220 = n4101 & n9506 ;
  assign n17221 = n17220 ^ n4156 ^ 1'b0 ;
  assign n17222 = n17221 ^ n3373 ^ 1'b0 ;
  assign n17223 = n17219 | n17222 ;
  assign n17224 = n17223 ^ n3889 ^ 1'b0 ;
  assign n17225 = n2063 & ~n2989 ;
  assign n17226 = n17225 ^ n6199 ^ 1'b0 ;
  assign n17227 = n6198 & ~n17226 ;
  assign n17228 = n8170 ^ n5569 ^ n4739 ;
  assign n17229 = n17228 ^ n5070 ^ 1'b0 ;
  assign n17230 = n740 & ~n17229 ;
  assign n17231 = n14352 ^ n11392 ^ 1'b0 ;
  assign n17232 = n17230 & ~n17231 ;
  assign n17233 = n16564 ^ n1178 ^ 1'b0 ;
  assign n17234 = n3189 & n17233 ;
  assign n17235 = ~n12779 & n17234 ;
  assign n17236 = n17235 ^ n3650 ^ 1'b0 ;
  assign n17237 = n1928 | n12866 ;
  assign n17238 = n17237 ^ n16501 ^ 1'b0 ;
  assign n17239 = n8740 | n17238 ;
  assign n17240 = n17239 ^ n14344 ^ 1'b0 ;
  assign n17241 = n8457 ^ n2703 ^ 1'b0 ;
  assign n17242 = n3865 & n17241 ;
  assign n17243 = n9327 & n17242 ;
  assign n17249 = n3582 ^ n1203 ^ 1'b0 ;
  assign n17244 = n4839 | n11953 ;
  assign n17245 = n8097 & ~n17244 ;
  assign n17246 = n7229 | n17245 ;
  assign n17247 = n1666 & ~n17246 ;
  assign n17248 = n1751 & n17247 ;
  assign n17250 = n17249 ^ n17248 ^ n2565 ;
  assign n17251 = n5078 ^ n3600 ^ n2423 ;
  assign n17252 = ~n4675 & n17251 ;
  assign n17253 = ( ~n9736 & n17250 ) | ( ~n9736 & n17252 ) | ( n17250 & n17252 ) ;
  assign n17254 = ~n508 & n2332 ;
  assign n17256 = n2243 & ~n8577 ;
  assign n17257 = ~n16807 & n17256 ;
  assign n17255 = n11004 ^ n6853 ^ n6283 ;
  assign n17258 = n17257 ^ n17255 ^ 1'b0 ;
  assign n17259 = n4830 & ~n6222 ;
  assign n17260 = ~n2654 & n17259 ;
  assign n17261 = n10318 | n12926 ;
  assign n17262 = n10770 & ~n17261 ;
  assign n17263 = ( n8938 & n17260 ) | ( n8938 & n17262 ) | ( n17260 & n17262 ) ;
  assign n17264 = n16443 ^ n12828 ^ n6859 ;
  assign n17265 = n17264 ^ n15468 ^ 1'b0 ;
  assign n17266 = n4904 ^ n2377 ^ n347 ;
  assign n17267 = ~n4025 & n5213 ;
  assign n17268 = n17266 & n17267 ;
  assign n17269 = n14541 ^ n5627 ^ 1'b0 ;
  assign n17270 = n2147 & ~n6140 ;
  assign n17271 = n3642 & n4949 ;
  assign n17272 = ( n8185 & n17270 ) | ( n8185 & n17271 ) | ( n17270 & n17271 ) ;
  assign n17273 = n15662 ^ n12771 ^ n2670 ;
  assign n17274 = n6275 & n7972 ;
  assign n17275 = ~n307 & n17274 ;
  assign n17276 = n10807 | n17275 ;
  assign n17277 = n8899 & ~n17276 ;
  assign n17278 = ( n4380 & ~n15183 ) | ( n4380 & n17277 ) | ( ~n15183 & n17277 ) ;
  assign n17279 = ~n8679 & n17278 ;
  assign n17285 = n1986 | n6807 ;
  assign n17286 = n17285 ^ n8721 ^ 1'b0 ;
  assign n17281 = n965 & ~n4516 ;
  assign n17282 = n17281 ^ n2810 ^ 1'b0 ;
  assign n17283 = n1306 | n17282 ;
  assign n17280 = ~n641 & n15053 ;
  assign n17284 = n17283 ^ n17280 ^ n7209 ;
  assign n17287 = n17286 ^ n17284 ^ 1'b0 ;
  assign n17288 = n17287 ^ n7233 ^ 1'b0 ;
  assign n17289 = n14617 ^ n4878 ^ 1'b0 ;
  assign n17290 = ~n15178 & n17289 ;
  assign n17291 = n17290 ^ n11002 ^ n3010 ;
  assign n17292 = ( ~n6873 & n15459 ) | ( ~n6873 & n17291 ) | ( n15459 & n17291 ) ;
  assign n17293 = n6838 & ~n9218 ;
  assign n17294 = ~n9913 & n17293 ;
  assign n17295 = ( n3228 & ~n7427 ) | ( n3228 & n17294 ) | ( ~n7427 & n17294 ) ;
  assign n17296 = ~n2231 & n7988 ;
  assign n17297 = ( n14622 & ~n16205 ) | ( n14622 & n17296 ) | ( ~n16205 & n17296 ) ;
  assign n17298 = n4356 ^ n2172 ^ 1'b0 ;
  assign n17299 = n11272 & ~n13452 ;
  assign n17300 = n17299 ^ n13158 ^ 1'b0 ;
  assign n17301 = n2766 ^ n1935 ^ 1'b0 ;
  assign n17302 = ( n6797 & n10832 ) | ( n6797 & n17301 ) | ( n10832 & n17301 ) ;
  assign n17303 = ~n3217 & n17302 ;
  assign n17304 = n2042 ^ n1480 ^ 1'b0 ;
  assign n17305 = n17304 ^ n6566 ^ n2733 ;
  assign n17306 = ( n1620 & n3493 ) | ( n1620 & n4645 ) | ( n3493 & n4645 ) ;
  assign n17307 = n7287 | n17306 ;
  assign n17308 = n17307 ^ n2152 ^ 1'b0 ;
  assign n17309 = ~n4029 & n6930 ;
  assign n17310 = n4221 ^ n2390 ^ n1870 ;
  assign n17311 = n17310 ^ n845 ^ 1'b0 ;
  assign n17312 = ~n9227 & n17311 ;
  assign n17313 = n17312 ^ n8677 ^ 1'b0 ;
  assign n17314 = n15963 & n17313 ;
  assign n17315 = ( n10158 & n15135 ) | ( n10158 & ~n17314 ) | ( n15135 & ~n17314 ) ;
  assign n17316 = n17315 ^ n15212 ^ n2061 ;
  assign n17317 = n6999 ^ n3610 ^ 1'b0 ;
  assign n17318 = ~n4308 & n17317 ;
  assign n17319 = ~n4215 & n17318 ;
  assign n17320 = ~n5347 & n17319 ;
  assign n17321 = n17320 ^ n8514 ^ 1'b0 ;
  assign n17322 = ~n5903 & n17321 ;
  assign n17323 = n14410 | n16360 ;
  assign n17324 = ( n505 & n2971 ) | ( n505 & ~n4713 ) | ( n2971 & ~n4713 ) ;
  assign n17325 = n17324 ^ n11196 ^ n2697 ;
  assign n17326 = n17325 ^ n1851 ^ 1'b0 ;
  assign n17327 = n9746 ^ n5742 ^ 1'b0 ;
  assign n17328 = n15053 ^ n10459 ^ 1'b0 ;
  assign n17329 = x21 & ~n17328 ;
  assign n17330 = n15551 ^ n5741 ^ 1'b0 ;
  assign n17331 = n1902 | n17330 ;
  assign n17332 = n17331 ^ n781 ^ 1'b0 ;
  assign n17333 = n13493 & ~n14082 ;
  assign n17334 = ( n6387 & ~n17332 ) | ( n6387 & n17333 ) | ( ~n17332 & n17333 ) ;
  assign n17335 = n9804 & ~n14624 ;
  assign n17336 = ~n5537 & n8909 ;
  assign n17337 = n6169 & n17336 ;
  assign n17338 = n9047 | n16316 ;
  assign n17340 = n827 | n3948 ;
  assign n17339 = n13425 ^ n5461 ^ 1'b0 ;
  assign n17341 = n17340 ^ n17339 ^ n7162 ;
  assign n17342 = ~n2139 & n9563 ;
  assign n17343 = ~n2072 & n17342 ;
  assign n17344 = ( n6328 & ~n12418 ) | ( n6328 & n17343 ) | ( ~n12418 & n17343 ) ;
  assign n17345 = n981 & n9698 ;
  assign n17346 = ~n6277 & n17345 ;
  assign n17347 = ~n11330 & n17346 ;
  assign n17348 = n14287 ^ n7096 ^ n5013 ;
  assign n17349 = n7999 & ~n11689 ;
  assign n17350 = n17348 & n17349 ;
  assign n17351 = n1176 & ~n2360 ;
  assign n17352 = n10191 | n17351 ;
  assign n17353 = n17350 & ~n17352 ;
  assign n17354 = ~n10343 & n12761 ;
  assign n17355 = n8415 & n17354 ;
  assign n17356 = n17355 ^ n8572 ^ 1'b0 ;
  assign n17357 = n3287 ^ n1962 ^ 1'b0 ;
  assign n17358 = n14157 ^ n13577 ^ n12827 ;
  assign n17359 = n13658 ^ n8822 ^ 1'b0 ;
  assign n17360 = n3178 & n17359 ;
  assign n17361 = ( ~n2894 & n3917 ) | ( ~n2894 & n5570 ) | ( n3917 & n5570 ) ;
  assign n17362 = n17361 ^ n5560 ^ 1'b0 ;
  assign n17363 = n6856 & n17362 ;
  assign n17364 = n7815 & n17363 ;
  assign n17365 = ~n4737 & n17364 ;
  assign n17366 = n5764 | n16408 ;
  assign n17367 = n12704 ^ n8006 ^ n7683 ;
  assign n17368 = n17367 ^ n13018 ^ 1'b0 ;
  assign n17369 = n17368 ^ n13896 ^ n9827 ;
  assign n17370 = n4022 ^ n1759 ^ 1'b0 ;
  assign n17371 = n17370 ^ n14445 ^ n1679 ;
  assign n17372 = n17371 ^ n13223 ^ 1'b0 ;
  assign n17373 = n16630 | n17372 ;
  assign n17375 = n7626 ^ n6211 ^ n4285 ;
  assign n17376 = n17375 ^ n3461 ^ n1175 ;
  assign n17374 = n3653 | n6036 ;
  assign n17377 = n17376 ^ n17374 ^ 1'b0 ;
  assign n17378 = ~n8623 & n12276 ;
  assign n17379 = n17378 ^ n11612 ^ n9284 ;
  assign n17380 = n2252 & n17379 ;
  assign n17381 = n17380 ^ n15130 ^ n10240 ;
  assign n17382 = n4131 ^ n3948 ^ n2072 ;
  assign n17383 = n16058 & ~n17382 ;
  assign n17384 = ( n2305 & n2872 ) | ( n2305 & n5831 ) | ( n2872 & n5831 ) ;
  assign n17385 = ~n8472 & n16843 ;
  assign n17386 = n17385 ^ n7926 ^ 1'b0 ;
  assign n17387 = n15064 ^ n6579 ^ n5482 ;
  assign n17388 = n6553 & ~n17387 ;
  assign n17389 = n15014 ^ n6726 ^ n2671 ;
  assign n17390 = n890 & n17389 ;
  assign n17391 = n17390 ^ n5303 ^ 1'b0 ;
  assign n17392 = n722 & n5261 ;
  assign n17393 = n1036 | n2524 ;
  assign n17394 = n17393 ^ n5491 ^ 1'b0 ;
  assign n17395 = n14496 & n17394 ;
  assign n17396 = n5261 & n17395 ;
  assign n17397 = n13227 ^ n1223 ^ 1'b0 ;
  assign n17398 = n11340 & n17397 ;
  assign n17399 = ~n1591 & n13062 ;
  assign n17400 = ~n4477 & n14597 ;
  assign n17401 = n17400 ^ n11746 ^ 1'b0 ;
  assign n17402 = ( n8480 & n13960 ) | ( n8480 & ~n17401 ) | ( n13960 & ~n17401 ) ;
  assign n17403 = ~n9511 & n14850 ;
  assign n17404 = n17403 ^ n8775 ^ 1'b0 ;
  assign n17405 = ( ~x16 & n15342 ) | ( ~x16 & n17404 ) | ( n15342 & n17404 ) ;
  assign n17406 = n16197 ^ n8198 ^ n2056 ;
  assign n17407 = ( ~n1153 & n2350 ) | ( ~n1153 & n7743 ) | ( n2350 & n7743 ) ;
  assign n17408 = ( n5861 & n17406 ) | ( n5861 & n17407 ) | ( n17406 & n17407 ) ;
  assign n17409 = ~n1558 & n17408 ;
  assign n17410 = n5396 ^ n2086 ^ 1'b0 ;
  assign n17411 = ~n17409 & n17410 ;
  assign n17412 = n10220 & ~n15442 ;
  assign n17413 = ~x93 & n17412 ;
  assign n17414 = n17413 ^ n9368 ^ 1'b0 ;
  assign n17415 = n17411 & n17414 ;
  assign n17416 = ( n14361 & n17405 ) | ( n14361 & n17415 ) | ( n17405 & n17415 ) ;
  assign n17418 = n8501 | n12684 ;
  assign n17417 = n7144 & n8090 ;
  assign n17419 = n17418 ^ n17417 ^ 1'b0 ;
  assign n17420 = ~n3398 & n9824 ;
  assign n17421 = n12752 ^ n8008 ^ 1'b0 ;
  assign n17422 = n5732 & ~n17421 ;
  assign n17423 = n17420 | n17422 ;
  assign n17424 = n17423 ^ n3374 ^ 1'b0 ;
  assign n17425 = n2232 & ~n2433 ;
  assign n17426 = n17425 ^ n12382 ^ 1'b0 ;
  assign n17427 = ~n1921 & n6082 ;
  assign n17428 = n17427 ^ n17070 ^ 1'b0 ;
  assign n17429 = n17428 ^ n8092 ^ n861 ;
  assign n17430 = n9657 ^ n1913 ^ n233 ;
  assign n17431 = ( n7153 & ~n11198 ) | ( n7153 & n17430 ) | ( ~n11198 & n17430 ) ;
  assign n17432 = n17431 ^ n9160 ^ 1'b0 ;
  assign n17434 = n6010 ^ n2522 ^ n1154 ;
  assign n17433 = n11524 & ~n13897 ;
  assign n17435 = n17434 ^ n17433 ^ 1'b0 ;
  assign n17436 = n11868 ^ n6133 ^ 1'b0 ;
  assign n17437 = n5451 | n17436 ;
  assign n17438 = ( n239 & n6083 ) | ( n239 & ~n17437 ) | ( n6083 & ~n17437 ) ;
  assign n17439 = ~n8323 & n17438 ;
  assign n17440 = ~n8269 & n17439 ;
  assign n17441 = n11112 & n17440 ;
  assign n17442 = ( n3848 & n6453 ) | ( n3848 & n9409 ) | ( n6453 & n9409 ) ;
  assign n17443 = n2498 & ~n17442 ;
  assign n17444 = n16956 ^ n12779 ^ n9485 ;
  assign n17445 = n12698 ^ n4030 ^ 1'b0 ;
  assign n17446 = n8133 | n17445 ;
  assign n17447 = ( ~n7835 & n14895 ) | ( ~n7835 & n17446 ) | ( n14895 & n17446 ) ;
  assign n17448 = n17447 ^ n9064 ^ 1'b0 ;
  assign n17449 = ( x38 & ~n11597 ) | ( x38 & n17448 ) | ( ~n11597 & n17448 ) ;
  assign n17450 = n15384 ^ n5004 ^ n4304 ;
  assign n17451 = n3825 ^ n1643 ^ n937 ;
  assign n17452 = ~n3433 & n17451 ;
  assign n17453 = n11151 ^ n4148 ^ 1'b0 ;
  assign n17454 = n5173 | n17453 ;
  assign n17455 = ~n2659 & n4706 ;
  assign n17456 = n17455 ^ n3642 ^ 1'b0 ;
  assign n17457 = n4905 ^ n3029 ^ n1754 ;
  assign n17458 = n4422 & ~n8842 ;
  assign n17459 = n777 & n17458 ;
  assign n17460 = n17459 ^ n12026 ^ 1'b0 ;
  assign n17461 = n3483 ^ x101 ^ 1'b0 ;
  assign n17462 = n9674 ^ n2964 ^ 1'b0 ;
  assign n17463 = ( n5131 & n6485 ) | ( n5131 & ~n17462 ) | ( n6485 & ~n17462 ) ;
  assign n17464 = x54 & ~n1514 ;
  assign n17465 = n17464 ^ n1784 ^ 1'b0 ;
  assign n17466 = n17465 ^ n14801 ^ 1'b0 ;
  assign n17467 = n3514 | n4059 ;
  assign n17468 = n10827 & n11329 ;
  assign n17469 = ~n4943 & n10982 ;
  assign n17470 = n3677 & ~n9860 ;
  assign n17471 = n17470 ^ n5578 ^ 1'b0 ;
  assign n17472 = n13479 ^ n1640 ^ 1'b0 ;
  assign n17473 = n17472 ^ n13168 ^ 1'b0 ;
  assign n17474 = n13979 & ~n17473 ;
  assign n17475 = n9762 ^ n5664 ^ n2031 ;
  assign n17476 = n917 & ~n17475 ;
  assign n17477 = ~n6799 & n17476 ;
  assign n17478 = ~n1223 & n17477 ;
  assign n17479 = ( n6075 & ~n7448 ) | ( n6075 & n10389 ) | ( ~n7448 & n10389 ) ;
  assign n17480 = n10109 ^ n6378 ^ 1'b0 ;
  assign n17481 = n14560 & n17480 ;
  assign n17482 = n17481 ^ n12297 ^ n2342 ;
  assign n17483 = n3792 & ~n8414 ;
  assign n17484 = n17483 ^ n5313 ^ 1'b0 ;
  assign n17485 = n17482 & ~n17484 ;
  assign n17486 = n17485 ^ n6976 ^ n2219 ;
  assign n17487 = n4825 | n14505 ;
  assign n17488 = n17487 ^ n13849 ^ 1'b0 ;
  assign n17489 = n11385 ^ n4950 ^ 1'b0 ;
  assign n17490 = n2295 | n17489 ;
  assign n17491 = n15216 | n17490 ;
  assign n17492 = n13060 ^ n12094 ^ 1'b0 ;
  assign n17493 = n17492 ^ n7830 ^ n1957 ;
  assign n17494 = n17493 ^ n6107 ^ 1'b0 ;
  assign n17495 = n6343 & n17494 ;
  assign n17496 = n866 & ~n5349 ;
  assign n17497 = n17496 ^ n15053 ^ 1'b0 ;
  assign n17498 = n17497 ^ n14926 ^ n3380 ;
  assign n17500 = n1656 | n6496 ;
  assign n17501 = n1438 & ~n17500 ;
  assign n17499 = n16288 ^ n4681 ^ 1'b0 ;
  assign n17502 = n17501 ^ n17499 ^ n7334 ;
  assign n17503 = n4111 ^ n1422 ^ 1'b0 ;
  assign n17504 = n11708 & n17503 ;
  assign n17505 = ~n13754 & n17504 ;
  assign n17506 = ~n8242 & n17505 ;
  assign n17507 = n2679 | n10258 ;
  assign n17508 = n8370 | n17507 ;
  assign n17509 = n3784 & ~n6593 ;
  assign n17510 = n17509 ^ n4606 ^ 1'b0 ;
  assign n17511 = n17510 ^ n6655 ^ 1'b0 ;
  assign n17512 = n6133 | n17511 ;
  assign n17513 = n3556 & n4181 ;
  assign n17514 = n17513 ^ n4928 ^ 1'b0 ;
  assign n17515 = n5381 & ~n8829 ;
  assign n17516 = ( n6376 & n14100 ) | ( n6376 & n16619 ) | ( n14100 & n16619 ) ;
  assign n17517 = n17516 ^ n14009 ^ 1'b0 ;
  assign n17518 = n4286 | n17517 ;
  assign n17519 = n6858 ^ n4984 ^ 1'b0 ;
  assign n17520 = n7526 & ~n17519 ;
  assign n17521 = n5730 ^ n4729 ^ 1'b0 ;
  assign n17526 = ( n3332 & n5579 ) | ( n3332 & n16346 ) | ( n5579 & n16346 ) ;
  assign n17525 = n582 & n14284 ;
  assign n17527 = n17526 ^ n17525 ^ 1'b0 ;
  assign n17524 = n5349 ^ n4099 ^ n3096 ;
  assign n17522 = n11061 ^ n2905 ^ 1'b0 ;
  assign n17523 = ~n4068 & n17522 ;
  assign n17528 = n17527 ^ n17524 ^ n17523 ;
  assign n17529 = n7574 & n9204 ;
  assign n17530 = ~n7928 & n17529 ;
  assign n17531 = n2980 & ~n9511 ;
  assign n17532 = n17531 ^ n8880 ^ 1'b0 ;
  assign n17533 = n14931 ^ n14140 ^ n1213 ;
  assign n17534 = n10910 ^ n9664 ^ 1'b0 ;
  assign n17535 = ~n2600 & n3732 ;
  assign n17536 = n13576 & n17535 ;
  assign n17537 = n5799 & ~n17536 ;
  assign n17538 = n6018 & ~n17537 ;
  assign n17539 = n5397 & ~n10255 ;
  assign n17540 = n17539 ^ n9999 ^ 1'b0 ;
  assign n17541 = ( ~n5221 & n6424 ) | ( ~n5221 & n11577 ) | ( n6424 & n11577 ) ;
  assign n17542 = n10926 ^ n5460 ^ 1'b0 ;
  assign n17543 = n8326 & n17542 ;
  assign n17544 = ~n17541 & n17543 ;
  assign n17545 = ~n17540 & n17544 ;
  assign n17547 = n4717 ^ n3134 ^ n159 ;
  assign n17548 = n17547 ^ n6993 ^ n1108 ;
  assign n17546 = n3961 | n5221 ;
  assign n17549 = n17548 ^ n17546 ^ 1'b0 ;
  assign n17550 = n14460 ^ n11790 ^ n1302 ;
  assign n17551 = n7913 ^ n3929 ^ n1352 ;
  assign n17552 = n4379 & ~n15723 ;
  assign n17553 = n17552 ^ n1918 ^ 1'b0 ;
  assign n17554 = n17553 ^ n6492 ^ 1'b0 ;
  assign n17555 = ~n9507 & n17554 ;
  assign n17556 = n17555 ^ n7711 ^ 1'b0 ;
  assign n17557 = ~n3831 & n7676 ;
  assign n17558 = ~n11465 & n17557 ;
  assign n17559 = ~n1903 & n16947 ;
  assign n17560 = n17559 ^ n3856 ^ 1'b0 ;
  assign n17561 = n14242 ^ n2636 ^ 1'b0 ;
  assign n17562 = ~n3072 & n17561 ;
  assign n17563 = n10564 & ~n17562 ;
  assign n17564 = ~n3905 & n17563 ;
  assign n17565 = n14083 ^ n9016 ^ 1'b0 ;
  assign n17566 = n1002 & n14683 ;
  assign n17567 = n17566 ^ n5216 ^ 1'b0 ;
  assign n17568 = ~n4336 & n9058 ;
  assign n17569 = n2282 | n17568 ;
  assign n17574 = ~n1390 & n5159 ;
  assign n17575 = ~n1554 & n17574 ;
  assign n17570 = n16715 ^ n5367 ^ n384 ;
  assign n17571 = n17570 ^ n2420 ^ 1'b0 ;
  assign n17572 = n9551 & n17571 ;
  assign n17573 = n7947 & n17572 ;
  assign n17576 = n17575 ^ n17573 ^ 1'b0 ;
  assign n17577 = n8168 ^ n5491 ^ 1'b0 ;
  assign n17578 = n7436 | n17577 ;
  assign n17579 = n17578 ^ n7908 ^ 1'b0 ;
  assign n17580 = n17576 & n17579 ;
  assign n17581 = ( ~n233 & n12235 ) | ( ~n233 & n17580 ) | ( n12235 & n17580 ) ;
  assign n17582 = ( ~n348 & n8440 ) | ( ~n348 & n11522 ) | ( n8440 & n11522 ) ;
  assign n17583 = ~n7112 & n17582 ;
  assign n17584 = n16327 ^ n2360 ^ 1'b0 ;
  assign n17585 = n7579 | n17584 ;
  assign n17586 = ( ~n723 & n4221 ) | ( ~n723 & n17585 ) | ( n4221 & n17585 ) ;
  assign n17587 = n17586 ^ n7933 ^ 1'b0 ;
  assign n17588 = ~n17583 & n17587 ;
  assign n17589 = ~n6059 & n16431 ;
  assign n17590 = n16737 ^ n4703 ^ 1'b0 ;
  assign n17592 = ( ~n2143 & n3132 ) | ( ~n2143 & n13893 ) | ( n3132 & n13893 ) ;
  assign n17591 = ( n1084 & ~n1302 ) | ( n1084 & n3374 ) | ( ~n1302 & n3374 ) ;
  assign n17593 = n17592 ^ n17591 ^ n2271 ;
  assign n17594 = n3632 & n17593 ;
  assign n17596 = n3738 & n10807 ;
  assign n17597 = n7910 & ~n17596 ;
  assign n17598 = n17597 ^ n11297 ^ 1'b0 ;
  assign n17595 = ( n3212 & n4986 ) | ( n3212 & n14235 ) | ( n4986 & n14235 ) ;
  assign n17599 = n17598 ^ n17595 ^ 1'b0 ;
  assign n17600 = ( n325 & ~n10264 ) | ( n325 & n17599 ) | ( ~n10264 & n17599 ) ;
  assign n17601 = n4501 ^ n500 ^ 1'b0 ;
  assign n17602 = n3279 & ~n8173 ;
  assign n17603 = ~n1851 & n17602 ;
  assign n17604 = n17603 ^ n12276 ^ 1'b0 ;
  assign n17605 = n17601 & ~n17604 ;
  assign n17608 = n871 & ~n1896 ;
  assign n17609 = ~n871 & n17608 ;
  assign n17610 = n292 & n9005 ;
  assign n17611 = n17609 & n17610 ;
  assign n17612 = n15946 ^ n4356 ^ 1'b0 ;
  assign n17613 = ( n10445 & n17611 ) | ( n10445 & ~n17612 ) | ( n17611 & ~n17612 ) ;
  assign n17606 = ( n3887 & n5690 ) | ( n3887 & ~n9901 ) | ( n5690 & ~n9901 ) ;
  assign n17607 = n740 & n17606 ;
  assign n17614 = n17613 ^ n17607 ^ 1'b0 ;
  assign n17615 = n5099 ^ n4203 ^ 1'b0 ;
  assign n17616 = n17614 & n17615 ;
  assign n17618 = n10160 & ~n11512 ;
  assign n17617 = ( n390 & n2237 ) | ( n390 & n8843 ) | ( n2237 & n8843 ) ;
  assign n17619 = n17618 ^ n17617 ^ 1'b0 ;
  assign n17620 = n7555 & ~n17619 ;
  assign n17621 = n8757 ^ n4902 ^ 1'b0 ;
  assign n17622 = n1546 | n3552 ;
  assign n17623 = n17622 ^ n17203 ^ 1'b0 ;
  assign n17624 = n17621 & n17623 ;
  assign n17625 = n17548 ^ n15296 ^ 1'b0 ;
  assign n17626 = ( ~n7225 & n8106 ) | ( ~n7225 & n9207 ) | ( n8106 & n9207 ) ;
  assign n17627 = n3169 ^ n2086 ^ n375 ;
  assign n17628 = ( n8409 & n17626 ) | ( n8409 & n17627 ) | ( n17626 & n17627 ) ;
  assign n17629 = n15801 ^ n13924 ^ n9106 ;
  assign n17630 = n17629 ^ n1066 ^ n548 ;
  assign n17631 = ~x107 & n290 ;
  assign n17632 = ~n13334 & n17631 ;
  assign n17633 = ( n672 & n7285 ) | ( n672 & n10619 ) | ( n7285 & n10619 ) ;
  assign n17634 = ( n2356 & ~n6032 ) | ( n2356 & n17633 ) | ( ~n6032 & n17633 ) ;
  assign n17635 = n10538 ^ n6134 ^ 1'b0 ;
  assign n17636 = n17635 ^ n2394 ^ n1921 ;
  assign n17637 = n11253 ^ n1087 ^ 1'b0 ;
  assign n17638 = ~n14461 & n17637 ;
  assign n17639 = ( n3334 & ~n10997 ) | ( n3334 & n14750 ) | ( ~n10997 & n14750 ) ;
  assign n17640 = n9348 ^ n6577 ^ n528 ;
  assign n17641 = n9330 ^ n3303 ^ n2342 ;
  assign n17642 = ( n5597 & ~n14689 ) | ( n5597 & n17641 ) | ( ~n14689 & n17641 ) ;
  assign n17643 = n16342 ^ n5922 ^ n3597 ;
  assign n17644 = n3128 & n7284 ;
  assign n17645 = n3346 & n14328 ;
  assign n17646 = n5925 ^ n2925 ^ 1'b0 ;
  assign n17647 = n4745 | n17646 ;
  assign n17648 = n15813 | n17647 ;
  assign n17650 = n7677 ^ n3326 ^ 1'b0 ;
  assign n17649 = n7647 & n15195 ;
  assign n17651 = n17650 ^ n17649 ^ 1'b0 ;
  assign n17652 = ( n9001 & n12722 ) | ( n9001 & ~n15729 ) | ( n12722 & ~n15729 ) ;
  assign n17653 = ( n8190 & ~n11665 ) | ( n8190 & n17652 ) | ( ~n11665 & n17652 ) ;
  assign n17654 = n6198 | n14742 ;
  assign n17655 = n5017 ^ n3202 ^ 1'b0 ;
  assign n17656 = ( n9597 & n11374 ) | ( n9597 & n14493 ) | ( n11374 & n14493 ) ;
  assign n17657 = n17656 ^ n14245 ^ n10795 ;
  assign n17658 = ( n4973 & ~n8170 ) | ( n4973 & n12928 ) | ( ~n8170 & n12928 ) ;
  assign n17659 = n12820 & ~n13949 ;
  assign n17660 = ( n7342 & ~n8474 ) | ( n7342 & n17659 ) | ( ~n8474 & n17659 ) ;
  assign n17661 = ( n7105 & n9639 ) | ( n7105 & n12001 ) | ( n9639 & n12001 ) ;
  assign n17662 = n17661 ^ n15299 ^ n4373 ;
  assign n17663 = n17662 ^ n9315 ^ n3070 ;
  assign n17664 = n15563 ^ n5176 ^ 1'b0 ;
  assign n17665 = ~n9505 & n17664 ;
  assign n17666 = n3796 & n6298 ;
  assign n17667 = ~n10704 & n17666 ;
  assign n17668 = n8748 ^ n908 ^ 1'b0 ;
  assign n17669 = ( n272 & n2985 ) | ( n272 & n4430 ) | ( n2985 & n4430 ) ;
  assign n17670 = n7214 & ~n17669 ;
  assign n17671 = n15639 & n17670 ;
  assign n17673 = n5535 ^ n1252 ^ 1'b0 ;
  assign n17672 = ( n173 & n7652 ) | ( n173 & ~n10904 ) | ( n7652 & ~n10904 ) ;
  assign n17674 = n17673 ^ n17672 ^ 1'b0 ;
  assign n17675 = n8359 | n17674 ;
  assign n17676 = n3325 ^ n207 ^ 1'b0 ;
  assign n17677 = n5423 ^ n2752 ^ 1'b0 ;
  assign n17678 = n1432 & n2728 ;
  assign n17679 = n9364 & n17678 ;
  assign n17680 = n8055 | n17679 ;
  assign n17681 = n17677 & ~n17680 ;
  assign n17682 = n10160 & ~n17681 ;
  assign n17683 = ~n9192 & n17682 ;
  assign n17684 = ~n5837 & n7072 ;
  assign n17685 = n7746 & n17684 ;
  assign n17686 = n10318 ^ n5600 ^ 1'b0 ;
  assign n17687 = n6451 ^ n1214 ^ 1'b0 ;
  assign n17688 = n10773 & n17687 ;
  assign n17689 = ~n17686 & n17688 ;
  assign n17690 = n17689 ^ n10309 ^ n1794 ;
  assign n17691 = n17690 ^ n2197 ^ 1'b0 ;
  assign n17692 = ( ~n1843 & n4613 ) | ( ~n1843 & n10066 ) | ( n4613 & n10066 ) ;
  assign n17693 = n13425 & ~n17692 ;
  assign n17694 = n17693 ^ n2681 ^ 1'b0 ;
  assign n17695 = n323 & ~n1220 ;
  assign n17696 = n12766 & ~n17695 ;
  assign n17697 = ~n4402 & n17696 ;
  assign n17698 = n7234 ^ n5189 ^ 1'b0 ;
  assign n17699 = n17252 & n17698 ;
  assign n17700 = n17699 ^ n6502 ^ 1'b0 ;
  assign n17701 = n7986 ^ n7031 ^ 1'b0 ;
  assign n17702 = n11437 & n17701 ;
  assign n17703 = n11131 & n17702 ;
  assign n17704 = ( n994 & n15826 ) | ( n994 & n17703 ) | ( n15826 & n17703 ) ;
  assign n17705 = n17369 ^ n11258 ^ 1'b0 ;
  assign n17706 = n11017 | n17705 ;
  assign n17707 = n8591 ^ n7456 ^ n3534 ;
  assign n17708 = n10393 & ~n17707 ;
  assign n17709 = n10882 ^ n6796 ^ 1'b0 ;
  assign n17710 = n17708 & n17709 ;
  assign n17711 = n6654 ^ n2069 ^ n906 ;
  assign n17712 = n197 | n17711 ;
  assign n17713 = n9336 | n17712 ;
  assign n17714 = n11595 ^ n1354 ^ 1'b0 ;
  assign n17715 = n17714 ^ n9225 ^ 1'b0 ;
  assign n17716 = n17713 & ~n17715 ;
  assign n17717 = n673 & ~n5311 ;
  assign n17718 = ~n17245 & n17329 ;
  assign n17719 = ~n12732 & n17718 ;
  assign n17720 = n17719 ^ n13367 ^ 1'b0 ;
  assign n17721 = n17151 | n17720 ;
  assign n17722 = n17721 ^ n1761 ^ n1435 ;
  assign n17723 = n2996 | n6737 ;
  assign n17724 = n3496 & ~n17723 ;
  assign n17725 = x106 & ~n16715 ;
  assign n17726 = n17724 & n17725 ;
  assign n17727 = n5795 & ~n17078 ;
  assign n17728 = n2224 & n10425 ;
  assign n17729 = n17728 ^ n1615 ^ 1'b0 ;
  assign n17730 = ( ~n2163 & n10251 ) | ( ~n2163 & n13034 ) | ( n10251 & n13034 ) ;
  assign n17731 = n4661 & ~n17730 ;
  assign n17732 = n17731 ^ n16433 ^ 1'b0 ;
  assign n17733 = n17729 | n17732 ;
  assign n17734 = ( ~n560 & n6357 ) | ( ~n560 & n8346 ) | ( n6357 & n8346 ) ;
  assign n17735 = ( n5593 & n15846 ) | ( n5593 & ~n17734 ) | ( n15846 & ~n17734 ) ;
  assign n17736 = n529 | n1015 ;
  assign n17737 = n17736 ^ n5699 ^ 1'b0 ;
  assign n17738 = n11471 & ~n17737 ;
  assign n17739 = ( n2908 & n3249 ) | ( n2908 & ~n17738 ) | ( n3249 & ~n17738 ) ;
  assign n17740 = n8109 & ~n16146 ;
  assign n17741 = n17740 ^ n16549 ^ n2718 ;
  assign n17742 = n17741 ^ n10643 ^ n7067 ;
  assign n17743 = n13267 ^ n8919 ^ 1'b0 ;
  assign n17744 = n3429 & ~n17743 ;
  assign n17745 = n9866 ^ n6896 ^ 1'b0 ;
  assign n17746 = n8487 ^ n7693 ^ 1'b0 ;
  assign n17747 = n17745 & n17746 ;
  assign n17748 = n17747 ^ n2163 ^ 1'b0 ;
  assign n17749 = n2014 & n11471 ;
  assign n17750 = n12250 ^ n3791 ^ n3025 ;
  assign n17751 = n17750 ^ n14550 ^ 1'b0 ;
  assign n17752 = ~n4469 & n17751 ;
  assign n17753 = n12347 & n17752 ;
  assign n17754 = n17749 & n17753 ;
  assign n17755 = ~n6281 & n12491 ;
  assign n17756 = n468 & n17755 ;
  assign n17757 = n174 & ~n6883 ;
  assign n17758 = ~n2015 & n17757 ;
  assign n17759 = n17758 ^ n9390 ^ n7819 ;
  assign n17760 = n1505 & n6528 ;
  assign n17761 = n11687 ^ n8284 ^ 1'b0 ;
  assign n17762 = n5609 ^ n1834 ^ 1'b0 ;
  assign n17763 = n17762 ^ n15181 ^ 1'b0 ;
  assign n17764 = ~n485 & n17763 ;
  assign n17765 = ( n2305 & n17761 ) | ( n2305 & ~n17764 ) | ( n17761 & ~n17764 ) ;
  assign n17766 = n9566 & n12829 ;
  assign n17767 = n17766 ^ n10304 ^ 1'b0 ;
  assign n17768 = n17185 ^ n1925 ^ 1'b0 ;
  assign n17769 = n16737 | n17768 ;
  assign n17770 = ~n4553 & n10050 ;
  assign n17771 = n11225 & n11820 ;
  assign n17772 = n12823 ^ n10668 ^ n4941 ;
  assign n17773 = n3162 ^ n646 ^ 1'b0 ;
  assign n17774 = ( n7092 & n9116 ) | ( n7092 & ~n17773 ) | ( n9116 & ~n17773 ) ;
  assign n17775 = n17371 ^ n12366 ^ n768 ;
  assign n17776 = n9403 ^ n3206 ^ n2469 ;
  assign n17777 = n17776 ^ n16301 ^ n1092 ;
  assign n17778 = n17777 ^ n7903 ^ n706 ;
  assign n17779 = n17778 ^ n8003 ^ 1'b0 ;
  assign n17780 = ( n3154 & n12273 ) | ( n3154 & n17779 ) | ( n12273 & n17779 ) ;
  assign n17781 = n16676 ^ n8273 ^ 1'b0 ;
  assign n17782 = ~n2115 & n17781 ;
  assign n17783 = ( n255 & n6866 ) | ( n255 & n13453 ) | ( n6866 & n13453 ) ;
  assign n17784 = n17783 ^ n4629 ^ n2621 ;
  assign n17785 = n17784 ^ n2460 ^ 1'b0 ;
  assign n17789 = n12812 | n16151 ;
  assign n17787 = n4329 & n7324 ;
  assign n17786 = n10249 ^ n4059 ^ 1'b0 ;
  assign n17788 = n17787 ^ n17786 ^ 1'b0 ;
  assign n17790 = n17789 ^ n17788 ^ 1'b0 ;
  assign n17791 = n951 & ~n4498 ;
  assign n17795 = ( n2426 & n4811 ) | ( n2426 & n9470 ) | ( n4811 & n9470 ) ;
  assign n17792 = n12803 ^ n1986 ^ 1'b0 ;
  assign n17793 = n9440 & ~n17792 ;
  assign n17794 = n8073 & n17793 ;
  assign n17796 = n17795 ^ n17794 ^ n6614 ;
  assign n17797 = n15479 ^ n7034 ^ n1765 ;
  assign n17798 = n17797 ^ n9187 ^ 1'b0 ;
  assign n17799 = ~n2612 & n11494 ;
  assign n17800 = n17799 ^ n10291 ^ 1'b0 ;
  assign n17801 = n3398 & n17800 ;
  assign n17802 = n17801 ^ n14980 ^ 1'b0 ;
  assign n17803 = n8653 ^ n5960 ^ 1'b0 ;
  assign n17804 = n17205 ^ n558 ^ n548 ;
  assign n17805 = n17804 ^ n4881 ^ 1'b0 ;
  assign n17806 = n13149 & ~n17805 ;
  assign n17807 = ( n2627 & n7951 ) | ( n2627 & n10880 ) | ( n7951 & n10880 ) ;
  assign n17808 = n7005 ^ n141 ^ 1'b0 ;
  assign n17809 = n10822 & n17808 ;
  assign n17810 = n15482 & n17809 ;
  assign n17811 = n7865 ^ n129 ^ 1'b0 ;
  assign n17812 = ( n16615 & n17810 ) | ( n16615 & n17811 ) | ( n17810 & n17811 ) ;
  assign n17813 = ( n1592 & n5246 ) | ( n1592 & n17472 ) | ( n5246 & n17472 ) ;
  assign n17814 = n17406 ^ n16117 ^ n4522 ;
  assign n17815 = n15325 ^ n7412 ^ n1830 ;
  assign n17816 = n17814 | n17815 ;
  assign n17817 = n17816 ^ n6297 ^ 1'b0 ;
  assign n17818 = ~n11391 & n17817 ;
  assign n17819 = ~n17813 & n17818 ;
  assign n17821 = n920 & ~n9472 ;
  assign n17822 = n17821 ^ n3560 ^ 1'b0 ;
  assign n17823 = n17822 ^ n8212 ^ n2609 ;
  assign n17820 = n5595 & ~n14536 ;
  assign n17824 = n17823 ^ n17820 ^ 1'b0 ;
  assign n17825 = n16468 ^ n6057 ^ 1'b0 ;
  assign n17826 = n12152 | n17825 ;
  assign n17827 = n3679 | n7806 ;
  assign n17828 = n3791 | n17827 ;
  assign n17829 = n13170 | n17828 ;
  assign n17830 = n10767 ^ n9023 ^ n8686 ;
  assign n17832 = n13003 ^ n3824 ^ n307 ;
  assign n17831 = ( n3879 & n5121 ) | ( n3879 & ~n6375 ) | ( n5121 & ~n6375 ) ;
  assign n17833 = n17832 ^ n17831 ^ n17182 ;
  assign n17834 = n14958 ^ n10663 ^ n3373 ;
  assign n17835 = n17834 ^ n4033 ^ 1'b0 ;
  assign n17836 = n4287 ^ n4111 ^ 1'b0 ;
  assign n17837 = n17836 ^ n17646 ^ 1'b0 ;
  assign n17838 = n17835 & n17837 ;
  assign n17839 = ( n2885 & n4359 ) | ( n2885 & n17337 ) | ( n4359 & n17337 ) ;
  assign n17840 = n439 & n761 ;
  assign n17841 = n17840 ^ n13575 ^ 1'b0 ;
  assign n17842 = n10489 ^ n5603 ^ n693 ;
  assign n17843 = n17842 ^ n2496 ^ 1'b0 ;
  assign n17844 = ~n5996 & n17843 ;
  assign n17845 = n9018 & n16077 ;
  assign n17846 = n7347 | n17845 ;
  assign n17847 = ( ~n2623 & n4723 ) | ( ~n2623 & n16870 ) | ( n4723 & n16870 ) ;
  assign n17848 = n10843 ^ n6169 ^ n2096 ;
  assign n17849 = n17848 ^ n4110 ^ 1'b0 ;
  assign n17850 = n13083 | n17849 ;
  assign n17851 = n12637 ^ n7080 ^ n281 ;
  assign n17852 = n17851 ^ n15639 ^ n12356 ;
  assign n17853 = n17852 ^ n10297 ^ n9120 ;
  assign n17854 = ( ~n5177 & n17850 ) | ( ~n5177 & n17853 ) | ( n17850 & n17853 ) ;
  assign n17855 = ~n1776 & n2288 ;
  assign n17856 = ( n3573 & ~n6765 ) | ( n3573 & n17855 ) | ( ~n6765 & n17855 ) ;
  assign n17857 = n9092 ^ n9089 ^ 1'b0 ;
  assign n17858 = ~n200 & n2542 ;
  assign n17859 = n16838 ^ n11080 ^ 1'b0 ;
  assign n17860 = n14041 ^ n6926 ^ n773 ;
  assign n17861 = n815 & ~n3832 ;
  assign n17862 = ( n1416 & ~n4341 ) | ( n1416 & n17861 ) | ( ~n4341 & n17861 ) ;
  assign n17863 = n11881 ^ n8220 ^ 1'b0 ;
  assign n17864 = n16787 ^ n2106 ^ 1'b0 ;
  assign n17865 = n6337 & ~n17864 ;
  assign n17866 = n13620 ^ n470 ^ 1'b0 ;
  assign n17867 = ~n576 & n17866 ;
  assign n17868 = n3322 & ~n13001 ;
  assign n17869 = n6171 | n17868 ;
  assign n17870 = n17869 ^ n17440 ^ 1'b0 ;
  assign n17871 = ( x77 & ~n12900 ) | ( x77 & n17870 ) | ( ~n12900 & n17870 ) ;
  assign n17872 = ( n2298 & n6701 ) | ( n2298 & n15608 ) | ( n6701 & n15608 ) ;
  assign n17873 = ( ~n4458 & n5396 ) | ( ~n4458 & n12045 ) | ( n5396 & n12045 ) ;
  assign n17879 = ( n612 & n5606 ) | ( n612 & ~n15698 ) | ( n5606 & ~n15698 ) ;
  assign n17874 = n5659 ^ n2399 ^ 1'b0 ;
  assign n17875 = n14094 | n17874 ;
  assign n17876 = n17875 ^ n3831 ^ 1'b0 ;
  assign n17877 = n17876 ^ n14961 ^ n14757 ;
  assign n17878 = ~n12813 & n17877 ;
  assign n17880 = n17879 ^ n17878 ^ 1'b0 ;
  assign n17881 = n17880 ^ n6169 ^ 1'b0 ;
  assign n17882 = n6906 & ~n17881 ;
  assign n17883 = n17882 ^ n3662 ^ n390 ;
  assign n17884 = ( x58 & n529 ) | ( x58 & n6361 ) | ( n529 & n6361 ) ;
  assign n17885 = n1762 & ~n17884 ;
  assign n17886 = n17172 ^ n10627 ^ n2194 ;
  assign n17887 = ~n11326 & n13615 ;
  assign n17888 = n10595 ^ n1886 ^ 1'b0 ;
  assign n17889 = n2500 | n11593 ;
  assign n17890 = n17889 ^ n3073 ^ 1'b0 ;
  assign n17891 = n3175 & ~n17890 ;
  assign n17892 = n17891 ^ n3188 ^ 1'b0 ;
  assign n17893 = n12501 ^ n2347 ^ 1'b0 ;
  assign n17894 = n323 & ~n17893 ;
  assign n17895 = ( n5474 & ~n15492 ) | ( n5474 & n17894 ) | ( ~n15492 & n17894 ) ;
  assign n17896 = ( n15295 & n15514 ) | ( n15295 & ~n15659 ) | ( n15514 & ~n15659 ) ;
  assign n17897 = n17896 ^ n14564 ^ n2603 ;
  assign n17898 = ( n248 & n15257 ) | ( n248 & ~n17897 ) | ( n15257 & ~n17897 ) ;
  assign n17899 = n14789 ^ n11465 ^ 1'b0 ;
  assign n17900 = n4246 & n17899 ;
  assign n17901 = n16229 ^ n6046 ^ n1219 ;
  assign n17902 = n15275 | n17901 ;
  assign n17903 = n1688 ^ n717 ^ 1'b0 ;
  assign n17904 = n8978 & ~n9434 ;
  assign n17905 = n3747 ^ n322 ^ 1'b0 ;
  assign n17906 = ~n1902 & n17905 ;
  assign n17907 = n15274 & n17906 ;
  assign n17908 = n17907 ^ n14097 ^ 1'b0 ;
  assign n17909 = n7112 ^ n3273 ^ 1'b0 ;
  assign n17910 = ( n1124 & ~n10445 ) | ( n1124 & n13109 ) | ( ~n10445 & n13109 ) ;
  assign n17911 = n11198 ^ n3367 ^ n1838 ;
  assign n17912 = n17911 ^ n2938 ^ 1'b0 ;
  assign n17913 = n17912 ^ n8588 ^ n3712 ;
  assign n17914 = n6362 ^ n3727 ^ 1'b0 ;
  assign n17915 = ~n8022 & n17914 ;
  assign n17916 = n17915 ^ n17614 ^ 1'b0 ;
  assign n17917 = ( ~n5180 & n10288 ) | ( ~n5180 & n17916 ) | ( n10288 & n17916 ) ;
  assign n17920 = ( n3498 & ~n3782 ) | ( n3498 & n17310 ) | ( ~n3782 & n17310 ) ;
  assign n17918 = n9573 & ~n12386 ;
  assign n17919 = ~n4081 & n17918 ;
  assign n17921 = n17920 ^ n17919 ^ 1'b0 ;
  assign n17922 = n14388 & ~n17396 ;
  assign n17923 = ~n13613 & n17922 ;
  assign n17924 = n10184 & ~n13188 ;
  assign n17925 = n13247 ^ n8775 ^ n8294 ;
  assign n17927 = ( n3751 & n17510 ) | ( n3751 & n17811 ) | ( n17510 & n17811 ) ;
  assign n17926 = ( n2339 & ~n6588 ) | ( n2339 & n10506 ) | ( ~n6588 & n10506 ) ;
  assign n17928 = n17927 ^ n17926 ^ n2595 ;
  assign n17931 = n293 | n11526 ;
  assign n17932 = n3005 | n17931 ;
  assign n17929 = ( ~n4938 & n7190 ) | ( ~n4938 & n10284 ) | ( n7190 & n10284 ) ;
  assign n17930 = n15615 & n17929 ;
  assign n17933 = n17932 ^ n17930 ^ 1'b0 ;
  assign n17934 = n2227 ^ n1993 ^ 1'b0 ;
  assign n17935 = n7726 ^ n930 ^ 1'b0 ;
  assign n17936 = n9242 ^ n5073 ^ n3644 ;
  assign n17937 = n1570 | n15854 ;
  assign n17938 = n6122 & ~n17937 ;
  assign n17939 = n3774 ^ n2563 ^ 1'b0 ;
  assign n17940 = ~n8130 & n17939 ;
  assign n17941 = n807 & n14543 ;
  assign n17942 = ( n12952 & ~n17940 ) | ( n12952 & n17941 ) | ( ~n17940 & n17941 ) ;
  assign n17943 = n12704 ^ n8416 ^ 1'b0 ;
  assign n17944 = n11855 | n17943 ;
  assign n17945 = n17944 ^ n8456 ^ n6283 ;
  assign n17946 = n17942 & n17945 ;
  assign n17947 = n17946 ^ n11059 ^ 1'b0 ;
  assign n17948 = ~n6303 & n11101 ;
  assign n17949 = n17948 ^ n3055 ^ 1'b0 ;
  assign n17950 = n7824 | n17949 ;
  assign n17951 = n17950 ^ n7827 ^ 1'b0 ;
  assign n17952 = n17951 ^ n6875 ^ 1'b0 ;
  assign n17953 = n3759 ^ n2561 ^ n696 ;
  assign n17954 = n17953 ^ n13612 ^ 1'b0 ;
  assign n17955 = n4956 ^ n2724 ^ 1'b0 ;
  assign n17958 = n13298 ^ n12425 ^ 1'b0 ;
  assign n17957 = n11889 ^ n9988 ^ n4124 ;
  assign n17956 = n4263 | n15773 ;
  assign n17959 = n17958 ^ n17957 ^ n17956 ;
  assign n17960 = n3576 & ~n17959 ;
  assign n17961 = n5180 & ~n9216 ;
  assign n17962 = n17961 ^ n151 ^ 1'b0 ;
  assign n17963 = n2178 & ~n13810 ;
  assign n17964 = n4980 | n17963 ;
  assign n17968 = n17355 ^ n9343 ^ 1'b0 ;
  assign n17965 = n5124 & n11262 ;
  assign n17966 = n6190 & n17965 ;
  assign n17967 = n17966 ^ n5563 ^ n4280 ;
  assign n17969 = n17968 ^ n17967 ^ 1'b0 ;
  assign n17970 = n10491 & ~n17969 ;
  assign n17971 = n17970 ^ n8616 ^ n7492 ;
  assign n17972 = n13355 ^ n8069 ^ n5178 ;
  assign n17973 = n3447 & ~n17972 ;
  assign n17974 = n6085 ^ n647 ^ 1'b0 ;
  assign n17975 = n17974 ^ n13834 ^ n6775 ;
  assign n17976 = n5259 | n17975 ;
  assign n17977 = ( x59 & n10242 ) | ( x59 & ~n17976 ) | ( n10242 & ~n17976 ) ;
  assign n17978 = n15281 & n17977 ;
  assign n17980 = n3996 ^ n3844 ^ 1'b0 ;
  assign n17981 = n17980 ^ n4331 ^ 1'b0 ;
  assign n17982 = n6879 | n17981 ;
  assign n17979 = n5320 | n8683 ;
  assign n17983 = n17982 ^ n17979 ^ 1'b0 ;
  assign n17984 = ( n3178 & n11009 ) | ( n3178 & ~n17983 ) | ( n11009 & ~n17983 ) ;
  assign n17985 = ( ~n1649 & n10580 ) | ( ~n1649 & n17984 ) | ( n10580 & n17984 ) ;
  assign n17986 = n14608 ^ n6963 ^ 1'b0 ;
  assign n17987 = n339 & ~n17986 ;
  assign n17988 = n4075 & ~n17987 ;
  assign n17989 = n15178 ^ n13288 ^ n7774 ;
  assign n17990 = n17989 ^ n6533 ^ n5905 ;
  assign n17991 = n17990 ^ n4367 ^ 1'b0 ;
  assign n17992 = n11339 ^ n1726 ^ 1'b0 ;
  assign n17993 = n3862 | n17992 ;
  assign n17994 = n16854 ^ n12611 ^ n8729 ;
  assign n17995 = ( n3394 & n7412 ) | ( n3394 & ~n9230 ) | ( n7412 & ~n9230 ) ;
  assign n17996 = n10360 ^ n3296 ^ n933 ;
  assign n17997 = n13130 ^ n9870 ^ n1794 ;
  assign n17998 = n2141 & n10558 ;
  assign n17999 = n6534 ^ n421 ^ 1'b0 ;
  assign n18000 = n17998 | n17999 ;
  assign n18001 = n14010 ^ n12001 ^ n6162 ;
  assign n18002 = n12487 & n18001 ;
  assign n18003 = n18002 ^ n10871 ^ 1'b0 ;
  assign n18004 = ~n3462 & n8039 ;
  assign n18005 = n10000 & n18004 ;
  assign n18006 = n246 & ~n18005 ;
  assign n18007 = n18006 ^ n8077 ^ 1'b0 ;
  assign n18008 = n5811 | n15930 ;
  assign n18009 = n14554 & ~n18008 ;
  assign n18010 = n14536 ^ n3923 ^ n2684 ;
  assign n18011 = ~n8514 & n18010 ;
  assign n18012 = ( ~n4048 & n8002 ) | ( ~n4048 & n16365 ) | ( n8002 & n16365 ) ;
  assign n18013 = n14926 ^ n4501 ^ 1'b0 ;
  assign n18015 = n4067 ^ n1921 ^ 1'b0 ;
  assign n18016 = n5234 ^ n4680 ^ 1'b0 ;
  assign n18017 = ( n15873 & n18015 ) | ( n15873 & ~n18016 ) | ( n18015 & ~n18016 ) ;
  assign n18014 = n10926 | n15219 ;
  assign n18018 = n18017 ^ n18014 ^ 1'b0 ;
  assign n18019 = ( ~n2776 & n3590 ) | ( ~n2776 & n8454 ) | ( n3590 & n8454 ) ;
  assign n18020 = ~n3585 & n18019 ;
  assign n18021 = n13279 & n18020 ;
  assign n18022 = ( n1882 & n8170 ) | ( n1882 & ~n8429 ) | ( n8170 & ~n8429 ) ;
  assign n18023 = n5533 & ~n18022 ;
  assign n18024 = n18023 ^ n3768 ^ n2019 ;
  assign n18025 = ~n7910 & n18024 ;
  assign n18026 = n877 & ~n4838 ;
  assign n18027 = n8437 & n18026 ;
  assign n18028 = ( n7325 & ~n12062 ) | ( n7325 & n18027 ) | ( ~n12062 & n18027 ) ;
  assign n18029 = ( n12328 & n13774 ) | ( n12328 & ~n15802 ) | ( n13774 & ~n15802 ) ;
  assign n18030 = n7647 ^ n2805 ^ 1'b0 ;
  assign n18031 = n14757 ^ n6945 ^ 1'b0 ;
  assign n18032 = ~n18030 & n18031 ;
  assign n18033 = n10872 & ~n17614 ;
  assign n18034 = ~n3411 & n13413 ;
  assign n18035 = ( n7914 & n11091 ) | ( n7914 & n18034 ) | ( n11091 & n18034 ) ;
  assign n18036 = ~n1541 & n2296 ;
  assign n18037 = n18036 ^ n4138 ^ 1'b0 ;
  assign n18038 = ~n14822 & n18037 ;
  assign n18039 = n7187 & ~n18038 ;
  assign n18043 = ~n2478 & n8938 ;
  assign n18044 = n6891 & n18043 ;
  assign n18040 = x26 & ~n5249 ;
  assign n18041 = n18040 ^ n5301 ^ 1'b0 ;
  assign n18042 = n16343 & n18041 ;
  assign n18045 = n18044 ^ n18042 ^ 1'b0 ;
  assign n18046 = ( ~n4711 & n17690 ) | ( ~n4711 & n18045 ) | ( n17690 & n18045 ) ;
  assign n18047 = x1 & n717 ;
  assign n18048 = n15990 & n18047 ;
  assign n18049 = n18048 ^ n6185 ^ n2323 ;
  assign n18050 = n8887 | n18049 ;
  assign n18051 = ( n1611 & n14216 ) | ( n1611 & ~n17242 ) | ( n14216 & ~n17242 ) ;
  assign n18052 = ~n5291 & n9748 ;
  assign n18053 = n18052 ^ n5120 ^ 1'b0 ;
  assign n18054 = n7267 & n18053 ;
  assign n18055 = n18051 & n18054 ;
  assign n18056 = n8451 ^ n5535 ^ 1'b0 ;
  assign n18057 = ( ~x19 & n7320 ) | ( ~x19 & n18056 ) | ( n7320 & n18056 ) ;
  assign n18058 = n18057 ^ n203 ^ 1'b0 ;
  assign n18059 = n2666 & n18058 ;
  assign n18060 = n8565 & n18059 ;
  assign n18061 = ~n18055 & n18060 ;
  assign n18062 = n6197 ^ n2457 ^ 1'b0 ;
  assign n18063 = ( ~n232 & n5266 ) | ( ~n232 & n10225 ) | ( n5266 & n10225 ) ;
  assign n18064 = n983 & ~n9082 ;
  assign n18065 = n18063 & n18064 ;
  assign n18066 = ~n5000 & n18065 ;
  assign n18067 = ( n12481 & ~n18062 ) | ( n12481 & n18066 ) | ( ~n18062 & n18066 ) ;
  assign n18068 = ( ~n12642 & n15026 ) | ( ~n12642 & n16672 ) | ( n15026 & n16672 ) ;
  assign n18070 = n9911 ^ n2157 ^ 1'b0 ;
  assign n18069 = n457 & n2056 ;
  assign n18071 = n18070 ^ n18069 ^ 1'b0 ;
  assign n18072 = n9728 ^ n4971 ^ 1'b0 ;
  assign n18073 = n6414 | n18072 ;
  assign n18074 = n672 & n4543 ;
  assign n18075 = n18073 & n18074 ;
  assign n18076 = n2010 ^ n479 ^ 1'b0 ;
  assign n18077 = n18075 | n18076 ;
  assign n18078 = ~n4427 & n9170 ;
  assign n18079 = ~n1862 & n18078 ;
  assign n18080 = ( n2730 & n3483 ) | ( n2730 & n8282 ) | ( n3483 & n8282 ) ;
  assign n18081 = n7930 ^ n6187 ^ 1'b0 ;
  assign n18082 = n1964 & n18081 ;
  assign n18083 = ~n4156 & n4315 ;
  assign n18084 = n18083 ^ n10285 ^ n7791 ;
  assign n18085 = ~n8710 & n18084 ;
  assign n18086 = ~n18082 & n18085 ;
  assign n18089 = n7203 ^ n4842 ^ 1'b0 ;
  assign n18090 = ~n6453 & n18089 ;
  assign n18091 = n4859 | n9660 ;
  assign n18092 = n18091 ^ n12690 ^ 1'b0 ;
  assign n18093 = ( n307 & n18090 ) | ( n307 & ~n18092 ) | ( n18090 & ~n18092 ) ;
  assign n18087 = ( ~n1292 & n7987 ) | ( ~n1292 & n11814 ) | ( n7987 & n11814 ) ;
  assign n18088 = n13755 & ~n18087 ;
  assign n18094 = n18093 ^ n18088 ^ 1'b0 ;
  assign n18095 = n7739 ^ n4469 ^ n1204 ;
  assign n18098 = n7503 | n8714 ;
  assign n18099 = n5932 & ~n18098 ;
  assign n18096 = n5353 ^ n2778 ^ n1821 ;
  assign n18097 = n11890 | n18096 ;
  assign n18100 = n18099 ^ n18097 ^ 1'b0 ;
  assign n18101 = n18095 | n18100 ;
  assign n18102 = ~n3008 & n6202 ;
  assign n18103 = ( ~n888 & n903 ) | ( ~n888 & n18102 ) | ( n903 & n18102 ) ;
  assign n18104 = n8354 ^ n4736 ^ 1'b0 ;
  assign n18105 = n7368 | n8936 ;
  assign n18106 = n18105 ^ n2163 ^ 1'b0 ;
  assign n18107 = n2729 & n18106 ;
  assign n18108 = n18104 & n18107 ;
  assign n18109 = n3599 | n18108 ;
  assign n18110 = n17399 & ~n18109 ;
  assign n18111 = ( n8298 & n18103 ) | ( n8298 & ~n18110 ) | ( n18103 & ~n18110 ) ;
  assign n18112 = ( ~n3588 & n9876 ) | ( ~n3588 & n10469 ) | ( n9876 & n10469 ) ;
  assign n18113 = n15855 ^ n2641 ^ 1'b0 ;
  assign n18114 = ~n4259 & n16796 ;
  assign n18115 = ~n18113 & n18114 ;
  assign n18116 = ~n9569 & n15482 ;
  assign n18117 = n4185 ^ n3826 ^ 1'b0 ;
  assign n18118 = ( ~n8101 & n16918 ) | ( ~n8101 & n18117 ) | ( n16918 & n18117 ) ;
  assign n18119 = n9928 ^ n3276 ^ 1'b0 ;
  assign n18120 = ~n18118 & n18119 ;
  assign n18121 = ( n1053 & n6136 ) | ( n1053 & ~n9349 ) | ( n6136 & ~n9349 ) ;
  assign n18122 = n18121 ^ n14260 ^ n11910 ;
  assign n18123 = n7966 | n8529 ;
  assign n18124 = ~n6754 & n15837 ;
  assign n18125 = n17653 & n18124 ;
  assign n18126 = n5905 & n8757 ;
  assign n18127 = ( n8724 & n10674 ) | ( n8724 & n17283 ) | ( n10674 & n17283 ) ;
  assign n18128 = n1980 ^ n1714 ^ 1'b0 ;
  assign n18130 = ( n976 & n1580 ) | ( n976 & ~n7542 ) | ( n1580 & ~n7542 ) ;
  assign n18131 = n18130 ^ n13283 ^ n6922 ;
  assign n18129 = n1033 & ~n3500 ;
  assign n18132 = n18131 ^ n18129 ^ 1'b0 ;
  assign n18133 = n6143 ^ n6139 ^ n471 ;
  assign n18134 = n18133 ^ n9921 ^ 1'b0 ;
  assign n18135 = n12073 & ~n18134 ;
  assign n18138 = x124 ^ x79 ^ 1'b0 ;
  assign n18139 = ~n4538 & n18138 ;
  assign n18136 = n1637 | n10481 ;
  assign n18137 = ( ~n3792 & n11357 ) | ( ~n3792 & n18136 ) | ( n11357 & n18136 ) ;
  assign n18140 = n18139 ^ n18137 ^ n12811 ;
  assign n18141 = n6665 ^ n3740 ^ n3185 ;
  assign n18142 = n4061 | n18141 ;
  assign n18143 = n18142 ^ n15707 ^ n1836 ;
  assign n18144 = n18143 ^ n4680 ^ n3173 ;
  assign n18145 = n15574 ^ n9205 ^ 1'b0 ;
  assign n18146 = n12248 & n18145 ;
  assign n18148 = n1683 ^ n334 ^ 1'b0 ;
  assign n18149 = n1626 & n18148 ;
  assign n18150 = ( n13567 & ~n15418 ) | ( n13567 & n18149 ) | ( ~n15418 & n18149 ) ;
  assign n18147 = n4101 & ~n6518 ;
  assign n18151 = n18150 ^ n18147 ^ 1'b0 ;
  assign n18152 = n6150 | n10993 ;
  assign n18153 = n18152 ^ n9664 ^ n4854 ;
  assign n18154 = n18153 ^ n12663 ^ n2578 ;
  assign n18155 = n15859 ^ n11820 ^ n9195 ;
  assign n18156 = ( n1990 & n2794 ) | ( n1990 & n10111 ) | ( n2794 & n10111 ) ;
  assign n18157 = ( n4502 & ~n8061 ) | ( n4502 & n17508 ) | ( ~n8061 & n17508 ) ;
  assign n18158 = n1830 | n11136 ;
  assign n18159 = n18158 ^ n14511 ^ n8166 ;
  assign n18160 = n2824 | n9079 ;
  assign n18161 = n5986 | n18160 ;
  assign n18162 = n6085 | n12712 ;
  assign n18163 = n18161 | n18162 ;
  assign n18164 = ( x113 & n11339 ) | ( x113 & ~n12722 ) | ( n11339 & ~n12722 ) ;
  assign n18165 = ( n2370 & n14245 ) | ( n2370 & n18164 ) | ( n14245 & n18164 ) ;
  assign n18166 = ( ~n905 & n1185 ) | ( ~n905 & n11487 ) | ( n1185 & n11487 ) ;
  assign n18167 = n8237 | n18166 ;
  assign n18168 = n5313 | n18167 ;
  assign n18169 = ( n3192 & n12491 ) | ( n3192 & ~n18168 ) | ( n12491 & ~n18168 ) ;
  assign n18170 = n15970 ^ n4332 ^ n2627 ;
  assign n18171 = n869 & n5891 ;
  assign n18172 = n12465 | n18171 ;
  assign n18173 = n8275 | n18172 ;
  assign n18175 = ~n1903 & n11804 ;
  assign n18176 = n18175 ^ n5302 ^ 1'b0 ;
  assign n18177 = n4727 | n14177 ;
  assign n18178 = n18176 & ~n18177 ;
  assign n18174 = n5322 & ~n7291 ;
  assign n18179 = n18178 ^ n18174 ^ 1'b0 ;
  assign n18181 = n9223 ^ n9016 ^ 1'b0 ;
  assign n18182 = ~n16323 & n18181 ;
  assign n18183 = ~n2931 & n18182 ;
  assign n18184 = n18183 ^ n11062 ^ 1'b0 ;
  assign n18180 = n890 & n8838 ;
  assign n18185 = n18184 ^ n18180 ^ 1'b0 ;
  assign n18190 = n9744 ^ n8322 ^ n5848 ;
  assign n18186 = n3721 ^ n3190 ^ 1'b0 ;
  assign n18187 = ( ~n5013 & n6967 ) | ( ~n5013 & n18186 ) | ( n6967 & n18186 ) ;
  assign n18188 = ~n1193 & n5819 ;
  assign n18189 = n18187 | n18188 ;
  assign n18191 = n18190 ^ n18189 ^ 1'b0 ;
  assign n18192 = n10320 ^ n2072 ^ 1'b0 ;
  assign n18193 = n3349 & ~n18192 ;
  assign n18194 = ( n6469 & n17583 ) | ( n6469 & ~n18193 ) | ( n17583 & ~n18193 ) ;
  assign n18195 = n12637 & n14098 ;
  assign n18196 = n3247 ^ n2209 ^ x49 ;
  assign n18198 = n4583 ^ n804 ^ 1'b0 ;
  assign n18197 = n16751 | n17739 ;
  assign n18199 = n18198 ^ n18197 ^ 1'b0 ;
  assign n18202 = n1673 ^ n1561 ^ n232 ;
  assign n18200 = n3555 ^ n2990 ^ 1'b0 ;
  assign n18201 = n8824 & n18200 ;
  assign n18203 = n18202 ^ n18201 ^ 1'b0 ;
  assign n18204 = n9902 ^ n1753 ^ 1'b0 ;
  assign n18205 = n4941 | n18204 ;
  assign n18206 = ( n11192 & ~n11357 ) | ( n11192 & n11712 ) | ( ~n11357 & n11712 ) ;
  assign n18207 = n18206 ^ n9460 ^ 1'b0 ;
  assign n18208 = n2487 & ~n18207 ;
  assign n18209 = n18208 ^ n12950 ^ 1'b0 ;
  assign n18210 = n6007 & n14872 ;
  assign n18211 = n8523 & n11801 ;
  assign n18212 = ( n506 & n2691 ) | ( n506 & n9715 ) | ( n2691 & n9715 ) ;
  assign n18213 = ( n3678 & n3950 ) | ( n3678 & n18212 ) | ( n3950 & n18212 ) ;
  assign n18214 = n18213 ^ n3176 ^ n1370 ;
  assign n18215 = ( n1840 & ~n15846 ) | ( n1840 & n18214 ) | ( ~n15846 & n18214 ) ;
  assign n18216 = n348 | n18215 ;
  assign n18217 = n12132 | n18216 ;
  assign n18218 = n1178 & ~n13281 ;
  assign n18219 = n12371 ^ n2264 ^ 1'b0 ;
  assign n18220 = n18219 ^ n7951 ^ 1'b0 ;
  assign n18221 = ~n4082 & n18220 ;
  assign n18222 = n767 | n10380 ;
  assign n18223 = ( ~n11815 & n18221 ) | ( ~n11815 & n18222 ) | ( n18221 & n18222 ) ;
  assign n18224 = n960 & ~n1793 ;
  assign n18225 = n9660 & n18224 ;
  assign n18226 = n18225 ^ n15733 ^ n7740 ;
  assign n18227 = n18226 ^ n1104 ^ 1'b0 ;
  assign n18228 = n8500 & ~n11694 ;
  assign n18229 = n2802 & ~n9965 ;
  assign n18230 = n18229 ^ n5369 ^ 1'b0 ;
  assign n18231 = n18230 ^ n18187 ^ n2013 ;
  assign n18232 = n5805 & n11967 ;
  assign n18233 = n18232 ^ n13212 ^ 1'b0 ;
  assign n18234 = ~n5875 & n11922 ;
  assign n18235 = ( n4475 & ~n6126 ) | ( n4475 & n9497 ) | ( ~n6126 & n9497 ) ;
  assign n18236 = ( n7136 & n11444 ) | ( n7136 & n18235 ) | ( n11444 & n18235 ) ;
  assign n18237 = n18236 ^ n13480 ^ 1'b0 ;
  assign n18238 = ~n4989 & n8256 ;
  assign n18239 = n18238 ^ n17350 ^ 1'b0 ;
  assign n18240 = ~n6026 & n18239 ;
  assign n18241 = n18240 ^ n2618 ^ 1'b0 ;
  assign n18242 = n17941 ^ n2326 ^ 1'b0 ;
  assign n18245 = ( n8530 & ~n11093 ) | ( n8530 & n13447 ) | ( ~n11093 & n13447 ) ;
  assign n18246 = n18245 ^ n14326 ^ x120 ;
  assign n18243 = n8521 | n8637 ;
  assign n18244 = n18149 & ~n18243 ;
  assign n18247 = n18246 ^ n18244 ^ n3803 ;
  assign n18248 = n15586 ^ n9949 ^ n7714 ;
  assign n18249 = n11737 ^ n6557 ^ n1527 ;
  assign n18250 = ( n3671 & ~n10080 ) | ( n3671 & n15824 ) | ( ~n10080 & n15824 ) ;
  assign n18251 = n18250 ^ n4850 ^ 1'b0 ;
  assign n18252 = n13708 & n18251 ;
  assign n18253 = n2360 & n18252 ;
  assign n18254 = ( ~n4131 & n7457 ) | ( ~n4131 & n8516 ) | ( n7457 & n8516 ) ;
  assign n18255 = n18254 ^ n580 ^ 1'b0 ;
  assign n18256 = ( ~n6491 & n12213 ) | ( ~n6491 & n18255 ) | ( n12213 & n18255 ) ;
  assign n18257 = ( n2401 & ~n2557 ) | ( n2401 & n12735 ) | ( ~n2557 & n12735 ) ;
  assign n18258 = ( ~n307 & n2059 ) | ( ~n307 & n18257 ) | ( n2059 & n18257 ) ;
  assign n18259 = n12382 ^ n5894 ^ 1'b0 ;
  assign n18261 = n4304 | n5632 ;
  assign n18262 = n9506 | n18261 ;
  assign n18260 = n9433 & n14441 ;
  assign n18263 = n18262 ^ n18260 ^ n15377 ;
  assign n18264 = ( ~n1548 & n1891 ) | ( ~n1548 & n7042 ) | ( n1891 & n7042 ) ;
  assign n18265 = n18264 ^ n663 ^ 1'b0 ;
  assign n18267 = n1208 & ~n2086 ;
  assign n18268 = n8037 & ~n18267 ;
  assign n18266 = n3757 | n5495 ;
  assign n18269 = n18268 ^ n18266 ^ 1'b0 ;
  assign n18270 = n18146 ^ n4451 ^ 1'b0 ;
  assign n18271 = n9850 ^ n3120 ^ 1'b0 ;
  assign n18272 = ( n3841 & ~n7646 ) | ( n3841 & n7913 ) | ( ~n7646 & n7913 ) ;
  assign n18273 = n14643 ^ n14629 ^ n1785 ;
  assign n18274 = ~n1779 & n15428 ;
  assign n18275 = ~n9331 & n18274 ;
  assign n18276 = ~n6903 & n18275 ;
  assign n18277 = n8019 | n13324 ;
  assign n18278 = n5629 | n18277 ;
  assign n18279 = n2328 | n5376 ;
  assign n18280 = n16735 | n18279 ;
  assign n18281 = ~n1580 & n18280 ;
  assign n18282 = ~n3162 & n4510 ;
  assign n18283 = ( ~n8456 & n14758 ) | ( ~n8456 & n18282 ) | ( n14758 & n18282 ) ;
  assign n18284 = ~n3073 & n12029 ;
  assign n18285 = n14320 | n18284 ;
  assign n18286 = n3461 & ~n10922 ;
  assign n18287 = n8410 ^ n7186 ^ n197 ;
  assign n18288 = n205 ^ n149 ^ 1'b0 ;
  assign n18289 = n2129 & n18288 ;
  assign n18290 = n8298 ^ n4831 ^ 1'b0 ;
  assign n18291 = n14911 & n18290 ;
  assign n18292 = n18291 ^ n13582 ^ n5954 ;
  assign n18293 = n5414 & n17631 ;
  assign n18294 = ( n6828 & ~n17852 ) | ( n6828 & n18293 ) | ( ~n17852 & n18293 ) ;
  assign n18297 = ( ~n5778 & n6042 ) | ( ~n5778 & n12429 ) | ( n6042 & n12429 ) ;
  assign n18295 = ( n429 & n1856 ) | ( n429 & n6860 ) | ( n1856 & n6860 ) ;
  assign n18296 = n18295 ^ n14689 ^ n5387 ;
  assign n18298 = n18297 ^ n18296 ^ n11612 ;
  assign n18299 = ( n10343 & ~n18294 ) | ( n10343 & n18298 ) | ( ~n18294 & n18298 ) ;
  assign n18300 = n7518 ^ n2146 ^ 1'b0 ;
  assign n18301 = ( n2621 & ~n11942 ) | ( n2621 & n18300 ) | ( ~n11942 & n18300 ) ;
  assign n18302 = n919 & n14154 ;
  assign n18303 = n18302 ^ n9281 ^ 1'b0 ;
  assign n18304 = ~n4185 & n13846 ;
  assign n18305 = n13244 & n18304 ;
  assign n18306 = ~n11297 & n18230 ;
  assign n18307 = n18306 ^ n2071 ^ 1'b0 ;
  assign n18308 = n1533 & ~n18307 ;
  assign n18309 = n18308 ^ n15763 ^ n2797 ;
  assign n18310 = n4155 & ~n12945 ;
  assign n18311 = n12782 & n18310 ;
  assign n18313 = ( n2404 & n5621 ) | ( n2404 & n10848 ) | ( n5621 & n10848 ) ;
  assign n18314 = n18313 ^ n9713 ^ n626 ;
  assign n18312 = n15531 & n17120 ;
  assign n18315 = n18314 ^ n18312 ^ 1'b0 ;
  assign n18316 = n18311 | n18315 ;
  assign n18318 = ~n13082 & n15094 ;
  assign n18319 = n18318 ^ n4885 ^ 1'b0 ;
  assign n18317 = ~n1314 & n12373 ;
  assign n18320 = n18319 ^ n18317 ^ 1'b0 ;
  assign n18321 = n8795 & n10556 ;
  assign n18322 = n12316 & n18321 ;
  assign n18323 = n3270 & ~n18322 ;
  assign n18324 = n6494 & ~n7360 ;
  assign n18325 = n7374 ^ n3569 ^ 1'b0 ;
  assign n18326 = n4193 & ~n18325 ;
  assign n18327 = n18326 ^ n1839 ^ n413 ;
  assign n18328 = ~n12081 & n15236 ;
  assign n18329 = n1458 & n2363 ;
  assign n18330 = ~n1354 & n18329 ;
  assign n18331 = n18330 ^ n16924 ^ 1'b0 ;
  assign n18332 = n8288 ^ n4344 ^ x83 ;
  assign n18333 = n14172 ^ n6088 ^ n2334 ;
  assign n18334 = n5021 & ~n18333 ;
  assign n18335 = ( n7422 & n11931 ) | ( n7422 & ~n18334 ) | ( n11931 & ~n18334 ) ;
  assign n18336 = n17921 ^ n8807 ^ 1'b0 ;
  assign n18337 = ~n3120 & n5350 ;
  assign n18338 = n2808 & n5844 ;
  assign n18339 = n11462 & n18338 ;
  assign n18340 = n18339 ^ n14492 ^ 1'b0 ;
  assign n18341 = ( n6158 & ~n8724 ) | ( n6158 & n18340 ) | ( ~n8724 & n18340 ) ;
  assign n18342 = n13977 ^ n11915 ^ n5837 ;
  assign n18343 = n1354 | n5351 ;
  assign n18344 = x101 | n18343 ;
  assign n18345 = n18344 ^ n3239 ^ 1'b0 ;
  assign n18346 = n2348 | n14927 ;
  assign n18347 = n1519 & n9605 ;
  assign n18348 = ( ~n6043 & n18346 ) | ( ~n6043 & n18347 ) | ( n18346 & n18347 ) ;
  assign n18349 = n5600 ^ x15 ^ 1'b0 ;
  assign n18350 = ( n9035 & n13737 ) | ( n9035 & n18349 ) | ( n13737 & n18349 ) ;
  assign n18351 = n18350 ^ n7806 ^ n987 ;
  assign n18352 = n18351 ^ n1696 ^ 1'b0 ;
  assign n18353 = n1550 & ~n18352 ;
  assign n18354 = n1402 ^ n1382 ^ 1'b0 ;
  assign n18355 = ( n1330 & n2407 ) | ( n1330 & n10724 ) | ( n2407 & n10724 ) ;
  assign n18356 = n9471 & n18355 ;
  assign n18357 = n18354 & n18356 ;
  assign n18358 = n667 | n10543 ;
  assign n18359 = n1104 | n18358 ;
  assign n18360 = ~n3222 & n10794 ;
  assign n18361 = ~n18359 & n18360 ;
  assign n18364 = ( n4970 & ~n8835 ) | ( n4970 & n10229 ) | ( ~n8835 & n10229 ) ;
  assign n18362 = n1585 & ~n4320 ;
  assign n18363 = n18362 ^ n447 ^ 1'b0 ;
  assign n18365 = n18364 ^ n18363 ^ n3297 ;
  assign n18366 = n6548 ^ n2114 ^ x33 ;
  assign n18367 = ~n15045 & n18366 ;
  assign n18370 = n14968 ^ n12091 ^ 1'b0 ;
  assign n18371 = ~n2231 & n18370 ;
  assign n18368 = n7471 & n8510 ;
  assign n18369 = n18368 ^ n6378 ^ 1'b0 ;
  assign n18372 = n18371 ^ n18369 ^ n4073 ;
  assign n18373 = ( n8061 & n8174 ) | ( n8061 & n16765 ) | ( n8174 & n16765 ) ;
  assign n18374 = n6343 & n9201 ;
  assign n18375 = n18374 ^ n12260 ^ 1'b0 ;
  assign n18376 = ( n6330 & n18373 ) | ( n6330 & n18375 ) | ( n18373 & n18375 ) ;
  assign n18377 = ~n4071 & n7450 ;
  assign n18378 = n18377 ^ n15759 ^ 1'b0 ;
  assign n18379 = ~n4741 & n10229 ;
  assign n18380 = n18379 ^ n15202 ^ 1'b0 ;
  assign n18381 = n6226 ^ n6169 ^ n4156 ;
  assign n18382 = n18381 ^ n16776 ^ 1'b0 ;
  assign n18383 = n2532 & ~n18382 ;
  assign n18384 = n429 & n1082 ;
  assign n18385 = n1456 & ~n10018 ;
  assign n18386 = n18385 ^ n9307 ^ 1'b0 ;
  assign n18387 = ( ~n6458 & n15483 ) | ( ~n6458 & n18386 ) | ( n15483 & n18386 ) ;
  assign n18388 = n15526 ^ n14289 ^ x83 ;
  assign n18389 = n14021 ^ n5305 ^ 1'b0 ;
  assign n18390 = n10247 & ~n18389 ;
  assign n18394 = n7749 ^ n4247 ^ n3798 ;
  assign n18395 = n18394 ^ n13124 ^ 1'b0 ;
  assign n18396 = n3614 | n18395 ;
  assign n18391 = n1319 & n2389 ;
  assign n18392 = ~n2839 & n18391 ;
  assign n18393 = n11008 & ~n18392 ;
  assign n18397 = n18396 ^ n18393 ^ 1'b0 ;
  assign n18398 = n2334 & ~n9176 ;
  assign n18399 = n12073 ^ n5370 ^ 1'b0 ;
  assign n18400 = x106 & n18399 ;
  assign n18401 = n18400 ^ n17209 ^ 1'b0 ;
  assign n18402 = n13058 | n18401 ;
  assign n18403 = n3508 & ~n7520 ;
  assign n18404 = n18403 ^ n7207 ^ 1'b0 ;
  assign n18405 = n2356 & n13613 ;
  assign n18406 = ( ~n3975 & n11289 ) | ( ~n3975 & n11443 ) | ( n11289 & n11443 ) ;
  assign n18407 = n18405 | n18406 ;
  assign n18408 = n18407 ^ n12503 ^ 1'b0 ;
  assign n18409 = n18408 ^ n16281 ^ 1'b0 ;
  assign n18410 = n3426 & ~n18409 ;
  assign n18411 = ( n16096 & n18404 ) | ( n16096 & n18410 ) | ( n18404 & n18410 ) ;
  assign n18412 = n18411 ^ n4618 ^ n3718 ;
  assign n18413 = n7180 ^ n5127 ^ n2138 ;
  assign n18414 = n14915 ^ x126 ^ 1'b0 ;
  assign n18415 = n1989 & n7085 ;
  assign n18416 = n14921 ^ n8883 ^ n6281 ;
  assign n18417 = n18416 ^ n4118 ^ 1'b0 ;
  assign n18418 = ~n18415 & n18417 ;
  assign n18419 = n16722 ^ n15600 ^ n3711 ;
  assign n18420 = n18419 ^ n6104 ^ 1'b0 ;
  assign n18421 = n12229 ^ n3448 ^ 1'b0 ;
  assign n18422 = n3449 | n18421 ;
  assign n18423 = ( n456 & n3947 ) | ( n456 & ~n9507 ) | ( n3947 & ~n9507 ) ;
  assign n18424 = ( ~n4177 & n13400 ) | ( ~n4177 & n14919 ) | ( n13400 & n14919 ) ;
  assign n18425 = ~n3321 & n4193 ;
  assign n18426 = n18117 & n18425 ;
  assign n18427 = n7866 & ~n15771 ;
  assign n18428 = n18427 ^ n13661 ^ 1'b0 ;
  assign n18429 = ( ~n6452 & n7746 ) | ( ~n6452 & n8691 ) | ( n7746 & n8691 ) ;
  assign n18430 = n5282 | n18429 ;
  assign n18431 = ( n4805 & ~n5952 ) | ( n4805 & n8629 ) | ( ~n5952 & n8629 ) ;
  assign n18432 = n9261 & n18431 ;
  assign n18433 = n4745 & n18432 ;
  assign n18434 = n7094 ^ n1654 ^ 1'b0 ;
  assign n18435 = n2589 & n18434 ;
  assign n18436 = ( n15212 & n17822 ) | ( n15212 & n18435 ) | ( n17822 & n18435 ) ;
  assign n18438 = ( n2278 & n8359 ) | ( n2278 & ~n12372 ) | ( n8359 & ~n12372 ) ;
  assign n18437 = ( n13871 & n16389 ) | ( n13871 & ~n17339 ) | ( n16389 & ~n17339 ) ;
  assign n18439 = n18438 ^ n18437 ^ n15754 ;
  assign n18440 = n8679 ^ n7900 ^ n3715 ;
  assign n18441 = n996 | n7531 ;
  assign n18442 = n18441 ^ n1835 ^ 1'b0 ;
  assign n18443 = n5156 ^ n1075 ^ 1'b0 ;
  assign n18444 = ~n2338 & n18443 ;
  assign n18445 = n13298 & ~n14609 ;
  assign n18446 = n6489 | n18445 ;
  assign n18447 = n428 | n18446 ;
  assign n18448 = ~n1076 & n2154 ;
  assign n18449 = n18448 ^ n14149 ^ 1'b0 ;
  assign n18450 = x92 & ~n15754 ;
  assign n18451 = ~n18449 & n18450 ;
  assign n18452 = ~n5351 & n10677 ;
  assign n18453 = n11625 ^ n11473 ^ n4121 ;
  assign n18454 = n18453 ^ n13434 ^ n7911 ;
  assign n18455 = n2941 | n13695 ;
  assign n18456 = n8529 & ~n18455 ;
  assign n18457 = ~n2881 & n9284 ;
  assign n18458 = ( n14985 & n18456 ) | ( n14985 & n18457 ) | ( n18456 & n18457 ) ;
  assign n18459 = n4874 ^ n4732 ^ 1'b0 ;
  assign n18460 = n12750 ^ n4266 ^ 1'b0 ;
  assign n18461 = n18459 & ~n18460 ;
  assign n18462 = n5224 & n18461 ;
  assign n18463 = n5384 | n5556 ;
  assign n18464 = n7367 & n15879 ;
  assign n18465 = n9931 ^ n6713 ^ n4819 ;
  assign n18466 = n10790 ^ n3784 ^ 1'b0 ;
  assign n18467 = n9928 & ~n18466 ;
  assign n18468 = n17786 ^ n9256 ^ 1'b0 ;
  assign n18469 = ~n8782 & n18468 ;
  assign n18470 = n17702 ^ n7636 ^ n7105 ;
  assign n18473 = n4609 & ~n12058 ;
  assign n18474 = n18473 ^ n3409 ^ 1'b0 ;
  assign n18471 = ~n3750 & n16735 ;
  assign n18472 = n18471 ^ x23 ^ 1'b0 ;
  assign n18475 = n18474 ^ n18472 ^ n13416 ;
  assign n18476 = n12275 ^ n4516 ^ 1'b0 ;
  assign n18477 = n18476 ^ n16676 ^ 1'b0 ;
  assign n18478 = n365 & ~n18477 ;
  assign n18479 = ( n5177 & ~n18475 ) | ( n5177 & n18478 ) | ( ~n18475 & n18478 ) ;
  assign n18480 = ~n18470 & n18479 ;
  assign n18481 = n18480 ^ n11080 ^ 1'b0 ;
  assign n18482 = n2386 | n16756 ;
  assign n18483 = n12793 | n18482 ;
  assign n18484 = n8482 ^ n6777 ^ n4821 ;
  assign n18485 = n18484 ^ n8239 ^ 1'b0 ;
  assign n18486 = n18483 & ~n18485 ;
  assign n18487 = n18486 ^ n12960 ^ 1'b0 ;
  assign n18489 = n10751 ^ n7415 ^ 1'b0 ;
  assign n18490 = n4075 & n18489 ;
  assign n18488 = n14273 & ~n16888 ;
  assign n18491 = n18490 ^ n18488 ^ n3164 ;
  assign n18492 = n13137 ^ n6079 ^ n4597 ;
  assign n18493 = ( n7314 & n9859 ) | ( n7314 & n13410 ) | ( n9859 & n13410 ) ;
  assign n18494 = ( n17750 & n18492 ) | ( n17750 & n18493 ) | ( n18492 & n18493 ) ;
  assign n18495 = n5729 & n9849 ;
  assign n18496 = n18495 ^ n5402 ^ 1'b0 ;
  assign n18497 = n18496 ^ n9609 ^ 1'b0 ;
  assign n18498 = n14353 ^ n11187 ^ n635 ;
  assign n18499 = ~n1939 & n15465 ;
  assign n18500 = n18499 ^ n14750 ^ 1'b0 ;
  assign n18501 = n18500 ^ n9254 ^ 1'b0 ;
  assign n18502 = n10534 | n18501 ;
  assign n18503 = n11931 ^ n5147 ^ n4005 ;
  assign n18504 = ( n4185 & ~n10443 ) | ( n4185 & n18503 ) | ( ~n10443 & n18503 ) ;
  assign n18505 = n1858 & ~n14966 ;
  assign n18506 = n18505 ^ n2698 ^ 1'b0 ;
  assign n18507 = n18506 ^ n3624 ^ n498 ;
  assign n18508 = ~n454 & n18507 ;
  assign n18509 = ~n9441 & n18508 ;
  assign n18510 = n296 | n18509 ;
  assign n18511 = n16527 ^ n10324 ^ 1'b0 ;
  assign n18512 = n18511 ^ n10529 ^ n10475 ;
  assign n18513 = n1188 & ~n11496 ;
  assign n18514 = ~n1534 & n18513 ;
  assign n18515 = n18514 ^ n12707 ^ n6554 ;
  assign n18516 = n18515 ^ n875 ^ 1'b0 ;
  assign n18517 = n2181 & ~n18516 ;
  assign n18519 = n8422 ^ n5702 ^ 1'b0 ;
  assign n18518 = ~n4905 & n12704 ;
  assign n18520 = n18519 ^ n18518 ^ 1'b0 ;
  assign n18521 = ( x18 & ~n11438 ) | ( x18 & n11982 ) | ( ~n11438 & n11982 ) ;
  assign n18522 = n18521 ^ n3696 ^ 1'b0 ;
  assign n18523 = ~n5096 & n18522 ;
  assign n18524 = n1853 | n2146 ;
  assign n18525 = n746 & n18524 ;
  assign n18526 = n15930 & ~n18525 ;
  assign n18527 = n9643 ^ n2481 ^ 1'b0 ;
  assign n18528 = n8071 | n17471 ;
  assign n18529 = n5431 & ~n5701 ;
  assign n18530 = n18529 ^ n2007 ^ 1'b0 ;
  assign n18531 = n9523 ^ n3166 ^ n1131 ;
  assign n18532 = n10896 & ~n18531 ;
  assign n18533 = n18532 ^ n10843 ^ 1'b0 ;
  assign n18534 = n9253 ^ n7379 ^ n1469 ;
  assign n18535 = n9491 & n18534 ;
  assign n18536 = n18535 ^ n9927 ^ 1'b0 ;
  assign n18537 = n14849 ^ n14522 ^ 1'b0 ;
  assign n18538 = ( n2834 & ~n5114 ) | ( n2834 & n5749 ) | ( ~n5114 & n5749 ) ;
  assign n18539 = n11909 & n18538 ;
  assign n18540 = n16447 ^ n2079 ^ n307 ;
  assign n18541 = n8908 ^ n8139 ^ n6140 ;
  assign n18542 = ( n458 & n2308 ) | ( n458 & n9909 ) | ( n2308 & n9909 ) ;
  assign n18543 = n699 & n18542 ;
  assign n18544 = n6566 & n18543 ;
  assign n18545 = ~n540 & n6558 ;
  assign n18546 = n1425 & n18545 ;
  assign n18547 = ( n3790 & ~n13305 ) | ( n3790 & n16841 ) | ( ~n13305 & n16841 ) ;
  assign n18548 = n10730 & n18547 ;
  assign n18549 = n16546 ^ n6893 ^ n5238 ;
  assign n18550 = n18549 ^ n721 ^ 1'b0 ;
  assign n18551 = ~n16962 & n18550 ;
  assign n18552 = n5165 & ~n7171 ;
  assign n18553 = n18552 ^ n5347 ^ 1'b0 ;
  assign n18554 = n18553 ^ n9857 ^ n7468 ;
  assign n18555 = n1484 | n3817 ;
  assign n18556 = n3817 & ~n18555 ;
  assign n18557 = n5867 & ~n13201 ;
  assign n18558 = n13201 & n18557 ;
  assign n18559 = n199 & ~n18558 ;
  assign n18560 = n18556 & n18559 ;
  assign n18561 = n10888 | n12719 ;
  assign n18562 = n18561 ^ n558 ^ 1'b0 ;
  assign n18563 = n15381 ^ n3975 ^ 1'b0 ;
  assign n18564 = n18563 ^ n12576 ^ n12322 ;
  assign n18565 = ( n1079 & n2958 ) | ( n1079 & ~n15190 ) | ( n2958 & ~n15190 ) ;
  assign n18566 = ( n4101 & ~n15086 ) | ( n4101 & n18565 ) | ( ~n15086 & n18565 ) ;
  assign n18568 = n2932 & n14664 ;
  assign n18569 = n18568 ^ n10946 ^ 1'b0 ;
  assign n18567 = n2177 & n18506 ;
  assign n18570 = n18569 ^ n18567 ^ n11314 ;
  assign n18571 = n18570 ^ n17211 ^ n11999 ;
  assign n18572 = n13562 ^ n12971 ^ 1'b0 ;
  assign n18573 = n12297 ^ n2562 ^ 1'b0 ;
  assign n18574 = n18573 ^ n18512 ^ 1'b0 ;
  assign n18575 = n16941 ^ n14081 ^ 1'b0 ;
  assign n18576 = n1754 | n18575 ;
  assign n18577 = n15408 & n16840 ;
  assign n18578 = ( ~n12330 & n16005 ) | ( ~n12330 & n16277 ) | ( n16005 & n16277 ) ;
  assign n18579 = n2011 & n14702 ;
  assign n18580 = n241 | n15395 ;
  assign n18581 = n3348 & n16748 ;
  assign n18585 = n1056 & n5082 ;
  assign n18582 = n8827 ^ n2798 ^ n1986 ;
  assign n18583 = n18582 ^ n3715 ^ n1213 ;
  assign n18584 = ( n763 & n16589 ) | ( n763 & n18583 ) | ( n16589 & n18583 ) ;
  assign n18586 = n18585 ^ n18584 ^ n13333 ;
  assign n18588 = n1302 | n8104 ;
  assign n18589 = n8577 | n18588 ;
  assign n18587 = ~n7968 & n10863 ;
  assign n18590 = n18589 ^ n18587 ^ 1'b0 ;
  assign n18591 = n6519 ^ n2507 ^ 1'b0 ;
  assign n18592 = ~n17677 & n18591 ;
  assign n18593 = x13 & n9902 ;
  assign n18594 = n7768 & n18593 ;
  assign n18595 = ( ~n11542 & n11915 ) | ( ~n11542 & n13416 ) | ( n11915 & n13416 ) ;
  assign n18596 = n12926 ^ n1204 ^ 1'b0 ;
  assign n18597 = ~n479 & n18596 ;
  assign n18598 = n18597 ^ n18212 ^ 1'b0 ;
  assign n18599 = n3218 | n4974 ;
  assign n18600 = n14643 & ~n18027 ;
  assign n18601 = n6249 & n18600 ;
  assign n18602 = n18599 & ~n18601 ;
  assign n18604 = ( ~n6800 & n7563 ) | ( ~n6800 & n10432 ) | ( n7563 & n10432 ) ;
  assign n18605 = n11369 ^ n8382 ^ n5878 ;
  assign n18606 = n2081 & ~n6954 ;
  assign n18607 = n7224 & n18606 ;
  assign n18608 = ( ~n18604 & n18605 ) | ( ~n18604 & n18607 ) | ( n18605 & n18607 ) ;
  assign n18603 = n7513 ^ n6773 ^ n4820 ;
  assign n18609 = n18608 ^ n18603 ^ 1'b0 ;
  assign n18610 = n16462 ^ n10049 ^ 1'b0 ;
  assign n18611 = ~n3917 & n18610 ;
  assign n18612 = n10731 & ~n11668 ;
  assign n18613 = n2524 & n18612 ;
  assign n18614 = n18143 ^ n5216 ^ 1'b0 ;
  assign n18615 = n9478 ^ n2893 ^ 1'b0 ;
  assign n18616 = ( n7572 & n10658 ) | ( n7572 & n12266 ) | ( n10658 & n12266 ) ;
  assign n18617 = n10616 | n18616 ;
  assign n18618 = n18615 | n18617 ;
  assign n18619 = ( n2919 & n3247 ) | ( n2919 & n5962 ) | ( n3247 & n5962 ) ;
  assign n18620 = n4984 | n18619 ;
  assign n18621 = n310 & ~n9363 ;
  assign n18622 = n18621 ^ n2113 ^ 1'b0 ;
  assign n18623 = n695 & n6689 ;
  assign n18624 = n18623 ^ n1829 ^ 1'b0 ;
  assign n18625 = n18624 ^ n3869 ^ 1'b0 ;
  assign n18626 = n12677 ^ n4336 ^ 1'b0 ;
  assign n18627 = ( ~n208 & n4653 ) | ( ~n208 & n5259 ) | ( n4653 & n5259 ) ;
  assign n18628 = n18627 ^ n8618 ^ 1'b0 ;
  assign n18629 = n11427 & n18628 ;
  assign n18630 = n16991 ^ n1833 ^ 1'b0 ;
  assign n18631 = n7492 & ~n18630 ;
  assign n18632 = n5179 & ~n18631 ;
  assign n18633 = n7842 | n10177 ;
  assign n18634 = n7232 ^ n2305 ^ n1601 ;
  assign n18635 = n18633 & n18634 ;
  assign n18636 = n4877 & ~n5432 ;
  assign n18637 = ~n2654 & n18636 ;
  assign n18638 = n1586 & ~n3688 ;
  assign n18639 = n8564 ^ n6368 ^ 1'b0 ;
  assign n18640 = n18639 ^ n2728 ^ 1'b0 ;
  assign n18641 = ( n18637 & n18638 ) | ( n18637 & ~n18640 ) | ( n18638 & ~n18640 ) ;
  assign n18642 = n1116 | n13047 ;
  assign n18643 = n2003 ^ n1966 ^ 1'b0 ;
  assign n18644 = n1057 & ~n4986 ;
  assign n18645 = n1870 | n18644 ;
  assign n18646 = n18645 ^ n6288 ^ n3838 ;
  assign n18647 = n4808 ^ n1292 ^ 1'b0 ;
  assign n18648 = ~n17446 & n18647 ;
  assign n18649 = n14835 ^ n8341 ^ n7984 ;
  assign n18650 = n4718 & ~n18649 ;
  assign n18651 = ( ~n15706 & n18648 ) | ( ~n15706 & n18650 ) | ( n18648 & n18650 ) ;
  assign n18652 = n11572 | n17967 ;
  assign n18653 = n18651 | n18652 ;
  assign n18654 = n12447 | n18212 ;
  assign n18655 = n5218 | n18654 ;
  assign n18656 = n508 & ~n18655 ;
  assign n18657 = n13033 & n17943 ;
  assign n18659 = ( ~n2978 & n8192 ) | ( ~n2978 & n14833 ) | ( n8192 & n14833 ) ;
  assign n18660 = n18659 ^ n6299 ^ 1'b0 ;
  assign n18661 = n18660 ^ n17442 ^ 1'b0 ;
  assign n18662 = ~n2891 & n18661 ;
  assign n18658 = n9179 & n11637 ;
  assign n18663 = n18662 ^ n18658 ^ 1'b0 ;
  assign n18667 = n2200 ^ n1498 ^ 1'b0 ;
  assign n18668 = n4179 & ~n18667 ;
  assign n18669 = n12928 & ~n18668 ;
  assign n18670 = ( ~n14044 & n14657 ) | ( ~n14044 & n18669 ) | ( n14657 & n18669 ) ;
  assign n18664 = n3055 ^ n320 ^ 1'b0 ;
  assign n18665 = n12359 & n18664 ;
  assign n18666 = n8380 | n18665 ;
  assign n18671 = n18670 ^ n18666 ^ 1'b0 ;
  assign n18672 = n5654 & ~n10955 ;
  assign n18673 = ~n17000 & n18672 ;
  assign n18674 = n12621 & n18673 ;
  assign n18675 = x2 & n18299 ;
  assign n18676 = n5990 ^ n3380 ^ n976 ;
  assign n18677 = ~n562 & n3796 ;
  assign n18678 = n18677 ^ n1431 ^ 1'b0 ;
  assign n18679 = n3686 & ~n18678 ;
  assign n18680 = ( ~n8293 & n18676 ) | ( ~n8293 & n18679 ) | ( n18676 & n18679 ) ;
  assign n18681 = n7270 ^ n4042 ^ 1'b0 ;
  assign n18682 = ~n9477 & n18681 ;
  assign n18683 = ( n3374 & n4999 ) | ( n3374 & ~n7591 ) | ( n4999 & ~n7591 ) ;
  assign n18684 = n18682 & ~n18683 ;
  assign n18685 = n8293 ^ n3118 ^ n2156 ;
  assign n18688 = n6862 & ~n14726 ;
  assign n18686 = n7395 & ~n7774 ;
  assign n18687 = n10443 & n18686 ;
  assign n18689 = n18688 ^ n18687 ^ 1'b0 ;
  assign n18690 = ~n18685 & n18689 ;
  assign n18691 = n826 | n13079 ;
  assign n18692 = n10469 & ~n18691 ;
  assign n18693 = ( n2958 & n13848 ) | ( n2958 & n18692 ) | ( n13848 & n18692 ) ;
  assign n18694 = n18693 ^ n3529 ^ 1'b0 ;
  assign n18695 = n1514 | n18694 ;
  assign n18696 = n10917 ^ n1364 ^ 1'b0 ;
  assign n18697 = n18696 ^ n11930 ^ 1'b0 ;
  assign n18698 = n6785 & n13422 ;
  assign n18699 = n18698 ^ n3072 ^ 1'b0 ;
  assign n18700 = n18699 ^ n12853 ^ n10721 ;
  assign n18701 = n11841 ^ n5108 ^ n4795 ;
  assign n18702 = n15872 | n18701 ;
  assign n18703 = n6079 ^ n1728 ^ 1'b0 ;
  assign n18704 = n541 & n18703 ;
  assign n18705 = ~n7611 & n18704 ;
  assign n18706 = n12331 ^ n11570 ^ n7043 ;
  assign n18707 = ( n1213 & n16816 ) | ( n1213 & n18706 ) | ( n16816 & n18706 ) ;
  assign n18711 = n2522 | n5904 ;
  assign n18712 = n18711 ^ n4642 ^ 1'b0 ;
  assign n18713 = n18712 ^ n5470 ^ 1'b0 ;
  assign n18714 = n15022 & n18713 ;
  assign n18708 = n6797 | n18639 ;
  assign n18709 = n3592 | n18708 ;
  assign n18710 = n18709 ^ n12457 ^ 1'b0 ;
  assign n18715 = n18714 ^ n18710 ^ n15654 ;
  assign n18716 = n1883 ^ n569 ^ 1'b0 ;
  assign n18717 = n3804 ^ n339 ^ 1'b0 ;
  assign n18718 = ~n1484 & n18717 ;
  assign n18719 = n18718 ^ n14650 ^ 1'b0 ;
  assign n18720 = n18719 ^ n5623 ^ 1'b0 ;
  assign n18721 = n18716 & ~n18720 ;
  assign n18722 = n7396 ^ n364 ^ 1'b0 ;
  assign n18723 = n16902 ^ n12058 ^ 1'b0 ;
  assign n18724 = n18723 ^ n5940 ^ 1'b0 ;
  assign n18725 = n18724 ^ n7682 ^ n3136 ;
  assign n18726 = n2160 ^ n319 ^ 1'b0 ;
  assign n18727 = n4259 | n11362 ;
  assign n18728 = n18727 ^ n6123 ^ 1'b0 ;
  assign n18729 = n18728 ^ n15096 ^ n3388 ;
  assign n18730 = n7845 & n18729 ;
  assign n18731 = n18730 ^ n10450 ^ 1'b0 ;
  assign n18732 = ( n1466 & ~n2500 ) | ( n1466 & n7726 ) | ( ~n2500 & n7726 ) ;
  assign n18733 = ~n12511 & n18732 ;
  assign n18734 = n18733 ^ n7229 ^ 1'b0 ;
  assign n18735 = n3950 ^ n3612 ^ 1'b0 ;
  assign n18736 = n588 & ~n18735 ;
  assign n18737 = n18736 ^ n15397 ^ x119 ;
  assign n18738 = n5328 & ~n9364 ;
  assign n18739 = n18738 ^ n17120 ^ n3533 ;
  assign n18740 = ( n7112 & n9678 ) | ( n7112 & ~n18739 ) | ( n9678 & ~n18739 ) ;
  assign n18741 = n3857 ^ n1860 ^ n597 ;
  assign n18742 = n4772 | n18741 ;
  assign n18743 = n8099 & ~n8183 ;
  assign n18744 = n17176 & n18743 ;
  assign n18746 = n3554 | n4775 ;
  assign n18747 = x93 | n18746 ;
  assign n18745 = n18438 ^ n13858 ^ 1'b0 ;
  assign n18748 = n18747 ^ n18745 ^ n6756 ;
  assign n18749 = ( ~n3986 & n10785 ) | ( ~n3986 & n18748 ) | ( n10785 & n18748 ) ;
  assign n18750 = ( n18742 & n18744 ) | ( n18742 & n18749 ) | ( n18744 & n18749 ) ;
  assign n18751 = n17100 ^ n8934 ^ n2100 ;
  assign n18752 = ~n3247 & n18751 ;
  assign n18753 = n12323 & n18752 ;
  assign n18754 = n18753 ^ n4176 ^ n1274 ;
  assign n18756 = n8785 ^ n1942 ^ 1'b0 ;
  assign n18757 = n18756 ^ n5371 ^ n4725 ;
  assign n18755 = n1927 | n10140 ;
  assign n18758 = n18757 ^ n18755 ^ n11605 ;
  assign n18759 = ( ~n12563 & n12970 ) | ( ~n12563 & n13591 ) | ( n12970 & n13591 ) ;
  assign n18760 = n16477 ^ n12345 ^ n3374 ;
  assign n18761 = n12347 ^ n1949 ^ 1'b0 ;
  assign n18762 = n18761 ^ n15773 ^ 1'b0 ;
  assign n18763 = n5962 | n18762 ;
  assign n18764 = n243 | n18763 ;
  assign n18765 = n4875 | n18764 ;
  assign n18766 = n15696 ^ n6231 ^ n2110 ;
  assign n18767 = ( n8660 & ~n8880 ) | ( n8660 & n17184 ) | ( ~n8880 & n17184 ) ;
  assign n18768 = n9419 & ~n9999 ;
  assign n18769 = n3540 & n18768 ;
  assign n18770 = ( n1600 & ~n2360 ) | ( n1600 & n18769 ) | ( ~n2360 & n18769 ) ;
  assign n18771 = ( n9279 & n11694 ) | ( n9279 & n18770 ) | ( n11694 & n18770 ) ;
  assign n18772 = n15074 ^ n10704 ^ n3948 ;
  assign n18773 = ~n5163 & n5209 ;
  assign n18774 = n18773 ^ n2038 ^ 1'b0 ;
  assign n18775 = n10951 ^ n8229 ^ n2303 ;
  assign n18776 = ( n344 & ~n1135 ) | ( n344 & n3188 ) | ( ~n1135 & n3188 ) ;
  assign n18777 = ( n12392 & n12812 ) | ( n12392 & ~n18776 ) | ( n12812 & ~n18776 ) ;
  assign n18783 = n14771 ^ n5097 ^ 1'b0 ;
  assign n18784 = n11691 & ~n18783 ;
  assign n18785 = ~n3337 & n10108 ;
  assign n18786 = ~n18784 & n18785 ;
  assign n18787 = n11647 ^ n714 ^ 1'b0 ;
  assign n18788 = n18786 | n18787 ;
  assign n18781 = n7190 & ~n9691 ;
  assign n18782 = n18781 ^ n12515 ^ 1'b0 ;
  assign n18778 = n7614 ^ n2900 ^ 1'b0 ;
  assign n18779 = ~n6858 & n18778 ;
  assign n18780 = ( n9867 & n12328 ) | ( n9867 & n18779 ) | ( n12328 & n18779 ) ;
  assign n18789 = n18788 ^ n18782 ^ n18780 ;
  assign n18790 = ~n6918 & n11357 ;
  assign n18791 = n18790 ^ n14172 ^ 1'b0 ;
  assign n18792 = n18791 ^ n14619 ^ n11578 ;
  assign n18795 = ( n1855 & n8580 ) | ( n1855 & n9123 ) | ( n8580 & n9123 ) ;
  assign n18793 = ~n3162 & n15992 ;
  assign n18794 = n18793 ^ n692 ^ 1'b0 ;
  assign n18796 = n18795 ^ n18794 ^ n3876 ;
  assign n18797 = n2792 & n4999 ;
  assign n18798 = n4567 & n18797 ;
  assign n18799 = n18798 ^ n1221 ^ 1'b0 ;
  assign n18800 = n7921 | n18799 ;
  assign n18801 = ~n5184 & n13836 ;
  assign n18802 = n18801 ^ n5077 ^ 1'b0 ;
  assign n18803 = n7869 | n18456 ;
  assign n18804 = n3923 ^ n1402 ^ 1'b0 ;
  assign n18805 = n8447 & ~n18804 ;
  assign n18806 = ~n15651 & n18805 ;
  assign n18807 = ~n10248 & n18806 ;
  assign n18808 = ( n5028 & ~n5430 ) | ( n5028 & n7378 ) | ( ~n5430 & n7378 ) ;
  assign n18811 = n3698 & n16757 ;
  assign n18809 = n12499 & ~n14773 ;
  assign n18810 = n18809 ^ n9857 ^ 1'b0 ;
  assign n18812 = n18811 ^ n18810 ^ n1590 ;
  assign n18813 = ( ~n9019 & n9220 ) | ( ~n9019 & n18812 ) | ( n9220 & n18812 ) ;
  assign n18815 = n5996 ^ n4874 ^ 1'b0 ;
  assign n18814 = n260 & ~n11566 ;
  assign n18816 = n18815 ^ n18814 ^ 1'b0 ;
  assign n18821 = n539 & ~n6272 ;
  assign n18817 = n5889 ^ n1758 ^ 1'b0 ;
  assign n18818 = ~n5825 & n9451 ;
  assign n18819 = n18818 ^ n13036 ^ 1'b0 ;
  assign n18820 = ~n18817 & n18819 ;
  assign n18822 = n18821 ^ n18820 ^ 1'b0 ;
  assign n18823 = n16526 ^ n8142 ^ 1'b0 ;
  assign n18824 = n6914 | n18823 ;
  assign n18825 = n2496 | n17477 ;
  assign n18826 = n18824 & ~n18825 ;
  assign n18827 = n4745 ^ n2350 ^ 1'b0 ;
  assign n18828 = ( n7195 & n9348 ) | ( n7195 & n16010 ) | ( n9348 & n16010 ) ;
  assign n18829 = ( n3561 & ~n18827 ) | ( n3561 & n18828 ) | ( ~n18827 & n18828 ) ;
  assign n18830 = n18829 ^ n15859 ^ n1799 ;
  assign n18831 = n10892 ^ n1771 ^ 1'b0 ;
  assign n18832 = n3149 & ~n18831 ;
  assign n18833 = ( n256 & n582 ) | ( n256 & ~n18832 ) | ( n582 & ~n18832 ) ;
  assign n18834 = ~n4098 & n11437 ;
  assign n18835 = n7622 | n18834 ;
  assign n18836 = n2475 & ~n18835 ;
  assign n18838 = n14812 ^ n8423 ^ n7116 ;
  assign n18839 = n18838 ^ n4208 ^ n1050 ;
  assign n18837 = ~n16968 & n17926 ;
  assign n18840 = n18839 ^ n18837 ^ 1'b0 ;
  assign n18841 = n12256 ^ n4588 ^ n4123 ;
  assign n18842 = ( ~n6627 & n11776 ) | ( ~n6627 & n18841 ) | ( n11776 & n18841 ) ;
  assign n18843 = x10 | n5527 ;
  assign n18844 = n18843 ^ n4647 ^ 1'b0 ;
  assign n18845 = n11804 ^ n8062 ^ 1'b0 ;
  assign n18846 = ~n1749 & n18845 ;
  assign n18847 = ( n4424 & n18844 ) | ( n4424 & ~n18846 ) | ( n18844 & ~n18846 ) ;
  assign n18848 = n11188 ^ n7411 ^ 1'b0 ;
  assign n18849 = ~n296 & n18848 ;
  assign n18850 = n18849 ^ n3419 ^ 1'b0 ;
  assign n18851 = n13646 | n18850 ;
  assign n18852 = ( ~n275 & n3780 ) | ( ~n275 & n18282 ) | ( n3780 & n18282 ) ;
  assign n18853 = n18852 ^ n1123 ^ 1'b0 ;
  assign n18857 = n635 ^ n454 ^ 1'b0 ;
  assign n18854 = n9761 ^ n1114 ^ 1'b0 ;
  assign n18855 = ~n17159 & n18854 ;
  assign n18856 = ~n7031 & n18855 ;
  assign n18858 = n18857 ^ n18856 ^ 1'b0 ;
  assign n18859 = ~n6864 & n10327 ;
  assign n18860 = n18859 ^ n7532 ^ 1'b0 ;
  assign n18861 = ~n4266 & n18860 ;
  assign n18862 = ( ~n1002 & n10024 ) | ( ~n1002 & n18861 ) | ( n10024 & n18861 ) ;
  assign n18863 = n18862 ^ n7375 ^ 1'b0 ;
  assign n18864 = n11120 ^ n7117 ^ n6504 ;
  assign n18865 = n3441 | n18864 ;
  assign n18866 = n13130 ^ n6740 ^ 1'b0 ;
  assign n18867 = n3346 & ~n18866 ;
  assign n18868 = n17355 ^ n2083 ^ 1'b0 ;
  assign n18869 = ~n1695 & n18868 ;
  assign n18870 = n11187 ^ n3574 ^ n2386 ;
  assign n18871 = ( n7284 & n9850 ) | ( n7284 & ~n13160 ) | ( n9850 & ~n13160 ) ;
  assign n18872 = ( n6151 & n10128 ) | ( n6151 & ~n17324 ) | ( n10128 & ~n17324 ) ;
  assign n18874 = ( ~n972 & n3617 ) | ( ~n972 & n5940 ) | ( n3617 & n5940 ) ;
  assign n18875 = ( n1363 & ~n14103 ) | ( n1363 & n18874 ) | ( ~n14103 & n18874 ) ;
  assign n18873 = n1383 & ~n18696 ;
  assign n18876 = n18875 ^ n18873 ^ 1'b0 ;
  assign n18877 = n10477 | n18876 ;
  assign n18878 = n18877 ^ n3333 ^ 1'b0 ;
  assign n18879 = n781 & n1713 ;
  assign n18880 = n18879 ^ n12735 ^ 1'b0 ;
  assign n18887 = ( n1456 & n2090 ) | ( n1456 & ~n4198 ) | ( n2090 & ~n4198 ) ;
  assign n18886 = n4976 & ~n7033 ;
  assign n18888 = n18887 ^ n18886 ^ 1'b0 ;
  assign n18881 = n4038 & n13232 ;
  assign n18882 = n11124 & n18881 ;
  assign n18883 = n18882 ^ n9757 ^ 1'b0 ;
  assign n18884 = n2211 | n18883 ;
  assign n18885 = n12201 | n18884 ;
  assign n18889 = n18888 ^ n18885 ^ 1'b0 ;
  assign n18890 = n7349 | n12043 ;
  assign n18891 = n12576 ^ n7850 ^ n2114 ;
  assign n18892 = n18891 ^ n9199 ^ 1'b0 ;
  assign n18893 = n1881 | n10911 ;
  assign n18894 = ( n5507 & n6498 ) | ( n5507 & n16266 ) | ( n6498 & n16266 ) ;
  assign n18895 = n18894 ^ n11519 ^ n3297 ;
  assign n18896 = n18895 ^ n11944 ^ 1'b0 ;
  assign n18897 = n9471 & ~n18896 ;
  assign n18900 = n3297 ^ n2254 ^ 1'b0 ;
  assign n18901 = n18732 & n18900 ;
  assign n18898 = n13908 ^ n12825 ^ 1'b0 ;
  assign n18899 = n11004 & ~n18898 ;
  assign n18902 = n18901 ^ n18899 ^ 1'b0 ;
  assign n18903 = n8355 & ~n18902 ;
  assign n18904 = n11128 ^ n6299 ^ n487 ;
  assign n18905 = n7600 ^ n2971 ^ 1'b0 ;
  assign n18906 = ~n18904 & n18905 ;
  assign n18907 = n3552 & ~n18906 ;
  assign n18908 = n2460 & n18907 ;
  assign n18909 = n9823 ^ n8019 ^ 1'b0 ;
  assign n18910 = n325 | n18909 ;
  assign n18911 = n11358 ^ n6271 ^ n3056 ;
  assign n18912 = ( ~n1533 & n1605 ) | ( ~n1533 & n2744 ) | ( n1605 & n2744 ) ;
  assign n18913 = ~n556 & n3422 ;
  assign n18914 = n18913 ^ n8351 ^ n5999 ;
  assign n18915 = n5049 & ~n10917 ;
  assign n18916 = n18914 & n18915 ;
  assign n18917 = ( n17848 & n18912 ) | ( n17848 & n18916 ) | ( n18912 & n18916 ) ;
  assign n18918 = n18917 ^ n11192 ^ n6448 ;
  assign n18919 = ~n10590 & n13370 ;
  assign n18920 = n13988 | n18919 ;
  assign n18921 = n18920 ^ n9375 ^ 1'b0 ;
  assign n18922 = ~n3812 & n5805 ;
  assign n18923 = n7612 ^ n5876 ^ 1'b0 ;
  assign n18924 = n18922 & n18923 ;
  assign n18927 = ( ~n1327 & n9043 ) | ( ~n1327 & n10913 ) | ( n9043 & n10913 ) ;
  assign n18925 = n13781 ^ n955 ^ 1'b0 ;
  assign n18926 = n2943 | n18925 ;
  assign n18928 = n18927 ^ n18926 ^ n13344 ;
  assign n18929 = ( n3037 & ~n6357 ) | ( n3037 & n12540 ) | ( ~n6357 & n12540 ) ;
  assign n18930 = n1292 & n2610 ;
  assign n18931 = n18929 & n18930 ;
  assign n18932 = ~n9841 & n18931 ;
  assign n18933 = n9594 | n15341 ;
  assign n18934 = n390 | n18933 ;
  assign n18935 = ( ~n1046 & n1578 ) | ( ~n1046 & n9224 ) | ( n1578 & n9224 ) ;
  assign n18936 = n1940 | n18935 ;
  assign n18937 = n18936 ^ n12243 ^ 1'b0 ;
  assign n18939 = n755 & ~n3696 ;
  assign n18940 = ~n5876 & n18939 ;
  assign n18938 = n13211 & n16114 ;
  assign n18941 = n18940 ^ n18938 ^ 1'b0 ;
  assign n18942 = ( n8271 & n13796 ) | ( n8271 & n18941 ) | ( n13796 & n18941 ) ;
  assign n18943 = n5430 | n6002 ;
  assign n18944 = n14743 ^ n7594 ^ 1'b0 ;
  assign n18949 = n880 ^ x59 ^ 1'b0 ;
  assign n18950 = n1058 & ~n18949 ;
  assign n18951 = ( n483 & n6449 ) | ( n483 & n18950 ) | ( n6449 & n18950 ) ;
  assign n18952 = n1764 & n18951 ;
  assign n18953 = n10506 & n18952 ;
  assign n18945 = n3376 & ~n10860 ;
  assign n18946 = n18945 ^ n3134 ^ 1'b0 ;
  assign n18947 = ~n13301 & n18946 ;
  assign n18948 = ~n11441 & n18947 ;
  assign n18954 = n18953 ^ n18948 ^ 1'b0 ;
  assign n18955 = n12208 ^ n9699 ^ 1'b0 ;
  assign n18956 = ~n3706 & n14721 ;
  assign n18957 = n6146 & n18956 ;
  assign n18958 = ( n5893 & ~n14506 ) | ( n5893 & n18957 ) | ( ~n14506 & n18957 ) ;
  assign n18959 = ~n5907 & n7788 ;
  assign n18960 = n18959 ^ n11433 ^ n4650 ;
  assign n18962 = n4602 | n13673 ;
  assign n18963 = n18962 ^ n6301 ^ 1'b0 ;
  assign n18961 = ( ~x102 & n2498 ) | ( ~x102 & n7848 ) | ( n2498 & n7848 ) ;
  assign n18964 = n18963 ^ n18961 ^ 1'b0 ;
  assign n18965 = n3573 & n4365 ;
  assign n18966 = n18965 ^ n4506 ^ 1'b0 ;
  assign n18967 = ( ~n3547 & n11769 ) | ( ~n3547 & n18966 ) | ( n11769 & n18966 ) ;
  assign n18968 = n1445 ^ n1176 ^ 1'b0 ;
  assign n18969 = n18968 ^ n12772 ^ n11644 ;
  assign n18970 = ~n3296 & n18969 ;
  assign n18971 = n7018 ^ n6330 ^ 1'b0 ;
  assign n18972 = n18971 ^ n12038 ^ n5076 ;
  assign n18973 = ( ~n7800 & n14612 ) | ( ~n7800 & n18972 ) | ( n14612 & n18972 ) ;
  assign n18974 = ( n527 & ~n2072 ) | ( n527 & n11808 ) | ( ~n2072 & n11808 ) ;
  assign n18975 = n18974 ^ n1860 ^ 1'b0 ;
  assign n18976 = n2701 & ~n12618 ;
  assign n18977 = ~n18975 & n18976 ;
  assign n18978 = n10634 ^ n6989 ^ 1'b0 ;
  assign n18979 = n2179 & n11119 ;
  assign n18980 = ~n18978 & n18979 ;
  assign n18982 = n17406 ^ n5272 ^ 1'b0 ;
  assign n18981 = n999 & ~n1333 ;
  assign n18983 = n18982 ^ n18981 ^ 1'b0 ;
  assign n18984 = n13675 | n14028 ;
  assign n18985 = n18984 ^ n10452 ^ 1'b0 ;
  assign n18986 = n11196 ^ n6965 ^ n1521 ;
  assign n18987 = n17020 ^ n16473 ^ 1'b0 ;
  assign n18988 = n14976 | n18987 ;
  assign n18989 = ~n5633 & n10182 ;
  assign n18990 = n18989 ^ n9639 ^ 1'b0 ;
  assign n18991 = n18990 ^ n6981 ^ n6951 ;
  assign n18992 = n16377 ^ n3974 ^ n1084 ;
  assign n18993 = n6624 ^ n1975 ^ 1'b0 ;
  assign n18994 = n394 & ~n18993 ;
  assign n18995 = n7780 | n11678 ;
  assign n18996 = ( n6700 & ~n9898 ) | ( n6700 & n15206 ) | ( ~n9898 & n15206 ) ;
  assign n18997 = ( n1364 & n5632 ) | ( n1364 & n8229 ) | ( n5632 & n8229 ) ;
  assign n18998 = n18997 ^ n5586 ^ 1'b0 ;
  assign n18999 = n18998 ^ n12764 ^ 1'b0 ;
  assign n19000 = n18999 ^ n16618 ^ n8910 ;
  assign n19001 = n3566 | n12948 ;
  assign n19002 = n19001 ^ n4234 ^ 1'b0 ;
  assign n19003 = n4915 & n19002 ;
  assign n19004 = n7945 ^ n141 ^ x113 ;
  assign n19005 = n4415 & n19004 ;
  assign n19006 = ~n7966 & n19005 ;
  assign n19007 = n1212 | n4131 ;
  assign n19008 = n2742 & ~n19007 ;
  assign n19009 = ( ~n8446 & n14835 ) | ( ~n8446 & n19008 ) | ( n14835 & n19008 ) ;
  assign n19010 = n2723 & n14066 ;
  assign n19011 = n9954 ^ n770 ^ 1'b0 ;
  assign n19012 = n6639 | n19011 ;
  assign n19013 = ( n1019 & n3098 ) | ( n1019 & ~n19012 ) | ( n3098 & ~n19012 ) ;
  assign n19014 = n19013 ^ n10991 ^ n4402 ;
  assign n19015 = n19014 ^ n10144 ^ 1'b0 ;
  assign n19016 = n10687 ^ n1170 ^ 1'b0 ;
  assign n19017 = n13146 ^ n1605 ^ 1'b0 ;
  assign n19018 = n19017 ^ n5316 ^ 1'b0 ;
  assign n19019 = n3864 & ~n19018 ;
  assign n19020 = n19016 & n19019 ;
  assign n19021 = n1236 & n6089 ;
  assign n19022 = ( n8182 & ~n9007 ) | ( n8182 & n16183 ) | ( ~n9007 & n16183 ) ;
  assign n19023 = ( n14492 & n19021 ) | ( n14492 & n19022 ) | ( n19021 & n19022 ) ;
  assign n19024 = n8868 & n19023 ;
  assign n19025 = n19020 & n19024 ;
  assign n19026 = n5436 ^ n1559 ^ 1'b0 ;
  assign n19027 = n11987 & ~n19026 ;
  assign n19028 = n8605 ^ n7673 ^ 1'b0 ;
  assign n19029 = n19028 ^ n13862 ^ 1'b0 ;
  assign n19030 = n4306 & n7499 ;
  assign n19031 = n19030 ^ n13973 ^ 1'b0 ;
  assign n19032 = n3375 & ~n19031 ;
  assign n19033 = ( ~n1973 & n8572 ) | ( ~n1973 & n19032 ) | ( n8572 & n19032 ) ;
  assign n19034 = x118 & n9115 ;
  assign n19035 = n19034 ^ n9198 ^ 1'b0 ;
  assign n19036 = n9556 ^ n7691 ^ n2539 ;
  assign n19037 = ~n7918 & n19036 ;
  assign n19038 = n18626 ^ n9563 ^ 1'b0 ;
  assign n19039 = n7325 | n8843 ;
  assign n19040 = n19039 ^ n452 ^ 1'b0 ;
  assign n19041 = ( n1998 & n2663 ) | ( n1998 & n16154 ) | ( n2663 & n16154 ) ;
  assign n19042 = n15996 & n19041 ;
  assign n19043 = n19042 ^ n9105 ^ n2296 ;
  assign n19044 = n5537 | n18054 ;
  assign n19045 = n7007 & n8393 ;
  assign n19046 = n12092 ^ n11377 ^ 1'b0 ;
  assign n19047 = n19046 ^ n4978 ^ 1'b0 ;
  assign n19048 = n4957 & n8921 ;
  assign n19049 = n19047 & n19048 ;
  assign n19050 = n19049 ^ n17102 ^ n343 ;
  assign n19052 = ( n11349 & n12930 ) | ( n11349 & n16241 ) | ( n12930 & n16241 ) ;
  assign n19051 = n10472 & n16246 ;
  assign n19053 = n19052 ^ n19051 ^ 1'b0 ;
  assign n19054 = n9061 | n9359 ;
  assign n19055 = n8473 | n19054 ;
  assign n19056 = ~n1914 & n5464 ;
  assign n19057 = ~n908 & n19056 ;
  assign n19061 = ( n6473 & n7314 ) | ( n6473 & ~n8471 ) | ( n7314 & ~n8471 ) ;
  assign n19058 = n6284 ^ n3897 ^ 1'b0 ;
  assign n19059 = ~n8714 & n19058 ;
  assign n19060 = n19059 ^ n18238 ^ 1'b0 ;
  assign n19062 = n19061 ^ n19060 ^ n11671 ;
  assign n19064 = n6711 ^ x107 ^ 1'b0 ;
  assign n19063 = n173 & n6773 ;
  assign n19065 = n19064 ^ n19063 ^ 1'b0 ;
  assign n19066 = ~n4539 & n19065 ;
  assign n19067 = n19066 ^ n10858 ^ n441 ;
  assign n19068 = n12727 ^ n8896 ^ 1'b0 ;
  assign n19069 = n15014 ^ n10098 ^ n1998 ;
  assign n19070 = ~n7219 & n19069 ;
  assign n19071 = n9785 ^ n6607 ^ 1'b0 ;
  assign n19077 = n270 & ~n3406 ;
  assign n19078 = ~n5704 & n19077 ;
  assign n19079 = n19078 ^ n2955 ^ 1'b0 ;
  assign n19080 = n5418 & n19079 ;
  assign n19076 = n11145 ^ n10425 ^ n7783 ;
  assign n19073 = ~n9942 & n12030 ;
  assign n19074 = n19073 ^ n8545 ^ 1'b0 ;
  assign n19072 = n16888 ^ n9896 ^ n9574 ;
  assign n19075 = n19074 ^ n19072 ^ 1'b0 ;
  assign n19081 = n19080 ^ n19076 ^ n19075 ;
  assign n19082 = ~n7933 & n17495 ;
  assign n19083 = n10116 & n19082 ;
  assign n19084 = ( ~n4655 & n5665 ) | ( ~n4655 & n7726 ) | ( n5665 & n7726 ) ;
  assign n19085 = n19084 ^ n13729 ^ n12735 ;
  assign n19086 = x69 | n6895 ;
  assign n19087 = n19086 ^ n16350 ^ n10341 ;
  assign n19088 = n18742 ^ n2263 ^ 1'b0 ;
  assign n19089 = ( n404 & n10048 ) | ( n404 & n19088 ) | ( n10048 & n19088 ) ;
  assign n19090 = n13033 ^ n13005 ^ n7313 ;
  assign n19091 = n5826 & ~n9953 ;
  assign n19092 = n7524 & n19091 ;
  assign n19093 = ~n6683 & n10414 ;
  assign n19094 = n13684 & n17626 ;
  assign n19095 = ~n19093 & n19094 ;
  assign n19096 = n13505 ^ n315 ^ 1'b0 ;
  assign n19097 = n19095 | n19096 ;
  assign n19098 = n15406 & ~n19097 ;
  assign n19099 = n12446 & n16156 ;
  assign n19100 = n11607 & n19099 ;
  assign n19101 = ( n366 & ~n8910 ) | ( n366 & n19100 ) | ( ~n8910 & n19100 ) ;
  assign n19102 = n7387 ^ n4949 ^ n4639 ;
  assign n19103 = ( n10093 & n19101 ) | ( n10093 & ~n19102 ) | ( n19101 & ~n19102 ) ;
  assign n19104 = n17711 ^ n17618 ^ n3069 ;
  assign n19105 = n18974 ^ n1227 ^ 1'b0 ;
  assign n19106 = n9277 & ~n19105 ;
  assign n19107 = ~n1652 & n19106 ;
  assign n19108 = n19107 ^ n8039 ^ 1'b0 ;
  assign n19109 = n1819 | n9639 ;
  assign n19110 = n5334 ^ n1643 ^ 1'b0 ;
  assign n19111 = ( n2911 & ~n8502 ) | ( n2911 & n19110 ) | ( ~n8502 & n19110 ) ;
  assign n19112 = ~n7597 & n19111 ;
  assign n19113 = n19112 ^ n7988 ^ 1'b0 ;
  assign n19114 = n19113 ^ n12276 ^ 1'b0 ;
  assign n19115 = n2087 & n8765 ;
  assign n19116 = n19115 ^ n498 ^ 1'b0 ;
  assign n19117 = ~n9472 & n19116 ;
  assign n19118 = ( n1074 & n3410 ) | ( n1074 & ~n19117 ) | ( n3410 & ~n19117 ) ;
  assign n19119 = ( n2756 & ~n12829 ) | ( n2756 & n19118 ) | ( ~n12829 & n19118 ) ;
  assign n19120 = ( n3246 & ~n8800 ) | ( n3246 & n15850 ) | ( ~n8800 & n15850 ) ;
  assign n19121 = n19120 ^ n3655 ^ 1'b0 ;
  assign n19122 = n7475 ^ n5749 ^ 1'b0 ;
  assign n19123 = n13896 | n19122 ;
  assign n19124 = ~n7304 & n19123 ;
  assign n19125 = n10315 & ~n15217 ;
  assign n19126 = n7963 ^ n531 ^ 1'b0 ;
  assign n19127 = n3841 & ~n19126 ;
  assign n19130 = n12361 ^ n4255 ^ n2929 ;
  assign n19131 = n3209 | n19130 ;
  assign n19128 = ( n176 & n1234 ) | ( n176 & n4458 ) | ( n1234 & n4458 ) ;
  assign n19129 = ( x39 & n940 ) | ( x39 & ~n19128 ) | ( n940 & ~n19128 ) ;
  assign n19132 = n19131 ^ n19129 ^ 1'b0 ;
  assign n19133 = n19132 ^ n17139 ^ n2642 ;
  assign n19134 = n13449 ^ n12289 ^ n4083 ;
  assign n19135 = n7424 ^ n3463 ^ 1'b0 ;
  assign n19136 = ~n14856 & n19135 ;
  assign n19137 = n15411 & n19136 ;
  assign n19138 = n19137 ^ n4576 ^ 1'b0 ;
  assign n19139 = n2874 ^ n2058 ^ 1'b0 ;
  assign n19140 = n6697 & ~n19139 ;
  assign n19141 = n19140 ^ n7192 ^ 1'b0 ;
  assign n19142 = n19141 ^ n10433 ^ 1'b0 ;
  assign n19143 = n19138 & ~n19142 ;
  assign n19144 = n3010 ^ n990 ^ n424 ;
  assign n19145 = ~n2737 & n19144 ;
  assign n19146 = n19145 ^ n6858 ^ 1'b0 ;
  assign n19147 = n11733 ^ n182 ^ 1'b0 ;
  assign n19148 = n19146 & ~n19147 ;
  assign n19149 = n12319 & n19148 ;
  assign n19150 = n15003 ^ n14092 ^ n4673 ;
  assign n19151 = n12222 ^ n6024 ^ 1'b0 ;
  assign n19152 = ~n9849 & n18648 ;
  assign n19153 = n12975 | n13764 ;
  assign n19154 = n6224 & ~n11193 ;
  assign n19155 = n19154 ^ n14807 ^ 1'b0 ;
  assign n19156 = n5891 ^ n5606 ^ 1'b0 ;
  assign n19157 = n17776 | n19156 ;
  assign n19158 = n19157 ^ n15645 ^ 1'b0 ;
  assign n19159 = n18788 ^ n7424 ^ 1'b0 ;
  assign n19160 = n1569 & ~n19159 ;
  assign n19161 = ~n8314 & n12008 ;
  assign n19162 = ~n10977 & n19161 ;
  assign n19163 = n2528 | n12788 ;
  assign n19164 = n19162 & ~n19163 ;
  assign n19165 = n174 & ~n13643 ;
  assign n19166 = n9766 ^ n5293 ^ n2222 ;
  assign n19167 = n19165 & n19166 ;
  assign n19168 = n13683 ^ n2443 ^ 1'b0 ;
  assign n19169 = n18678 ^ n296 ^ 1'b0 ;
  assign n19170 = ( n4145 & n9920 ) | ( n4145 & n19169 ) | ( n9920 & n19169 ) ;
  assign n19171 = n10164 | n11117 ;
  assign n19172 = ~n3604 & n6561 ;
  assign n19175 = n13810 ^ n2229 ^ n1458 ;
  assign n19173 = n1202 & n2842 ;
  assign n19174 = n19173 ^ n9937 ^ n6055 ;
  assign n19176 = n19175 ^ n19174 ^ 1'b0 ;
  assign n19177 = n2329 ^ n2041 ^ 1'b0 ;
  assign n19178 = n2467 & ~n2673 ;
  assign n19179 = ~n19177 & n19178 ;
  assign n19180 = ( n5963 & n9158 ) | ( n5963 & n14155 ) | ( n9158 & n14155 ) ;
  assign n19181 = ( ~n6173 & n19179 ) | ( ~n6173 & n19180 ) | ( n19179 & n19180 ) ;
  assign n19182 = n10647 & n19181 ;
  assign n19183 = n11433 & n11642 ;
  assign n19184 = n10584 & ~n12078 ;
  assign n19185 = n19184 ^ n6319 ^ 1'b0 ;
  assign n19186 = n7878 ^ n5641 ^ 1'b0 ;
  assign n19187 = n11421 ^ n6092 ^ 1'b0 ;
  assign n19188 = n10062 ^ n2297 ^ 1'b0 ;
  assign n19189 = n19187 & n19188 ;
  assign n19190 = n19189 ^ n6896 ^ n5161 ;
  assign n19191 = n17010 ^ n3383 ^ 1'b0 ;
  assign n19192 = n2903 & n19191 ;
  assign n19193 = n19192 ^ n6987 ^ 1'b0 ;
  assign n19194 = ~n11012 & n19193 ;
  assign n19195 = n15513 ^ n1754 ^ 1'b0 ;
  assign n19196 = n19194 & ~n19195 ;
  assign n19197 = n7469 | n10580 ;
  assign n19198 = ( n1920 & ~n3628 ) | ( n1920 & n4719 ) | ( ~n3628 & n4719 ) ;
  assign n19199 = n2420 & ~n12968 ;
  assign n19200 = ~n19198 & n19199 ;
  assign n19201 = n19200 ^ n13375 ^ 1'b0 ;
  assign n19202 = n12375 ^ n9446 ^ n1418 ;
  assign n19203 = ( n2762 & n10240 ) | ( n2762 & n17320 ) | ( n10240 & n17320 ) ;
  assign n19204 = n3519 ^ n368 ^ 1'b0 ;
  assign n19205 = n1271 & n2282 ;
  assign n19206 = n5403 & n19205 ;
  assign n19207 = n8845 | n19206 ;
  assign n19208 = n19207 ^ n11544 ^ 1'b0 ;
  assign n19209 = n15644 & ~n19208 ;
  assign n19210 = ~n1462 & n19209 ;
  assign n19211 = n10554 | n17677 ;
  assign n19212 = n11150 & ~n19211 ;
  assign n19213 = ( n3160 & n3753 ) | ( n3160 & ~n8265 ) | ( n3753 & ~n8265 ) ;
  assign n19214 = n17842 ^ n10722 ^ n994 ;
  assign n19215 = n19214 ^ n17394 ^ 1'b0 ;
  assign n19216 = n3847 | n8722 ;
  assign n19217 = n19216 ^ n7197 ^ n3118 ;
  assign n19218 = n19217 ^ n4424 ^ 1'b0 ;
  assign n19219 = n2275 ^ n2031 ^ 1'b0 ;
  assign n19220 = ( ~n8432 & n10376 ) | ( ~n8432 & n11698 ) | ( n10376 & n11698 ) ;
  assign n19221 = n19220 ^ n14043 ^ n10529 ;
  assign n19222 = ( n2000 & n3165 ) | ( n2000 & ~n7659 ) | ( n3165 & ~n7659 ) ;
  assign n19223 = n6633 | n19222 ;
  assign n19224 = n5996 ^ n5523 ^ n1050 ;
  assign n19225 = ( n1894 & ~n8660 ) | ( n1894 & n17384 ) | ( ~n8660 & n17384 ) ;
  assign n19229 = n10105 ^ n937 ^ 1'b0 ;
  assign n19226 = n6392 ^ n3044 ^ 1'b0 ;
  assign n19227 = ~n4133 & n19226 ;
  assign n19228 = n19227 ^ n7832 ^ n2772 ;
  assign n19230 = n19229 ^ n19228 ^ n1411 ;
  assign n19231 = n18246 ^ n2571 ^ 1'b0 ;
  assign n19232 = n19231 ^ n8780 ^ 1'b0 ;
  assign n19233 = ( n908 & ~n7242 ) | ( n908 & n10314 ) | ( ~n7242 & n10314 ) ;
  assign n19234 = ~n1145 & n10156 ;
  assign n19235 = ~n5286 & n19234 ;
  assign n19236 = ( ~n5940 & n13505 ) | ( ~n5940 & n19235 ) | ( n13505 & n19235 ) ;
  assign n19237 = n9605 ^ n5127 ^ 1'b0 ;
  assign n19238 = n8495 | n19237 ;
  assign n19239 = n19238 ^ n13813 ^ 1'b0 ;
  assign n19244 = n2746 ^ n2147 ^ n1704 ;
  assign n19243 = n492 & ~n11984 ;
  assign n19245 = n19244 ^ n19243 ^ 1'b0 ;
  assign n19240 = n9184 ^ n5818 ^ 1'b0 ;
  assign n19241 = n4475 & n19240 ;
  assign n19242 = n2632 | n19241 ;
  assign n19246 = n19245 ^ n19242 ^ 1'b0 ;
  assign n19247 = n1406 & ~n4572 ;
  assign n19248 = ~n2985 & n19247 ;
  assign n19249 = ( n270 & n5527 ) | ( n270 & ~n19248 ) | ( n5527 & ~n19248 ) ;
  assign n19250 = n19249 ^ n15691 ^ n2116 ;
  assign n19251 = ~n6254 & n19250 ;
  assign n19252 = n11211 ^ n7565 ^ 1'b0 ;
  assign n19253 = ( n2535 & n5966 ) | ( n2535 & ~n5995 ) | ( n5966 & ~n5995 ) ;
  assign n19254 = n19253 ^ n7052 ^ n4226 ;
  assign n19255 = ~n2682 & n8928 ;
  assign n19256 = n9230 ^ n2938 ^ 1'b0 ;
  assign n19257 = n8301 & ~n19256 ;
  assign n19258 = n7545 & n18852 ;
  assign n19259 = ~n4580 & n19258 ;
  assign n19260 = ( n9172 & n9467 ) | ( n9172 & ~n10331 ) | ( n9467 & ~n10331 ) ;
  assign n19261 = n16876 ^ n921 ^ 1'b0 ;
  assign n19263 = n2326 ^ n228 ^ 1'b0 ;
  assign n19262 = n1780 | n9427 ;
  assign n19264 = n19263 ^ n19262 ^ 1'b0 ;
  assign n19265 = ~n8690 & n10263 ;
  assign n19266 = n19265 ^ n12297 ^ 1'b0 ;
  assign n19267 = n19264 & ~n19266 ;
  assign n19268 = n7940 & n19267 ;
  assign n19269 = n4799 ^ n4390 ^ n4353 ;
  assign n19270 = n13545 & n19269 ;
  assign n19271 = n9937 & ~n18262 ;
  assign n19272 = n16102 ^ n8140 ^ n2217 ;
  assign n19273 = ~n7365 & n19063 ;
  assign n19274 = n19273 ^ n10234 ^ 1'b0 ;
  assign n19275 = n10581 & n19274 ;
  assign n19277 = n13733 ^ n6794 ^ n4297 ;
  assign n19276 = n3154 & ~n9081 ;
  assign n19278 = n19277 ^ n19276 ^ n7365 ;
  assign n19279 = n19278 ^ n3763 ^ 1'b0 ;
  assign n19280 = ~n4116 & n19279 ;
  assign n19281 = n5766 ^ n4237 ^ 1'b0 ;
  assign n19282 = n19281 ^ n11292 ^ n1288 ;
  assign n19283 = n19282 ^ n9024 ^ n2780 ;
  assign n19284 = ( n2564 & ~n4534 ) | ( n2564 & n6860 ) | ( ~n4534 & n6860 ) ;
  assign n19285 = ~n19283 & n19284 ;
  assign n19286 = n10450 ^ n9608 ^ 1'b0 ;
  assign n19287 = n3398 & ~n19286 ;
  assign n19288 = n18751 ^ n14925 ^ n12892 ;
  assign n19289 = ( n2163 & n19287 ) | ( n2163 & ~n19288 ) | ( n19287 & ~n19288 ) ;
  assign n19290 = n16212 ^ n2127 ^ n1733 ;
  assign n19291 = n4251 & ~n19290 ;
  assign n19292 = n19291 ^ n15475 ^ n7105 ;
  assign n19293 = ( ~n5265 & n6811 ) | ( ~n5265 & n16128 ) | ( n6811 & n16128 ) ;
  assign n19294 = n19293 ^ n13673 ^ 1'b0 ;
  assign n19295 = n2283 & n19294 ;
  assign n19296 = n4448 & ~n12067 ;
  assign n19297 = n19296 ^ n2889 ^ 1'b0 ;
  assign n19298 = n11337 ^ n3206 ^ 1'b0 ;
  assign n19299 = n19297 | n19298 ;
  assign n19300 = n3349 & n12035 ;
  assign n19301 = ( n7986 & ~n13407 ) | ( n7986 & n19300 ) | ( ~n13407 & n19300 ) ;
  assign n19302 = n6275 | n19301 ;
  assign n19303 = n4962 & n12481 ;
  assign n19304 = n19303 ^ n8605 ^ 1'b0 ;
  assign n19305 = n19304 ^ n2292 ^ 1'b0 ;
  assign n19306 = n4335 & n19305 ;
  assign n19307 = n19306 ^ n16954 ^ 1'b0 ;
  assign n19308 = ~n11722 & n16929 ;
  assign n19309 = n8283 ^ n316 ^ 1'b0 ;
  assign n19310 = n15606 & n19309 ;
  assign n19311 = n17446 ^ n12256 ^ n11939 ;
  assign n19312 = ( n6399 & ~n7743 ) | ( n6399 & n19311 ) | ( ~n7743 & n19311 ) ;
  assign n19313 = n11783 | n16806 ;
  assign n19314 = n19313 ^ n5371 ^ 1'b0 ;
  assign n19316 = n3297 ^ n2440 ^ 1'b0 ;
  assign n19317 = n8922 & ~n19316 ;
  assign n19315 = ( n831 & ~n9822 ) | ( n831 & n15879 ) | ( ~n9822 & n15879 ) ;
  assign n19318 = n19317 ^ n19315 ^ 1'b0 ;
  assign n19319 = n11890 ^ n8503 ^ 1'b0 ;
  assign n19320 = n19319 ^ n9351 ^ n4986 ;
  assign n19321 = n5753 & n8436 ;
  assign n19322 = n19321 ^ n16158 ^ 1'b0 ;
  assign n19323 = n4639 & n15860 ;
  assign n19324 = ~n19322 & n19323 ;
  assign n19325 = n11768 & ~n12678 ;
  assign n19326 = ~n3103 & n9053 ;
  assign n19327 = n8320 | n19326 ;
  assign n19328 = n2608 & n16302 ;
  assign n19329 = n19328 ^ n12513 ^ 1'b0 ;
  assign n19330 = n19329 ^ n10249 ^ n2871 ;
  assign n19331 = ( n6306 & ~n7119 ) | ( n6306 & n12291 ) | ( ~n7119 & n12291 ) ;
  assign n19332 = n6590 & n19331 ;
  assign n19333 = ( n3958 & ~n15986 ) | ( n3958 & n19332 ) | ( ~n15986 & n19332 ) ;
  assign n19335 = n15723 ^ n238 ^ 1'b0 ;
  assign n19334 = n7820 & n15664 ;
  assign n19336 = n19335 ^ n19334 ^ 1'b0 ;
  assign n19337 = n2316 | n6842 ;
  assign n19338 = n19337 ^ n291 ^ 1'b0 ;
  assign n19339 = ( n3746 & n5274 ) | ( n3746 & ~n5373 ) | ( n5274 & ~n5373 ) ;
  assign n19340 = n19339 ^ n11648 ^ 1'b0 ;
  assign n19344 = n13367 ^ n11844 ^ n893 ;
  assign n19341 = n11147 & ~n19110 ;
  assign n19342 = n19341 ^ n7934 ^ 1'b0 ;
  assign n19343 = n19342 ^ n8598 ^ n1113 ;
  assign n19345 = n19344 ^ n19343 ^ n4129 ;
  assign n19346 = ~n6475 & n7966 ;
  assign n19347 = n5774 | n15128 ;
  assign n19348 = n5528 ^ n3076 ^ n850 ;
  assign n19349 = n6951 & n19348 ;
  assign n19350 = n19349 ^ n3405 ^ 1'b0 ;
  assign n19351 = n4892 & n19350 ;
  assign n19352 = n19351 ^ n12745 ^ 1'b0 ;
  assign n19353 = n18862 & n19352 ;
  assign n19354 = ~n18045 & n19353 ;
  assign n19355 = ( ~n5590 & n9948 ) | ( ~n5590 & n10934 ) | ( n9948 & n10934 ) ;
  assign n19356 = n19355 ^ n5151 ^ 1'b0 ;
  assign n19357 = n8379 | n10449 ;
  assign n19358 = n2724 | n19357 ;
  assign n19359 = n19358 ^ n14287 ^ n13579 ;
  assign n19360 = n12481 & ~n19359 ;
  assign n19361 = n6183 | n14149 ;
  assign n19362 = n3724 & ~n19361 ;
  assign n19363 = n875 & n5865 ;
  assign n19364 = n7156 & n19363 ;
  assign n19365 = n3510 ^ n2361 ^ 1'b0 ;
  assign n19366 = n5448 ^ n1732 ^ 1'b0 ;
  assign n19367 = ~n11115 & n19366 ;
  assign n19368 = n19367 ^ n18041 ^ 1'b0 ;
  assign n19369 = n971 & ~n2296 ;
  assign n19370 = n19369 ^ n1646 ^ n915 ;
  assign n19371 = n19370 ^ n319 ^ 1'b0 ;
  assign n19372 = n11419 & n19371 ;
  assign n19373 = ~n19368 & n19372 ;
  assign n19374 = n18232 ^ n3975 ^ 1'b0 ;
  assign n19375 = n12715 ^ n10297 ^ 1'b0 ;
  assign n19376 = ~n5443 & n19375 ;
  assign n19377 = n13160 ^ n5131 ^ 1'b0 ;
  assign n19378 = n14865 ^ n4441 ^ 1'b0 ;
  assign n19379 = n18311 ^ n12053 ^ 1'b0 ;
  assign n19380 = n2254 & n4991 ;
  assign n19381 = n19380 ^ n1283 ^ 1'b0 ;
  assign n19382 = n19381 ^ n1105 ^ 1'b0 ;
  assign n19389 = n14713 ^ n8124 ^ 1'b0 ;
  assign n19390 = n1754 & n19389 ;
  assign n19383 = ( ~x12 & n8398 ) | ( ~x12 & n9193 ) | ( n8398 & n9193 ) ;
  assign n19384 = n14260 & ~n19383 ;
  assign n19385 = n19384 ^ n2178 ^ 1'b0 ;
  assign n19386 = n2125 & ~n19385 ;
  assign n19387 = n9512 & n19386 ;
  assign n19388 = n6621 | n19387 ;
  assign n19391 = n19390 ^ n19388 ^ 1'b0 ;
  assign n19392 = n1867 | n4971 ;
  assign n19393 = n19392 ^ n4972 ^ n834 ;
  assign n19394 = n3136 | n19393 ;
  assign n19395 = n18232 ^ n10981 ^ 1'b0 ;
  assign n19396 = n19394 & n19395 ;
  assign n19397 = n16833 ^ n15921 ^ n5405 ;
  assign n19398 = n4984 | n7916 ;
  assign n19399 = n14908 & ~n19398 ;
  assign n19400 = n550 | n9511 ;
  assign n19401 = n2989 & n19400 ;
  assign n19402 = n19401 ^ n2350 ^ 1'b0 ;
  assign n19403 = n10846 ^ n2523 ^ 1'b0 ;
  assign n19404 = n509 & n19403 ;
  assign n19405 = n19404 ^ n6099 ^ n5706 ;
  assign n19406 = ~n9402 & n19405 ;
  assign n19407 = n19406 ^ n5922 ^ 1'b0 ;
  assign n19408 = ( n4406 & n7481 ) | ( n4406 & n8879 ) | ( n7481 & n8879 ) ;
  assign n19410 = n16651 ^ n9552 ^ n1670 ;
  assign n19409 = n10422 & n11879 ;
  assign n19411 = n19410 ^ n19409 ^ 1'b0 ;
  assign n19412 = ( n5522 & n19408 ) | ( n5522 & ~n19411 ) | ( n19408 & ~n19411 ) ;
  assign n19413 = n10033 | n11688 ;
  assign n19414 = n15999 ^ n11215 ^ n6060 ;
  assign n19415 = x101 & n13467 ;
  assign n19416 = n19414 & n19415 ;
  assign n19417 = n10474 ^ n808 ^ 1'b0 ;
  assign n19418 = ~n19416 & n19417 ;
  assign n19419 = n8140 | n10843 ;
  assign n19420 = n2125 & ~n6469 ;
  assign n19421 = ~n19419 & n19420 ;
  assign n19422 = n15263 | n17621 ;
  assign n19423 = n10199 ^ n3761 ^ 1'b0 ;
  assign n19424 = n3807 & ~n19423 ;
  assign n19425 = n11491 ^ n7271 ^ 1'b0 ;
  assign n19426 = n19425 ^ n7229 ^ n1972 ;
  assign n19427 = n8035 & n13003 ;
  assign n19428 = n13201 ^ n3279 ^ 1'b0 ;
  assign n19429 = ~n5323 & n19428 ;
  assign n19430 = ( x101 & ~n2768 ) | ( x101 & n19429 ) | ( ~n2768 & n19429 ) ;
  assign n19431 = ( n4526 & n19427 ) | ( n4526 & ~n19430 ) | ( n19427 & ~n19430 ) ;
  assign n19432 = n1275 & n4237 ;
  assign n19433 = n19432 ^ n6421 ^ 1'b0 ;
  assign n19434 = n19433 ^ n2514 ^ 1'b0 ;
  assign n19435 = ( ~n3823 & n11972 ) | ( ~n3823 & n19434 ) | ( n11972 & n19434 ) ;
  assign n19436 = n19435 ^ n16258 ^ 1'b0 ;
  assign n19437 = ~n17846 & n19436 ;
  assign n19438 = ( n744 & ~n6888 ) | ( n744 & n12080 ) | ( ~n6888 & n12080 ) ;
  assign n19439 = ~n2244 & n3281 ;
  assign n19440 = n19439 ^ n1889 ^ 1'b0 ;
  assign n19441 = n5490 & ~n19440 ;
  assign n19442 = ~n1055 & n1455 ;
  assign n19443 = n19442 ^ n1320 ^ 1'b0 ;
  assign n19444 = ( n9580 & ~n17030 ) | ( n9580 & n19443 ) | ( ~n17030 & n19443 ) ;
  assign n19445 = n19444 ^ n5535 ^ 1'b0 ;
  assign n19446 = n9253 & ~n19445 ;
  assign n19447 = ( n5014 & n19441 ) | ( n5014 & ~n19446 ) | ( n19441 & ~n19446 ) ;
  assign n19448 = n16482 ^ n6633 ^ 1'b0 ;
  assign n19449 = n1312 | n19448 ;
  assign n19450 = n19449 ^ n1918 ^ 1'b0 ;
  assign n19451 = n19450 ^ n522 ^ 1'b0 ;
  assign n19452 = n14427 ^ n10538 ^ n3533 ;
  assign n19453 = n19452 ^ n5060 ^ n3968 ;
  assign n19455 = n11782 ^ n9172 ^ 1'b0 ;
  assign n19454 = n7763 & n16289 ;
  assign n19456 = n19455 ^ n19454 ^ 1'b0 ;
  assign n19457 = n17714 ^ n13738 ^ 1'b0 ;
  assign n19458 = n3677 & ~n5724 ;
  assign n19459 = n3459 | n4448 ;
  assign n19460 = ( n2124 & ~n5380 ) | ( n2124 & n7079 ) | ( ~n5380 & n7079 ) ;
  assign n19461 = ( n19458 & n19459 ) | ( n19458 & n19460 ) | ( n19459 & n19460 ) ;
  assign n19462 = n15022 & n19154 ;
  assign n19463 = n8040 ^ n7504 ^ 1'b0 ;
  assign n19464 = n19462 | n19463 ;
  assign n19465 = ( n11086 & n19461 ) | ( n11086 & n19464 ) | ( n19461 & n19464 ) ;
  assign n19466 = n5248 ^ n2141 ^ n419 ;
  assign n19467 = ( n2354 & n7854 ) | ( n2354 & ~n15681 ) | ( n7854 & ~n15681 ) ;
  assign n19468 = n5913 ^ n4786 ^ 1'b0 ;
  assign n19469 = n19468 ^ n5774 ^ 1'b0 ;
  assign n19470 = n12821 & n19469 ;
  assign n19471 = ~n545 & n13555 ;
  assign n19474 = n2558 & n10915 ;
  assign n19473 = n4999 & ~n7407 ;
  assign n19475 = n19474 ^ n19473 ^ 1'b0 ;
  assign n19472 = n15096 & n16921 ;
  assign n19476 = n19475 ^ n19472 ^ n3644 ;
  assign n19477 = ( n7156 & n19471 ) | ( n7156 & n19476 ) | ( n19471 & n19476 ) ;
  assign n19478 = n19477 ^ n10413 ^ 1'b0 ;
  assign n19479 = n5004 | n19478 ;
  assign n19480 = n5940 | n9015 ;
  assign n19481 = ( n11235 & n13168 ) | ( n11235 & ~n19480 ) | ( n13168 & ~n19480 ) ;
  assign n19482 = n7634 | n19481 ;
  assign n19483 = n19482 ^ n11050 ^ 1'b0 ;
  assign n19484 = ( n10940 & n16394 ) | ( n10940 & ~n19036 ) | ( n16394 & ~n19036 ) ;
  assign n19485 = ( n7725 & n8770 ) | ( n7725 & ~n11730 ) | ( n8770 & ~n11730 ) ;
  assign n19486 = n19485 ^ n19339 ^ n4735 ;
  assign n19487 = ~n2515 & n5764 ;
  assign n19488 = ~n2399 & n19487 ;
  assign n19489 = ~n4980 & n19488 ;
  assign n19490 = ( ~n1295 & n3641 ) | ( ~n1295 & n9368 ) | ( n3641 & n9368 ) ;
  assign n19491 = n6572 & ~n19490 ;
  assign n19492 = x107 & ~n12117 ;
  assign n19493 = ~n19491 & n19492 ;
  assign n19494 = n19489 & ~n19493 ;
  assign n19495 = ( n8949 & n10667 ) | ( n8949 & n11777 ) | ( n10667 & n11777 ) ;
  assign n19496 = n11710 & ~n18117 ;
  assign n19497 = ~n19495 & n19496 ;
  assign n19498 = n12491 ^ n6173 ^ n149 ;
  assign n19499 = n19498 ^ n17278 ^ n13219 ;
  assign n19500 = n1843 & ~n19499 ;
  assign n19506 = n4628 & n11282 ;
  assign n19507 = ~n16146 & n19506 ;
  assign n19508 = n19507 ^ n10467 ^ n4722 ;
  assign n19501 = ( x90 & n1949 ) | ( x90 & n12963 ) | ( n1949 & n12963 ) ;
  assign n19502 = n19501 ^ n6436 ^ n1124 ;
  assign n19503 = n19502 ^ n4164 ^ 1'b0 ;
  assign n19504 = ~n14839 & n19503 ;
  assign n19505 = n15685 & n19504 ;
  assign n19509 = n19508 ^ n19505 ^ 1'b0 ;
  assign n19510 = ~n3035 & n8020 ;
  assign n19511 = n10993 | n19510 ;
  assign n19513 = n11795 ^ n2624 ^ n597 ;
  assign n19512 = n965 & n17926 ;
  assign n19514 = n19513 ^ n19512 ^ n5400 ;
  assign n19515 = n451 & ~n6074 ;
  assign n19516 = n4124 ^ n1385 ^ 1'b0 ;
  assign n19517 = n13127 & n19516 ;
  assign n19518 = ~n3630 & n19517 ;
  assign n19519 = n19515 & ~n19518 ;
  assign n19520 = ~n9362 & n10330 ;
  assign n19521 = n13614 ^ n8844 ^ 1'b0 ;
  assign n19522 = ( ~n3224 & n5463 ) | ( ~n3224 & n8508 ) | ( n5463 & n8508 ) ;
  assign n19523 = n16036 | n19522 ;
  assign n19524 = ( ~n1647 & n13019 ) | ( ~n1647 & n17734 ) | ( n13019 & n17734 ) ;
  assign n19525 = n19524 ^ n7301 ^ 1'b0 ;
  assign n19526 = ~n18308 & n19525 ;
  assign n19527 = n9587 ^ n8273 ^ 1'b0 ;
  assign n19528 = n7935 | n19527 ;
  assign n19537 = n761 & n9559 ;
  assign n19538 = ~n9087 & n19537 ;
  assign n19529 = n5498 ^ n1605 ^ 1'b0 ;
  assign n19533 = n14461 ^ n12460 ^ 1'b0 ;
  assign n19534 = ~n7033 & n19533 ;
  assign n19530 = n14176 ^ n6334 ^ 1'b0 ;
  assign n19531 = ~n1515 & n19530 ;
  assign n19532 = n15833 | n19531 ;
  assign n19535 = n19534 ^ n19532 ^ n13421 ;
  assign n19536 = ( n12554 & n19529 ) | ( n12554 & n19535 ) | ( n19529 & n19535 ) ;
  assign n19539 = n19538 ^ n19536 ^ n9953 ;
  assign n19540 = n8874 ^ x27 ^ 1'b0 ;
  assign n19541 = n13141 & n19540 ;
  assign n19542 = n6793 | n7579 ;
  assign n19543 = n4970 & ~n19542 ;
  assign n19544 = n4376 | n4770 ;
  assign n19545 = n19544 ^ n10564 ^ 1'b0 ;
  assign n19546 = ( n13135 & ~n19543 ) | ( n13135 & n19545 ) | ( ~n19543 & n19545 ) ;
  assign n19547 = n6067 & n19546 ;
  assign n19548 = n3994 & n5133 ;
  assign n19549 = n3862 & n19548 ;
  assign n19550 = ~n930 & n8493 ;
  assign n19551 = n7116 | n13110 ;
  assign n19552 = n10123 ^ n3137 ^ 1'b0 ;
  assign n19553 = ~n3610 & n19552 ;
  assign n19554 = n19553 ^ n14905 ^ 1'b0 ;
  assign n19555 = ( n6890 & n19551 ) | ( n6890 & ~n19554 ) | ( n19551 & ~n19554 ) ;
  assign n19556 = ( ~n7994 & n10831 ) | ( ~n7994 & n16979 ) | ( n10831 & n16979 ) ;
  assign n19557 = n10062 | n19556 ;
  assign n19558 = n19557 ^ n11730 ^ n4645 ;
  assign n19559 = n19558 ^ n16915 ^ n7103 ;
  assign n19560 = n8883 ^ n8777 ^ 1'b0 ;
  assign n19561 = ~n13965 & n14952 ;
  assign n19562 = ~n652 & n19561 ;
  assign n19563 = n12724 & ~n19562 ;
  assign n19564 = ~n19560 & n19563 ;
  assign n19565 = n8092 & ~n13885 ;
  assign n19566 = ~n6699 & n7724 ;
  assign n19567 = n19566 ^ n6899 ^ 1'b0 ;
  assign n19568 = n11362 & ~n12147 ;
  assign n19569 = n4327 | n19568 ;
  assign n19570 = n3366 | n19569 ;
  assign n19571 = n2925 | n13696 ;
  assign n19572 = n2647 | n19571 ;
  assign n19573 = ( n19567 & n19570 ) | ( n19567 & ~n19572 ) | ( n19570 & ~n19572 ) ;
  assign n19574 = ~n294 & n1445 ;
  assign n19575 = n19574 ^ n5078 ^ 1'b0 ;
  assign n19576 = n1548 & n19575 ;
  assign n19582 = n18027 ^ n5164 ^ 1'b0 ;
  assign n19583 = n1739 & n19582 ;
  assign n19577 = n3465 & n7085 ;
  assign n19578 = n19577 ^ n4176 ^ 1'b0 ;
  assign n19579 = n19578 ^ n5711 ^ 1'b0 ;
  assign n19580 = n3111 & ~n19579 ;
  assign n19581 = ~n6779 & n19580 ;
  assign n19584 = n19583 ^ n19581 ^ n6922 ;
  assign n19585 = n7346 & ~n14179 ;
  assign n19586 = n19585 ^ n17911 ^ n12657 ;
  assign n19587 = n2152 | n14813 ;
  assign n19590 = ~n3215 & n11632 ;
  assign n19588 = ( ~n7434 & n9076 ) | ( ~n7434 & n12654 ) | ( n9076 & n12654 ) ;
  assign n19589 = n19588 ^ n16214 ^ n4661 ;
  assign n19591 = n19590 ^ n19589 ^ 1'b0 ;
  assign n19593 = n5097 ^ n4202 ^ 1'b0 ;
  assign n19594 = ~n13079 & n19593 ;
  assign n19592 = n12864 ^ n5821 ^ n1511 ;
  assign n19595 = n19594 ^ n19592 ^ n4779 ;
  assign n19596 = n7907 ^ n6605 ^ n1637 ;
  assign n19597 = n15265 ^ n13685 ^ 1'b0 ;
  assign n19598 = n12494 | n19597 ;
  assign n19599 = n2860 | n10017 ;
  assign n19600 = n865 & ~n3509 ;
  assign n19601 = n19600 ^ n15081 ^ 1'b0 ;
  assign n19602 = n8458 ^ n7357 ^ 1'b0 ;
  assign n19603 = n19601 | n19602 ;
  assign n19604 = n706 & n4232 ;
  assign n19605 = n19604 ^ n9762 ^ 1'b0 ;
  assign n19606 = n19605 ^ n15859 ^ 1'b0 ;
  assign n19607 = n17879 ^ n14775 ^ n2336 ;
  assign n19608 = n582 & ~n1439 ;
  assign n19609 = n1587 & n19608 ;
  assign n19610 = ( ~n12139 & n18760 ) | ( ~n12139 & n19609 ) | ( n18760 & n19609 ) ;
  assign n19611 = n5674 & n10916 ;
  assign n19612 = n19611 ^ n3035 ^ 1'b0 ;
  assign n19613 = n13684 ^ n4174 ^ 1'b0 ;
  assign n19614 = n2639 ^ n495 ^ 1'b0 ;
  assign n19615 = ~n6325 & n19614 ;
  assign n19616 = n19393 & n19615 ;
  assign n19617 = n19616 ^ n9121 ^ 1'b0 ;
  assign n19618 = n19617 ^ n16725 ^ 1'b0 ;
  assign n19619 = n18782 ^ n16004 ^ n4969 ;
  assign n19620 = ( n12465 & n15146 ) | ( n12465 & n17901 ) | ( n15146 & n17901 ) ;
  assign n19622 = n1264 & n2715 ;
  assign n19621 = n17482 ^ n2404 ^ 1'b0 ;
  assign n19623 = n19622 ^ n19621 ^ n17944 ;
  assign n19624 = n1598 & n2937 ;
  assign n19625 = ~n10122 & n19624 ;
  assign n19626 = n18817 & ~n19625 ;
  assign n19627 = x49 & n10467 ;
  assign n19628 = ( ~n12139 & n13649 ) | ( ~n12139 & n19627 ) | ( n13649 & n19627 ) ;
  assign n19629 = ( n1277 & ~n2679 ) | ( n1277 & n7848 ) | ( ~n2679 & n7848 ) ;
  assign n19630 = n19629 ^ n9938 ^ n4415 ;
  assign n19631 = n5173 ^ n3973 ^ n1188 ;
  assign n19632 = n7682 | n19631 ;
  assign n19633 = n9948 ^ n8987 ^ 1'b0 ;
  assign n19634 = n19632 & n19633 ;
  assign n19635 = n6210 & n6451 ;
  assign n19636 = n4157 ^ n2939 ^ n1384 ;
  assign n19637 = n19635 & n19636 ;
  assign n19638 = n11027 ^ n5822 ^ 1'b0 ;
  assign n19639 = ( n1779 & n9899 ) | ( n1779 & n19638 ) | ( n9899 & n19638 ) ;
  assign n19640 = n19639 ^ n5762 ^ 1'b0 ;
  assign n19641 = n8055 ^ x113 ^ 1'b0 ;
  assign n19642 = n267 & ~n3235 ;
  assign n19643 = ( ~n4465 & n5387 ) | ( ~n4465 & n19642 ) | ( n5387 & n19642 ) ;
  assign n19644 = n1543 & ~n16306 ;
  assign n19645 = ~n2663 & n19644 ;
  assign n19646 = ( n4414 & n13278 ) | ( n4414 & n19645 ) | ( n13278 & n19645 ) ;
  assign n19648 = n4091 ^ n2232 ^ 1'b0 ;
  assign n19647 = n13005 ^ n1494 ^ 1'b0 ;
  assign n19649 = n19648 ^ n19647 ^ 1'b0 ;
  assign n19650 = n19649 ^ n10552 ^ 1'b0 ;
  assign n19651 = n6439 ^ n1537 ^ 1'b0 ;
  assign n19652 = n969 | n13777 ;
  assign n19653 = ( ~n3607 & n19651 ) | ( ~n3607 & n19652 ) | ( n19651 & n19652 ) ;
  assign n19654 = n19653 ^ n6298 ^ 1'b0 ;
  assign n19655 = n13754 | n15757 ;
  assign n19656 = n15496 & ~n19655 ;
  assign n19657 = n11481 | n19656 ;
  assign n19658 = n19657 ^ n4956 ^ 1'b0 ;
  assign n19659 = n2013 | n9015 ;
  assign n19660 = x7 | n19659 ;
  assign n19661 = n16208 ^ n5139 ^ 1'b0 ;
  assign n19662 = n5673 & ~n16595 ;
  assign n19663 = ( n250 & n3218 ) | ( n250 & n9402 ) | ( n3218 & n9402 ) ;
  assign n19670 = x100 & ~n971 ;
  assign n19671 = n19670 ^ n2596 ^ 1'b0 ;
  assign n19672 = ( ~n964 & n1262 ) | ( ~n964 & n19671 ) | ( n1262 & n19671 ) ;
  assign n19666 = n5891 ^ n4105 ^ n2214 ;
  assign n19667 = n19666 ^ n18092 ^ n7127 ;
  assign n19668 = n19667 ^ n8571 ^ n6817 ;
  assign n19669 = ( n1543 & ~n2336 ) | ( n1543 & n19668 ) | ( ~n2336 & n19668 ) ;
  assign n19664 = n5322 & ~n10273 ;
  assign n19665 = n19664 ^ n723 ^ 1'b0 ;
  assign n19673 = n19672 ^ n19669 ^ n19665 ;
  assign n19674 = n9957 ^ n9403 ^ n8441 ;
  assign n19675 = n2205 & n15452 ;
  assign n19676 = n3247 & n19675 ;
  assign n19677 = ~n8530 & n14899 ;
  assign n19678 = n12204 & n19677 ;
  assign n19679 = ~n11646 & n17865 ;
  assign n19680 = ~n526 & n3010 ;
  assign n19681 = ~n3319 & n14465 ;
  assign n19682 = n5609 & n7951 ;
  assign n19683 = ( n5702 & ~n8341 ) | ( n5702 & n19682 ) | ( ~n8341 & n19682 ) ;
  assign n19684 = ( n7105 & n8371 ) | ( n7105 & n10915 ) | ( n8371 & n10915 ) ;
  assign n19685 = n17434 & n19684 ;
  assign n19686 = ~n3788 & n7954 ;
  assign n19687 = n19686 ^ n7254 ^ 1'b0 ;
  assign n19688 = n19687 ^ n13135 ^ n7907 ;
  assign n19689 = ~n9472 & n16738 ;
  assign n19690 = ~n1592 & n19689 ;
  assign n19691 = n13391 & n19690 ;
  assign n19692 = n19691 ^ n16277 ^ n4949 ;
  assign n19693 = ( n2304 & n17212 ) | ( n2304 & ~n19639 ) | ( n17212 & ~n19639 ) ;
  assign n19694 = ( n2302 & ~n5995 ) | ( n2302 & n17107 ) | ( ~n5995 & n17107 ) ;
  assign n19695 = n8271 ^ n8242 ^ 1'b0 ;
  assign n19696 = n17120 & ~n19695 ;
  assign n19697 = n5996 | n14310 ;
  assign n19698 = n19697 ^ n6187 ^ 1'b0 ;
  assign n19699 = ~n12380 & n19698 ;
  assign n19700 = n7467 & n19699 ;
  assign n19701 = n19700 ^ n3799 ^ 1'b0 ;
  assign n19705 = n8582 & ~n14827 ;
  assign n19702 = n12051 ^ n6256 ^ n911 ;
  assign n19703 = n16483 ^ n13005 ^ n3296 ;
  assign n19704 = ( n2377 & n19702 ) | ( n2377 & n19703 ) | ( n19702 & n19703 ) ;
  assign n19706 = n19705 ^ n19704 ^ n6951 ;
  assign n19707 = n637 & ~n1753 ;
  assign n19708 = ~n637 & n19707 ;
  assign n19709 = ~n8354 & n19708 ;
  assign n19710 = n1387 & n19709 ;
  assign n19711 = n1283 & n19710 ;
  assign n19712 = n19711 ^ n2255 ^ 1'b0 ;
  assign n19713 = ( ~n3573 & n11698 ) | ( ~n3573 & n19712 ) | ( n11698 & n19712 ) ;
  assign n19714 = n1553 & ~n4859 ;
  assign n19715 = n2799 | n19714 ;
  assign n19716 = ~n1922 & n14664 ;
  assign n19717 = n5465 ^ n406 ^ 1'b0 ;
  assign n19718 = n12560 ^ n4465 ^ 1'b0 ;
  assign n19719 = n13678 & ~n19718 ;
  assign n19720 = n19719 ^ n7412 ^ n924 ;
  assign n19721 = ( n7299 & ~n9463 ) | ( n7299 & n14887 ) | ( ~n9463 & n14887 ) ;
  assign n19722 = ~n5392 & n5894 ;
  assign n19723 = n13396 ^ n12663 ^ n8723 ;
  assign n19724 = ( n6068 & ~n8131 ) | ( n6068 & n19723 ) | ( ~n8131 & n19723 ) ;
  assign n19725 = n16081 ^ n4857 ^ 1'b0 ;
  assign n19726 = ~n19724 & n19725 ;
  assign n19727 = n508 & n4082 ;
  assign n19728 = n19698 | n19727 ;
  assign n19729 = n12501 ^ n12446 ^ n6128 ;
  assign n19730 = n11150 ^ n8928 ^ n4042 ;
  assign n19731 = n5126 ^ n3496 ^ 1'b0 ;
  assign n19732 = n4708 & n19731 ;
  assign n19733 = n3367 & n19732 ;
  assign n19734 = ~n19730 & n19733 ;
  assign n19735 = n17865 ^ n9256 ^ 1'b0 ;
  assign n19736 = n13634 & ~n19735 ;
  assign n19737 = ( ~n19729 & n19734 ) | ( ~n19729 & n19736 ) | ( n19734 & n19736 ) ;
  assign n19738 = n4004 | n10048 ;
  assign n19739 = n955 & n12982 ;
  assign n19740 = ( n5241 & ~n14029 ) | ( n5241 & n19739 ) | ( ~n14029 & n19739 ) ;
  assign n19741 = n1466 & n5370 ;
  assign n19742 = n3503 & n19741 ;
  assign n19743 = ( n11027 & n15795 ) | ( n11027 & n19742 ) | ( n15795 & n19742 ) ;
  assign n19744 = n19740 & n19743 ;
  assign n19745 = n13334 | n19744 ;
  assign n19746 = n5815 | n19745 ;
  assign n19747 = ( n4874 & n5083 ) | ( n4874 & n9830 ) | ( n5083 & n9830 ) ;
  assign n19748 = n11560 & ~n19747 ;
  assign n19749 = n14463 ^ n13158 ^ n9673 ;
  assign n19750 = n7572 | n16762 ;
  assign n19751 = ( n5670 & n18137 ) | ( n5670 & ~n19750 ) | ( n18137 & ~n19750 ) ;
  assign n19752 = n19751 ^ n11841 ^ 1'b0 ;
  assign n19753 = n7243 ^ n6565 ^ 1'b0 ;
  assign n19754 = n19753 ^ n15112 ^ 1'b0 ;
  assign n19755 = ~n17369 & n19754 ;
  assign n19756 = ~n5231 & n19755 ;
  assign n19757 = ~n6210 & n7945 ;
  assign n19758 = n8833 & ~n19757 ;
  assign n19759 = n2567 & n19758 ;
  assign n19760 = n11668 ^ n5301 ^ 1'b0 ;
  assign n19761 = n10095 ^ n7542 ^ 1'b0 ;
  assign n19762 = n19760 & n19761 ;
  assign n19764 = n137 & ~n11404 ;
  assign n19765 = n3845 & n7863 ;
  assign n19766 = n19765 ^ n19072 ^ 1'b0 ;
  assign n19767 = n9547 & n19766 ;
  assign n19768 = ( n7025 & n14463 ) | ( n7025 & ~n14784 ) | ( n14463 & ~n14784 ) ;
  assign n19769 = ( n19764 & ~n19767 ) | ( n19764 & n19768 ) | ( ~n19767 & n19768 ) ;
  assign n19763 = n14245 | n14297 ;
  assign n19770 = n19769 ^ n19763 ^ n13673 ;
  assign n19771 = ( n1559 & n2998 ) | ( n1559 & ~n10458 ) | ( n2998 & ~n10458 ) ;
  assign n19772 = n174 & ~n13685 ;
  assign n19773 = n19772 ^ n10400 ^ 1'b0 ;
  assign n19774 = n9342 ^ n4684 ^ n4025 ;
  assign n19775 = n14273 ^ n9460 ^ n9374 ;
  assign n19776 = ~n2797 & n8273 ;
  assign n19777 = ~n7954 & n19776 ;
  assign n19778 = ( n7190 & ~n9102 ) | ( n7190 & n19777 ) | ( ~n9102 & n19777 ) ;
  assign n19779 = n15992 ^ n10327 ^ 1'b0 ;
  assign n19780 = n3232 & n19779 ;
  assign n19781 = n19780 ^ n5180 ^ 1'b0 ;
  assign n19782 = n17596 ^ n14711 ^ n4691 ;
  assign n19783 = ( n694 & n7053 ) | ( n694 & n8512 ) | ( n7053 & n8512 ) ;
  assign n19784 = n19783 ^ n10368 ^ 1'b0 ;
  assign n19785 = ~n1704 & n2279 ;
  assign n19786 = ~n19408 & n19785 ;
  assign n19787 = n2601 & ~n7022 ;
  assign n19788 = ~n8175 & n19787 ;
  assign n19789 = n8075 & n19788 ;
  assign n19791 = ( n669 & ~n2513 ) | ( n669 & n10074 ) | ( ~n2513 & n10074 ) ;
  assign n19792 = ( x115 & ~n2522 ) | ( x115 & n6322 ) | ( ~n2522 & n6322 ) ;
  assign n19793 = n10250 ^ n6353 ^ 1'b0 ;
  assign n19794 = ~n5396 & n19793 ;
  assign n19795 = n19794 ^ n7733 ^ 1'b0 ;
  assign n19796 = n6049 & n19795 ;
  assign n19797 = ( ~n11518 & n19792 ) | ( ~n11518 & n19796 ) | ( n19792 & n19796 ) ;
  assign n19798 = n926 & n19797 ;
  assign n19799 = n19791 & n19798 ;
  assign n19790 = n1017 | n18835 ;
  assign n19800 = n19799 ^ n19790 ^ 1'b0 ;
  assign n19801 = ~n2042 & n8341 ;
  assign n19802 = n19801 ^ n17832 ^ 1'b0 ;
  assign n19803 = n7136 | n9855 ;
  assign n19804 = ~n15275 & n19803 ;
  assign n19805 = n1918 | n9658 ;
  assign n19806 = n1952 | n19805 ;
  assign n19807 = n19806 ^ n13065 ^ n2163 ;
  assign n19808 = ( n3553 & n6700 ) | ( n3553 & n10963 ) | ( n6700 & n10963 ) ;
  assign n19809 = ( n5858 & n15859 ) | ( n5858 & n16067 ) | ( n15859 & n16067 ) ;
  assign n19810 = n19809 ^ n9801 ^ n2074 ;
  assign n19811 = n16324 ^ n6184 ^ 1'b0 ;
  assign n19812 = n14441 & ~n19811 ;
  assign n19813 = n19812 ^ n1003 ^ 1'b0 ;
  assign n19814 = n2559 ^ n2282 ^ 1'b0 ;
  assign n19815 = n2257 | n19814 ;
  assign n19816 = n2204 & ~n19815 ;
  assign n19817 = n3677 & ~n19816 ;
  assign n19818 = n5925 & n6046 ;
  assign n19819 = n19818 ^ n7012 ^ 1'b0 ;
  assign n19820 = n19819 ^ n6399 ^ n4743 ;
  assign n19821 = n10193 & n10993 ;
  assign n19822 = n6676 & ~n19821 ;
  assign n19823 = n4772 & n19822 ;
  assign n19824 = n7839 ^ n2077 ^ n2060 ;
  assign n19825 = n16168 ^ n8839 ^ 1'b0 ;
  assign n19826 = ~n19824 & n19825 ;
  assign n19827 = ( n804 & n11720 ) | ( n804 & n18887 ) | ( n11720 & n18887 ) ;
  assign n19828 = ~n8552 & n12345 ;
  assign n19829 = n17568 ^ n14668 ^ n2310 ;
  assign n19830 = n19829 ^ n13623 ^ n2008 ;
  assign n19831 = n5013 | n18112 ;
  assign n19832 = n19831 ^ n13104 ^ 1'b0 ;
  assign n19834 = n13480 & ~n16929 ;
  assign n19835 = n19834 ^ n7886 ^ 1'b0 ;
  assign n19836 = ~n366 & n6477 ;
  assign n19837 = n9386 & n19836 ;
  assign n19838 = ~n19835 & n19837 ;
  assign n19833 = n14091 ^ n398 ^ 1'b0 ;
  assign n19839 = n19838 ^ n19833 ^ n2058 ;
  assign n19840 = ( n1385 & n4508 ) | ( n1385 & n11326 ) | ( n4508 & n11326 ) ;
  assign n19841 = n14216 ^ n12503 ^ n5706 ;
  assign n19842 = ( ~n8206 & n19840 ) | ( ~n8206 & n19841 ) | ( n19840 & n19841 ) ;
  assign n19843 = n19842 ^ n13119 ^ 1'b0 ;
  assign n19844 = ( ~n8159 & n15586 ) | ( ~n8159 & n19843 ) | ( n15586 & n19843 ) ;
  assign n19845 = n2955 | n4430 ;
  assign n19846 = n7654 | n19845 ;
  assign n19847 = ( ~n4991 & n6848 ) | ( ~n4991 & n18254 ) | ( n6848 & n18254 ) ;
  assign n19848 = ~n7890 & n19847 ;
  assign n19849 = n16241 | n19848 ;
  assign n19850 = n19849 ^ n7897 ^ 1'b0 ;
  assign n19851 = n19846 & ~n19850 ;
  assign n19852 = n3322 | n15018 ;
  assign n19853 = n19852 ^ n4410 ^ 1'b0 ;
  assign n19854 = n18678 ^ n15211 ^ 1'b0 ;
  assign n19855 = ( ~n5862 & n6796 ) | ( ~n5862 & n19854 ) | ( n6796 & n19854 ) ;
  assign n19856 = n19855 ^ n16275 ^ n4344 ;
  assign n19857 = ~n9321 & n12938 ;
  assign n19858 = n19857 ^ n9775 ^ 1'b0 ;
  assign n19859 = n19858 ^ n16932 ^ 1'b0 ;
  assign n19860 = ~n571 & n12787 ;
  assign n19861 = n17283 & n19860 ;
  assign n19862 = n7612 ^ n6565 ^ 1'b0 ;
  assign n19863 = n18095 & n19862 ;
  assign n19864 = ( ~n3281 & n6714 ) | ( ~n3281 & n19732 ) | ( n6714 & n19732 ) ;
  assign n19865 = ~n325 & n4179 ;
  assign n19866 = n5132 & n19865 ;
  assign n19867 = n19864 & ~n19866 ;
  assign n19868 = ~n12938 & n19867 ;
  assign n19869 = n12569 & ~n17580 ;
  assign n19872 = n11164 ^ n8052 ^ 1'b0 ;
  assign n19873 = n14106 & n19872 ;
  assign n19870 = n3062 & n4022 ;
  assign n19871 = n9469 & n19870 ;
  assign n19874 = n19873 ^ n19871 ^ 1'b0 ;
  assign n19875 = n19671 ^ n850 ^ 1'b0 ;
  assign n19876 = n19875 ^ n5063 ^ 1'b0 ;
  assign n19877 = ~n153 & n19876 ;
  assign n19878 = n8117 & n16342 ;
  assign n19879 = n13244 & n19878 ;
  assign n19880 = n7306 ^ n3499 ^ 1'b0 ;
  assign n19881 = ~n19879 & n19880 ;
  assign n19882 = ~n19877 & n19881 ;
  assign n19883 = n4199 ^ n2098 ^ 1'b0 ;
  assign n19884 = n6344 | n19883 ;
  assign n19885 = n2087 | n19884 ;
  assign n19886 = n848 & ~n19885 ;
  assign n19887 = n19886 ^ n16728 ^ n687 ;
  assign n19888 = n14493 & ~n14709 ;
  assign n19889 = ~n3202 & n19888 ;
  assign n19891 = n16945 ^ n7339 ^ n4410 ;
  assign n19890 = n7986 ^ n603 ^ 1'b0 ;
  assign n19892 = n19891 ^ n19890 ^ n5316 ;
  assign n19893 = ( n19887 & ~n19889 ) | ( n19887 & n19892 ) | ( ~n19889 & n19892 ) ;
  assign n19894 = ~n1794 & n4564 ;
  assign n19895 = n11678 & n19894 ;
  assign n19896 = ( ~n12135 & n19322 ) | ( ~n12135 & n19895 ) | ( n19322 & n19895 ) ;
  assign n19897 = ( ~n7820 & n10587 ) | ( ~n7820 & n14098 ) | ( n10587 & n14098 ) ;
  assign n19898 = n17828 ^ n15272 ^ n334 ;
  assign n19899 = ( ~n3777 & n15551 ) | ( ~n3777 & n19366 ) | ( n15551 & n19366 ) ;
  assign n19900 = ( n19897 & n19898 ) | ( n19897 & ~n19899 ) | ( n19898 & ~n19899 ) ;
  assign n19901 = n16803 & ~n17376 ;
  assign n19903 = n2451 & n4666 ;
  assign n19904 = n19903 ^ n11308 ^ 1'b0 ;
  assign n19902 = n6170 ^ n2781 ^ n1056 ;
  assign n19905 = n19904 ^ n19902 ^ n2172 ;
  assign n19906 = n19901 | n19905 ;
  assign n19907 = n3346 & n3432 ;
  assign n19908 = ~n693 & n19907 ;
  assign n19909 = n19796 ^ n8360 ^ 1'b0 ;
  assign n19910 = ~n19908 & n19909 ;
  assign n19911 = n1072 & ~n1535 ;
  assign n19912 = n19911 ^ n13209 ^ 1'b0 ;
  assign n19913 = ~n17956 & n19912 ;
  assign n19914 = n19913 ^ n11893 ^ 1'b0 ;
  assign n19915 = n1607 | n6371 ;
  assign n19916 = n18584 & ~n19915 ;
  assign n19917 = n16499 ^ n3002 ^ n1968 ;
  assign n19918 = ( n1819 & ~n13353 ) | ( n1819 & n19917 ) | ( ~n13353 & n19917 ) ;
  assign n19919 = n9521 ^ n7422 ^ 1'b0 ;
  assign n19920 = ~n13219 & n19919 ;
  assign n19921 = n2215 & n19920 ;
  assign n19922 = ( n505 & ~n5417 ) | ( n505 & n13764 ) | ( ~n5417 & n13764 ) ;
  assign n19923 = n19551 & ~n19922 ;
  assign n19924 = n10668 ^ n7875 ^ n6370 ;
  assign n19925 = ( ~n18212 & n19838 ) | ( ~n18212 & n19924 ) | ( n19838 & n19924 ) ;
  assign n19926 = n19925 ^ n14901 ^ n1456 ;
  assign n19927 = n15458 & n19149 ;
  assign n19928 = n15661 & n19927 ;
  assign n19929 = ( n596 & n4741 ) | ( n596 & n11094 ) | ( n4741 & n11094 ) ;
  assign n19930 = n2671 | n19929 ;
  assign n19931 = ( n3984 & ~n4630 ) | ( n3984 & n4854 ) | ( ~n4630 & n4854 ) ;
  assign n19932 = n6159 & ~n19931 ;
  assign n19933 = n19932 ^ n4891 ^ 1'b0 ;
  assign n19935 = n6330 & n8997 ;
  assign n19934 = n16919 ^ n5263 ^ 1'b0 ;
  assign n19936 = n19935 ^ n19934 ^ 1'b0 ;
  assign n19937 = ~n6287 & n8011 ;
  assign n19938 = ~n628 & n661 ;
  assign n19939 = n19938 ^ n11826 ^ 1'b0 ;
  assign n19940 = n19937 & n19939 ;
  assign n19941 = ( ~n12631 & n18293 ) | ( ~n12631 & n19940 ) | ( n18293 & n19940 ) ;
  assign n19942 = n692 | n17422 ;
  assign n19943 = n7076 ^ n2906 ^ 1'b0 ;
  assign n19944 = n16765 & ~n19943 ;
  assign n19945 = n17312 ^ n11030 ^ 1'b0 ;
  assign n19946 = n19944 & n19945 ;
  assign n19947 = n19946 ^ n2593 ^ 1'b0 ;
  assign n19948 = n3174 & ~n4390 ;
  assign n19949 = n6750 & ~n19723 ;
  assign n19950 = n14788 ^ n3864 ^ n2480 ;
  assign n19951 = n19950 ^ n12104 ^ 1'b0 ;
  assign n19952 = n11007 & n19951 ;
  assign n19953 = n1510 | n1574 ;
  assign n19954 = ( ~n2501 & n7968 ) | ( ~n2501 & n14190 ) | ( n7968 & n14190 ) ;
  assign n19955 = ( n10535 & ~n19953 ) | ( n10535 & n19954 ) | ( ~n19953 & n19954 ) ;
  assign n19956 = n12680 ^ n12425 ^ n1590 ;
  assign n19957 = n3272 | n19956 ;
  assign n19958 = n19955 & ~n19957 ;
  assign n19959 = n9860 ^ n1794 ^ 1'b0 ;
  assign n19960 = n19959 ^ n4482 ^ 1'b0 ;
  assign n19961 = n5463 | n11453 ;
  assign n19962 = n19961 ^ n1921 ^ 1'b0 ;
  assign n19963 = n12800 ^ n3074 ^ 1'b0 ;
  assign n19964 = n19962 | n19963 ;
  assign n19965 = n10174 | n19964 ;
  assign n19966 = n19965 ^ n2541 ^ 1'b0 ;
  assign n19967 = n15924 ^ n2150 ^ n422 ;
  assign n19968 = ~n2682 & n19967 ;
  assign n19969 = ( n13216 & ~n19966 ) | ( n13216 & n19968 ) | ( ~n19966 & n19968 ) ;
  assign n19970 = n3181 ^ n248 ^ 1'b0 ;
  assign n19971 = n4834 & ~n19970 ;
  assign n19972 = n19971 ^ n6586 ^ 1'b0 ;
  assign n19973 = n5639 & ~n10748 ;
  assign n19974 = n19973 ^ n10963 ^ 1'b0 ;
  assign n19975 = n8658 ^ n7505 ^ n6109 ;
  assign n19976 = n14858 ^ n1478 ^ 1'b0 ;
  assign n19977 = ( n458 & n6684 ) | ( n458 & n11105 ) | ( n6684 & n11105 ) ;
  assign n19978 = n17633 ^ n12269 ^ n1541 ;
  assign n19979 = n14711 & n19978 ;
  assign n19980 = ~n7014 & n19979 ;
  assign n19981 = x44 & ~n3694 ;
  assign n19982 = n19981 ^ n14497 ^ 1'b0 ;
  assign n19983 = x74 & ~n5369 ;
  assign n19984 = n19934 & n19983 ;
  assign n19985 = n1541 & ~n7516 ;
  assign n19986 = n7343 & n19985 ;
  assign n19987 = n9841 & n19986 ;
  assign n19989 = n9937 ^ n8960 ^ 1'b0 ;
  assign n19990 = n1843 & ~n19989 ;
  assign n19988 = ~n1533 & n6839 ;
  assign n19991 = n19990 ^ n19988 ^ 1'b0 ;
  assign n19992 = n19991 ^ n11206 ^ 1'b0 ;
  assign n19993 = ~n11362 & n19992 ;
  assign n19994 = n19993 ^ n14904 ^ n13705 ;
  assign n19995 = n19271 ^ n15150 ^ 1'b0 ;
  assign n19996 = ( n926 & ~n1120 ) | ( n926 & n5219 ) | ( ~n1120 & n5219 ) ;
  assign n19997 = n196 | n9971 ;
  assign n19998 = n19997 ^ n776 ^ 1'b0 ;
  assign n19999 = ( n3524 & ~n19996 ) | ( n3524 & n19998 ) | ( ~n19996 & n19998 ) ;
  assign n20000 = n19999 ^ n13223 ^ x118 ;
  assign n20004 = ~n477 & n1016 ;
  assign n20005 = n20004 ^ n4307 ^ 1'b0 ;
  assign n20001 = n3617 ^ n2689 ^ 1'b0 ;
  assign n20002 = n2114 | n20001 ;
  assign n20003 = n16142 | n20002 ;
  assign n20006 = n20005 ^ n20003 ^ 1'b0 ;
  assign n20007 = n13467 ^ n1558 ^ 1'b0 ;
  assign n20008 = n5351 & n17602 ;
  assign n20009 = ~n1678 & n20008 ;
  assign n20010 = n20009 ^ n13714 ^ n2162 ;
  assign n20011 = ~n260 & n1781 ;
  assign n20012 = n6752 | n18607 ;
  assign n20013 = n14822 & ~n20012 ;
  assign n20023 = n11791 ^ n9316 ^ 1'b0 ;
  assign n20024 = n1643 & n20023 ;
  assign n20025 = ( ~n2398 & n13337 ) | ( ~n2398 & n20024 ) | ( n13337 & n20024 ) ;
  assign n20014 = n4630 & ~n9001 ;
  assign n20015 = n6616 & n20014 ;
  assign n20016 = n852 & ~n16778 ;
  assign n20017 = n850 | n11651 ;
  assign n20018 = n20017 ^ n12437 ^ 1'b0 ;
  assign n20019 = n20016 | n20018 ;
  assign n20020 = n20015 & ~n20019 ;
  assign n20021 = ~n4421 & n6382 ;
  assign n20022 = n20020 & n20021 ;
  assign n20026 = n20025 ^ n20022 ^ n6331 ;
  assign n20027 = n1052 & ~n17541 ;
  assign n20028 = ~n9582 & n20027 ;
  assign n20029 = ( n17189 & n17283 ) | ( n17189 & n20028 ) | ( n17283 & n20028 ) ;
  assign n20030 = ( x77 & ~n1346 ) | ( x77 & n4349 ) | ( ~n1346 & n4349 ) ;
  assign n20031 = n20030 ^ n1292 ^ 1'b0 ;
  assign n20032 = n842 & ~n20031 ;
  assign n20033 = n4858 & n8109 ;
  assign n20034 = ( n5114 & ~n9964 ) | ( n5114 & n20033 ) | ( ~n9964 & n20033 ) ;
  assign n20035 = n20034 ^ n6940 ^ 1'b0 ;
  assign n20036 = n2637 & ~n7524 ;
  assign n20037 = n16581 & n18349 ;
  assign n20038 = ~n8708 & n20037 ;
  assign n20039 = ( n5512 & ~n19452 ) | ( n5512 & n20038 ) | ( ~n19452 & n20038 ) ;
  assign n20041 = ~n6485 & n11964 ;
  assign n20042 = n20041 ^ x99 ^ 1'b0 ;
  assign n20043 = ~n5616 & n14812 ;
  assign n20044 = n20043 ^ n1996 ^ 1'b0 ;
  assign n20045 = n20042 | n20044 ;
  assign n20046 = ( n9740 & n14619 ) | ( n9740 & n20045 ) | ( n14619 & n20045 ) ;
  assign n20040 = ( n5073 & n14575 ) | ( n5073 & n17578 ) | ( n14575 & n17578 ) ;
  assign n20047 = n20046 ^ n20040 ^ n2660 ;
  assign n20048 = n6818 ^ n1853 ^ 1'b0 ;
  assign n20049 = n10828 & ~n20048 ;
  assign n20050 = n8493 ^ n3364 ^ 1'b0 ;
  assign n20051 = n9067 & ~n20050 ;
  assign n20052 = ~n3803 & n20051 ;
  assign n20053 = ~n2883 & n20052 ;
  assign n20054 = ( n3766 & n6261 ) | ( n3766 & n6702 ) | ( n6261 & n6702 ) ;
  assign n20055 = n20054 ^ n7913 ^ 1'b0 ;
  assign n20056 = n8626 & ~n20055 ;
  assign n20057 = n19507 ^ n12522 ^ 1'b0 ;
  assign n20058 = n20057 ^ n3189 ^ 1'b0 ;
  assign n20059 = n20056 & n20058 ;
  assign n20060 = ( ~n2359 & n20053 ) | ( ~n2359 & n20059 ) | ( n20053 & n20059 ) ;
  assign n20061 = n16441 ^ n8073 ^ 1'b0 ;
  assign n20062 = n20060 & ~n20061 ;
  assign n20063 = n4341 & n12642 ;
  assign n20064 = ( n2626 & n4819 ) | ( n2626 & ~n11452 ) | ( n4819 & ~n11452 ) ;
  assign n20065 = ( n2402 & n10190 ) | ( n2402 & ~n20064 ) | ( n10190 & ~n20064 ) ;
  assign n20066 = n12457 ^ n3546 ^ 1'b0 ;
  assign n20067 = n20066 ^ n8702 ^ n8073 ;
  assign n20068 = n20067 ^ n14514 ^ 1'b0 ;
  assign n20069 = ( n11701 & ~n20065 ) | ( n11701 & n20068 ) | ( ~n20065 & n20068 ) ;
  assign n20070 = n6163 ^ n5682 ^ 1'b0 ;
  assign n20071 = n1743 & n20070 ;
  assign n20072 = n17024 ^ x32 ^ 1'b0 ;
  assign n20073 = n9092 ^ n4334 ^ n2937 ;
  assign n20074 = n11027 | n19238 ;
  assign n20075 = n16215 & n20074 ;
  assign n20076 = ~n20073 & n20075 ;
  assign n20077 = ( n20071 & ~n20072 ) | ( n20071 & n20076 ) | ( ~n20072 & n20076 ) ;
  assign n20078 = ( n2802 & n7015 ) | ( n2802 & ~n11117 ) | ( n7015 & ~n11117 ) ;
  assign n20079 = n1234 | n20078 ;
  assign n20080 = n1820 & ~n9132 ;
  assign n20081 = ~n10710 & n20080 ;
  assign n20082 = ~n20079 & n20081 ;
  assign n20083 = ~n9501 & n10803 ;
  assign n20084 = ~n7206 & n20083 ;
  assign n20085 = n1337 & n19762 ;
  assign n20086 = n12971 ^ n5410 ^ 1'b0 ;
  assign n20087 = n20086 ^ n11623 ^ n5618 ;
  assign n20088 = ( ~n1114 & n3986 ) | ( ~n1114 & n20087 ) | ( n3986 & n20087 ) ;
  assign n20089 = n2867 & n20088 ;
  assign n20090 = ( n11312 & ~n14282 ) | ( n11312 & n15149 ) | ( ~n14282 & n15149 ) ;
  assign n20091 = n6461 ^ n1987 ^ 1'b0 ;
  assign n20092 = n6683 | n20091 ;
  assign n20093 = n7053 | n20092 ;
  assign n20094 = n20093 ^ n6410 ^ 1'b0 ;
  assign n20095 = ( n4836 & n10066 ) | ( n4836 & n20094 ) | ( n10066 & n20094 ) ;
  assign n20096 = ( n2564 & n4615 ) | ( n2564 & ~n20095 ) | ( n4615 & ~n20095 ) ;
  assign n20097 = ( ~n11176 & n17831 ) | ( ~n11176 & n20096 ) | ( n17831 & n20096 ) ;
  assign n20098 = ( ~n3816 & n5098 ) | ( ~n3816 & n20097 ) | ( n5098 & n20097 ) ;
  assign n20099 = n13695 ^ n8179 ^ 1'b0 ;
  assign n20100 = n1304 | n20099 ;
  assign n20101 = n4484 & ~n20100 ;
  assign n20102 = n20101 ^ n18005 ^ 1'b0 ;
  assign n20103 = n545 & ~n5479 ;
  assign n20104 = ~n246 & n20103 ;
  assign n20105 = ( n1397 & n10593 ) | ( n1397 & n20104 ) | ( n10593 & n20104 ) ;
  assign n20106 = n14258 & n20105 ;
  assign n20107 = n17875 ^ n7343 ^ 1'b0 ;
  assign n20108 = n8587 ^ n898 ^ n341 ;
  assign n20109 = n17828 ^ n13207 ^ 1'b0 ;
  assign n20110 = n20108 & ~n20109 ;
  assign n20111 = n12245 ^ n7855 ^ 1'b0 ;
  assign n20112 = n4023 | n20111 ;
  assign n20113 = ( ~n647 & n16625 ) | ( ~n647 & n20112 ) | ( n16625 & n20112 ) ;
  assign n20114 = n2222 & n20113 ;
  assign n20115 = n11382 ^ n8441 ^ 1'b0 ;
  assign n20116 = n2134 | n20115 ;
  assign n20117 = n20116 ^ n4400 ^ n486 ;
  assign n20118 = n703 | n4400 ;
  assign n20119 = n6993 | n20118 ;
  assign n20120 = n20119 ^ n18079 ^ n1059 ;
  assign n20121 = ~n2396 & n20120 ;
  assign n20122 = ~n1723 & n18164 ;
  assign n20123 = ( n12992 & n19229 ) | ( n12992 & ~n20122 ) | ( n19229 & ~n20122 ) ;
  assign n20124 = n7188 ^ n5960 ^ 1'b0 ;
  assign n20125 = n2826 ^ n1961 ^ 1'b0 ;
  assign n20126 = n19455 ^ n7928 ^ n227 ;
  assign n20127 = n20126 ^ n13661 ^ 1'b0 ;
  assign n20128 = n4377 & n20127 ;
  assign n20129 = ( n636 & n5679 ) | ( n636 & ~n20128 ) | ( n5679 & ~n20128 ) ;
  assign n20134 = n12752 ^ n10140 ^ n4067 ;
  assign n20130 = n4073 & n4956 ;
  assign n20131 = n3774 | n5806 ;
  assign n20132 = n20130 & ~n20131 ;
  assign n20133 = n18931 & ~n20132 ;
  assign n20135 = n20134 ^ n20133 ^ n2640 ;
  assign n20136 = n14834 ^ n1079 ^ 1'b0 ;
  assign n20137 = ( n1429 & n10854 ) | ( n1429 & ~n20136 ) | ( n10854 & ~n20136 ) ;
  assign n20138 = ( n7289 & ~n10443 ) | ( n7289 & n20137 ) | ( ~n10443 & n20137 ) ;
  assign n20139 = n11314 ^ n7039 ^ 1'b0 ;
  assign n20140 = n7369 | n7484 ;
  assign n20141 = n5173 & ~n20140 ;
  assign n20142 = ~n9910 & n10000 ;
  assign n20143 = n5480 & n18507 ;
  assign n20144 = ~n20142 & n20143 ;
  assign n20145 = n20141 | n20144 ;
  assign n20146 = n8929 | n14026 ;
  assign n20147 = ( n4904 & n14407 ) | ( n4904 & n20146 ) | ( n14407 & n20146 ) ;
  assign n20148 = n20141 ^ n19444 ^ n5237 ;
  assign n20149 = ~n2220 & n9445 ;
  assign n20150 = ~n18689 & n20149 ;
  assign n20151 = n15802 ^ n13047 ^ 1'b0 ;
  assign n20152 = ~n20150 & n20151 ;
  assign n20153 = n13721 & ~n17923 ;
  assign n20154 = ~n20152 & n20153 ;
  assign n20155 = ~n1134 & n9552 ;
  assign n20156 = n15771 ^ n13367 ^ n2820 ;
  assign n20157 = n4197 ^ n3813 ^ n3677 ;
  assign n20158 = ~n4952 & n16521 ;
  assign n20159 = n20158 ^ n13945 ^ n13427 ;
  assign n20160 = n18639 ^ n4811 ^ 1'b0 ;
  assign n20161 = n2131 & n20160 ;
  assign n20162 = ( n1352 & n1683 ) | ( n1352 & ~n20161 ) | ( n1683 & ~n20161 ) ;
  assign n20163 = n20162 ^ n17653 ^ 1'b0 ;
  assign n20164 = ( n2751 & n3913 ) | ( n2751 & n16067 ) | ( n3913 & n16067 ) ;
  assign n20165 = n6034 ^ n1476 ^ 1'b0 ;
  assign n20166 = n2516 & ~n20165 ;
  assign n20167 = ~n12503 & n20166 ;
  assign n20168 = ~n4198 & n20167 ;
  assign n20169 = n3277 & ~n20168 ;
  assign n20170 = n948 & n20169 ;
  assign n20171 = n3369 & n20170 ;
  assign n20172 = n5844 | n20171 ;
  assign n20173 = n20172 ^ n14103 ^ 1'b0 ;
  assign n20174 = n20173 ^ n18736 ^ 1'b0 ;
  assign n20175 = ~n612 & n7810 ;
  assign n20176 = ( n4633 & n7374 ) | ( n4633 & n20175 ) | ( n7374 & n20175 ) ;
  assign n20177 = n20176 ^ n11831 ^ n9757 ;
  assign n20178 = ( ~n4733 & n12463 ) | ( ~n4733 & n20177 ) | ( n12463 & n20177 ) ;
  assign n20179 = n6767 ^ n1720 ^ 1'b0 ;
  assign n20181 = n2271 & n7497 ;
  assign n20180 = n306 & n9919 ;
  assign n20182 = n20181 ^ n20180 ^ 1'b0 ;
  assign n20183 = n20182 ^ n2140 ^ n1681 ;
  assign n20184 = n19501 ^ n7233 ^ 1'b0 ;
  assign n20185 = n7771 & ~n9526 ;
  assign n20186 = ( n1769 & n5547 ) | ( n1769 & n5903 ) | ( n5547 & n5903 ) ;
  assign n20187 = n8758 | n20186 ;
  assign n20188 = n7077 & ~n20187 ;
  assign n20189 = n1348 | n4836 ;
  assign n20190 = n2165 | n20189 ;
  assign n20191 = ( n7883 & n19326 ) | ( n7883 & ~n20190 ) | ( n19326 & ~n20190 ) ;
  assign n20192 = n20191 ^ n14971 ^ n3701 ;
  assign n20193 = ( n20185 & n20188 ) | ( n20185 & n20192 ) | ( n20188 & n20192 ) ;
  assign n20194 = n7062 | n11137 ;
  assign n20195 = n20194 ^ n1481 ^ 1'b0 ;
  assign n20196 = n6976 | n20195 ;
  assign n20197 = n10908 | n13642 ;
  assign n20198 = n20197 ^ n5037 ^ 1'b0 ;
  assign n20199 = n20198 ^ n14721 ^ 1'b0 ;
  assign n20200 = n4684 | n7958 ;
  assign n20201 = n4714 | n20200 ;
  assign n20202 = n20201 ^ n6990 ^ 1'b0 ;
  assign n20203 = n19656 ^ n14391 ^ n3617 ;
  assign n20204 = n19753 ^ n9385 ^ 1'b0 ;
  assign n20205 = n14009 & ~n20204 ;
  assign n20206 = n18763 ^ n11431 ^ 1'b0 ;
  assign n20207 = n13078 | n20206 ;
  assign n20208 = n694 & ~n7762 ;
  assign n20209 = n8749 & n20208 ;
  assign n20210 = ( n5524 & ~n9770 ) | ( n5524 & n16601 ) | ( ~n9770 & n16601 ) ;
  assign n20211 = n11948 ^ n5225 ^ 1'b0 ;
  assign n20212 = n15514 ^ n8748 ^ n1302 ;
  assign n20213 = n12620 ^ n979 ^ 1'b0 ;
  assign n20214 = n6275 & ~n20213 ;
  assign n20215 = ( ~n16168 & n20212 ) | ( ~n16168 & n20214 ) | ( n20212 & n20214 ) ;
  assign n20219 = ( n1628 & n5054 ) | ( n1628 & n11779 ) | ( n5054 & n11779 ) ;
  assign n20216 = ~n806 & n6811 ;
  assign n20217 = n15490 & n20216 ;
  assign n20218 = n4275 & ~n20217 ;
  assign n20220 = n20219 ^ n20218 ^ 1'b0 ;
  assign n20221 = n3410 & ~n19884 ;
  assign n20222 = n6484 & n8346 ;
  assign n20223 = n20222 ^ n19510 ^ n11502 ;
  assign n20224 = ( n5603 & ~n16123 ) | ( n5603 & n20223 ) | ( ~n16123 & n20223 ) ;
  assign n20225 = n6970 ^ n3351 ^ 1'b0 ;
  assign n20226 = ~n8651 & n20225 ;
  assign n20227 = n20226 ^ n5122 ^ n898 ;
  assign n20228 = n752 & n20227 ;
  assign n20229 = ~n8302 & n20228 ;
  assign n20230 = ~n3684 & n3804 ;
  assign n20231 = n1027 & n20230 ;
  assign n20232 = n5349 ^ n196 ^ 1'b0 ;
  assign n20233 = ~n20231 & n20232 ;
  assign n20234 = n7521 ^ n3031 ^ n2115 ;
  assign n20235 = ( n7959 & n20233 ) | ( n7959 & ~n20234 ) | ( n20233 & ~n20234 ) ;
  assign n20236 = n20235 ^ n17673 ^ n319 ;
  assign n20237 = n3575 & ~n14641 ;
  assign n20238 = n20237 ^ n1555 ^ 1'b0 ;
  assign n20239 = n2671 & ~n20238 ;
  assign n20240 = n4956 ^ n1357 ^ 1'b0 ;
  assign n20241 = n6283 & n20240 ;
  assign n20243 = n13325 ^ n7357 ^ n1330 ;
  assign n20242 = n390 & ~n14865 ;
  assign n20244 = n20243 ^ n20242 ^ 1'b0 ;
  assign n20245 = ( n10779 & n18670 ) | ( n10779 & n20244 ) | ( n18670 & n20244 ) ;
  assign n20246 = ( n2356 & n4714 ) | ( n2356 & ~n13997 ) | ( n4714 & ~n13997 ) ;
  assign n20247 = ( ~n328 & n3419 ) | ( ~n328 & n9334 ) | ( n3419 & n9334 ) ;
  assign n20248 = n7300 & ~n20247 ;
  assign n20249 = ( n12008 & n20246 ) | ( n12008 & n20248 ) | ( n20246 & n20248 ) ;
  assign n20250 = n2011 & ~n10291 ;
  assign n20251 = n4917 & n20250 ;
  assign n20252 = n4684 | n20251 ;
  assign n20253 = n7002 | n20252 ;
  assign n20254 = n20253 ^ n2960 ^ 1'b0 ;
  assign n20255 = n20254 ^ n16086 ^ n10195 ;
  assign n20256 = n474 & n973 ;
  assign n20257 = n4714 & n20256 ;
  assign n20258 = n3945 | n13288 ;
  assign n20259 = n20258 ^ n9539 ^ 1'b0 ;
  assign n20260 = n2300 | n6079 ;
  assign n20261 = n339 | n20260 ;
  assign n20262 = n11733 & ~n20261 ;
  assign n20263 = n7415 ^ n6838 ^ n6250 ;
  assign n20264 = ( n9913 & ~n20262 ) | ( n9913 & n20263 ) | ( ~n20262 & n20263 ) ;
  assign n20265 = n20264 ^ n5254 ^ n934 ;
  assign n20266 = n11646 & n20265 ;
  assign n20267 = n3393 & ~n5106 ;
  assign n20268 = n20267 ^ n12489 ^ n6382 ;
  assign n20269 = ~n3915 & n20268 ;
  assign n20270 = n3013 & n20269 ;
  assign n20271 = ~n318 & n5919 ;
  assign n20272 = ( n7317 & n15842 ) | ( n7317 & ~n17284 ) | ( n15842 & ~n17284 ) ;
  assign n20273 = n20271 | n20272 ;
  assign n20274 = ~n1523 & n3494 ;
  assign n20275 = n20274 ^ n7627 ^ 1'b0 ;
  assign n20276 = n20275 ^ n14379 ^ 1'b0 ;
  assign n20277 = n1837 & n10199 ;
  assign n20278 = n14011 & n19304 ;
  assign n20279 = ~n14406 & n20278 ;
  assign n20280 = n373 | n6830 ;
  assign n20281 = n20279 & n20280 ;
  assign n20282 = n20281 ^ n10410 ^ 1'b0 ;
  assign n20283 = n3844 & ~n12911 ;
  assign n20284 = n15723 ^ n9780 ^ 1'b0 ;
  assign n20285 = n14592 | n20284 ;
  assign n20286 = n5759 | n7146 ;
  assign n20287 = n20286 ^ n17227 ^ 1'b0 ;
  assign n20288 = n3324 & n8080 ;
  assign n20289 = n13924 ^ n12633 ^ n2296 ;
  assign n20290 = n16029 ^ n14898 ^ n3970 ;
  assign n20291 = n15155 ^ n3183 ^ 1'b0 ;
  assign n20292 = n3334 | n13898 ;
  assign n20293 = n17054 & ~n20292 ;
  assign n20294 = x81 & ~n17997 ;
  assign n20295 = n1704 | n20294 ;
  assign n20296 = n986 & n4232 ;
  assign n20297 = n20296 ^ n8134 ^ 1'b0 ;
  assign n20298 = ( n3022 & n13903 ) | ( n3022 & ~n20297 ) | ( n13903 & ~n20297 ) ;
  assign n20299 = ( n3365 & n4158 ) | ( n3365 & ~n13266 ) | ( n4158 & ~n13266 ) ;
  assign n20300 = ~n164 & n1223 ;
  assign n20301 = ~n10029 & n20300 ;
  assign n20302 = n9561 & ~n20301 ;
  assign n20303 = n20302 ^ n7784 ^ 1'b0 ;
  assign n20304 = ( n7168 & n10759 ) | ( n7168 & ~n18496 ) | ( n10759 & ~n18496 ) ;
  assign n20305 = ~n1383 & n10997 ;
  assign n20306 = ( n5289 & n12723 ) | ( n5289 & n20305 ) | ( n12723 & n20305 ) ;
  assign n20307 = n2481 ^ n248 ^ 1'b0 ;
  assign n20308 = x18 & n12345 ;
  assign n20309 = ~n20307 & n20308 ;
  assign n20310 = n20309 ^ n7753 ^ n7407 ;
  assign n20311 = n3612 & n5474 ;
  assign n20312 = n2623 ^ n1279 ^ 1'b0 ;
  assign n20313 = n20312 ^ n7710 ^ 1'b0 ;
  assign n20314 = n7306 & ~n20313 ;
  assign n20315 = n14289 ^ n8860 ^ 1'b0 ;
  assign n20316 = ~n18166 & n20315 ;
  assign n20317 = n20316 ^ n2917 ^ 1'b0 ;
  assign n20318 = n16665 ^ n4059 ^ 1'b0 ;
  assign n20319 = n12218 | n20318 ;
  assign n20320 = n334 & ~n3476 ;
  assign n20321 = n1343 & n9473 ;
  assign n20322 = n18149 ^ n13841 ^ n4592 ;
  assign n20323 = ~n20321 & n20322 ;
  assign n20324 = n12625 ^ n365 ^ 1'b0 ;
  assign n20325 = ( n2752 & n3398 ) | ( n2752 & n12449 ) | ( n3398 & n12449 ) ;
  assign n20326 = n20248 & n20325 ;
  assign n20327 = n20305 ^ x18 ^ 1'b0 ;
  assign n20328 = ~n831 & n20327 ;
  assign n20330 = n17695 ^ n3101 ^ 1'b0 ;
  assign n20331 = n5848 & ~n20330 ;
  assign n20329 = ~n1698 & n10391 ;
  assign n20332 = n20331 ^ n20329 ^ 1'b0 ;
  assign n20333 = n8904 | n11928 ;
  assign n20334 = n12543 ^ n9370 ^ 1'b0 ;
  assign n20341 = n9186 ^ n3403 ^ 1'b0 ;
  assign n20340 = n13212 & ~n15404 ;
  assign n20335 = ( ~n992 & n5673 ) | ( ~n992 & n9249 ) | ( n5673 & n9249 ) ;
  assign n20336 = ~n984 & n20335 ;
  assign n20337 = n844 & n20336 ;
  assign n20338 = n13346 ^ n3797 ^ 1'b0 ;
  assign n20339 = n20337 | n20338 ;
  assign n20342 = n20341 ^ n20340 ^ n20339 ;
  assign n20343 = n15053 ^ n7207 ^ n2420 ;
  assign n20344 = n5859 & n20343 ;
  assign n20345 = n4210 | n20344 ;
  assign n20346 = n20345 ^ n10793 ^ 1'b0 ;
  assign n20347 = ~n3569 & n20346 ;
  assign n20348 = n20347 ^ n12287 ^ 1'b0 ;
  assign n20349 = n5807 ^ n689 ^ 1'b0 ;
  assign n20350 = n10289 ^ n9458 ^ n4503 ;
  assign n20351 = n17256 | n20350 ;
  assign n20352 = ~n1876 & n15639 ;
  assign n20353 = ( ~n1218 & n1602 ) | ( ~n1218 & n5543 ) | ( n1602 & n5543 ) ;
  assign n20354 = n680 & ~n20353 ;
  assign n20355 = ~n565 & n20354 ;
  assign n20356 = ~n4543 & n20355 ;
  assign n20357 = n20352 | n20356 ;
  assign n20358 = ~n984 & n9559 ;
  assign n20359 = ~n20357 & n20358 ;
  assign n20360 = n3907 | n9423 ;
  assign n20361 = n12257 | n20360 ;
  assign n20362 = ~n2485 & n3450 ;
  assign n20363 = n20362 ^ n4735 ^ 1'b0 ;
  assign n20364 = n8003 ^ n7606 ^ 1'b0 ;
  assign n20365 = n20364 ^ n14028 ^ n4000 ;
  assign n20366 = n6311 | n11997 ;
  assign n20367 = n14522 & ~n20366 ;
  assign n20368 = ( n2199 & ~n4269 ) | ( n2199 & n20367 ) | ( ~n4269 & n20367 ) ;
  assign n20369 = n20368 ^ n3063 ^ 1'b0 ;
  assign n20370 = n11925 & ~n20369 ;
  assign n20372 = n5800 ^ n4073 ^ 1'b0 ;
  assign n20373 = n7508 | n20372 ;
  assign n20371 = n9513 | n11040 ;
  assign n20374 = n20373 ^ n20371 ^ 1'b0 ;
  assign n20375 = n14094 ^ n714 ^ 1'b0 ;
  assign n20376 = n6637 | n20375 ;
  assign n20377 = n20376 ^ n10118 ^ n1940 ;
  assign n20378 = ~n565 & n20377 ;
  assign n20379 = n20374 & n20378 ;
  assign n20380 = ( n10202 & n13605 ) | ( n10202 & ~n19177 ) | ( n13605 & ~n19177 ) ;
  assign n20381 = n20380 ^ n9609 ^ n7460 ;
  assign n20382 = n19074 ^ n9842 ^ 1'b0 ;
  assign n20385 = ( ~n2561 & n12936 ) | ( ~n2561 & n19937 ) | ( n12936 & n19937 ) ;
  assign n20383 = n6092 | n6954 ;
  assign n20384 = n2138 | n20383 ;
  assign n20386 = n20385 ^ n20384 ^ n9065 ;
  assign n20387 = ( ~n5301 & n20382 ) | ( ~n5301 & n20386 ) | ( n20382 & n20386 ) ;
  assign n20388 = n8603 ^ n8214 ^ 1'b0 ;
  assign n20389 = ~n14354 & n20388 ;
  assign n20390 = n17530 | n18503 ;
  assign n20391 = ( n2616 & n8029 ) | ( n2616 & n8752 ) | ( n8029 & n8752 ) ;
  assign n20392 = ( n2785 & ~n8297 ) | ( n2785 & n15490 ) | ( ~n8297 & n15490 ) ;
  assign n20393 = n10236 | n20392 ;
  assign n20394 = ( ~n2870 & n11963 ) | ( ~n2870 & n20393 ) | ( n11963 & n20393 ) ;
  assign n20395 = n19840 & n20394 ;
  assign n20396 = ~n20391 & n20395 ;
  assign n20397 = n2295 | n13744 ;
  assign n20398 = n15770 | n20397 ;
  assign n20399 = n17019 ^ n1125 ^ 1'b0 ;
  assign n20400 = n9011 ^ n4491 ^ n4192 ;
  assign n20401 = ( n703 & ~n10898 ) | ( n703 & n15344 ) | ( ~n10898 & n15344 ) ;
  assign n20402 = n6770 & ~n20401 ;
  assign n20403 = ( ~n3497 & n4477 ) | ( ~n3497 & n20402 ) | ( n4477 & n20402 ) ;
  assign n20404 = n17682 ^ n4644 ^ n2600 ;
  assign n20405 = n8116 | n12005 ;
  assign n20406 = ( n356 & n11427 ) | ( n356 & n20405 ) | ( n11427 & n20405 ) ;
  assign n20408 = n10820 | n11722 ;
  assign n20407 = n3710 & n7574 ;
  assign n20409 = n20408 ^ n20407 ^ 1'b0 ;
  assign n20410 = n9160 ^ n8283 ^ n6392 ;
  assign n20411 = n20409 & ~n20410 ;
  assign n20412 = n6908 & ~n8777 ;
  assign n20413 = ( n1716 & n1774 ) | ( n1716 & ~n7022 ) | ( n1774 & ~n7022 ) ;
  assign n20414 = n16690 ^ n13022 ^ n11381 ;
  assign n20415 = n5078 ^ n2906 ^ 1'b0 ;
  assign n20416 = n3624 | n20415 ;
  assign n20417 = n20416 ^ n7986 ^ 1'b0 ;
  assign n20418 = n5041 | n12108 ;
  assign n20419 = ( n1203 & n20417 ) | ( n1203 & ~n20418 ) | ( n20417 & ~n20418 ) ;
  assign n20420 = n3049 & n14794 ;
  assign n20421 = n20420 ^ n9096 ^ 1'b0 ;
  assign n20422 = n3968 & n9306 ;
  assign n20423 = n20422 ^ n2511 ^ 1'b0 ;
  assign n20424 = ~n951 & n2476 ;
  assign n20425 = n18187 ^ n14389 ^ n10240 ;
  assign n20426 = n20425 ^ n12875 ^ n11665 ;
  assign n20427 = ~n2326 & n14650 ;
  assign n20428 = ( n1157 & ~n2782 ) | ( n1157 & n2799 ) | ( ~n2782 & n2799 ) ;
  assign n20429 = n2660 ^ n1550 ^ n525 ;
  assign n20430 = n20429 ^ n15212 ^ 1'b0 ;
  assign n20431 = n20428 & n20430 ;
  assign n20432 = n6075 & n10537 ;
  assign n20433 = n10642 & n20432 ;
  assign n20434 = n3194 | n4955 ;
  assign n20435 = ( n10763 & ~n11374 ) | ( n10763 & n20434 ) | ( ~n11374 & n20434 ) ;
  assign n20436 = n20435 ^ n19506 ^ 1'b0 ;
  assign n20437 = n11599 & ~n20436 ;
  assign n20438 = n20433 & n20437 ;
  assign n20439 = n20438 ^ n15677 ^ n8931 ;
  assign n20440 = n11258 & n13120 ;
  assign n20441 = n20440 ^ n12589 ^ 1'b0 ;
  assign n20442 = n19586 ^ n5449 ^ 1'b0 ;
  assign n20443 = ~n20441 & n20442 ;
  assign n20444 = ( ~n1798 & n2675 ) | ( ~n1798 & n14100 ) | ( n2675 & n14100 ) ;
  assign n20445 = n2774 & n6040 ;
  assign n20446 = n20444 & n20445 ;
  assign n20447 = n19884 ^ n4642 ^ 1'b0 ;
  assign n20448 = ( n2029 & ~n8258 ) | ( n2029 & n17652 ) | ( ~n8258 & n17652 ) ;
  assign n20451 = ~n3879 & n7701 ;
  assign n20452 = ~n1548 & n20451 ;
  assign n20449 = n18712 ^ n10678 ^ n8105 ;
  assign n20450 = ( n2726 & ~n10240 ) | ( n2726 & n20449 ) | ( ~n10240 & n20449 ) ;
  assign n20453 = n20452 ^ n20450 ^ n18829 ;
  assign n20454 = n19858 ^ n1212 ^ 1'b0 ;
  assign n20455 = n15406 ^ n4862 ^ 1'b0 ;
  assign n20456 = n15667 & n20455 ;
  assign n20457 = n1160 & ~n2156 ;
  assign n20458 = n7113 & n20457 ;
  assign n20459 = n20458 ^ n6168 ^ 1'b0 ;
  assign n20460 = n6628 ^ n3322 ^ 1'b0 ;
  assign n20461 = n675 & n4357 ;
  assign n20462 = ~n20460 & n20461 ;
  assign n20463 = n20462 ^ n14630 ^ 1'b0 ;
  assign n20464 = n20463 ^ n8712 ^ n2114 ;
  assign n20465 = n9230 & n20464 ;
  assign n20466 = n20465 ^ n19954 ^ 1'b0 ;
  assign n20467 = n1357 | n6974 ;
  assign n20468 = n20467 ^ n2817 ^ n2399 ;
  assign n20469 = ~n19095 & n20468 ;
  assign n20470 = n9146 ^ n5050 ^ n4964 ;
  assign n20471 = n20470 ^ n9824 ^ 1'b0 ;
  assign n20472 = n9958 & n19429 ;
  assign n20473 = n517 | n20472 ;
  assign n20474 = ~n7353 & n10205 ;
  assign n20475 = ~n3457 & n20474 ;
  assign n20476 = n5814 ^ n5461 ^ 1'b0 ;
  assign n20477 = ~n465 & n17775 ;
  assign n20478 = n20476 & n20477 ;
  assign n20479 = n6267 ^ n4530 ^ 1'b0 ;
  assign n20480 = n18479 & ~n20479 ;
  assign n20481 = ~n18633 & n20480 ;
  assign n20482 = ~n10494 & n17456 ;
  assign n20483 = n3694 & n20482 ;
  assign n20484 = n17575 ^ n11685 ^ n1350 ;
  assign n20485 = ( n1041 & n2353 ) | ( n1041 & n7776 ) | ( n2353 & n7776 ) ;
  assign n20486 = ~n20484 & n20485 ;
  assign n20487 = ( n1851 & n3790 ) | ( n1851 & n20486 ) | ( n3790 & n20486 ) ;
  assign n20488 = n1952 & ~n3630 ;
  assign n20489 = n20488 ^ n18133 ^ n1114 ;
  assign n20490 = n9669 ^ n1571 ^ n1349 ;
  assign n20491 = n15924 ^ n8601 ^ 1'b0 ;
  assign n20492 = ~n5616 & n20491 ;
  assign n20493 = ( n3384 & n20490 ) | ( n3384 & ~n20492 ) | ( n20490 & ~n20492 ) ;
  assign n20494 = n15103 ^ n4105 ^ 1'b0 ;
  assign n20495 = n20494 ^ n13052 ^ 1'b0 ;
  assign n20496 = n16621 & ~n20495 ;
  assign n20497 = ~n466 & n620 ;
  assign n20498 = n14340 & ~n14342 ;
  assign n20499 = ~n949 & n20498 ;
  assign n20500 = ( n12361 & ~n12691 ) | ( n12361 & n20499 ) | ( ~n12691 & n20499 ) ;
  assign n20501 = n2831 & ~n19609 ;
  assign n20502 = ~n1213 & n20501 ;
  assign n20507 = n11004 ^ n8000 ^ 1'b0 ;
  assign n20503 = n18238 ^ n196 ^ 1'b0 ;
  assign n20504 = n16895 & n20503 ;
  assign n20505 = n5144 & n20504 ;
  assign n20506 = ~n11626 & n20505 ;
  assign n20508 = n20507 ^ n20506 ^ 1'b0 ;
  assign n20509 = ~n12185 & n20508 ;
  assign n20510 = n3131 | n8212 ;
  assign n20511 = n20510 ^ n3441 ^ 1'b0 ;
  assign n20512 = ~n403 & n20511 ;
  assign n20513 = n20512 ^ n13493 ^ 1'b0 ;
  assign n20514 = n16697 ^ n11371 ^ 1'b0 ;
  assign n20515 = n1194 & n20514 ;
  assign n20516 = n1769 | n9539 ;
  assign n20517 = n12975 | n20516 ;
  assign n20518 = ( n4164 & ~n4957 ) | ( n4164 & n20517 ) | ( ~n4957 & n20517 ) ;
  assign n20520 = n8240 ^ n4500 ^ 1'b0 ;
  assign n20521 = n3796 & n20520 ;
  assign n20519 = n1385 & ~n4461 ;
  assign n20522 = n20521 ^ n20519 ^ n2929 ;
  assign n20523 = n1646 ^ x74 ^ 1'b0 ;
  assign n20524 = n5743 & n20523 ;
  assign n20525 = n20524 ^ n8437 ^ n8079 ;
  assign n20526 = n11927 ^ n5495 ^ 1'b0 ;
  assign n20527 = n10238 | n20526 ;
  assign n20528 = n20527 ^ n6899 ^ 1'b0 ;
  assign n20529 = n20525 | n20528 ;
  assign n20530 = n1410 | n10642 ;
  assign n20531 = n14393 & ~n20530 ;
  assign n20532 = n6109 & n20531 ;
  assign n20533 = ~n3538 & n14432 ;
  assign n20534 = n6752 & n20533 ;
  assign n20535 = n1070 | n20534 ;
  assign n20536 = ~n847 & n5745 ;
  assign n20537 = n20536 ^ n19326 ^ n6968 ;
  assign n20538 = n12599 ^ n2770 ^ 1'b0 ;
  assign n20539 = n20538 ^ n8074 ^ 1'b0 ;
  assign n20540 = n20537 | n20539 ;
  assign n20541 = n2547 | n16051 ;
  assign n20542 = n20541 ^ n12616 ^ x125 ;
  assign n20543 = n11790 ^ n8859 ^ 1'b0 ;
  assign n20545 = n8776 ^ n1018 ^ 1'b0 ;
  assign n20546 = n1894 & ~n2147 ;
  assign n20547 = ~n20545 & n20546 ;
  assign n20544 = ~n4004 & n5732 ;
  assign n20548 = n20547 ^ n20544 ^ 1'b0 ;
  assign n20549 = ( n20357 & n20543 ) | ( n20357 & ~n20548 ) | ( n20543 & ~n20548 ) ;
  assign n20551 = n9662 ^ n6451 ^ 1'b0 ;
  assign n20552 = n8309 & ~n20551 ;
  assign n20550 = n16971 & ~n20116 ;
  assign n20553 = n20552 ^ n20550 ^ 1'b0 ;
  assign n20554 = n5728 & n7727 ;
  assign n20555 = ~n12046 & n20554 ;
  assign n20556 = n19751 ^ n12812 ^ x19 ;
  assign n20557 = ~n2106 & n20556 ;
  assign n20558 = n19732 ^ n11341 ^ 1'b0 ;
  assign n20559 = n10364 & ~n11531 ;
  assign n20560 = n6495 & n20559 ;
  assign n20561 = n1973 ^ n612 ^ 1'b0 ;
  assign n20562 = n14381 & n20561 ;
  assign n20563 = n20562 ^ n371 ^ 1'b0 ;
  assign n20564 = ( n4743 & ~n16673 ) | ( n4743 & n20563 ) | ( ~n16673 & n20563 ) ;
  assign n20565 = n20564 ^ n13400 ^ 1'b0 ;
  assign n20566 = ~n20560 & n20565 ;
  assign n20567 = n4028 ^ n812 ^ 1'b0 ;
  assign n20568 = n7536 & n20567 ;
  assign n20569 = ~n20566 & n20568 ;
  assign n20570 = ~x112 & n4811 ;
  assign n20571 = ~n10529 & n20570 ;
  assign n20572 = n2945 & n20571 ;
  assign n20573 = n20572 ^ n12752 ^ n2006 ;
  assign n20574 = n6101 ^ n3232 ^ 1'b0 ;
  assign n20575 = ~n2025 & n20574 ;
  assign n20576 = n20575 ^ n3952 ^ 1'b0 ;
  assign n20577 = n18063 ^ n5963 ^ 1'b0 ;
  assign n20578 = n19835 ^ n7407 ^ 1'b0 ;
  assign n20579 = n7219 ^ n6105 ^ 1'b0 ;
  assign n20584 = n2744 & n2842 ;
  assign n20585 = n20584 ^ n2740 ^ 1'b0 ;
  assign n20583 = n14673 & ~n16154 ;
  assign n20586 = n20585 ^ n20583 ^ 1'b0 ;
  assign n20587 = ~n1761 & n20586 ;
  assign n20580 = n6892 & n8298 ;
  assign n20581 = n20580 ^ n8255 ^ 1'b0 ;
  assign n20582 = n20581 ^ n1896 ^ n1274 ;
  assign n20588 = n20587 ^ n20582 ^ n2884 ;
  assign n20589 = ~n162 & n2547 ;
  assign n20590 = n5277 & n20589 ;
  assign n20591 = ~n6199 & n20590 ;
  assign n20592 = ( n3095 & n3631 ) | ( n3095 & n20591 ) | ( n3631 & n20591 ) ;
  assign n20593 = ~n727 & n7819 ;
  assign n20594 = ~n16730 & n20593 ;
  assign n20596 = n1894 & n10127 ;
  assign n20597 = ~n3394 & n20596 ;
  assign n20598 = n20597 ^ n14235 ^ n3756 ;
  assign n20595 = n2223 & n5928 ;
  assign n20599 = n20598 ^ n20595 ^ 1'b0 ;
  assign n20600 = n14755 ^ n9984 ^ 1'b0 ;
  assign n20601 = n9804 & n20600 ;
  assign n20602 = ~n16751 & n20601 ;
  assign n20604 = n4867 & n20562 ;
  assign n20603 = n3120 | n6026 ;
  assign n20605 = n20604 ^ n20603 ^ n6392 ;
  assign n20606 = n6235 | n11421 ;
  assign n20607 = n20606 ^ n13885 ^ 1'b0 ;
  assign n20610 = n9913 ^ n2413 ^ 1'b0 ;
  assign n20609 = n7469 & n7972 ;
  assign n20611 = n20610 ^ n20609 ^ 1'b0 ;
  assign n20612 = n2513 & n20611 ;
  assign n20608 = ( n3254 & n5502 ) | ( n3254 & ~n7999 ) | ( n5502 & ~n7999 ) ;
  assign n20613 = n20612 ^ n20608 ^ 1'b0 ;
  assign n20614 = n20613 ^ n4325 ^ 1'b0 ;
  assign n20615 = n20607 & ~n20614 ;
  assign n20616 = ( ~n9081 & n20605 ) | ( ~n9081 & n20615 ) | ( n20605 & n20615 ) ;
  assign n20617 = n20616 ^ n5632 ^ 1'b0 ;
  assign n20618 = ( n3617 & n6557 ) | ( n3617 & n16954 ) | ( n6557 & n16954 ) ;
  assign n20619 = ( n3146 & ~n12916 ) | ( n3146 & n20618 ) | ( ~n12916 & n20618 ) ;
  assign n20620 = n14257 ^ n7104 ^ 1'b0 ;
  assign n20621 = ~n6867 & n7396 ;
  assign n20622 = n7392 & n20621 ;
  assign n20623 = n20136 ^ n11722 ^ n3500 ;
  assign n20624 = n20538 | n20623 ;
  assign n20625 = n19131 ^ n10986 ^ n3403 ;
  assign n20626 = n20625 ^ n1530 ^ 1'b0 ;
  assign n20627 = ~n13823 & n17918 ;
  assign n20628 = n8130 | n11138 ;
  assign n20629 = ( n4055 & n10346 ) | ( n4055 & ~n15517 ) | ( n10346 & ~n15517 ) ;
  assign n20630 = n20629 ^ n4727 ^ 1'b0 ;
  assign n20631 = n4630 & n20630 ;
  assign n20632 = n6010 & n6231 ;
  assign n20633 = n1546 & n9914 ;
  assign n20634 = n10178 | n20633 ;
  assign n20635 = n20634 ^ n11319 ^ 1'b0 ;
  assign n20636 = n18268 ^ n5566 ^ 1'b0 ;
  assign n20637 = n8699 | n20636 ;
  assign n20638 = n20637 ^ n7701 ^ 1'b0 ;
  assign n20639 = n7244 | n15295 ;
  assign n20640 = ( n2331 & n8451 ) | ( n2331 & ~n20639 ) | ( n8451 & ~n20639 ) ;
  assign n20641 = ~n6085 & n12346 ;
  assign n20642 = n20641 ^ n5899 ^ n5248 ;
  assign n20643 = ( n1431 & n19277 ) | ( n1431 & ~n20228 ) | ( n19277 & ~n20228 ) ;
  assign n20644 = n7132 ^ n399 ^ 1'b0 ;
  assign n20645 = n4508 | n20644 ;
  assign n20646 = n20645 ^ n1226 ^ 1'b0 ;
  assign n20647 = n7617 | n20646 ;
  assign n20648 = ( n771 & n6374 ) | ( n771 & ~n8076 ) | ( n6374 & ~n8076 ) ;
  assign n20649 = ( n8238 & ~n10957 ) | ( n8238 & n20648 ) | ( ~n10957 & n20648 ) ;
  assign n20650 = n17626 ^ n213 ^ 1'b0 ;
  assign n20651 = n8163 ^ n6607 ^ 1'b0 ;
  assign n20652 = n13194 & n20651 ;
  assign n20653 = n20652 ^ n19858 ^ n2295 ;
  assign n20654 = ( n4391 & ~n7152 ) | ( n4391 & n16027 ) | ( ~n7152 & n16027 ) ;
  assign n20655 = ~n8685 & n17142 ;
  assign n20656 = n11737 ^ n8541 ^ n5495 ;
  assign n20657 = n20656 ^ n17941 ^ n15736 ;
  assign n20658 = n20657 ^ n1650 ^ 1'b0 ;
  assign n20659 = n8915 | n20658 ;
  assign n20660 = n819 & ~n7354 ;
  assign n20661 = n4100 | n16891 ;
  assign n20662 = n10765 ^ n10258 ^ 1'b0 ;
  assign n20665 = n439 & n4407 ;
  assign n20664 = n8025 ^ n643 ^ 1'b0 ;
  assign n20663 = n5011 ^ n4392 ^ x108 ;
  assign n20666 = n20665 ^ n20664 ^ n20663 ;
  assign n20667 = n2773 ^ x25 ^ 1'b0 ;
  assign n20668 = n20667 ^ n18029 ^ n320 ;
  assign n20669 = ~n12256 & n14292 ;
  assign n20670 = n15176 & n20669 ;
  assign n20671 = n20670 ^ n10880 ^ n1137 ;
  assign n20672 = n1198 & ~n9521 ;
  assign n20673 = n20672 ^ n8643 ^ 1'b0 ;
  assign n20674 = n7490 | n13201 ;
  assign n20675 = n12468 & ~n20674 ;
  assign n20676 = ( n2447 & n14271 ) | ( n2447 & n16810 ) | ( n14271 & n16810 ) ;
  assign n20677 = n20676 ^ n3894 ^ 1'b0 ;
  assign n20678 = ~n7366 & n20677 ;
  assign n20679 = n2165 | n14198 ;
  assign n20680 = n16356 ^ n6446 ^ x57 ;
  assign n20681 = n1329 & ~n13832 ;
  assign n20682 = n8882 | n13890 ;
  assign n20683 = n2652 & ~n7492 ;
  assign n20684 = n2712 | n20683 ;
  assign n20685 = ~n11572 & n20684 ;
  assign n20687 = ( ~n8411 & n10368 ) | ( ~n8411 & n16611 ) | ( n10368 & n16611 ) ;
  assign n20686 = n3784 & n14601 ;
  assign n20688 = n20687 ^ n20686 ^ 1'b0 ;
  assign n20689 = n3533 | n8634 ;
  assign n20690 = ( n3808 & ~n6376 ) | ( n3808 & n10360 ) | ( ~n6376 & n10360 ) ;
  assign n20691 = n13744 ^ n13580 ^ n4684 ;
  assign n20692 = ( n5890 & n6572 ) | ( n5890 & n16183 ) | ( n6572 & n16183 ) ;
  assign n20693 = n3118 ^ n1832 ^ 1'b0 ;
  assign n20694 = n20692 & n20693 ;
  assign n20695 = n3214 | n17982 ;
  assign n20696 = n20695 ^ n15373 ^ 1'b0 ;
  assign n20697 = n6488 | n7484 ;
  assign n20698 = n3283 & n20697 ;
  assign n20699 = n18665 & n20698 ;
  assign n20700 = ~n4157 & n20656 ;
  assign n20702 = n4313 ^ n1568 ^ 1'b0 ;
  assign n20701 = n13158 ^ n13109 ^ n12489 ;
  assign n20703 = n20702 ^ n20701 ^ n7793 ;
  assign n20704 = n17031 ^ n3267 ^ n2023 ;
  assign n20705 = n20704 ^ n5093 ^ n412 ;
  assign n20706 = ( ~n491 & n1635 ) | ( ~n491 & n12603 ) | ( n1635 & n12603 ) ;
  assign n20707 = n6196 ^ n3477 ^ 1'b0 ;
  assign n20708 = n1805 & ~n20707 ;
  assign n20709 = n3721 & n3738 ;
  assign n20710 = n1901 & n7309 ;
  assign n20711 = n20710 ^ n16251 ^ 1'b0 ;
  assign n20712 = ~n14619 & n20711 ;
  assign n20713 = n14609 ^ n4742 ^ 1'b0 ;
  assign n20714 = n20712 | n20713 ;
  assign n20715 = ( n8334 & ~n20709 ) | ( n8334 & n20714 ) | ( ~n20709 & n20714 ) ;
  assign n20716 = ~n1225 & n5755 ;
  assign n20718 = n5719 ^ n141 ^ 1'b0 ;
  assign n20717 = ~n1990 & n10780 ;
  assign n20719 = n20718 ^ n20717 ^ 1'b0 ;
  assign n20720 = n20716 | n20719 ;
  assign n20721 = n5805 & ~n20720 ;
  assign n20722 = ( ~n12426 & n16091 ) | ( ~n12426 & n20721 ) | ( n16091 & n20721 ) ;
  assign n20723 = n4591 ^ n307 ^ 1'b0 ;
  assign n20724 = n4137 & n20723 ;
  assign n20725 = n12159 ^ n7494 ^ 1'b0 ;
  assign n20726 = ( ~n3595 & n20724 ) | ( ~n3595 & n20725 ) | ( n20724 & n20725 ) ;
  assign n20727 = ( n11272 & ~n15465 ) | ( n11272 & n18059 ) | ( ~n15465 & n18059 ) ;
  assign n20728 = n8610 | n14908 ;
  assign n20729 = n20728 ^ n11335 ^ 1'b0 ;
  assign n20730 = ( n13783 & n20727 ) | ( n13783 & n20729 ) | ( n20727 & n20729 ) ;
  assign n20731 = n16717 ^ n5709 ^ 1'b0 ;
  assign n20732 = n18841 & n19727 ;
  assign n20733 = ~n6847 & n20732 ;
  assign n20734 = ( n11357 & ~n15253 ) | ( n11357 & n20733 ) | ( ~n15253 & n20733 ) ;
  assign n20735 = n4347 | n13511 ;
  assign n20736 = ( n10817 & n12768 ) | ( n10817 & ~n20735 ) | ( n12768 & ~n20735 ) ;
  assign n20737 = n3262 & ~n16220 ;
  assign n20738 = n20737 ^ n11988 ^ 1'b0 ;
  assign n20739 = n8864 ^ n5140 ^ 1'b0 ;
  assign n20740 = n9194 & n20739 ;
  assign n20741 = n16280 ^ n13145 ^ n12522 ;
  assign n20742 = n10842 ^ n4681 ^ n1339 ;
  assign n20743 = n20742 ^ n7496 ^ n3437 ;
  assign n20744 = n13664 ^ n5461 ^ 1'b0 ;
  assign n20745 = n20560 ^ n18834 ^ x55 ;
  assign n20746 = ( n11984 & ~n20744 ) | ( n11984 & n20745 ) | ( ~n20744 & n20745 ) ;
  assign n20747 = ~n4237 & n10808 ;
  assign n20748 = n20747 ^ n4364 ^ n1681 ;
  assign n20749 = ~n6520 & n9143 ;
  assign n20750 = n20749 ^ n16302 ^ 1'b0 ;
  assign n20751 = n14298 | n14578 ;
  assign n20752 = ( n8280 & n8714 ) | ( n8280 & ~n20639 ) | ( n8714 & ~n20639 ) ;
  assign n20753 = n3003 & n6350 ;
  assign n20754 = n20753 ^ n7314 ^ 1'b0 ;
  assign n20758 = n6053 & n10764 ;
  assign n20756 = ~n1086 & n10548 ;
  assign n20757 = n2167 & n20756 ;
  assign n20759 = n20758 ^ n20757 ^ n18862 ;
  assign n20755 = n856 & ~n19086 ;
  assign n20760 = n20759 ^ n20755 ^ 1'b0 ;
  assign n20761 = n4441 & n13971 ;
  assign n20762 = ~n9102 & n20761 ;
  assign n20763 = ( n2222 & n3354 ) | ( n2222 & n3955 ) | ( n3354 & n3955 ) ;
  assign n20764 = n11122 ^ n2136 ^ 1'b0 ;
  assign n20765 = n14313 ^ n9220 ^ 1'b0 ;
  assign n20766 = n5525 & ~n20765 ;
  assign n20767 = n20766 ^ n14389 ^ n14069 ;
  assign n20768 = n20764 & n20767 ;
  assign n20769 = n20763 & n20768 ;
  assign n20770 = n18902 ^ n10990 ^ 1'b0 ;
  assign n20771 = n12739 ^ n474 ^ 1'b0 ;
  assign n20772 = n16917 | n17066 ;
  assign n20773 = n863 | n20772 ;
  assign n20774 = n10819 ^ n6988 ^ 1'b0 ;
  assign n20775 = n912 & n9409 ;
  assign n20776 = n20775 ^ n3303 ^ 1'b0 ;
  assign n20777 = n3808 & n10944 ;
  assign n20778 = n20142 & n20777 ;
  assign n20779 = n20344 & n20778 ;
  assign n20780 = n17729 ^ n11270 ^ 1'b0 ;
  assign n20781 = n730 | n20780 ;
  assign n20782 = n442 | n2389 ;
  assign n20783 = n10452 ^ n7071 ^ 1'b0 ;
  assign n20784 = ~n19046 & n20783 ;
  assign n20785 = n20784 ^ n12849 ^ 1'b0 ;
  assign n20786 = n20785 ^ n590 ^ 1'b0 ;
  assign n20787 = n20782 & n20786 ;
  assign n20788 = n18686 ^ n4878 ^ 1'b0 ;
  assign n20789 = n20788 ^ n11368 ^ n4726 ;
  assign n20790 = n18326 ^ n15150 ^ n12668 ;
  assign n20791 = n9869 ^ n8080 ^ 1'b0 ;
  assign n20792 = n1540 | n20181 ;
  assign n20793 = ~n1803 & n2420 ;
  assign n20794 = ~n4180 & n20793 ;
  assign n20799 = n2670 ^ n2165 ^ 1'b0 ;
  assign n20800 = n6611 & ~n20799 ;
  assign n20795 = n6422 ^ n3481 ^ 1'b0 ;
  assign n20796 = n20795 ^ n11650 ^ 1'b0 ;
  assign n20797 = n17420 ^ n815 ^ 1'b0 ;
  assign n20798 = n20796 | n20797 ;
  assign n20801 = n20800 ^ n20798 ^ 1'b0 ;
  assign n20802 = n17677 ^ n10017 ^ 1'b0 ;
  assign n20803 = n16772 ^ n9870 ^ 1'b0 ;
  assign n20804 = n4862 | n5479 ;
  assign n20805 = n10343 & ~n20804 ;
  assign n20806 = n8605 ^ n4417 ^ 1'b0 ;
  assign n20807 = n1027 | n20806 ;
  assign n20808 = ( x13 & n20805 ) | ( x13 & ~n20807 ) | ( n20805 & ~n20807 ) ;
  assign n20809 = ( ~n650 & n2165 ) | ( ~n650 & n6083 ) | ( n2165 & n6083 ) ;
  assign n20810 = ( n1921 & n6598 ) | ( n1921 & ~n20809 ) | ( n6598 & ~n20809 ) ;
  assign n20811 = n20810 ^ n5436 ^ 1'b0 ;
  assign n20812 = n2681 & ~n8890 ;
  assign n20813 = ~n15483 & n20812 ;
  assign n20814 = n20813 ^ n6146 ^ 1'b0 ;
  assign n20815 = n1377 & n7536 ;
  assign n20816 = n15464 & n20815 ;
  assign n20817 = n11746 & n19495 ;
  assign n20818 = ~n2131 & n20817 ;
  assign n20819 = ( n7819 & n8911 ) | ( n7819 & ~n13461 ) | ( n8911 & ~n13461 ) ;
  assign n20820 = ~n17600 & n20819 ;
  assign n20821 = ~n3524 & n20820 ;
  assign n20822 = n3921 & n13594 ;
  assign n20823 = n6838 & ~n20822 ;
  assign n20824 = n12550 | n20823 ;
  assign n20825 = ( n982 & ~n9111 ) | ( n982 & n20824 ) | ( ~n9111 & n20824 ) ;
  assign n20826 = ~n2242 & n2273 ;
  assign n20827 = n13499 ^ n8795 ^ 1'b0 ;
  assign n20828 = n20826 & ~n20827 ;
  assign n20829 = n4815 ^ n4789 ^ n4777 ;
  assign n20830 = n20829 ^ n14185 ^ 1'b0 ;
  assign n20831 = n20828 & ~n20830 ;
  assign n20832 = n4733 & ~n17497 ;
  assign n20833 = ~n9790 & n20832 ;
  assign n20834 = ~n6824 & n15608 ;
  assign n20835 = ( n13965 & ~n19777 ) | ( n13965 & n20834 ) | ( ~n19777 & n20834 ) ;
  assign n20836 = n19890 ^ n19685 ^ 1'b0 ;
  assign n20837 = ~n9155 & n20836 ;
  assign n20838 = n9331 ^ x93 ^ 1'b0 ;
  assign n20839 = ~n6370 & n20838 ;
  assign n20840 = n3666 & ~n5633 ;
  assign n20841 = ~n6008 & n20840 ;
  assign n20842 = ( n12811 & ~n18034 ) | ( n12811 & n20841 ) | ( ~n18034 & n20841 ) ;
  assign n20843 = n20842 ^ n1771 ^ 1'b0 ;
  assign n20846 = n7485 ^ n584 ^ 1'b0 ;
  assign n20847 = n5914 | n20846 ;
  assign n20844 = n17129 ^ n5788 ^ 1'b0 ;
  assign n20845 = n16067 & ~n20844 ;
  assign n20848 = n20847 ^ n20845 ^ n2038 ;
  assign n20849 = n6772 & ~n8117 ;
  assign n20850 = n3333 ^ n146 ^ 1'b0 ;
  assign n20851 = n5873 & n20850 ;
  assign n20852 = n4252 & ~n20851 ;
  assign n20854 = n4433 | n8697 ;
  assign n20855 = n20854 ^ n2112 ^ 1'b0 ;
  assign n20856 = ~n3565 & n20855 ;
  assign n20857 = n14886 & n20856 ;
  assign n20853 = n1867 & ~n16612 ;
  assign n20858 = n20857 ^ n20853 ^ 1'b0 ;
  assign n20859 = n13220 | n15579 ;
  assign n20860 = ~n241 & n14450 ;
  assign n20861 = n855 & n20860 ;
  assign n20862 = n6717 | n20861 ;
  assign n20863 = n714 | n13279 ;
  assign n20864 = n1209 & ~n20863 ;
  assign n20865 = n9024 ^ n8923 ^ n1357 ;
  assign n20866 = ( ~n1617 & n4681 ) | ( ~n1617 & n13642 ) | ( n4681 & n13642 ) ;
  assign n20867 = ( ~x103 & n12510 ) | ( ~x103 & n20866 ) | ( n12510 & n20866 ) ;
  assign n20868 = n10875 | n20867 ;
  assign n20869 = n13817 | n20868 ;
  assign n20875 = ( n265 & n7816 ) | ( n265 & n13043 ) | ( n7816 & n13043 ) ;
  assign n20870 = n13764 ^ n5384 ^ 1'b0 ;
  assign n20871 = n977 | n8623 ;
  assign n20872 = n20871 ^ n6452 ^ n2879 ;
  assign n20873 = n20872 ^ n1974 ^ 1'b0 ;
  assign n20874 = n20870 & n20873 ;
  assign n20876 = n20875 ^ n20874 ^ 1'b0 ;
  assign n20877 = n20876 ^ n7571 ^ n6261 ;
  assign n20878 = ( n20212 & n20869 ) | ( n20212 & ~n20877 ) | ( n20869 & ~n20877 ) ;
  assign n20879 = n659 | n10135 ;
  assign n20880 = n3109 & ~n20879 ;
  assign n20881 = n6888 ^ n4516 ^ 1'b0 ;
  assign n20882 = ~n19568 & n20881 ;
  assign n20883 = n4135 | n14207 ;
  assign n20884 = n6289 ^ n1230 ^ 1'b0 ;
  assign n20885 = ~n13253 & n20884 ;
  assign n20886 = n4869 & n20885 ;
  assign n20887 = n20886 ^ n11442 ^ 1'b0 ;
  assign n20888 = n2184 & ~n20887 ;
  assign n20889 = ~n10991 & n14077 ;
  assign n20890 = ( n17835 & ~n20888 ) | ( n17835 & n20889 ) | ( ~n20888 & n20889 ) ;
  assign n20891 = n9090 ^ n3707 ^ n1611 ;
  assign n20892 = n17219 ^ n7211 ^ n3742 ;
  assign n20893 = ~n1192 & n5960 ;
  assign n20894 = n6890 & n20893 ;
  assign n20895 = n1813 | n20894 ;
  assign n20896 = n9393 & ~n20895 ;
  assign n20897 = n9396 | n19114 ;
  assign n20898 = n14961 & n17093 ;
  assign n20899 = n20898 ^ n10286 ^ n2219 ;
  assign n20900 = n6769 ^ n3508 ^ 1'b0 ;
  assign n20901 = ~n7482 & n20900 ;
  assign n20902 = n20901 ^ n12076 ^ 1'b0 ;
  assign n20903 = n19742 | n20902 ;
  assign n20904 = n3811 ^ x107 ^ 1'b0 ;
  assign n20905 = n20904 ^ n6410 ^ 1'b0 ;
  assign n20906 = ( n20899 & n20903 ) | ( n20899 & ~n20905 ) | ( n20903 & ~n20905 ) ;
  assign n20907 = n4311 ^ n2095 ^ 1'b0 ;
  assign n20908 = n1327 & ~n20907 ;
  assign n20909 = ( ~n8342 & n10846 ) | ( ~n8342 & n20908 ) | ( n10846 & n20908 ) ;
  assign n20910 = n8415 & n10095 ;
  assign n20911 = ( x101 & n12348 ) | ( x101 & ~n17430 ) | ( n12348 & ~n17430 ) ;
  assign n20912 = n8957 ^ n6016 ^ n182 ;
  assign n20913 = ~n550 & n20912 ;
  assign n20914 = n20913 ^ n4465 ^ 1'b0 ;
  assign n20916 = n1282 | n15574 ;
  assign n20917 = n3235 | n20916 ;
  assign n20915 = ~n2763 & n10299 ;
  assign n20918 = n20917 ^ n20915 ^ 1'b0 ;
  assign n20919 = n9473 | n20918 ;
  assign n20920 = ( n8645 & n18810 ) | ( n8645 & n18876 ) | ( n18810 & n18876 ) ;
  assign n20921 = ( n3643 & ~n10092 ) | ( n3643 & n10190 ) | ( ~n10092 & n10190 ) ;
  assign n20922 = n16780 ^ n10213 ^ n6461 ;
  assign n20923 = ( n383 & ~n2816 ) | ( n383 & n6138 ) | ( ~n2816 & n6138 ) ;
  assign n20924 = n8984 ^ n6749 ^ 1'b0 ;
  assign n20925 = ~n20629 & n20924 ;
  assign n20926 = n20925 ^ n8446 ^ 1'b0 ;
  assign n20927 = n20923 | n20926 ;
  assign n20928 = n11505 ^ n10175 ^ 1'b0 ;
  assign n20929 = n10440 & ~n20928 ;
  assign n20930 = n11465 & n20929 ;
  assign n20931 = n20930 ^ n18041 ^ 1'b0 ;
  assign n20932 = n211 | n5681 ;
  assign n20933 = n19656 & ~n20932 ;
  assign n20934 = n8370 ^ n1153 ^ 1'b0 ;
  assign n20935 = ~n11015 & n20934 ;
  assign n20936 = ( ~n6974 & n11820 ) | ( ~n6974 & n20935 ) | ( n11820 & n20935 ) ;
  assign n20940 = ( n7362 & n9910 ) | ( n7362 & ~n15475 ) | ( n9910 & ~n15475 ) ;
  assign n20937 = ~n2869 & n9798 ;
  assign n20938 = n20937 ^ n12963 ^ n8801 ;
  assign n20939 = n8081 | n20938 ;
  assign n20941 = n20940 ^ n20939 ^ n19146 ;
  assign n20942 = n4527 ^ n3580 ^ 1'b0 ;
  assign n20943 = n13893 & ~n15525 ;
  assign n20944 = n20943 ^ n11181 ^ 1'b0 ;
  assign n20945 = ~n2396 & n2838 ;
  assign n20946 = n17970 ^ n842 ^ 1'b0 ;
  assign n20947 = n17998 ^ n8827 ^ n7232 ;
  assign n20948 = ( n7911 & ~n11718 ) | ( n7911 & n12477 ) | ( ~n11718 & n12477 ) ;
  assign n20949 = n20948 ^ n11576 ^ 1'b0 ;
  assign n20950 = ~n20947 & n20949 ;
  assign n20951 = n4060 & n7869 ;
  assign n20952 = ~n7423 & n20951 ;
  assign n20953 = ~n10659 & n16067 ;
  assign n20954 = n20953 ^ n13629 ^ 1'b0 ;
  assign n20955 = ( n6921 & n13079 ) | ( n6921 & ~n20954 ) | ( n13079 & ~n20954 ) ;
  assign n20956 = n20955 ^ n8287 ^ n239 ;
  assign n20957 = ~n2364 & n11371 ;
  assign n20958 = n6208 & n20957 ;
  assign n20959 = n10043 | n20958 ;
  assign n20960 = n11958 ^ n10418 ^ 1'b0 ;
  assign n20961 = n5235 & n16289 ;
  assign n20962 = ~n5251 & n20961 ;
  assign n20963 = ~n8687 & n20962 ;
  assign n20964 = n20963 ^ n11692 ^ 1'b0 ;
  assign n20965 = n15680 ^ n6649 ^ 1'b0 ;
  assign n20966 = n20965 ^ n12668 ^ 1'b0 ;
  assign n20967 = n10843 & n20966 ;
  assign n20968 = n8307 & n14428 ;
  assign n20969 = n983 ^ n379 ^ 1'b0 ;
  assign n20970 = ( n2433 & n4123 ) | ( n2433 & n20969 ) | ( n4123 & n20969 ) ;
  assign n20971 = ( ~n8265 & n12319 ) | ( ~n8265 & n20970 ) | ( n12319 & n20970 ) ;
  assign n20972 = n10986 ^ n2449 ^ n1664 ;
  assign n20973 = n2572 | n20972 ;
  assign n20974 = n16010 & ~n20973 ;
  assign n20975 = n20974 ^ n11286 ^ 1'b0 ;
  assign n20976 = n2281 | n3077 ;
  assign n20977 = n13534 & ~n20976 ;
  assign n20980 = n8409 ^ n6336 ^ n1412 ;
  assign n20979 = n889 & n5661 ;
  assign n20981 = n20980 ^ n20979 ^ 1'b0 ;
  assign n20978 = ~n5638 & n14170 ;
  assign n20982 = n20981 ^ n20978 ^ 1'b0 ;
  assign n20983 = ( n13515 & n20977 ) | ( n13515 & ~n20982 ) | ( n20977 & ~n20982 ) ;
  assign n20984 = x21 & ~n6495 ;
  assign n20985 = ~n3398 & n20984 ;
  assign n20986 = n20136 ^ n7760 ^ n2009 ;
  assign n20987 = n8170 & n20986 ;
  assign n20988 = n885 & n20987 ;
  assign n20989 = n20988 ^ n928 ^ 1'b0 ;
  assign n20990 = n20989 ^ n9617 ^ n3169 ;
  assign n20991 = n10809 & n14151 ;
  assign n20992 = ~n4840 & n20991 ;
  assign n20993 = x123 & n13961 ;
  assign n20994 = n7306 ^ n2273 ^ n1077 ;
  assign n20995 = n20994 ^ n10137 ^ 1'b0 ;
  assign n20996 = n8134 & n14297 ;
  assign n20997 = n5259 & n20996 ;
  assign n20998 = n12966 & n16607 ;
  assign n20999 = n257 & ~n1138 ;
  assign n21000 = n8665 ^ n6409 ^ 1'b0 ;
  assign n21001 = n20999 & n21000 ;
  assign n21002 = n18219 & n21001 ;
  assign n21003 = n21002 ^ n8603 ^ 1'b0 ;
  assign n21004 = ( n493 & n15287 ) | ( n493 & n20141 ) | ( n15287 & n20141 ) ;
  assign n21005 = ( n1730 & ~n2102 ) | ( n1730 & n3948 ) | ( ~n2102 & n3948 ) ;
  assign n21006 = n21005 ^ n3612 ^ 1'b0 ;
  assign n21007 = ~n21004 & n21006 ;
  assign n21008 = ( n2043 & n15872 ) | ( n2043 & n17686 ) | ( n15872 & n17686 ) ;
  assign n21009 = n12954 ^ n1431 ^ 1'b0 ;
  assign n21010 = n6995 ^ n6807 ^ n4341 ;
  assign n21011 = n21010 ^ n19698 ^ n11030 ;
  assign n21012 = n349 & ~n5570 ;
  assign n21013 = n1608 | n10297 ;
  assign n21014 = n21013 ^ n13758 ^ 1'b0 ;
  assign n21015 = n4857 & ~n8770 ;
  assign n21016 = n21014 & n21015 ;
  assign n21017 = ( n3704 & n4145 ) | ( n3704 & ~n4686 ) | ( n4145 & ~n4686 ) ;
  assign n21018 = n21017 ^ n18678 ^ n7762 ;
  assign n21019 = ~n16980 & n20611 ;
  assign n21020 = n21019 ^ n12611 ^ 1'b0 ;
  assign n21021 = ( ~n5886 & n21018 ) | ( ~n5886 & n21020 ) | ( n21018 & n21020 ) ;
  assign n21024 = n7318 & ~n9804 ;
  assign n21022 = ( n1910 & n4334 ) | ( n1910 & n7562 ) | ( n4334 & n7562 ) ;
  assign n21023 = ( n1745 & ~n17510 ) | ( n1745 & n21022 ) | ( ~n17510 & n21022 ) ;
  assign n21025 = n21024 ^ n21023 ^ n12928 ;
  assign n21026 = n1942 & n21025 ;
  assign n21027 = ~n21021 & n21026 ;
  assign n21029 = n13827 ^ n7228 ^ 1'b0 ;
  assign n21028 = ~n6881 & n11300 ;
  assign n21030 = n21029 ^ n21028 ^ 1'b0 ;
  assign n21031 = ( n8281 & n9811 ) | ( n8281 & ~n18202 ) | ( n9811 & ~n18202 ) ;
  assign n21032 = n10224 ^ n4157 ^ 1'b0 ;
  assign n21033 = n10460 & ~n21032 ;
  assign n21034 = ( ~n4669 & n15078 ) | ( ~n4669 & n21033 ) | ( n15078 & n21033 ) ;
  assign n21035 = ( n17896 & ~n21031 ) | ( n17896 & n21034 ) | ( ~n21031 & n21034 ) ;
  assign n21038 = ~n3192 & n5629 ;
  assign n21039 = n681 | n21038 ;
  assign n21040 = n7835 & ~n21039 ;
  assign n21036 = n168 & n341 ;
  assign n21037 = n21036 ^ n4577 ^ 1'b0 ;
  assign n21041 = n21040 ^ n21037 ^ n13848 ;
  assign n21042 = n14350 | n19208 ;
  assign n21043 = n3200 | n21042 ;
  assign n21044 = ( ~n8187 & n8281 ) | ( ~n8187 & n8634 ) | ( n8281 & n8634 ) ;
  assign n21045 = n12270 ^ n10417 ^ n8240 ;
  assign n21046 = n6104 | n18212 ;
  assign n21047 = n21045 & ~n21046 ;
  assign n21048 = n21044 | n21047 ;
  assign n21049 = n21048 ^ n18328 ^ n13063 ;
  assign n21050 = n11597 | n12218 ;
  assign n21051 = n13234 & ~n21050 ;
  assign n21052 = n7224 ^ n6005 ^ 1'b0 ;
  assign n21053 = n4619 & ~n21052 ;
  assign n21054 = ( n3534 & ~n4307 ) | ( n3534 & n7574 ) | ( ~n4307 & n7574 ) ;
  assign n21055 = n21054 ^ n539 ^ 1'b0 ;
  assign n21056 = n21053 & ~n21055 ;
  assign n21057 = n16738 ^ n12795 ^ x22 ;
  assign n21058 = ~n7350 & n14735 ;
  assign n21059 = n21058 ^ n12858 ^ 1'b0 ;
  assign n21060 = n777 & n21056 ;
  assign n21061 = n21060 ^ n10634 ^ 1'b0 ;
  assign n21062 = n1818 & ~n2092 ;
  assign n21063 = n21062 ^ n15274 ^ n1793 ;
  assign n21064 = n474 & n21063 ;
  assign n21065 = n10025 & n21064 ;
  assign n21066 = x77 & ~n21065 ;
  assign n21067 = n5334 & n21066 ;
  assign n21069 = n8991 ^ n3024 ^ n2115 ;
  assign n21072 = n3634 ^ n3185 ^ n2426 ;
  assign n21071 = n13997 ^ n11888 ^ 1'b0 ;
  assign n21073 = n21072 ^ n21071 ^ n3555 ;
  assign n21070 = x113 & n12589 ;
  assign n21074 = n21073 ^ n21070 ^ 1'b0 ;
  assign n21075 = ~n21069 & n21074 ;
  assign n21068 = n2821 & n20133 ;
  assign n21076 = n21075 ^ n21068 ^ 1'b0 ;
  assign n21078 = n829 | n4187 ;
  assign n21077 = n20051 ^ x65 ^ 1'b0 ;
  assign n21079 = n21078 ^ n21077 ^ n5133 ;
  assign n21083 = n18186 ^ n14908 ^ n405 ;
  assign n21084 = n11889 & ~n21083 ;
  assign n21080 = ( n8365 & n10380 ) | ( n8365 & n12756 ) | ( n10380 & n12756 ) ;
  assign n21081 = n5271 | n21080 ;
  assign n21082 = n11840 | n21081 ;
  assign n21085 = n21084 ^ n21082 ^ n18386 ;
  assign n21086 = n14875 ^ n12881 ^ 1'b0 ;
  assign n21087 = n8478 & ~n21086 ;
  assign n21088 = n6072 | n6319 ;
  assign n21089 = ~n8765 & n11328 ;
  assign n21090 = ~n18154 & n21089 ;
  assign n21091 = ( n7401 & n13160 ) | ( n7401 & n15564 ) | ( n13160 & n15564 ) ;
  assign n21092 = n21091 ^ n6646 ^ n2711 ;
  assign n21093 = n3272 & ~n14865 ;
  assign n21094 = n13863 | n18062 ;
  assign n21095 = ~n20857 & n21094 ;
  assign n21096 = ~n17652 & n21095 ;
  assign n21097 = n5992 & ~n18210 ;
  assign n21098 = n21097 ^ n12212 ^ 1'b0 ;
  assign n21099 = ~n13354 & n19317 ;
  assign n21100 = n14249 & n21099 ;
  assign n21101 = n16136 ^ n1705 ^ 1'b0 ;
  assign n21102 = ~n6566 & n21101 ;
  assign n21103 = n20507 ^ n7067 ^ 1'b0 ;
  assign n21104 = n16483 & n21103 ;
  assign n21105 = ( n13678 & n20981 ) | ( n13678 & ~n21104 ) | ( n20981 & ~n21104 ) ;
  assign n21106 = ( n4078 & ~n12077 ) | ( n4078 & n19729 ) | ( ~n12077 & n19729 ) ;
  assign n21107 = n21106 ^ n9675 ^ 1'b0 ;
  assign n21108 = n4440 ^ n2869 ^ n1149 ;
  assign n21109 = ( x112 & n12204 ) | ( x112 & n17124 ) | ( n12204 & n17124 ) ;
  assign n21110 = ( n1989 & n9097 ) | ( n1989 & n19216 ) | ( n9097 & n19216 ) ;
  assign n21111 = ( ~n153 & n5326 ) | ( ~n153 & n21110 ) | ( n5326 & n21110 ) ;
  assign n21112 = ~n17797 & n21111 ;
  assign n21117 = n1632 ^ n1302 ^ 1'b0 ;
  assign n21118 = n11388 & n21117 ;
  assign n21113 = n11337 | n13002 ;
  assign n21114 = n6551 & ~n21113 ;
  assign n21115 = ( ~n2568 & n5596 ) | ( ~n2568 & n21114 ) | ( n5596 & n21114 ) ;
  assign n21116 = n10562 & ~n21115 ;
  assign n21119 = n21118 ^ n21116 ^ 1'b0 ;
  assign n21120 = n3419 ^ n164 ^ 1'b0 ;
  assign n21121 = n16279 & n21120 ;
  assign n21122 = ( n6541 & n8434 ) | ( n6541 & ~n21121 ) | ( n8434 & ~n21121 ) ;
  assign n21123 = n21122 ^ n9790 ^ 1'b0 ;
  assign n21124 = ( ~n5470 & n11491 ) | ( ~n5470 & n13904 ) | ( n11491 & n13904 ) ;
  assign n21125 = n5142 ^ n5113 ^ 1'b0 ;
  assign n21126 = ( n11135 & n20870 ) | ( n11135 & ~n21125 ) | ( n20870 & ~n21125 ) ;
  assign n21127 = n1274 & ~n11905 ;
  assign n21128 = n17786 ^ n368 ^ 1'b0 ;
  assign n21129 = n21127 | n21128 ;
  assign n21130 = n2444 & n6674 ;
  assign n21131 = ~n9460 & n21130 ;
  assign n21132 = n21131 ^ n3220 ^ 1'b0 ;
  assign n21133 = n4633 | n5711 ;
  assign n21134 = n20875 & ~n21133 ;
  assign n21135 = ~n4272 & n13220 ;
  assign n21136 = n10650 & n21135 ;
  assign n21137 = ~n283 & n21136 ;
  assign n21138 = n17792 ^ n16691 ^ n6150 ;
  assign n21139 = n9815 ^ n3837 ^ 1'b0 ;
  assign n21141 = n4561 | n5952 ;
  assign n21142 = n14785 & ~n21141 ;
  assign n21140 = ( n2363 & n4195 ) | ( n2363 & n4204 ) | ( n4195 & n4204 ) ;
  assign n21143 = n21142 ^ n21140 ^ n5402 ;
  assign n21144 = n722 & n12003 ;
  assign n21145 = n21144 ^ n12008 ^ 1'b0 ;
  assign n21146 = n1883 & ~n6719 ;
  assign n21147 = n17583 & n21146 ;
  assign n21148 = ( n3325 & n3637 ) | ( n3325 & ~n11188 ) | ( n3637 & ~n11188 ) ;
  assign n21149 = n21148 ^ n196 ^ 1'b0 ;
  assign n21150 = n3766 | n21149 ;
  assign n21151 = n12646 & ~n13611 ;
  assign n21152 = n21151 ^ n18779 ^ n6350 ;
  assign n21153 = n21152 ^ x68 ^ 1'b0 ;
  assign n21154 = n18250 & ~n21153 ;
  assign n21155 = n12719 ^ n5375 ^ n2372 ;
  assign n21156 = ( ~n3095 & n4052 ) | ( ~n3095 & n21155 ) | ( n4052 & n21155 ) ;
  assign n21157 = ( ~n10348 & n11109 ) | ( ~n10348 & n21156 ) | ( n11109 & n21156 ) ;
  assign n21158 = n13576 ^ n6239 ^ 1'b0 ;
  assign n21159 = n3293 & n21158 ;
  assign n21160 = ~n12248 & n21159 ;
  assign n21161 = n7141 & n16902 ;
  assign n21162 = x22 & ~n20521 ;
  assign n21163 = n11031 ^ n6926 ^ 1'b0 ;
  assign n21164 = n1052 ^ x106 ^ 1'b0 ;
  assign n21165 = n21163 & n21164 ;
  assign n21166 = n16590 & n20948 ;
  assign n21167 = n3463 ^ n1898 ^ 1'b0 ;
  assign n21168 = n21167 ^ n13034 ^ 1'b0 ;
  assign n21169 = n12116 ^ n8450 ^ n2315 ;
  assign n21170 = ( n1059 & n1671 ) | ( n1059 & n1686 ) | ( n1671 & n1686 ) ;
  assign n21171 = n14055 & ~n21170 ;
  assign n21172 = ( ~n250 & n349 ) | ( ~n250 & n1382 ) | ( n349 & n1382 ) ;
  assign n21173 = n13413 & n21172 ;
  assign n21174 = ( ~n11685 & n21171 ) | ( ~n11685 & n21173 ) | ( n21171 & n21173 ) ;
  assign n21178 = n9552 ^ n619 ^ 1'b0 ;
  assign n21179 = n14003 & ~n21178 ;
  assign n21176 = ( ~n12822 & n15759 ) | ( ~n12822 & n16805 ) | ( n15759 & n16805 ) ;
  assign n21175 = n4825 ^ n2587 ^ 1'b0 ;
  assign n21177 = n21176 ^ n21175 ^ n8132 ;
  assign n21180 = n21179 ^ n21177 ^ n6125 ;
  assign n21181 = n21180 ^ n19304 ^ 1'b0 ;
  assign n21182 = n15955 ^ n15502 ^ 1'b0 ;
  assign n21183 = n15296 & n21182 ;
  assign n21184 = n11036 & n21183 ;
  assign n21185 = ~n14540 & n21184 ;
  assign n21186 = n21185 ^ n18141 ^ n6128 ;
  assign n21188 = ( n2091 & n9602 ) | ( n2091 & n10674 ) | ( n9602 & n10674 ) ;
  assign n21187 = n6976 & ~n7365 ;
  assign n21189 = n21188 ^ n21187 ^ n17135 ;
  assign n21190 = n21189 ^ n4880 ^ 1'b0 ;
  assign n21191 = n13113 & ~n21190 ;
  assign n21192 = n15785 ^ n10420 ^ n4706 ;
  assign n21193 = n9664 ^ n9657 ^ n8077 ;
  assign n21194 = n17612 ^ n15166 ^ n9497 ;
  assign n21195 = ( n4740 & n5222 ) | ( n4740 & n16368 ) | ( n5222 & n16368 ) ;
  assign n21196 = n15486 ^ n7635 ^ n6668 ;
  assign n21197 = n21196 ^ n5233 ^ 1'b0 ;
  assign n21198 = n16310 ^ n8758 ^ 1'b0 ;
  assign n21199 = n10349 & ~n21198 ;
  assign n21202 = n10611 ^ n6714 ^ n3416 ;
  assign n21203 = ( n6520 & n10205 ) | ( n6520 & ~n21202 ) | ( n10205 & ~n21202 ) ;
  assign n21201 = ~n6824 & n17629 ;
  assign n21204 = n21203 ^ n21201 ^ 1'b0 ;
  assign n21200 = n16174 & n18249 ;
  assign n21205 = n21204 ^ n21200 ^ 1'b0 ;
  assign n21206 = n5982 ^ n1009 ^ 1'b0 ;
  assign n21207 = n2311 & ~n21206 ;
  assign n21208 = ~n8422 & n13620 ;
  assign n21209 = ( x60 & ~n21207 ) | ( x60 & n21208 ) | ( ~n21207 & n21208 ) ;
  assign n21210 = ~n954 & n8361 ;
  assign n21211 = n21210 ^ n18935 ^ n13492 ;
  assign n21212 = ( n2497 & n6171 ) | ( n2497 & n19033 ) | ( n6171 & n19033 ) ;
  assign n21213 = ~n10324 & n12861 ;
  assign n21214 = ~n20190 & n21213 ;
  assign n21215 = ( n312 & n8552 ) | ( n312 & ~n21214 ) | ( n8552 & ~n21214 ) ;
  assign n21217 = x83 & ~n15486 ;
  assign n21216 = n9875 & ~n17477 ;
  assign n21218 = n21217 ^ n21216 ^ 1'b0 ;
  assign n21219 = ~n3448 & n21218 ;
  assign n21220 = n21219 ^ n6312 ^ 1'b0 ;
  assign n21221 = n12368 ^ n5954 ^ 1'b0 ;
  assign n21222 = n7011 & n21221 ;
  assign n21223 = ~n7488 & n21222 ;
  assign n21224 = n14266 ^ n8012 ^ 1'b0 ;
  assign n21225 = n8601 | n15746 ;
  assign n21226 = n20463 & ~n21225 ;
  assign n21227 = n1348 | n21226 ;
  assign n21228 = ( ~n3951 & n21224 ) | ( ~n3951 & n21227 ) | ( n21224 & n21227 ) ;
  assign n21229 = n21228 ^ n11745 ^ 1'b0 ;
  assign n21230 = n21229 ^ n5056 ^ 1'b0 ;
  assign n21235 = n1964 & n7171 ;
  assign n21236 = n21235 ^ n5403 ^ n3930 ;
  assign n21231 = n6211 & ~n8138 ;
  assign n21232 = ~n2811 & n21231 ;
  assign n21233 = n14404 ^ n12798 ^ 1'b0 ;
  assign n21234 = ~n21232 & n21233 ;
  assign n21237 = n21236 ^ n21234 ^ 1'b0 ;
  assign n21240 = ( n144 & n1570 ) | ( n144 & n3883 ) | ( n1570 & n3883 ) ;
  assign n21241 = n5511 | n21240 ;
  assign n21242 = n5211 | n21241 ;
  assign n21238 = n2152 & ~n13963 ;
  assign n21239 = n1571 & n21238 ;
  assign n21243 = n21242 ^ n21239 ^ 1'b0 ;
  assign n21244 = n19959 ^ n3590 ^ 1'b0 ;
  assign n21246 = ( ~n2267 & n6247 ) | ( ~n2267 & n8619 ) | ( n6247 & n8619 ) ;
  assign n21245 = n7284 | n14536 ;
  assign n21247 = n21246 ^ n21245 ^ n10297 ;
  assign n21248 = n7332 ^ n2726 ^ 1'b0 ;
  assign n21249 = n6777 | n21248 ;
  assign n21250 = ~n3004 & n21249 ;
  assign n21251 = ( n9418 & n13119 ) | ( n9418 & n16168 ) | ( n13119 & n16168 ) ;
  assign n21252 = n21251 ^ n579 ^ n314 ;
  assign n21253 = ( ~n4203 & n4754 ) | ( ~n4203 & n18649 ) | ( n4754 & n18649 ) ;
  assign n21254 = n3703 | n5665 ;
  assign n21255 = n19996 ^ n17492 ^ n11745 ;
  assign n21256 = n11308 ^ n5311 ^ n3221 ;
  assign n21257 = n8571 ^ n766 ^ 1'b0 ;
  assign n21258 = n5873 & n8466 ;
  assign n21259 = n7934 & n21258 ;
  assign n21260 = n21257 & n21259 ;
  assign n21262 = n7197 | n8029 ;
  assign n21263 = n1330 | n21262 ;
  assign n21261 = ~n1572 & n17391 ;
  assign n21264 = n21263 ^ n21261 ^ 1'b0 ;
  assign n21265 = ~n6592 & n6847 ;
  assign n21266 = n7618 ^ n171 ^ 1'b0 ;
  assign n21267 = n10989 & n21266 ;
  assign n21268 = n12109 ^ n7526 ^ n2949 ;
  assign n21269 = n11930 & n21268 ;
  assign n21270 = n11502 | n15213 ;
  assign n21271 = n21270 ^ n19063 ^ n11557 ;
  assign n21272 = n18051 ^ n2189 ^ 1'b0 ;
  assign n21273 = n2810 | n21272 ;
  assign n21274 = ( x27 & n7822 ) | ( x27 & n19754 ) | ( n7822 & n19754 ) ;
  assign n21275 = ( ~n12928 & n21273 ) | ( ~n12928 & n21274 ) | ( n21273 & n21274 ) ;
  assign n21276 = n2516 & n16279 ;
  assign n21277 = n21276 ^ n1609 ^ 1'b0 ;
  assign n21278 = ( n1704 & n11391 ) | ( n1704 & ~n21277 ) | ( n11391 & ~n21277 ) ;
  assign n21279 = n21278 ^ n15481 ^ n11632 ;
  assign n21280 = n13114 ^ n12041 ^ 1'b0 ;
  assign n21281 = n2468 | n15924 ;
  assign n21282 = n3992 & ~n21281 ;
  assign n21283 = n5714 | n17177 ;
  assign n21284 = ( ~n3862 & n21282 ) | ( ~n3862 & n21283 ) | ( n21282 & n21283 ) ;
  assign n21285 = n16810 | n21284 ;
  assign n21286 = ~n8890 & n20601 ;
  assign n21287 = n21286 ^ n14545 ^ 1'b0 ;
  assign n21288 = ( n3542 & ~n12425 ) | ( n3542 & n20417 ) | ( ~n12425 & n20417 ) ;
  assign n21289 = n21288 ^ n12481 ^ n8269 ;
  assign n21290 = n18295 ^ n2730 ^ n2156 ;
  assign n21291 = n21290 ^ n11382 ^ n7496 ;
  assign n21292 = n15030 ^ n10880 ^ n1467 ;
  assign n21293 = n20092 ^ n1152 ^ 1'b0 ;
  assign n21294 = ~n5682 & n21293 ;
  assign n21295 = n21294 ^ n8457 ^ 1'b0 ;
  assign n21296 = n10746 ^ n4234 ^ 1'b0 ;
  assign n21297 = ~n4941 & n21296 ;
  assign n21298 = n2842 ^ n2832 ^ 1'b0 ;
  assign n21299 = n6214 ^ n5411 ^ n5157 ;
  assign n21300 = ( n3655 & n4299 ) | ( n3655 & ~n6283 ) | ( n4299 & ~n6283 ) ;
  assign n21301 = ( n1054 & n13029 ) | ( n1054 & n21300 ) | ( n13029 & n21300 ) ;
  assign n21302 = ( n597 & n3027 ) | ( n597 & ~n19998 ) | ( n3027 & ~n19998 ) ;
  assign n21303 = n6668 ^ n6233 ^ n917 ;
  assign n21304 = n2853 | n21303 ;
  assign n21305 = ~n7409 & n17974 ;
  assign n21306 = n9342 & n21305 ;
  assign n21307 = n17639 ^ n1682 ^ 1'b0 ;
  assign n21308 = n10152 ^ n5889 ^ 1'b0 ;
  assign n21309 = n5228 | n21308 ;
  assign n21310 = n12355 & ~n21309 ;
  assign n21311 = n4299 & n21310 ;
  assign n21312 = n17280 ^ n11108 ^ n7234 ;
  assign n21313 = n19141 ^ n7578 ^ 1'b0 ;
  assign n21316 = n1511 | n17174 ;
  assign n21314 = n9515 ^ n5122 ^ x107 ;
  assign n21315 = n1369 | n21314 ;
  assign n21317 = n21316 ^ n21315 ^ 1'b0 ;
  assign n21318 = n15242 ^ n8961 ^ 1'b0 ;
  assign n21319 = ( x81 & n12170 ) | ( x81 & ~n21318 ) | ( n12170 & ~n21318 ) ;
  assign n21320 = ( ~n13716 & n20392 ) | ( ~n13716 & n21319 ) | ( n20392 & n21319 ) ;
  assign n21321 = ( n5056 & ~n9403 ) | ( n5056 & n13881 ) | ( ~n9403 & n13881 ) ;
  assign n21322 = n9968 ^ n2359 ^ 1'b0 ;
  assign n21323 = n5597 & ~n21322 ;
  assign n21324 = n6848 & ~n17303 ;
  assign n21325 = n4062 & n21324 ;
  assign n21326 = n1406 & ~n3467 ;
  assign n21327 = n4083 & n21326 ;
  assign n21328 = ~n5961 & n11038 ;
  assign n21329 = n21328 ^ n343 ^ 1'b0 ;
  assign n21330 = ( n3352 & ~n8366 ) | ( n3352 & n11771 ) | ( ~n8366 & n11771 ) ;
  assign n21331 = n7753 & ~n21330 ;
  assign n21332 = ~n21329 & n21331 ;
  assign n21333 = ( n5109 & n14904 ) | ( n5109 & ~n21332 ) | ( n14904 & ~n21332 ) ;
  assign n21334 = ( n4733 & n5053 ) | ( n4733 & ~n17582 ) | ( n5053 & ~n17582 ) ;
  assign n21335 = ( n3763 & n17256 ) | ( n3763 & ~n21334 ) | ( n17256 & ~n21334 ) ;
  assign n21336 = n14058 & ~n19103 ;
  assign n21337 = n21336 ^ n11288 ^ 1'b0 ;
  assign n21338 = n20100 ^ n4502 ^ 1'b0 ;
  assign n21339 = n11190 ^ n1034 ^ 1'b0 ;
  assign n21340 = n18278 ^ n1586 ^ 1'b0 ;
  assign n21341 = n21339 | n21340 ;
  assign n21342 = n4553 & n21341 ;
  assign n21344 = n266 & n7675 ;
  assign n21345 = n12368 | n21344 ;
  assign n21346 = n15449 | n21345 ;
  assign n21343 = n16239 | n16641 ;
  assign n21347 = n21346 ^ n21343 ^ 1'b0 ;
  assign n21348 = n10459 ^ n7251 ^ 1'b0 ;
  assign n21349 = ( ~n11629 & n11777 ) | ( ~n11629 & n21348 ) | ( n11777 & n21348 ) ;
  assign n21350 = n21349 ^ n13499 ^ 1'b0 ;
  assign n21351 = n18665 ^ n10812 ^ 1'b0 ;
  assign n21352 = n573 | n17817 ;
  assign n21353 = n18371 ^ n12075 ^ 1'b0 ;
  assign n21354 = ~n2697 & n21353 ;
  assign n21355 = n11444 ^ n5993 ^ 1'b0 ;
  assign n21356 = ~n1738 & n21355 ;
  assign n21357 = ~n14098 & n21356 ;
  assign n21358 = n17301 ^ n11406 ^ n9749 ;
  assign n21359 = n7424 | n10721 ;
  assign n21360 = ( n8777 & n21358 ) | ( n8777 & ~n21359 ) | ( n21358 & ~n21359 ) ;
  assign n21361 = ( ~n6131 & n7070 ) | ( ~n6131 & n21360 ) | ( n7070 & n21360 ) ;
  assign n21362 = ~n1520 & n10432 ;
  assign n21363 = ~n6947 & n21362 ;
  assign n21364 = n695 | n17686 ;
  assign n21365 = n21364 ^ n3713 ^ 1'b0 ;
  assign n21366 = n21363 & n21365 ;
  assign n21367 = ( ~n831 & n5228 ) | ( ~n831 & n11120 ) | ( n5228 & n11120 ) ;
  assign n21368 = n9848 | n21367 ;
  assign n21369 = ~n4602 & n5799 ;
  assign n21370 = ( n17562 & ~n18708 ) | ( n17562 & n21369 ) | ( ~n18708 & n21369 ) ;
  assign n21371 = n15649 ^ n8223 ^ 1'b0 ;
  assign n21372 = n9268 & n21371 ;
  assign n21373 = n9860 ^ n3980 ^ 1'b0 ;
  assign n21374 = ~n10295 & n21373 ;
  assign n21375 = n21374 ^ n10304 ^ 1'b0 ;
  assign n21376 = n11074 & n21375 ;
  assign n21377 = ( n1448 & ~n3274 ) | ( n1448 & n4658 ) | ( ~n3274 & n4658 ) ;
  assign n21378 = n19998 & ~n21152 ;
  assign n21379 = n3825 ^ n689 ^ 1'b0 ;
  assign n21380 = n19141 & n21379 ;
  assign n21381 = n2149 & ~n2706 ;
  assign n21382 = n21381 ^ n6564 ^ n4461 ;
  assign n21383 = ( n21378 & n21380 ) | ( n21378 & n21382 ) | ( n21380 & n21382 ) ;
  assign n21384 = n12457 ^ n5858 ^ 1'b0 ;
  assign n21385 = n2141 | n2796 ;
  assign n21386 = n21385 ^ n8789 ^ x30 ;
  assign n21387 = ( n7425 & n21384 ) | ( n7425 & n21386 ) | ( n21384 & n21386 ) ;
  assign n21391 = n4434 | n6866 ;
  assign n21392 = n16909 & ~n21391 ;
  assign n21388 = n9359 ^ n5355 ^ 1'b0 ;
  assign n21389 = n20585 | n21388 ;
  assign n21390 = n19063 | n21389 ;
  assign n21393 = n21392 ^ n21390 ^ n7757 ;
  assign n21394 = n3905 & n20324 ;
  assign n21395 = n21394 ^ n7627 ^ 1'b0 ;
  assign n21396 = n1566 | n14072 ;
  assign n21399 = n8314 ^ n318 ^ 1'b0 ;
  assign n21400 = ( n11570 & n15566 ) | ( n11570 & n21399 ) | ( n15566 & n21399 ) ;
  assign n21397 = ~n4986 & n19390 ;
  assign n21398 = ~n8936 & n21397 ;
  assign n21401 = n21400 ^ n21398 ^ 1'b0 ;
  assign n21402 = n2051 | n17271 ;
  assign n21403 = ( n403 & n9414 ) | ( n403 & ~n21402 ) | ( n9414 & ~n21402 ) ;
  assign n21404 = n21403 ^ n3971 ^ 1'b0 ;
  assign n21405 = ( n652 & ~n3742 ) | ( n652 & n18631 ) | ( ~n3742 & n18631 ) ;
  assign n21406 = n15823 ^ n12644 ^ n11867 ;
  assign n21407 = n16047 & ~n16053 ;
  assign n21408 = n10820 ^ n8349 ^ 1'b0 ;
  assign n21409 = ~n5281 & n21408 ;
  assign n21410 = n21409 ^ n11134 ^ n4703 ;
  assign n21411 = ( n7375 & ~n11955 ) | ( n7375 & n12606 ) | ( ~n11955 & n12606 ) ;
  assign n21412 = n12341 & ~n17262 ;
  assign n21413 = n21412 ^ n8887 ^ 1'b0 ;
  assign n21417 = n12284 ^ n9338 ^ n7347 ;
  assign n21414 = n8997 ^ n3828 ^ 1'b0 ;
  assign n21415 = n21414 ^ n8444 ^ 1'b0 ;
  assign n21416 = n12657 & n21415 ;
  assign n21418 = n21417 ^ n21416 ^ 1'b0 ;
  assign n21419 = n20100 ^ n3595 ^ n452 ;
  assign n21420 = n5497 & ~n7488 ;
  assign n21421 = n5604 | n10724 ;
  assign n21422 = n21421 ^ n5510 ^ 1'b0 ;
  assign n21423 = n10084 ^ n8392 ^ 1'b0 ;
  assign n21424 = ~n11849 & n21423 ;
  assign n21425 = n21424 ^ n11910 ^ 1'b0 ;
  assign n21426 = n3396 ^ n2436 ^ n506 ;
  assign n21427 = n21426 ^ n9427 ^ 1'b0 ;
  assign n21428 = n14342 | n21427 ;
  assign n21437 = n6599 & ~n10829 ;
  assign n21438 = n21437 ^ n6706 ^ 1'b0 ;
  assign n21439 = ( ~n2910 & n9580 ) | ( ~n2910 & n21438 ) | ( n9580 & n21438 ) ;
  assign n21435 = n4222 & ~n7197 ;
  assign n21436 = n21435 ^ n14949 ^ 1'b0 ;
  assign n21430 = ~n8579 & n9878 ;
  assign n21431 = n10306 & n21430 ;
  assign n21429 = n1342 | n15281 ;
  assign n21432 = n21431 ^ n21429 ^ 1'b0 ;
  assign n21433 = n14721 & ~n21432 ;
  assign n21434 = n21433 ^ n10920 ^ 1'b0 ;
  assign n21440 = n21439 ^ n21436 ^ n21434 ;
  assign n21442 = n1427 & ~n1695 ;
  assign n21441 = n5118 ^ n4083 ^ n153 ;
  assign n21443 = n21442 ^ n21441 ^ n4147 ;
  assign n21444 = n16541 ^ n12088 ^ 1'b0 ;
  assign n21445 = ( n1267 & n6483 ) | ( n1267 & n16024 ) | ( n6483 & n16024 ) ;
  assign n21446 = n2074 | n21445 ;
  assign n21447 = n12404 ^ n1656 ^ x65 ;
  assign n21448 = n8670 & ~n21447 ;
  assign n21449 = n21448 ^ n11140 ^ 1'b0 ;
  assign n21450 = n3244 & n9591 ;
  assign n21455 = n20615 ^ n2279 ^ 1'b0 ;
  assign n21456 = ~n4684 & n21455 ;
  assign n21451 = n3596 & n9561 ;
  assign n21452 = ~n2419 & n21451 ;
  assign n21453 = n21452 ^ n11653 ^ 1'b0 ;
  assign n21454 = n11776 & n21453 ;
  assign n21457 = n21456 ^ n21454 ^ 1'b0 ;
  assign n21458 = n11235 ^ n8502 ^ 1'b0 ;
  assign n21459 = ( n7597 & ~n20475 ) | ( n7597 & n20538 ) | ( ~n20475 & n20538 ) ;
  assign n21460 = n2663 & ~n12907 ;
  assign n21461 = n21460 ^ n13614 ^ n2631 ;
  assign n21462 = n15612 ^ n13769 ^ n4440 ;
  assign n21464 = n3999 ^ n3965 ^ 1'b0 ;
  assign n21463 = n14508 ^ n11689 ^ 1'b0 ;
  assign n21465 = n21464 ^ n21463 ^ n7737 ;
  assign n21466 = n8749 ^ n2975 ^ 1'b0 ;
  assign n21467 = n10065 & n21466 ;
  assign n21468 = ( n2558 & n7754 ) | ( n2558 & n21467 ) | ( n7754 & n21467 ) ;
  assign n21469 = ( n1745 & n3126 ) | ( n1745 & ~n7007 ) | ( n3126 & ~n7007 ) ;
  assign n21470 = ( n10197 & n21468 ) | ( n10197 & ~n21469 ) | ( n21468 & ~n21469 ) ;
  assign n21471 = n4176 ^ n2188 ^ n815 ;
  assign n21472 = n20777 & n21471 ;
  assign n21474 = ( ~n2528 & n2689 ) | ( ~n2528 & n4142 ) | ( n2689 & n4142 ) ;
  assign n21473 = n5472 & n16840 ;
  assign n21475 = n21474 ^ n21473 ^ 1'b0 ;
  assign n21476 = ( n994 & n8399 ) | ( n994 & ~n10688 ) | ( n8399 & ~n10688 ) ;
  assign n21477 = ( n1268 & n10713 ) | ( n1268 & ~n11465 ) | ( n10713 & ~n11465 ) ;
  assign n21478 = n21476 | n21477 ;
  assign n21479 = n4318 & n21478 ;
  assign n21480 = n9938 ^ n6779 ^ 1'b0 ;
  assign n21481 = n1858 & ~n5958 ;
  assign n21482 = n21480 | n21481 ;
  assign n21483 = n21482 ^ n14432 ^ 1'b0 ;
  assign n21484 = n5131 & ~n21483 ;
  assign n21485 = n21484 ^ n1687 ^ 1'b0 ;
  assign n21486 = ( n5704 & ~n17324 ) | ( n5704 & n17811 ) | ( ~n17324 & n17811 ) ;
  assign n21487 = n11241 ^ n5341 ^ 1'b0 ;
  assign n21488 = n7367 & n9127 ;
  assign n21489 = ~n3232 & n21488 ;
  assign n21490 = n15250 & ~n20857 ;
  assign n21491 = n810 & n21490 ;
  assign n21492 = n21491 ^ n5941 ^ 1'b0 ;
  assign n21493 = ~n1073 & n21492 ;
  assign n21494 = ( n2868 & n4800 ) | ( n2868 & n6347 ) | ( n4800 & n6347 ) ;
  assign n21495 = ( n5174 & n9677 ) | ( n5174 & ~n21494 ) | ( n9677 & ~n21494 ) ;
  assign n21496 = n18363 ^ n17523 ^ n5652 ;
  assign n21497 = n20258 ^ n19796 ^ 1'b0 ;
  assign n21498 = n7070 & n10688 ;
  assign n21499 = n21498 ^ n2729 ^ 1'b0 ;
  assign n21500 = n12747 | n21499 ;
  assign n21501 = n21500 ^ n4931 ^ 1'b0 ;
  assign n21502 = ~n12945 & n21501 ;
  assign n21503 = n6230 ^ n2254 ^ 1'b0 ;
  assign n21504 = n6903 ^ n6419 ^ n4287 ;
  assign n21505 = n21504 ^ n3104 ^ 1'b0 ;
  assign n21506 = ( n3266 & n14147 ) | ( n3266 & ~n20262 ) | ( n14147 & ~n20262 ) ;
  assign n21508 = n1236 & ~n9664 ;
  assign n21509 = ~n14162 & n21508 ;
  assign n21507 = ~n4446 & n11019 ;
  assign n21510 = n21509 ^ n21507 ^ 1'b0 ;
  assign n21511 = n1160 & ~n17122 ;
  assign n21512 = ~n18288 & n21511 ;
  assign n21513 = n12105 ^ n3334 ^ 1'b0 ;
  assign n21514 = n21513 ^ n15872 ^ 1'b0 ;
  assign n21515 = n17302 | n21514 ;
  assign n21516 = n16214 ^ n9319 ^ 1'b0 ;
  assign n21517 = n8018 ^ n6866 ^ 1'b0 ;
  assign n21518 = x88 & n2665 ;
  assign n21519 = n21518 ^ n10624 ^ n7871 ;
  assign n21520 = ~n8056 & n21519 ;
  assign n21521 = n13865 & n19649 ;
  assign n21522 = n19966 ^ n10175 ^ 1'b0 ;
  assign n21523 = n10926 | n21522 ;
  assign n21524 = n12151 ^ n9179 ^ 1'b0 ;
  assign n21525 = n21524 ^ n17073 ^ n9979 ;
  assign n21527 = n3167 & ~n14005 ;
  assign n21528 = ~n17886 & n21527 ;
  assign n21526 = n3198 & ~n16065 ;
  assign n21529 = n21528 ^ n21526 ^ 1'b0 ;
  assign n21530 = n6817 | n9958 ;
  assign n21531 = n3548 | n4498 ;
  assign n21532 = n16114 | n21531 ;
  assign n21533 = ~n6971 & n21532 ;
  assign n21534 = n21533 ^ n16969 ^ 1'b0 ;
  assign n21540 = n3411 & ~n7813 ;
  assign n21539 = n9173 & n11057 ;
  assign n21537 = n12330 ^ n2173 ^ 1'b0 ;
  assign n21535 = ~n3854 & n20101 ;
  assign n21536 = n9339 | n21535 ;
  assign n21538 = n21537 ^ n21536 ^ 1'b0 ;
  assign n21541 = n21540 ^ n21539 ^ n21538 ;
  assign n21542 = ( n3188 & n6393 ) | ( n3188 & n17966 ) | ( n6393 & n17966 ) ;
  assign n21543 = n6652 ^ n3661 ^ 1'b0 ;
  assign n21544 = ( n14055 & ~n16968 ) | ( n14055 & n21543 ) | ( ~n16968 & n21543 ) ;
  assign n21545 = n18171 ^ n1929 ^ 1'b0 ;
  assign n21546 = n2899 ^ n2849 ^ 1'b0 ;
  assign n21547 = ~n21545 & n21546 ;
  assign n21548 = ( ~n1357 & n5616 ) | ( ~n1357 & n11615 ) | ( n5616 & n11615 ) ;
  assign n21549 = n10817 ^ n479 ^ 1'b0 ;
  assign n21550 = ~n21548 & n21549 ;
  assign n21551 = n6437 & n6901 ;
  assign n21552 = ~n9922 & n21551 ;
  assign n21553 = n8143 & n9059 ;
  assign n21554 = n14901 | n21553 ;
  assign n21555 = n21552 & ~n21554 ;
  assign n21556 = n255 & n3723 ;
  assign n21557 = n6391 & n21556 ;
  assign n21558 = n4696 & n21557 ;
  assign n21560 = n12948 ^ n10023 ^ n4789 ;
  assign n21559 = ~n2934 & n5655 ;
  assign n21561 = n21560 ^ n21559 ^ 1'b0 ;
  assign n21562 = ( n3970 & n19310 ) | ( n3970 & n21561 ) | ( n19310 & n21561 ) ;
  assign n21563 = n8326 ^ n6751 ^ 1'b0 ;
  assign n21565 = n2925 | n6391 ;
  assign n21564 = ~n1345 & n4493 ;
  assign n21566 = n21565 ^ n21564 ^ 1'b0 ;
  assign n21567 = ( n2079 & n7523 ) | ( n2079 & n21566 ) | ( n7523 & n21566 ) ;
  assign n21568 = n13818 ^ n7141 ^ n5979 ;
  assign n21569 = n1171 | n21071 ;
  assign n21570 = ~n1806 & n1883 ;
  assign n21571 = n1990 & n21570 ;
  assign n21572 = n21571 ^ n8217 ^ 1'b0 ;
  assign n21573 = ( n3635 & n4993 ) | ( n3635 & ~n7945 ) | ( n4993 & ~n7945 ) ;
  assign n21574 = n5179 & ~n21573 ;
  assign n21575 = ~n6263 & n21574 ;
  assign n21576 = n8073 ^ n6732 ^ 1'b0 ;
  assign n21577 = n21576 ^ n3007 ^ 1'b0 ;
  assign n21578 = n2163 & ~n5844 ;
  assign n21579 = n21578 ^ n347 ^ 1'b0 ;
  assign n21580 = ( n1984 & ~n10352 ) | ( n1984 & n21579 ) | ( ~n10352 & n21579 ) ;
  assign n21581 = n6215 & n21580 ;
  assign n21582 = n21581 ^ x28 ^ 1'b0 ;
  assign n21583 = n8773 ^ n7521 ^ 1'b0 ;
  assign n21584 = ( n2897 & n6587 ) | ( n2897 & n21583 ) | ( n6587 & n21583 ) ;
  assign n21585 = n21584 ^ n19331 ^ n12680 ;
  assign n21586 = n14815 ^ n13718 ^ n10415 ;
  assign n21587 = n10626 & ~n17277 ;
  assign n21588 = n21587 ^ n7524 ^ n5513 ;
  assign n21589 = n5342 | n14812 ;
  assign n21590 = n21589 ^ n9799 ^ 1'b0 ;
  assign n21591 = ( ~n5405 & n18842 ) | ( ~n5405 & n21590 ) | ( n18842 & n21590 ) ;
  assign n21592 = n1531 & ~n2779 ;
  assign n21593 = n21592 ^ n2879 ^ 1'b0 ;
  assign n21594 = n9822 & ~n20392 ;
  assign n21595 = n21594 ^ n20476 ^ 1'b0 ;
  assign n21596 = ~n18916 & n21595 ;
  assign n21597 = n21593 & n21596 ;
  assign n21599 = n8477 ^ n1664 ^ 1'b0 ;
  assign n21598 = n4148 | n17471 ;
  assign n21600 = n21599 ^ n21598 ^ 1'b0 ;
  assign n21602 = n6977 ^ n5259 ^ 1'b0 ;
  assign n21601 = ~n4839 & n20267 ;
  assign n21603 = n21602 ^ n21601 ^ n5778 ;
  assign n21604 = n15136 & ~n17600 ;
  assign n21605 = n21604 ^ n20797 ^ 1'b0 ;
  assign n21606 = n14026 ^ n1909 ^ 1'b0 ;
  assign n21607 = ~n6853 & n19937 ;
  assign n21611 = ( ~n1769 & n12642 ) | ( ~n1769 & n16182 ) | ( n12642 & n16182 ) ;
  assign n21608 = n5963 & ~n9654 ;
  assign n21609 = n21608 ^ n774 ^ 1'b0 ;
  assign n21610 = ( ~n8447 & n20908 ) | ( ~n8447 & n21609 ) | ( n20908 & n21609 ) ;
  assign n21612 = n21611 ^ n21610 ^ 1'b0 ;
  assign n21613 = n16435 ^ n13534 ^ 1'b0 ;
  assign n21614 = n654 ^ n577 ^ 1'b0 ;
  assign n21615 = n20078 ^ n12389 ^ 1'b0 ;
  assign n21616 = n21614 | n21615 ;
  assign n21617 = n10858 ^ n7468 ^ 1'b0 ;
  assign n21618 = n6351 & n21617 ;
  assign n21619 = n10098 | n15131 ;
  assign n21620 = n21619 ^ n6668 ^ 1'b0 ;
  assign n21621 = ~n5510 & n21620 ;
  assign n21622 = n21621 ^ n9793 ^ 1'b0 ;
  assign n21623 = ~n12887 & n21622 ;
  assign n21624 = n6619 | n9935 ;
  assign n21625 = n8519 & ~n21624 ;
  assign n21626 = n21625 ^ n9932 ^ 1'b0 ;
  assign n21627 = ~n3662 & n17673 ;
  assign n21628 = n21627 ^ n18071 ^ n1292 ;
  assign n21629 = n2681 | n4592 ;
  assign n21630 = n21629 ^ n10951 ^ n5469 ;
  assign n21631 = n19757 ^ n6502 ^ 1'b0 ;
  assign n21632 = n13301 ^ n5254 ^ n139 ;
  assign n21633 = n21385 ^ n9475 ^ 1'b0 ;
  assign n21634 = n17465 | n21633 ;
  assign n21635 = n12919 | n21634 ;
  assign n21636 = n21635 ^ n14089 ^ 1'b0 ;
  assign n21637 = n5498 & ~n14232 ;
  assign n21638 = n21637 ^ n21282 ^ 1'b0 ;
  assign n21640 = n360 & ~n12782 ;
  assign n21641 = n4939 & ~n21640 ;
  assign n21639 = n7172 | n18222 ;
  assign n21642 = n21641 ^ n21639 ^ 1'b0 ;
  assign n21643 = n10645 ^ n3742 ^ n2824 ;
  assign n21644 = n2898 | n4351 ;
  assign n21645 = n21643 | n21644 ;
  assign n21646 = ~n12723 & n12828 ;
  assign n21647 = ( n6960 & ~n9662 ) | ( n6960 & n11360 ) | ( ~n9662 & n11360 ) ;
  assign n21648 = n21647 ^ n9546 ^ 1'b0 ;
  assign n21649 = n8479 & ~n11288 ;
  assign n21650 = ~n3411 & n5079 ;
  assign n21651 = n21650 ^ n14846 ^ 1'b0 ;
  assign n21652 = ~n12172 & n12778 ;
  assign n21653 = n21652 ^ n17580 ^ 1'b0 ;
  assign n21654 = n18225 ^ n11292 ^ n8706 ;
  assign n21655 = ~n5094 & n19803 ;
  assign n21656 = n13832 ^ n9956 ^ 1'b0 ;
  assign n21657 = ~n4859 & n21656 ;
  assign n21658 = n21657 ^ n18297 ^ n3532 ;
  assign n21659 = n2274 & n7062 ;
  assign n21660 = ( n8636 & n11999 ) | ( n8636 & ~n21659 ) | ( n11999 & ~n21659 ) ;
  assign n21661 = n21660 ^ n1038 ^ 1'b0 ;
  assign n21662 = n13251 & ~n20553 ;
  assign n21663 = ~n7698 & n21662 ;
  assign n21664 = ( n9511 & ~n14022 ) | ( n9511 & n21304 ) | ( ~n14022 & n21304 ) ;
  assign n21665 = n15039 ^ n9295 ^ n6236 ;
  assign n21666 = n20884 ^ n9649 ^ 1'b0 ;
  assign n21667 = n10394 ^ n1466 ^ 1'b0 ;
  assign n21668 = ~n18699 & n21667 ;
  assign n21669 = n2600 & n11733 ;
  assign n21670 = n21668 & n21669 ;
  assign n21671 = n13411 & ~n17992 ;
  assign n21672 = n17870 & n21671 ;
  assign n21673 = n17944 ^ x96 ^ 1'b0 ;
  assign n21674 = n21673 ^ n14473 ^ 1'b0 ;
  assign n21675 = ( n7589 & ~n10497 ) | ( n7589 & n16190 ) | ( ~n10497 & n16190 ) ;
  assign n21676 = n5188 ^ n2046 ^ 1'b0 ;
  assign n21677 = n21676 ^ n14972 ^ x98 ;
  assign n21678 = n21677 ^ n13701 ^ n1581 ;
  assign n21679 = n5795 ^ n1609 ^ 1'b0 ;
  assign n21680 = n14381 & n21679 ;
  assign n21681 = n21680 ^ n20449 ^ 1'b0 ;
  assign n21682 = n21227 ^ n4864 ^ 1'b0 ;
  assign n21685 = ( n566 & ~n5133 ) | ( n566 & n6402 ) | ( ~n5133 & n6402 ) ;
  assign n21686 = ~n1253 & n21685 ;
  assign n21683 = n4928 | n10456 ;
  assign n21684 = n8618 | n21683 ;
  assign n21687 = n21686 ^ n21684 ^ 1'b0 ;
  assign n21688 = ( n511 & n9656 ) | ( n511 & n14432 ) | ( n9656 & n14432 ) ;
  assign n21689 = ~n15144 & n16699 ;
  assign n21690 = n5739 | n9938 ;
  assign n21691 = n21690 ^ n16735 ^ 1'b0 ;
  assign n21692 = n21691 ^ n13140 ^ n6497 ;
  assign n21693 = n3190 & ~n11886 ;
  assign n21694 = n15180 & ~n19238 ;
  assign n21695 = n21694 ^ n968 ^ 1'b0 ;
  assign n21696 = n18206 ^ n4461 ^ 1'b0 ;
  assign n21697 = n4784 | n15804 ;
  assign n21698 = n16408 & ~n21697 ;
  assign n21699 = ~n9021 & n21698 ;
  assign n21700 = n5136 ^ n2898 ^ 1'b0 ;
  assign n21701 = n4356 & ~n21700 ;
  assign n21702 = n21701 ^ n20527 ^ 1'b0 ;
  assign n21703 = ~n7473 & n21702 ;
  assign n21704 = ( n7108 & n11419 ) | ( n7108 & ~n14055 ) | ( n11419 & ~n14055 ) ;
  assign n21705 = ~n7417 & n16516 ;
  assign n21706 = n18902 ^ n13858 ^ 1'b0 ;
  assign n21707 = n2641 & n21706 ;
  assign n21708 = n1287 ^ n259 ^ 1'b0 ;
  assign n21709 = n21708 ^ n10663 ^ 1'b0 ;
  assign n21710 = n203 & ~n7368 ;
  assign n21711 = ~n21709 & n21710 ;
  assign n21712 = n752 & ~n3338 ;
  assign n21713 = n21712 ^ n18596 ^ 1'b0 ;
  assign n21714 = n1456 & n4089 ;
  assign n21715 = ~n1801 & n21714 ;
  assign n21716 = ( n468 & n7948 ) | ( n468 & n21715 ) | ( n7948 & n21715 ) ;
  assign n21717 = n16167 ^ n5093 ^ 1'b0 ;
  assign n21718 = n19392 ^ n14257 ^ n11093 ;
  assign n21719 = n11669 & ~n20809 ;
  assign n21720 = n21719 ^ n12662 ^ 1'b0 ;
  assign n21721 = n8832 ^ n7313 ^ n323 ;
  assign n21722 = ~n2813 & n8733 ;
  assign n21723 = n21722 ^ n10730 ^ 1'b0 ;
  assign n21724 = n21723 ^ n11538 ^ n11531 ;
  assign n21725 = n21724 ^ n12290 ^ x73 ;
  assign n21726 = n421 & ~n21725 ;
  assign n21727 = n21721 & n21726 ;
  assign n21728 = n15376 ^ n6632 ^ 1'b0 ;
  assign n21729 = n16827 ^ n3436 ^ x63 ;
  assign n21730 = ~n2937 & n8060 ;
  assign n21731 = n6759 | n6892 ;
  assign n21732 = n5645 & n21731 ;
  assign n21733 = n21732 ^ n13802 ^ 1'b0 ;
  assign n21734 = ~n7188 & n21733 ;
  assign n21735 = n8338 ^ n2681 ^ 1'b0 ;
  assign n21736 = n21734 & n21735 ;
  assign n21737 = ~n20018 & n20684 ;
  assign n21738 = n19545 ^ n11068 ^ 1'b0 ;
  assign n21739 = ~n2815 & n21738 ;
  assign n21740 = ~n8279 & n11944 ;
  assign n21741 = n21257 ^ n3561 ^ 1'b0 ;
  assign n21742 = ~n21740 & n21741 ;
  assign n21743 = n21742 ^ n7002 ^ x70 ;
  assign n21744 = n7284 & n15480 ;
  assign n21745 = n21579 ^ x48 ^ 1'b0 ;
  assign n21746 = ( n7180 & n10854 ) | ( n7180 & ~n18945 ) | ( n10854 & ~n18945 ) ;
  assign n21747 = n4334 & n5826 ;
  assign n21748 = ~n10991 & n21747 ;
  assign n21749 = ( n16834 & n19068 ) | ( n16834 & ~n21748 ) | ( n19068 & ~n21748 ) ;
  assign n21750 = n7633 ^ n4825 ^ 1'b0 ;
  assign n21751 = n923 & ~n16634 ;
  assign n21752 = ~n3357 & n21751 ;
  assign n21753 = n21752 ^ n15956 ^ 1'b0 ;
  assign n21754 = n15976 & n21753 ;
  assign n21755 = n21754 ^ n12686 ^ x123 ;
  assign n21756 = n9492 | n12327 ;
  assign n21757 = n3612 | n13902 ;
  assign n21758 = n21757 ^ n2833 ^ 1'b0 ;
  assign n21759 = ~n631 & n21758 ;
  assign n21760 = n21759 ^ n354 ^ 1'b0 ;
  assign n21761 = n3276 | n11222 ;
  assign n21762 = n3337 & ~n21761 ;
  assign n21763 = n21762 ^ n12388 ^ 1'b0 ;
  assign n21764 = ( n1410 & ~n8785 ) | ( n1410 & n21763 ) | ( ~n8785 & n21763 ) ;
  assign n21765 = ( ~n6799 & n8490 ) | ( ~n6799 & n21764 ) | ( n8490 & n21764 ) ;
  assign n21766 = ( n15131 & n18057 ) | ( n15131 & n21765 ) | ( n18057 & n21765 ) ;
  assign n21767 = n21766 ^ n9608 ^ 1'b0 ;
  assign n21768 = ( x77 & n1426 ) | ( x77 & n16730 ) | ( n1426 & n16730 ) ;
  assign n21769 = n2701 | n7521 ;
  assign n21770 = n8803 | n17375 ;
  assign n21771 = ( n17359 & ~n21769 ) | ( n17359 & n21770 ) | ( ~n21769 & n21770 ) ;
  assign n21772 = n1743 & n21771 ;
  assign n21773 = n12829 ^ n11849 ^ 1'b0 ;
  assign n21774 = n14954 ^ n13706 ^ 1'b0 ;
  assign n21775 = ~n3491 & n21774 ;
  assign n21776 = ~n12037 & n21775 ;
  assign n21777 = n9093 | n13769 ;
  assign n21778 = n1927 & ~n21777 ;
  assign n21779 = n16923 | n21778 ;
  assign n21780 = n21779 ^ n13939 ^ 1'b0 ;
  assign n21781 = n1519 | n4321 ;
  assign n21782 = n21780 & ~n21781 ;
  assign n21783 = n11473 ^ n9482 ^ n9295 ;
  assign n21784 = n3808 | n7433 ;
  assign n21785 = n21784 ^ n16954 ^ n5248 ;
  assign n21786 = n4778 & n21785 ;
  assign n21787 = ( ~n8702 & n10754 ) | ( ~n8702 & n19271 ) | ( n10754 & n19271 ) ;
  assign n21788 = ~n12432 & n14972 ;
  assign n21789 = n13818 & n17808 ;
  assign n21790 = ~n3120 & n4177 ;
  assign n21791 = n998 & ~n21551 ;
  assign n21795 = n16117 ^ n752 ^ 1'b0 ;
  assign n21796 = n7987 & ~n21795 ;
  assign n21792 = n8143 ^ n1405 ^ 1'b0 ;
  assign n21793 = n306 & n3095 ;
  assign n21794 = n21792 & n21793 ;
  assign n21797 = n21796 ^ n21794 ^ 1'b0 ;
  assign n21798 = n21545 ^ n19817 ^ 1'b0 ;
  assign n21799 = n15546 & n21798 ;
  assign n21800 = n7121 & n7976 ;
  assign n21801 = n2654 & ~n8514 ;
  assign n21802 = n7354 & n21801 ;
  assign n21803 = n17166 & ~n21802 ;
  assign n21804 = ~n21053 & n21803 ;
  assign n21805 = n9441 ^ n6438 ^ 1'b0 ;
  assign n21806 = n1058 & ~n21805 ;
  assign n21807 = n5938 ^ n1959 ^ 1'b0 ;
  assign n21808 = ( n1843 & n3467 ) | ( n1843 & ~n18262 ) | ( n3467 & ~n18262 ) ;
  assign n21809 = n21807 & ~n21808 ;
  assign n21810 = n21809 ^ n5953 ^ 1'b0 ;
  assign n21811 = ( n15920 & n20348 ) | ( n15920 & n21810 ) | ( n20348 & n21810 ) ;
  assign n21812 = n20373 ^ n19515 ^ n15196 ;
  assign n21813 = n21812 ^ n20235 ^ n19912 ;
  assign n21814 = n16769 ^ n12995 ^ n7863 ;
  assign n21815 = n12572 | n21814 ;
  assign n21816 = n2665 & n18333 ;
  assign n21817 = n21483 ^ n17804 ^ n4520 ;
  assign n21818 = n21817 ^ n4201 ^ 1'b0 ;
  assign n21819 = n21818 ^ n15288 ^ 1'b0 ;
  assign n21820 = n21816 & n21819 ;
  assign n21826 = n9034 ^ n4160 ^ n1199 ;
  assign n21822 = n17776 ^ n3461 ^ 1'b0 ;
  assign n21823 = n746 | n21822 ;
  assign n21824 = n3364 & ~n21823 ;
  assign n21825 = n21824 ^ n4308 ^ n3842 ;
  assign n21821 = n15746 ^ n10949 ^ n3065 ;
  assign n21827 = n21826 ^ n21825 ^ n21821 ;
  assign n21828 = n5137 ^ n740 ^ 1'b0 ;
  assign n21829 = n21828 ^ n21822 ^ n11071 ;
  assign n21830 = n2619 & ~n21829 ;
  assign n21831 = n7230 ^ n5975 ^ n5104 ;
  assign n21832 = n8991 & ~n20020 ;
  assign n21833 = n8744 & n19664 ;
  assign n21834 = n21833 ^ n7360 ^ 1'b0 ;
  assign n21835 = ( n744 & n11677 ) | ( n744 & n21834 ) | ( n11677 & n21834 ) ;
  assign n21836 = n10417 | n21835 ;
  assign n21837 = ~n2352 & n18947 ;
  assign n21838 = ~x37 & n21837 ;
  assign n21839 = ~n8699 & n16676 ;
  assign n21840 = n21839 ^ n5719 ^ 1'b0 ;
  assign n21841 = ~n3696 & n5739 ;
  assign n21842 = n21841 ^ n1043 ^ 1'b0 ;
  assign n21843 = ~n1608 & n21842 ;
  assign n21844 = ( n6672 & n13181 ) | ( n6672 & ~n17324 ) | ( n13181 & ~n17324 ) ;
  assign n21845 = n9805 ^ n6475 ^ 1'b0 ;
  assign n21846 = n15946 ^ n12715 ^ n4889 ;
  assign n21847 = ~n1132 & n3874 ;
  assign n21848 = ~n7659 & n21847 ;
  assign n21849 = n21846 & n21848 ;
  assign n21850 = n8516 | n16304 ;
  assign n21851 = n20718 ^ n8501 ^ n7891 ;
  assign n21852 = ~n4990 & n11649 ;
  assign n21853 = n16641 & n21852 ;
  assign n21854 = ~n7280 & n16555 ;
  assign n21855 = ( n17673 & n21853 ) | ( n17673 & n21854 ) | ( n21853 & n21854 ) ;
  assign n21856 = ( n861 & n13152 ) | ( n861 & n14641 ) | ( n13152 & n14641 ) ;
  assign n21857 = n17626 ^ n2428 ^ 1'b0 ;
  assign n21858 = ~n5749 & n21857 ;
  assign n21859 = ( n5824 & n21856 ) | ( n5824 & n21858 ) | ( n21856 & n21858 ) ;
  assign n21861 = n7076 ^ n2237 ^ 1'b0 ;
  assign n21862 = ~n1824 & n21861 ;
  assign n21860 = n14015 | n21553 ;
  assign n21863 = n21862 ^ n21860 ^ 1'b0 ;
  assign n21864 = n11397 ^ n4875 ^ 1'b0 ;
  assign n21865 = n19489 | n21864 ;
  assign n21866 = n21865 ^ n9862 ^ 1'b0 ;
  assign n21867 = n11925 & ~n14702 ;
  assign n21868 = n17974 ^ n16410 ^ n5398 ;
  assign n21869 = n4690 & ~n5991 ;
  assign n21870 = n3118 & ~n9544 ;
  assign n21871 = n5147 & n21870 ;
  assign n21872 = n10439 ^ n5915 ^ n390 ;
  assign n21873 = n18429 | n21872 ;
  assign n21874 = n9928 | n17953 ;
  assign n21875 = n2018 | n21874 ;
  assign n21876 = n16852 & n21875 ;
  assign n21877 = n6639 & n21876 ;
  assign n21878 = n13507 ^ x92 ^ 1'b0 ;
  assign n21879 = n4468 & ~n7501 ;
  assign n21880 = n1135 & n21879 ;
  assign n21881 = n5579 & ~n11674 ;
  assign n21882 = n2558 & ~n21881 ;
  assign n21883 = ( n5787 & n21880 ) | ( n5787 & ~n21882 ) | ( n21880 & ~n21882 ) ;
  assign n21884 = n1418 ^ x85 ^ 1'b0 ;
  assign n21885 = n6249 ^ n3056 ^ n2263 ;
  assign n21886 = n4377 & ~n6657 ;
  assign n21887 = n21885 & n21886 ;
  assign n21888 = n21887 ^ n4735 ^ 1'b0 ;
  assign n21889 = ( ~n17815 & n21884 ) | ( ~n17815 & n21888 ) | ( n21884 & n21888 ) ;
  assign n21890 = n21176 ^ n4346 ^ 1'b0 ;
  assign n21891 = n8899 | n21890 ;
  assign n21893 = n3942 ^ n3612 ^ 1'b0 ;
  assign n21894 = n21893 ^ n1794 ^ 1'b0 ;
  assign n21895 = ~n7792 & n21894 ;
  assign n21892 = n10512 & ~n14156 ;
  assign n21896 = n21895 ^ n21892 ^ 1'b0 ;
  assign n21897 = n18171 ^ n2388 ^ 1'b0 ;
  assign n21901 = n9035 ^ n6330 ^ n442 ;
  assign n21899 = n6279 | n9539 ;
  assign n21900 = n350 | n21899 ;
  assign n21902 = n21901 ^ n21900 ^ n9984 ;
  assign n21898 = n9977 & ~n10077 ;
  assign n21903 = n21902 ^ n21898 ^ 1'b0 ;
  assign n21906 = n349 & n1912 ;
  assign n21905 = ( n5237 & ~n6046 ) | ( n5237 & n19400 ) | ( ~n6046 & n19400 ) ;
  assign n21904 = n5283 ^ n4914 ^ 1'b0 ;
  assign n21907 = n21906 ^ n21905 ^ n21904 ;
  assign n21908 = n15233 ^ n13929 ^ n11875 ;
  assign n21909 = n21908 ^ n7943 ^ n4270 ;
  assign n21910 = n21909 ^ n10179 ^ 1'b0 ;
  assign n21911 = n15237 ^ n14752 ^ 1'b0 ;
  assign n21912 = x42 & ~n3276 ;
  assign n21913 = ~n1236 & n21912 ;
  assign n21914 = n8948 & n21657 ;
  assign n21915 = ( n1501 & n21913 ) | ( n1501 & n21914 ) | ( n21913 & n21914 ) ;
  assign n21916 = n5798 | n21915 ;
  assign n21917 = n21916 ^ n6201 ^ 1'b0 ;
  assign n21918 = n12680 & n15070 ;
  assign n21919 = n21918 ^ n8456 ^ 1'b0 ;
  assign n21920 = n7903 & ~n15087 ;
  assign n21921 = n21919 & n21920 ;
  assign n21922 = n12001 ^ n7508 ^ 1'b0 ;
  assign n21927 = n16762 ^ n5573 ^ 1'b0 ;
  assign n21923 = n2100 | n10185 ;
  assign n21924 = n21923 ^ n6493 ^ 1'b0 ;
  assign n21925 = n20486 ^ n11932 ^ 1'b0 ;
  assign n21926 = n21924 & n21925 ;
  assign n21928 = n21927 ^ n21926 ^ 1'b0 ;
  assign n21929 = ( n20321 & n21922 ) | ( n20321 & ~n21928 ) | ( n21922 & ~n21928 ) ;
  assign n21930 = n9369 ^ n5365 ^ 1'b0 ;
  assign n21931 = n404 & n21930 ;
  assign n21932 = n7783 ^ n4240 ^ 1'b0 ;
  assign n21933 = ~n5889 & n21932 ;
  assign n21934 = n1835 & n16258 ;
  assign n21935 = n21934 ^ n12593 ^ 1'b0 ;
  assign n21936 = ~n21933 & n21935 ;
  assign n21937 = ~n5840 & n21936 ;
  assign n21938 = ~n6233 & n21937 ;
  assign n21939 = n21938 ^ n9488 ^ n5353 ;
  assign n21940 = n3001 & n12328 ;
  assign n21941 = ~n16662 & n21940 ;
  assign n21942 = n11875 ^ n6093 ^ 1'b0 ;
  assign n21943 = n13874 & ~n21942 ;
  assign n21944 = n6438 & ~n18744 ;
  assign n21945 = n12147 ^ n10688 ^ 1'b0 ;
  assign n21946 = n9105 & n21945 ;
  assign n21947 = ( n10799 & n14005 ) | ( n10799 & n18044 ) | ( n14005 & n18044 ) ;
  assign n21948 = ( n2121 & n9268 ) | ( n2121 & n9715 ) | ( n9268 & n9715 ) ;
  assign n21949 = n8821 & n19366 ;
  assign n21955 = ~n9811 & n10846 ;
  assign n21956 = n8610 & n21955 ;
  assign n21950 = n18096 & ~n20158 ;
  assign n21951 = ~n3701 & n21950 ;
  assign n21952 = n10304 & ~n21951 ;
  assign n21953 = n21952 ^ n7015 ^ 1'b0 ;
  assign n21954 = n6804 & ~n21953 ;
  assign n21957 = n21956 ^ n21954 ^ 1'b0 ;
  assign n21958 = n7905 ^ n5475 ^ n5215 ;
  assign n21959 = n9163 & ~n21958 ;
  assign n21960 = n7049 & n8399 ;
  assign n21961 = ( n8174 & n8467 ) | ( n8174 & n13078 ) | ( n8467 & n13078 ) ;
  assign n21962 = ~n7790 & n13416 ;
  assign n21963 = ~n11600 & n17526 ;
  assign n21964 = n8672 & ~n18205 ;
  assign n21965 = n21964 ^ n852 ^ 1'b0 ;
  assign n21966 = n9595 ^ n1758 ^ 1'b0 ;
  assign n21967 = ( n4285 & n4605 ) | ( n4285 & ~n13012 ) | ( n4605 & ~n13012 ) ;
  assign n21968 = ~n21966 & n21967 ;
  assign n21969 = n11812 ^ n1569 ^ 1'b0 ;
  assign n21970 = ~n5506 & n10945 ;
  assign n21971 = n12825 & n21825 ;
  assign n21972 = n21971 ^ n10613 ^ 1'b0 ;
  assign n21973 = ~n11032 & n18585 ;
  assign n21974 = n17880 ^ n5714 ^ 1'b0 ;
  assign n21975 = n4774 & n13865 ;
  assign n21976 = n21975 ^ n1628 ^ 1'b0 ;
  assign n21977 = n6830 & ~n21976 ;
  assign n21978 = ~n4188 & n20623 ;
  assign n21979 = n5596 & ~n9824 ;
  assign n21980 = n21979 ^ n6656 ^ 1'b0 ;
  assign n21981 = ~n5832 & n19430 ;
  assign n21982 = ~n19953 & n21981 ;
  assign n21983 = n14013 ^ n1700 ^ 1'b0 ;
  assign n21984 = n2031 & ~n21983 ;
  assign n21985 = n1110 & n21071 ;
  assign n21986 = n1100 ^ n1055 ^ 1'b0 ;
  assign n21987 = n18431 ^ n2163 ^ n1154 ;
  assign n21988 = n21987 ^ n383 ^ 1'b0 ;
  assign n21989 = n21986 | n21988 ;
  assign n21991 = n17561 ^ n10780 ^ n8621 ;
  assign n21990 = n2607 & ~n17228 ;
  assign n21992 = n21991 ^ n21990 ^ 1'b0 ;
  assign n21993 = n20813 | n21992 ;
  assign n21994 = n6382 | n21993 ;
  assign n21995 = ~n10496 & n21994 ;
  assign n21996 = ( n4727 & ~n10677 ) | ( n4727 & n12248 ) | ( ~n10677 & n12248 ) ;
  assign n21997 = ~n511 & n8259 ;
  assign n21998 = ~n21996 & n21997 ;
  assign n21999 = ( n6553 & n13933 ) | ( n6553 & ~n21998 ) | ( n13933 & ~n21998 ) ;
  assign n22000 = ~n2430 & n12642 ;
  assign n22002 = n1619 | n14447 ;
  assign n22003 = n12123 | n22002 ;
  assign n22001 = n4615 & ~n7116 ;
  assign n22004 = n22003 ^ n22001 ^ 1'b0 ;
  assign n22005 = ~n5529 & n13111 ;
  assign n22006 = n22005 ^ n2298 ^ 1'b0 ;
  assign n22007 = x75 & n22006 ;
  assign n22008 = n867 & n22007 ;
  assign n22009 = ( n2174 & n6817 ) | ( n2174 & n7115 ) | ( n6817 & n7115 ) ;
  assign n22010 = n7772 ^ n5887 ^ n5664 ;
  assign n22011 = ~n22009 & n22010 ;
  assign n22012 = ~n428 & n22011 ;
  assign n22013 = n20497 ^ n3267 ^ n2592 ;
  assign n22014 = n19647 ^ n1427 ^ 1'b0 ;
  assign n22015 = n5289 & ~n7205 ;
  assign n22016 = n1669 & n22015 ;
  assign n22017 = ~n10030 & n22016 ;
  assign n22018 = ~n2420 & n16053 ;
  assign n22019 = n17174 ^ n15492 ^ 1'b0 ;
  assign n22020 = n4511 & n11910 ;
  assign n22021 = n22019 & ~n22020 ;
  assign n22022 = n721 & ~n14033 ;
  assign n22024 = n11190 ^ n9588 ^ 1'b0 ;
  assign n22023 = n9295 ^ n5202 ^ 1'b0 ;
  assign n22025 = n22024 ^ n22023 ^ x40 ;
  assign n22028 = n2173 & n21426 ;
  assign n22029 = ~n3553 & n22028 ;
  assign n22026 = n18634 ^ n14388 ^ 1'b0 ;
  assign n22027 = n1962 & ~n22026 ;
  assign n22030 = n22029 ^ n22027 ^ 1'b0 ;
  assign n22036 = n586 | n6155 ;
  assign n22037 = n20470 & ~n22036 ;
  assign n22032 = n5325 & n7374 ;
  assign n22033 = n22032 ^ n1634 ^ 1'b0 ;
  assign n22031 = ~n3793 & n13194 ;
  assign n22034 = n22033 ^ n22031 ^ 1'b0 ;
  assign n22035 = n14143 & ~n22034 ;
  assign n22038 = n22037 ^ n22035 ^ 1'b0 ;
  assign n22039 = n7924 & ~n12681 ;
  assign n22040 = ~n17958 & n22039 ;
  assign n22041 = n22040 ^ n14521 ^ n4506 ;
  assign n22042 = n22041 ^ n18355 ^ 1'b0 ;
  assign n22043 = ~n10506 & n16671 ;
  assign n22044 = n22043 ^ n4857 ^ 1'b0 ;
  assign n22045 = ~n514 & n10784 ;
  assign n22046 = n22045 ^ n3277 ^ 1'b0 ;
  assign n22047 = n21189 ^ n13615 ^ n10872 ;
  assign n22048 = n7291 ^ n3611 ^ 1'b0 ;
  assign n22049 = n13797 & n22048 ;
  assign n22050 = n12919 | n13724 ;
  assign n22051 = n22050 ^ x98 ^ 1'b0 ;
  assign n22052 = n16455 ^ n7617 ^ 1'b0 ;
  assign n22053 = ~n15891 & n22052 ;
  assign n22054 = ~n4148 & n10232 ;
  assign n22055 = n1591 & ~n22054 ;
  assign n22056 = n22055 ^ n13154 ^ 1'b0 ;
  assign n22057 = ~n390 & n22056 ;
  assign n22058 = ~n4022 & n22057 ;
  assign n22059 = n2206 & n5110 ;
  assign n22060 = ~n8502 & n22059 ;
  assign n22061 = n22060 ^ n15068 ^ n6101 ;
  assign n22062 = n9887 ^ n6947 ^ n6170 ;
  assign n22063 = n16303 ^ n8562 ^ 1'b0 ;
  assign n22064 = n22063 ^ n13468 ^ n12715 ;
  assign n22065 = n22064 ^ n12501 ^ 1'b0 ;
  assign n22066 = n3658 & n22065 ;
  assign n22067 = n378 | n2659 ;
  assign n22068 = n19934 ^ n8816 ^ 1'b0 ;
  assign n22069 = ~n7330 & n22068 ;
  assign n22070 = ~n1182 & n7499 ;
  assign n22071 = n22070 ^ n9949 ^ 1'b0 ;
  assign n22072 = ( n14683 & n16879 ) | ( n14683 & ~n22071 ) | ( n16879 & ~n22071 ) ;
  assign n22073 = n22072 ^ n16499 ^ 1'b0 ;
  assign n22075 = n17604 ^ n6371 ^ n2378 ;
  assign n22074 = n12883 ^ n6130 ^ n3816 ;
  assign n22076 = n22075 ^ n22074 ^ n9945 ;
  assign n22077 = n12235 & ~n12899 ;
  assign n22078 = n22077 ^ n13759 ^ n11478 ;
  assign n22082 = ( n798 & n3502 ) | ( n798 & ~n8342 ) | ( n3502 & ~n8342 ) ;
  assign n22083 = n2886 & ~n10547 ;
  assign n22084 = ( n1283 & n22082 ) | ( n1283 & ~n22083 ) | ( n22082 & ~n22083 ) ;
  assign n22079 = n5937 & n12229 ;
  assign n22080 = n22079 ^ n310 ^ 1'b0 ;
  assign n22081 = ( n3527 & ~n9846 ) | ( n3527 & n22080 ) | ( ~n9846 & n22080 ) ;
  assign n22085 = n22084 ^ n22081 ^ n3463 ;
  assign n22086 = n7871 & n15221 ;
  assign n22087 = n7175 & n22086 ;
  assign n22088 = n12123 & ~n13865 ;
  assign n22089 = ~n824 & n22088 ;
  assign n22090 = ~n9464 & n22089 ;
  assign n22092 = n10880 ^ n6362 ^ 1'b0 ;
  assign n22093 = n7531 & ~n22092 ;
  assign n22091 = n18761 ^ n13045 ^ 1'b0 ;
  assign n22094 = n22093 ^ n22091 ^ n2231 ;
  assign n22095 = n7351 & ~n11988 ;
  assign n22096 = n5307 & n22095 ;
  assign n22097 = ( n2033 & n14548 ) | ( n2033 & ~n22096 ) | ( n14548 & ~n22096 ) ;
  assign n22098 = n22097 ^ n16598 ^ n3134 ;
  assign n22099 = ( n6060 & n11997 ) | ( n6060 & ~n16396 ) | ( n11997 & ~n16396 ) ;
  assign n22100 = ~n289 & n2168 ;
  assign n22101 = n436 & n20473 ;
  assign n22102 = n22101 ^ n15892 ^ 1'b0 ;
  assign n22103 = n7641 & n21977 ;
  assign n22104 = ~n10970 & n22103 ;
  assign n22105 = n9984 ^ n2636 ^ 1'b0 ;
  assign n22106 = n10929 & n11210 ;
  assign n22107 = ( n2019 & n4739 ) | ( n2019 & ~n20417 ) | ( n4739 & ~n20417 ) ;
  assign n22108 = n3296 ^ n2165 ^ 1'b0 ;
  assign n22109 = ~n3470 & n12747 ;
  assign n22110 = n2929 | n14975 ;
  assign n22111 = n20335 | n22110 ;
  assign n22112 = n10164 ^ n4582 ^ 1'b0 ;
  assign n22113 = n13931 & n22112 ;
  assign n22114 = ~n9145 & n22113 ;
  assign n22115 = ~n6644 & n11300 ;
  assign n22116 = n16275 ^ n9203 ^ 1'b0 ;
  assign n22117 = n22115 & ~n22116 ;
  assign n22118 = n17064 ^ n7257 ^ 1'b0 ;
  assign n22119 = n22117 & n22118 ;
  assign n22120 = ( n971 & n10842 ) | ( n971 & n11646 ) | ( n10842 & n11646 ) ;
  assign n22121 = n5798 ^ n4377 ^ n2125 ;
  assign n22122 = n22121 ^ n14177 ^ n11239 ;
  assign n22123 = n15211 ^ n14149 ^ 1'b0 ;
  assign n22124 = n13873 & n22123 ;
  assign n22125 = n22124 ^ n20283 ^ 1'b0 ;
  assign n22126 = ~n10183 & n13222 ;
  assign n22127 = n9323 & n13550 ;
  assign n22128 = ~n12234 & n22127 ;
  assign n22129 = ~n15319 & n16162 ;
  assign n22130 = n21214 & n22129 ;
  assign n22131 = n22130 ^ n9556 ^ 1'b0 ;
  assign n22132 = ( n855 & ~n19115 ) | ( n855 & n19180 ) | ( ~n19115 & n19180 ) ;
  assign n22133 = ~n20150 & n20364 ;
  assign n22134 = ~n849 & n13706 ;
  assign n22136 = n8568 | n16811 ;
  assign n22137 = n1341 & ~n22136 ;
  assign n22135 = n4365 & n17154 ;
  assign n22138 = n22137 ^ n22135 ^ 1'b0 ;
  assign n22139 = n8779 & n15303 ;
  assign n22140 = n14096 ^ n12593 ^ 1'b0 ;
  assign n22141 = n17941 & n22140 ;
  assign n22142 = n13600 ^ n9406 ^ 1'b0 ;
  assign n22143 = n16337 | n22142 ;
  assign n22144 = ~n5954 & n6252 ;
  assign n22145 = n22144 ^ n369 ^ 1'b0 ;
  assign n22146 = ( n10448 & ~n16062 ) | ( n10448 & n22145 ) | ( ~n16062 & n22145 ) ;
  assign n22147 = n22146 ^ n16870 ^ n13202 ;
  assign n22148 = n21844 ^ n635 ^ 1'b0 ;
  assign n22149 = ~n8239 & n20490 ;
  assign n22150 = n19996 & n22149 ;
  assign n22152 = n18861 ^ n6233 ^ 1'b0 ;
  assign n22151 = ~x89 & n5212 ;
  assign n22153 = n22152 ^ n22151 ^ n16373 ;
  assign n22154 = n22153 ^ n12097 ^ n8274 ;
  assign n22155 = ( ~n4653 & n13406 ) | ( ~n4653 & n20954 ) | ( n13406 & n20954 ) ;
  assign n22156 = n22154 | n22155 ;
  assign n22157 = ( n1942 & ~n2175 ) | ( n1942 & n15168 ) | ( ~n2175 & n15168 ) ;
  assign n22159 = n10098 | n19269 ;
  assign n22158 = n2317 | n19665 ;
  assign n22160 = n22159 ^ n22158 ^ n3750 ;
  assign n22161 = n16747 & ~n18300 ;
  assign n22162 = ~n13117 & n22161 ;
  assign n22163 = ( n9931 & n10139 ) | ( n9931 & ~n22088 ) | ( n10139 & ~n22088 ) ;
  assign n22164 = n14591 ^ n7855 ^ n2387 ;
  assign n22165 = ~n4315 & n15940 ;
  assign n22166 = n9746 & n22165 ;
  assign n22167 = n8406 | n22166 ;
  assign n22168 = n22167 ^ n15499 ^ 1'b0 ;
  assign n22169 = n22164 & n22168 ;
  assign n22170 = ( n11209 & n22163 ) | ( n11209 & n22169 ) | ( n22163 & n22169 ) ;
  assign n22171 = n7618 & n8447 ;
  assign n22172 = n22171 ^ n17778 ^ 1'b0 ;
  assign n22173 = ~n376 & n2836 ;
  assign n22174 = n2338 & n22173 ;
  assign n22175 = n22174 ^ n11457 ^ 1'b0 ;
  assign n22176 = n21507 | n22175 ;
  assign n22177 = n9155 ^ n7990 ^ n1617 ;
  assign n22178 = n22177 ^ x79 ^ 1'b0 ;
  assign n22179 = ~n22176 & n22178 ;
  assign n22180 = ~n18803 & n22179 ;
  assign n22181 = ~n22172 & n22180 ;
  assign n22182 = n10947 | n19329 ;
  assign n22183 = ~n2006 & n13894 ;
  assign n22184 = n5023 | n22183 ;
  assign n22185 = n22184 ^ n11199 ^ 1'b0 ;
  assign n22186 = ~n11701 & n22019 ;
  assign n22187 = n10562 ^ n7998 ^ n4285 ;
  assign n22188 = ( n1429 & n8809 ) | ( n1429 & n22187 ) | ( n8809 & n22187 ) ;
  assign n22189 = n2751 & n22188 ;
  assign n22190 = n22189 ^ n6969 ^ 1'b0 ;
  assign n22191 = n9273 ^ n5746 ^ n1480 ;
  assign n22192 = ~n4970 & n9331 ;
  assign n22193 = ~n22191 & n22192 ;
  assign n22194 = n22193 ^ n11573 ^ n5449 ;
  assign n22195 = n13605 & n14086 ;
  assign n22196 = n22195 ^ n1327 ^ 1'b0 ;
  assign n22197 = n22196 ^ n6960 ^ 1'b0 ;
  assign n22199 = x20 & ~n2097 ;
  assign n22198 = n13060 & ~n16514 ;
  assign n22200 = n22199 ^ n22198 ^ 1'b0 ;
  assign n22201 = n22200 ^ n16053 ^ 1'b0 ;
  assign n22202 = n5714 | n10334 ;
  assign n22203 = n22202 ^ n16358 ^ 1'b0 ;
  assign n22204 = ( n12924 & n17369 ) | ( n12924 & n22203 ) | ( n17369 & n22203 ) ;
  assign n22205 = n22204 ^ n8931 ^ 1'b0 ;
  assign n22208 = n5859 & ~n19575 ;
  assign n22206 = n21979 ^ n11002 ^ 1'b0 ;
  assign n22207 = n22206 ^ n15996 ^ n1530 ;
  assign n22209 = n22208 ^ n22207 ^ n18729 ;
  assign n22210 = n21232 ^ n2149 ^ 1'b0 ;
  assign n22214 = n5965 ^ n3835 ^ n3668 ;
  assign n22215 = n3169 & ~n22214 ;
  assign n22211 = n6304 ^ n615 ^ 1'b0 ;
  assign n22212 = n1530 | n22211 ;
  assign n22213 = n2091 & ~n22212 ;
  assign n22216 = n22215 ^ n22213 ^ 1'b0 ;
  assign n22217 = n22216 ^ n11412 ^ 1'b0 ;
  assign n22218 = ~n696 & n22217 ;
  assign n22219 = n21593 & n22218 ;
  assign n22220 = n6493 | n13378 ;
  assign n22221 = n22220 ^ n13891 ^ 1'b0 ;
  assign n22222 = ( ~n12108 & n21460 ) | ( ~n12108 & n22221 ) | ( n21460 & n22221 ) ;
  assign n22223 = n20247 ^ n14643 ^ 1'b0 ;
  assign n22224 = ~n15482 & n22223 ;
  assign n22225 = n22224 ^ n13614 ^ 1'b0 ;
  assign n22226 = n22222 & n22225 ;
  assign n22228 = ~n5086 & n11680 ;
  assign n22229 = n22228 ^ n8587 ^ 1'b0 ;
  assign n22230 = n1338 & n22229 ;
  assign n22231 = n390 & n22230 ;
  assign n22227 = n171 & n607 ;
  assign n22232 = n22231 ^ n22227 ^ 1'b0 ;
  assign n22234 = ( ~n6665 & n6819 ) | ( ~n6665 & n7972 ) | ( n6819 & n7972 ) ;
  assign n22233 = n15583 ^ n11565 ^ n6809 ;
  assign n22235 = n22234 ^ n22233 ^ n672 ;
  assign n22236 = ( x9 & n16495 ) | ( x9 & n22235 ) | ( n16495 & n22235 ) ;
  assign n22242 = ~n576 & n3556 ;
  assign n22237 = n576 | n5711 ;
  assign n22238 = n5690 | n22237 ;
  assign n22239 = n22238 ^ n12347 ^ 1'b0 ;
  assign n22240 = n22239 ^ n5776 ^ n615 ;
  assign n22241 = n22240 ^ n14482 ^ n486 ;
  assign n22243 = n22242 ^ n22241 ^ n18935 ;
  assign n22244 = n19264 ^ n10419 ^ n7591 ;
  assign n22245 = n1609 & ~n19455 ;
  assign n22246 = ~n11883 & n22245 ;
  assign n22247 = n4217 | n22246 ;
  assign n22248 = n22247 ^ n2031 ^ 1'b0 ;
  assign n22249 = n22248 ^ n16429 ^ 1'b0 ;
  assign n22250 = ~n1918 & n5782 ;
  assign n22251 = n22250 ^ n3089 ^ 1'b0 ;
  assign n22252 = n4354 ^ n1343 ^ n205 ;
  assign n22253 = n3542 & n8920 ;
  assign n22254 = ~n22252 & n22253 ;
  assign n22255 = ( ~n628 & n19812 ) | ( ~n628 & n22254 ) | ( n19812 & n22254 ) ;
  assign n22256 = n1272 | n12344 ;
  assign n22257 = ( ~n7744 & n8592 ) | ( ~n7744 & n22256 ) | ( n8592 & n22256 ) ;
  assign n22258 = n6398 & n9116 ;
  assign n22259 = n19093 ^ n11143 ^ n7048 ;
  assign n22260 = ( n21376 & n22258 ) | ( n21376 & ~n22259 ) | ( n22258 & ~n22259 ) ;
  assign n22261 = ( n1159 & n11206 ) | ( n1159 & ~n17541 ) | ( n11206 & ~n17541 ) ;
  assign n22262 = n10954 ^ n10917 ^ n3904 ;
  assign n22263 = n22262 ^ n16467 ^ 1'b0 ;
  assign n22264 = n7320 & ~n22263 ;
  assign n22265 = n7782 & n22264 ;
  assign n22266 = n5724 ^ n1679 ^ 1'b0 ;
  assign n22267 = ~n22265 & n22266 ;
  assign n22268 = n22267 ^ n4961 ^ 1'b0 ;
  assign n22273 = n4837 & n13477 ;
  assign n22274 = n22273 ^ n911 ^ 1'b0 ;
  assign n22275 = n22274 ^ n17117 ^ 1'b0 ;
  assign n22269 = n9701 ^ n7098 ^ n5110 ;
  assign n22270 = n8058 & n22269 ;
  assign n22271 = ~n15549 & n22270 ;
  assign n22272 = n239 & ~n22271 ;
  assign n22276 = n22275 ^ n22272 ^ 1'b0 ;
  assign n22277 = n6420 & ~n16025 ;
  assign n22278 = n22277 ^ n17177 ^ 1'b0 ;
  assign n22279 = n22278 ^ n19557 ^ n196 ;
  assign n22280 = n22279 ^ n4628 ^ 1'b0 ;
  assign n22283 = n7784 | n10650 ;
  assign n22284 = n8619 & ~n22283 ;
  assign n22285 = n727 | n3614 ;
  assign n22286 = n2383 & n22285 ;
  assign n22287 = n3551 | n22286 ;
  assign n22288 = ~n22284 & n22287 ;
  assign n22281 = n15850 & ~n20494 ;
  assign n22282 = n5590 | n22281 ;
  assign n22289 = n22288 ^ n22282 ^ 1'b0 ;
  assign n22290 = ( n7521 & n8701 ) | ( n7521 & ~n11982 ) | ( n8701 & ~n11982 ) ;
  assign n22291 = n18529 ^ n10161 ^ 1'b0 ;
  assign n22292 = n2833 & n4956 ;
  assign n22293 = n5302 | n9949 ;
  assign n22294 = ( ~n5850 & n8558 ) | ( ~n5850 & n9370 ) | ( n8558 & n9370 ) ;
  assign n22295 = ~n9179 & n16516 ;
  assign n22296 = n22294 & n22295 ;
  assign n22297 = n4489 & ~n5448 ;
  assign n22298 = ~n5167 & n12375 ;
  assign n22299 = n5654 | n18690 ;
  assign n22300 = n22299 ^ n13639 ^ 1'b0 ;
  assign n22301 = n22300 ^ n16873 ^ 1'b0 ;
  assign n22302 = n18542 & ~n18627 ;
  assign n22303 = n22302 ^ n13551 ^ 1'b0 ;
  assign n22304 = ( n2296 & ~n5601 ) | ( n2296 & n9473 ) | ( ~n5601 & n9473 ) ;
  assign n22305 = n22304 ^ n7360 ^ 1'b0 ;
  assign n22306 = n12328 ^ n10316 ^ 1'b0 ;
  assign n22307 = n22305 & n22306 ;
  assign n22308 = n19962 ^ n6350 ^ 1'b0 ;
  assign n22309 = n22308 ^ n20528 ^ n2781 ;
  assign n22310 = ( n933 & n1696 ) | ( n933 & ~n10413 ) | ( n1696 & ~n10413 ) ;
  assign n22311 = n22310 ^ n16245 ^ 1'b0 ;
  assign n22312 = ( n1309 & n3857 ) | ( n1309 & ~n14687 ) | ( n3857 & ~n14687 ) ;
  assign n22313 = n4182 & ~n20579 ;
  assign n22314 = ~n1615 & n20825 ;
  assign n22315 = n3402 & n22314 ;
  assign n22318 = n3483 ^ n470 ^ 1'b0 ;
  assign n22319 = n1077 & ~n22318 ;
  assign n22316 = n7271 | n20352 ;
  assign n22317 = n22316 ^ n15757 ^ 1'b0 ;
  assign n22320 = n22319 ^ n22317 ^ n13212 ;
  assign n22321 = n10157 ^ n6530 ^ 1'b0 ;
  assign n22322 = ~n13124 & n22321 ;
  assign n22323 = n22320 & n22322 ;
  assign n22324 = n21880 ^ n6213 ^ x50 ;
  assign n22325 = n905 & ~n6331 ;
  assign n22326 = n22325 ^ n3176 ^ 1'b0 ;
  assign n22327 = n4907 | n22326 ;
  assign n22328 = n22327 ^ n22006 ^ 1'b0 ;
  assign n22329 = ~n2561 & n3177 ;
  assign n22330 = ~n22328 & n22329 ;
  assign n22331 = n13343 & n21900 ;
  assign n22332 = n22331 ^ n3321 ^ 1'b0 ;
  assign n22333 = n22332 ^ n2404 ^ 1'b0 ;
  assign n22334 = n22330 | n22333 ;
  assign n22335 = n22324 | n22334 ;
  assign n22336 = n22335 ^ n7468 ^ 1'b0 ;
  assign n22337 = n136 & n859 ;
  assign n22338 = ( ~n970 & n1836 ) | ( ~n970 & n22337 ) | ( n1836 & n22337 ) ;
  assign n22339 = n3440 ^ n838 ^ 1'b0 ;
  assign n22340 = n22338 & ~n22339 ;
  assign n22341 = n10672 ^ n2416 ^ n1213 ;
  assign n22342 = n1511 | n22341 ;
  assign n22343 = n19864 | n22342 ;
  assign n22344 = n17112 ^ n13837 ^ 1'b0 ;
  assign n22345 = ~n5569 & n8423 ;
  assign n22346 = ( n2969 & ~n5083 ) | ( n2969 & n22345 ) | ( ~n5083 & n22345 ) ;
  assign n22347 = n2901 ^ n980 ^ 1'b0 ;
  assign n22348 = ( n2569 & n5006 ) | ( n2569 & ~n12958 ) | ( n5006 & ~n12958 ) ;
  assign n22349 = n6972 & n7614 ;
  assign n22350 = ~n759 & n10595 ;
  assign n22351 = ~n7145 & n22350 ;
  assign n22352 = n16845 ^ n2597 ^ 1'b0 ;
  assign n22353 = n1843 & ~n2389 ;
  assign n22354 = ( ~n3527 & n10349 ) | ( ~n3527 & n12788 ) | ( n10349 & n12788 ) ;
  assign n22355 = n2565 | n3548 ;
  assign n22356 = n8468 & ~n22355 ;
  assign n22357 = n18214 ^ n15245 ^ n3625 ;
  assign n22358 = ( n210 & n5954 ) | ( n210 & ~n9869 ) | ( n5954 & ~n9869 ) ;
  assign n22359 = ( n21685 & n22357 ) | ( n21685 & ~n22358 ) | ( n22357 & ~n22358 ) ;
  assign n22360 = n22356 | n22359 ;
  assign n22361 = n22360 ^ n16205 ^ 1'b0 ;
  assign n22362 = ~n22354 & n22361 ;
  assign n22363 = n22353 & n22362 ;
  assign n22364 = n2057 & n20312 ;
  assign n22365 = n13134 & n22364 ;
  assign n22366 = ( n16944 & ~n19215 ) | ( n16944 & n22365 ) | ( ~n19215 & n22365 ) ;
  assign n22367 = n8393 & n17069 ;
  assign n22368 = n22367 ^ n6275 ^ 1'b0 ;
  assign n22369 = ( ~n3217 & n21491 ) | ( ~n3217 & n22368 ) | ( n21491 & n22368 ) ;
  assign n22370 = ( ~n2717 & n20511 ) | ( ~n2717 & n21740 ) | ( n20511 & n21740 ) ;
  assign n22371 = n21059 ^ n1484 ^ 1'b0 ;
  assign n22372 = n8106 ^ n1475 ^ 1'b0 ;
  assign n22373 = n3008 & ~n22372 ;
  assign n22374 = n9249 ^ n4157 ^ n2720 ;
  assign n22375 = n9053 & ~n22374 ;
  assign n22376 = ~n22373 & n22375 ;
  assign n22377 = n9282 | n16225 ;
  assign n22378 = n12657 ^ n10816 ^ 1'b0 ;
  assign n22379 = n9348 ^ n6759 ^ 1'b0 ;
  assign n22380 = ( n6260 & n20667 ) | ( n6260 & n22379 ) | ( n20667 & n22379 ) ;
  assign n22381 = n22380 ^ n12832 ^ n307 ;
  assign n22382 = n9813 ^ n2131 ^ 1'b0 ;
  assign n22383 = ( ~n1316 & n7673 ) | ( ~n1316 & n10976 ) | ( n7673 & n10976 ) ;
  assign n22384 = n22383 ^ n18329 ^ n17440 ;
  assign n22385 = n9916 ^ n3639 ^ 1'b0 ;
  assign n22386 = n2811 ^ x77 ^ 1'b0 ;
  assign n22387 = n3338 ^ n692 ^ 1'b0 ;
  assign n22388 = ~n683 & n22387 ;
  assign n22389 = n22386 & n22388 ;
  assign n22390 = ~n12491 & n22389 ;
  assign n22391 = n3980 ^ n1240 ^ 1'b0 ;
  assign n22392 = ~n7476 & n22391 ;
  assign n22393 = n22392 ^ n1545 ^ 1'b0 ;
  assign n22394 = n307 & ~n7174 ;
  assign n22395 = ~n307 & n22394 ;
  assign n22396 = n22395 ^ n3383 ^ 1'b0 ;
  assign n22397 = n20102 & n22396 ;
  assign n22398 = ~n22396 & n22397 ;
  assign n22399 = n5049 & n10128 ;
  assign n22400 = n11633 & n12245 ;
  assign n22401 = n5986 & n8744 ;
  assign n22402 = n22401 ^ n8262 ^ 1'b0 ;
  assign n22403 = n22402 ^ n18073 ^ n14589 ;
  assign n22404 = n10619 ^ n2205 ^ n1202 ;
  assign n22405 = n16601 ^ n4900 ^ 1'b0 ;
  assign n22406 = n4754 & ~n22405 ;
  assign n22407 = n22406 ^ n17378 ^ n7972 ;
  assign n22408 = n22404 & ~n22407 ;
  assign n22409 = n6035 ^ n3862 ^ 1'b0 ;
  assign n22410 = n12815 & ~n22409 ;
  assign n22411 = ~n4762 & n22410 ;
  assign n22412 = n161 & n17886 ;
  assign n22413 = ~n1658 & n22412 ;
  assign n22414 = x32 & n5390 ;
  assign n22415 = ~n5774 & n22414 ;
  assign n22416 = ~n16173 & n22415 ;
  assign n22417 = n4304 & ~n5434 ;
  assign n22418 = n22417 ^ n18876 ^ n5350 ;
  assign n22421 = ~n5850 & n21385 ;
  assign n22422 = n22421 ^ n5407 ^ 1'b0 ;
  assign n22420 = n8713 ^ n3815 ^ 1'b0 ;
  assign n22423 = n22422 ^ n22420 ^ n12503 ;
  assign n22419 = n11059 & n14627 ;
  assign n22424 = n22423 ^ n22419 ^ n20917 ;
  assign n22425 = n22424 ^ n17629 ^ n13201 ;
  assign n22426 = n21175 ^ n4454 ^ n1599 ;
  assign n22427 = n22426 ^ n5056 ^ n1915 ;
  assign n22428 = n22427 ^ n13927 ^ n10640 ;
  assign n22429 = n22428 ^ n20126 ^ n3390 ;
  assign n22430 = n22429 ^ n10120 ^ n3688 ;
  assign n22431 = n9972 ^ n6446 ^ n6399 ;
  assign n22432 = ~n7338 & n17940 ;
  assign n22433 = n6936 & n22432 ;
  assign n22434 = ( n1076 & n2041 ) | ( n1076 & n22433 ) | ( n2041 & n22433 ) ;
  assign n22435 = n22434 ^ n13949 ^ 1'b0 ;
  assign n22436 = n22210 & n22435 ;
  assign n22437 = n18483 ^ n13939 ^ 1'b0 ;
  assign n22438 = n8341 & n17713 ;
  assign n22439 = n22438 ^ n5314 ^ 1'b0 ;
  assign n22440 = n22439 ^ n16805 ^ 1'b0 ;
  assign n22441 = n16188 ^ n6805 ^ n6180 ;
  assign n22442 = ~n9613 & n14591 ;
  assign n22443 = n20536 ^ n12755 ^ 1'b0 ;
  assign n22444 = n11930 & n22443 ;
  assign n22445 = ( ~n9053 & n22442 ) | ( ~n9053 & n22444 ) | ( n22442 & n22444 ) ;
  assign n22446 = n4571 & ~n5787 ;
  assign n22447 = n22446 ^ n6416 ^ 1'b0 ;
  assign n22448 = ( n6489 & n16553 ) | ( n6489 & n22447 ) | ( n16553 & n22447 ) ;
  assign n22449 = n6841 & n13903 ;
  assign n22450 = ~n754 & n4933 ;
  assign n22451 = n22450 ^ n3270 ^ 1'b0 ;
  assign n22452 = n22451 ^ n19781 ^ 1'b0 ;
  assign n22453 = n22449 & ~n22452 ;
  assign n22454 = n9621 | n13966 ;
  assign n22455 = n2625 ^ n1877 ^ 1'b0 ;
  assign n22456 = n6987 & n22455 ;
  assign n22457 = n379 & ~n927 ;
  assign n22458 = n22457 ^ n14474 ^ n3911 ;
  assign n22459 = n22456 & ~n22458 ;
  assign n22461 = n1100 & n2905 ;
  assign n22462 = n22461 ^ n2768 ^ n1943 ;
  assign n22460 = n10549 & n15317 ;
  assign n22463 = n22462 ^ n22460 ^ n3232 ;
  assign n22464 = ( n1952 & n18738 ) | ( n1952 & ~n22463 ) | ( n18738 & ~n22463 ) ;
  assign n22465 = n11420 ^ n7560 ^ 1'b0 ;
  assign n22466 = ( ~n15556 & n15824 ) | ( ~n15556 & n22465 ) | ( n15824 & n22465 ) ;
  assign n22467 = n22466 ^ n18619 ^ n476 ;
  assign n22471 = n21494 ^ n5603 ^ 1'b0 ;
  assign n22472 = n17277 | n22471 ;
  assign n22469 = ( n13219 & n15306 ) | ( n13219 & ~n17906 ) | ( n15306 & ~n17906 ) ;
  assign n22470 = ( ~n15536 & n22191 ) | ( ~n15536 & n22469 ) | ( n22191 & n22469 ) ;
  assign n22468 = ( n3206 & ~n15023 ) | ( n3206 & n18066 ) | ( ~n15023 & n18066 ) ;
  assign n22473 = n22472 ^ n22470 ^ n22468 ;
  assign n22474 = n6431 ^ n4010 ^ 1'b0 ;
  assign n22475 = n22474 ^ n14721 ^ n2366 ;
  assign n22479 = ~n364 & n14182 ;
  assign n22476 = ~n4492 & n12758 ;
  assign n22477 = n22476 ^ n21590 ^ 1'b0 ;
  assign n22478 = n448 & ~n22477 ;
  assign n22480 = n22479 ^ n22478 ^ 1'b0 ;
  assign n22481 = n16915 & n18921 ;
  assign n22482 = n22481 ^ n12494 ^ 1'b0 ;
  assign n22483 = n22482 ^ n10238 ^ n3986 ;
  assign n22484 = n22483 ^ n4520 ^ 1'b0 ;
  assign n22485 = n19884 ^ n18747 ^ n8018 ;
  assign n22486 = ( n2698 & ~n15625 ) | ( n2698 & n22485 ) | ( ~n15625 & n22485 ) ;
  assign n22487 = n5857 ^ n2432 ^ 1'b0 ;
  assign n22488 = ( n1319 & n16668 ) | ( n1319 & n22487 ) | ( n16668 & n22487 ) ;
  assign n22489 = n22488 ^ n19480 ^ n2751 ;
  assign n22490 = n8567 ^ n8445 ^ 1'b0 ;
  assign n22491 = n11919 & n22490 ;
  assign n22492 = ( n1117 & n2537 ) | ( n1117 & n8188 ) | ( n2537 & n8188 ) ;
  assign n22493 = ~n4529 & n22492 ;
  assign n22494 = n12208 & n22008 ;
  assign n22495 = n4323 ^ n1879 ^ x53 ;
  assign n22496 = x59 & n22495 ;
  assign n22499 = ( n4712 & n11100 ) | ( n4712 & n12874 ) | ( n11100 & n12874 ) ;
  assign n22497 = n4292 & ~n4385 ;
  assign n22498 = n22497 ^ n3921 ^ 1'b0 ;
  assign n22500 = n22499 ^ n22498 ^ n1065 ;
  assign n22501 = ( n7528 & n10440 ) | ( n7528 & ~n15892 ) | ( n10440 & ~n15892 ) ;
  assign n22502 = n1754 & n3631 ;
  assign n22503 = ~n10794 & n22502 ;
  assign n22504 = ~n2466 & n5768 ;
  assign n22505 = n1576 & ~n15334 ;
  assign n22506 = n22505 ^ n17425 ^ 1'b0 ;
  assign n22507 = n11937 ^ n8711 ^ n6672 ;
  assign n22508 = n15485 ^ n178 ^ 1'b0 ;
  assign n22509 = n22507 & n22508 ;
  assign n22511 = n4274 ^ n2868 ^ n1262 ;
  assign n22510 = n16121 ^ n3548 ^ 1'b0 ;
  assign n22512 = n22511 ^ n22510 ^ n4501 ;
  assign n22513 = ( n756 & n6284 ) | ( n756 & n22512 ) | ( n6284 & n22512 ) ;
  assign n22514 = ~n3134 & n13490 ;
  assign n22515 = n22514 ^ n10187 ^ 1'b0 ;
  assign n22516 = n16035 ^ n1576 ^ 1'b0 ;
  assign n22517 = ~n5142 & n22516 ;
  assign n22518 = n22517 ^ n3288 ^ 1'b0 ;
  assign n22519 = n595 & ~n22518 ;
  assign n22520 = n10433 & ~n22519 ;
  assign n22521 = n6477 & ~n7979 ;
  assign n22522 = ( n3523 & n6823 ) | ( n3523 & n21683 ) | ( n6823 & n21683 ) ;
  assign n22523 = n14660 & ~n22522 ;
  assign n22524 = n22523 ^ n2081 ^ 1'b0 ;
  assign n22525 = n22524 ^ n14068 ^ 1'b0 ;
  assign n22526 = n9343 ^ n9146 ^ 1'b0 ;
  assign n22527 = n22526 ^ n11088 ^ n7346 ;
  assign n22533 = n7165 | n19794 ;
  assign n22532 = ( ~n1992 & n12938 ) | ( ~n1992 & n14237 ) | ( n12938 & n14237 ) ;
  assign n22529 = n2279 ^ n2199 ^ n516 ;
  assign n22530 = n22529 ^ n15563 ^ 1'b0 ;
  assign n22528 = ~n3517 & n3777 ;
  assign n22531 = n22530 ^ n22528 ^ 1'b0 ;
  assign n22534 = n22533 ^ n22532 ^ n22531 ;
  assign n22535 = ( n11782 & ~n16360 ) | ( n11782 & n22163 ) | ( ~n16360 & n22163 ) ;
  assign n22536 = n4574 | n15886 ;
  assign n22537 = n22536 ^ n8028 ^ 1'b0 ;
  assign n22538 = n7914 & n22537 ;
  assign n22539 = ~n2014 & n22538 ;
  assign n22540 = n22539 ^ n2489 ^ 1'b0 ;
  assign n22541 = n2835 & n9746 ;
  assign n22542 = ( n5544 & ~n7545 ) | ( n5544 & n20045 ) | ( ~n7545 & n20045 ) ;
  assign n22543 = n386 & ~n6821 ;
  assign n22544 = n22542 & n22543 ;
  assign n22545 = n9054 ^ n2897 ^ 1'b0 ;
  assign n22546 = n16282 ^ n8752 ^ 1'b0 ;
  assign n22547 = ( n1485 & n1562 ) | ( n1485 & n6678 ) | ( n1562 & n6678 ) ;
  assign n22548 = n17142 ^ n474 ^ 1'b0 ;
  assign n22549 = n15233 | n22548 ;
  assign n22550 = n771 | n16353 ;
  assign n22551 = n7144 ^ n131 ^ 1'b0 ;
  assign n22552 = n188 & n7748 ;
  assign n22553 = n22552 ^ n18997 ^ 1'b0 ;
  assign n22554 = n6145 | n22553 ;
  assign n22555 = ( n3106 & ~n12608 ) | ( n3106 & n16619 ) | ( ~n12608 & n16619 ) ;
  assign n22556 = n8636 ^ n826 ^ 1'b0 ;
  assign n22557 = n13354 ^ n7237 ^ 1'b0 ;
  assign n22558 = n6590 & n22557 ;
  assign n22565 = n18741 ^ n7985 ^ 1'b0 ;
  assign n22559 = n8018 ^ n7560 ^ 1'b0 ;
  assign n22560 = ~n4172 & n22559 ;
  assign n22561 = n22560 ^ n20586 ^ n13848 ;
  assign n22562 = ~n11829 & n22145 ;
  assign n22563 = ~n4538 & n22562 ;
  assign n22564 = ~n22561 & n22563 ;
  assign n22566 = n22565 ^ n22564 ^ n15736 ;
  assign n22567 = ~n1417 & n7489 ;
  assign n22568 = ~n17138 & n22567 ;
  assign n22569 = n19554 & n21646 ;
  assign n22570 = n17896 & n22569 ;
  assign n22571 = ( ~n834 & n3510 ) | ( ~n834 & n6338 ) | ( n3510 & n6338 ) ;
  assign n22572 = ~n19827 & n22571 ;
  assign n22573 = n22572 ^ n537 ^ 1'b0 ;
  assign n22574 = ( n8052 & ~n10136 ) | ( n8052 & n16362 ) | ( ~n10136 & n16362 ) ;
  assign n22575 = n4429 & ~n22574 ;
  assign n22576 = n12891 & ~n20114 ;
  assign n22577 = n4025 & n22576 ;
  assign n22578 = ( n6201 & ~n22575 ) | ( n6201 & n22577 ) | ( ~n22575 & n22577 ) ;
  assign n22579 = n5604 ^ n2093 ^ 1'b0 ;
  assign n22580 = n22579 ^ n1966 ^ 1'b0 ;
  assign n22581 = ~n141 & n7542 ;
  assign n22582 = n3062 ^ n2263 ^ 1'b0 ;
  assign n22583 = n8985 | n17040 ;
  assign n22584 = n22582 | n22583 ;
  assign n22585 = n5525 ^ n1745 ^ 1'b0 ;
  assign n22586 = ( n3788 & n10668 ) | ( n3788 & ~n22585 ) | ( n10668 & ~n22585 ) ;
  assign n22587 = n22586 ^ n12721 ^ n4154 ;
  assign n22588 = x113 & n22587 ;
  assign n22589 = ( n10698 & n13955 ) | ( n10698 & ~n18678 ) | ( n13955 & ~n18678 ) ;
  assign n22590 = n10660 ^ n7441 ^ 1'b0 ;
  assign n22591 = n22590 ^ n19560 ^ n1282 ;
  assign n22592 = n22591 ^ n15785 ^ n11226 ;
  assign n22593 = ( n4494 & n9324 ) | ( n4494 & n15499 ) | ( n9324 & n15499 ) ;
  assign n22594 = ( ~n11628 & n19425 ) | ( ~n11628 & n19502 ) | ( n19425 & n19502 ) ;
  assign n22595 = n19862 | n20106 ;
  assign n22596 = ~n7268 & n9651 ;
  assign n22597 = n22596 ^ n9442 ^ 1'b0 ;
  assign n22598 = n16760 & n22597 ;
  assign n22601 = n11694 ^ n8242 ^ 1'b0 ;
  assign n22602 = ~n21348 & n22601 ;
  assign n22599 = n8796 & ~n13818 ;
  assign n22600 = ~n2173 & n22599 ;
  assign n22603 = n22602 ^ n22600 ^ n13138 ;
  assign n22604 = n22603 ^ n2896 ^ 1'b0 ;
  assign n22605 = n12009 & ~n22604 ;
  assign n22606 = n14645 ^ n11210 ^ n2679 ;
  assign n22607 = n9914 & n19796 ;
  assign n22608 = ( n5739 & ~n12431 ) | ( n5739 & n19538 ) | ( ~n12431 & n19538 ) ;
  assign n22609 = n14736 ^ n8508 ^ n6490 ;
  assign n22610 = ( n8436 & n20954 ) | ( n8436 & n22117 ) | ( n20954 & n22117 ) ;
  assign n22611 = ~n9298 & n14460 ;
  assign n22612 = n7175 ^ n5276 ^ 1'b0 ;
  assign n22613 = n214 & n22612 ;
  assign n22614 = n4999 & n7079 ;
  assign n22615 = ~n19117 & n22614 ;
  assign n22616 = n14326 ^ n4595 ^ 1'b0 ;
  assign n22617 = n22615 | n22616 ;
  assign n22618 = ( ~n17815 & n22613 ) | ( ~n17815 & n22617 ) | ( n22613 & n22617 ) ;
  assign n22619 = n22618 ^ n9574 ^ 1'b0 ;
  assign n22620 = n22611 & n22619 ;
  assign n22621 = n8349 ^ n7776 ^ 1'b0 ;
  assign n22622 = n14037 ^ n6008 ^ 1'b0 ;
  assign n22623 = ( n3476 & n13758 ) | ( n3476 & n19588 ) | ( n13758 & n19588 ) ;
  assign n22624 = n22623 ^ n6140 ^ 1'b0 ;
  assign n22625 = ( ~n3376 & n4878 ) | ( ~n3376 & n22071 ) | ( n4878 & n22071 ) ;
  assign n22626 = n22625 ^ n12858 ^ 1'b0 ;
  assign n22627 = n10449 | n15206 ;
  assign n22628 = n22627 ^ n10647 ^ 1'b0 ;
  assign n22629 = n8894 ^ n3776 ^ 1'b0 ;
  assign n22630 = n14807 ^ n3819 ^ 1'b0 ;
  assign n22631 = n16558 ^ n15667 ^ n10765 ;
  assign n22632 = n22631 ^ n17420 ^ n8097 ;
  assign n22633 = n7149 ^ n1568 ^ n398 ;
  assign n22634 = ( ~n6637 & n7335 ) | ( ~n6637 & n11815 ) | ( n7335 & n11815 ) ;
  assign n22635 = n22634 ^ n4073 ^ 1'b0 ;
  assign n22636 = n7513 & n14335 ;
  assign n22637 = n18769 & n22636 ;
  assign n22638 = ~n6455 & n10231 ;
  assign n22639 = n22638 ^ n2745 ^ 1'b0 ;
  assign n22640 = n924 & n7776 ;
  assign n22641 = n15752 ^ n12266 ^ n6480 ;
  assign n22642 = n16919 ^ n8660 ^ 1'b0 ;
  assign n22643 = n22642 ^ n11184 ^ n2981 ;
  assign n22646 = n14875 ^ n14557 ^ n13337 ;
  assign n22644 = n4287 & ~n19120 ;
  assign n22645 = n22644 ^ n9649 ^ 1'b0 ;
  assign n22647 = n22646 ^ n22645 ^ 1'b0 ;
  assign n22648 = n4718 | n9634 ;
  assign n22649 = n4836 & ~n22648 ;
  assign n22650 = n12475 ^ n10380 ^ n4814 ;
  assign n22651 = ( n294 & n9537 ) | ( n294 & ~n22650 ) | ( n9537 & ~n22650 ) ;
  assign n22652 = n22651 ^ n14380 ^ 1'b0 ;
  assign n22653 = ~n19131 & n22652 ;
  assign n22654 = ~n2804 & n2831 ;
  assign n22655 = ~n3337 & n5498 ;
  assign n22656 = ~n22654 & n22655 ;
  assign n22657 = ~n2129 & n22656 ;
  assign n22658 = n3042 & n9672 ;
  assign n22659 = n4418 & ~n6710 ;
  assign n22660 = n9622 ^ n5786 ^ n1789 ;
  assign n22661 = n10370 ^ n4851 ^ n3572 ;
  assign n22662 = n22661 ^ n20897 ^ n9828 ;
  assign n22665 = n6120 ^ n4691 ^ n1253 ;
  assign n22666 = n9265 & ~n22665 ;
  assign n22663 = ( n11582 & n15928 ) | ( n11582 & n21691 ) | ( n15928 & n21691 ) ;
  assign n22664 = n22663 ^ n3321 ^ 1'b0 ;
  assign n22667 = n22666 ^ n22664 ^ n5906 ;
  assign n22668 = n4563 & n12125 ;
  assign n22669 = ~n12185 & n22668 ;
  assign n22670 = n356 & ~n6890 ;
  assign n22671 = n22670 ^ n11791 ^ 1'b0 ;
  assign n22672 = n15595 & n22671 ;
  assign n22673 = n2371 & n22672 ;
  assign n22674 = n17008 ^ n11837 ^ n7913 ;
  assign n22675 = n4915 & ~n21392 ;
  assign n22676 = n8148 ^ n7958 ^ 1'b0 ;
  assign n22677 = n20253 ^ n19385 ^ n9664 ;
  assign n22678 = ~n3761 & n4578 ;
  assign n22679 = n14500 & n22678 ;
  assign n22680 = ~n22677 & n22679 ;
  assign n22681 = ( n4029 & ~n18963 ) | ( n4029 & n22680 ) | ( ~n18963 & n22680 ) ;
  assign n22682 = ( n1104 & n3422 ) | ( n1104 & ~n22519 ) | ( n3422 & ~n22519 ) ;
  assign n22683 = n8012 | n17275 ;
  assign n22684 = n22683 ^ n3858 ^ 1'b0 ;
  assign n22685 = n21030 & ~n22684 ;
  assign n22686 = n12144 ^ n1011 ^ 1'b0 ;
  assign n22687 = n20701 ^ n917 ^ 1'b0 ;
  assign n22688 = n3360 | n22687 ;
  assign n22689 = n10590 ^ n8301 ^ x96 ;
  assign n22690 = ( ~n6055 & n22688 ) | ( ~n6055 & n22689 ) | ( n22688 & n22689 ) ;
  assign n22691 = ~n10521 & n22690 ;
  assign n22692 = n22686 & n22691 ;
  assign n22693 = x26 & ~n12449 ;
  assign n22694 = n18073 & n22693 ;
  assign n22695 = n22694 ^ n16586 ^ 1'b0 ;
  assign n22696 = n1816 & ~n22695 ;
  assign n22697 = n15850 ^ n5213 ^ n5145 ;
  assign n22698 = n13700 ^ n12460 ^ 1'b0 ;
  assign n22699 = n22697 & n22698 ;
  assign n22700 = n6755 ^ n3588 ^ 1'b0 ;
  assign n22701 = n8215 & ~n22700 ;
  assign n22702 = ( ~n2663 & n5077 ) | ( ~n2663 & n22701 ) | ( n5077 & n22701 ) ;
  assign n22703 = n22702 ^ n16741 ^ n14745 ;
  assign n22704 = n22703 ^ n7633 ^ 1'b0 ;
  assign n22705 = n14512 & ~n22704 ;
  assign n22706 = n8422 ^ n5684 ^ 1'b0 ;
  assign n22707 = ( n4740 & n17060 ) | ( n4740 & ~n22706 ) | ( n17060 & ~n22706 ) ;
  assign n22708 = n305 & ~n3104 ;
  assign n22709 = n12573 & n22708 ;
  assign n22710 = n1411 & ~n22709 ;
  assign n22711 = n10792 ^ n7966 ^ 1'b0 ;
  assign n22712 = n22710 & n22711 ;
  assign n22713 = n16683 ^ n12563 ^ 1'b0 ;
  assign n22714 = ( n14486 & ~n17580 ) | ( n14486 & n22713 ) | ( ~n17580 & n22713 ) ;
  assign n22715 = n16791 ^ n5077 ^ 1'b0 ;
  assign n22716 = ( n9713 & n10564 ) | ( n9713 & n10601 ) | ( n10564 & n10601 ) ;
  assign n22717 = ( n10645 & n22715 ) | ( n10645 & ~n22716 ) | ( n22715 & ~n22716 ) ;
  assign n22718 = n6847 ^ n3246 ^ 1'b0 ;
  assign n22721 = n3542 & ~n8043 ;
  assign n22722 = n13764 & n22721 ;
  assign n22719 = n5468 ^ n2253 ^ 1'b0 ;
  assign n22720 = n17242 & n22719 ;
  assign n22723 = n22722 ^ n22720 ^ 1'b0 ;
  assign n22724 = n5095 & ~n9216 ;
  assign n22725 = n13255 ^ n7724 ^ n5297 ;
  assign n22726 = ( n676 & n986 ) | ( n676 & n22725 ) | ( n986 & n22725 ) ;
  assign n22727 = n22724 & n22726 ;
  assign n22728 = n16680 | n17139 ;
  assign n22729 = n22728 ^ n8471 ^ 1'b0 ;
  assign n22730 = ( n2062 & n12258 ) | ( n2062 & n22729 ) | ( n12258 & n22729 ) ;
  assign n22731 = n7606 ^ n4955 ^ 1'b0 ;
  assign n22732 = ~n829 & n9998 ;
  assign n22733 = n3462 & n22732 ;
  assign n22734 = n22733 ^ n21382 ^ n13242 ;
  assign n22735 = n22666 ^ n500 ^ 1'b0 ;
  assign n22736 = n12685 & n22735 ;
  assign n22737 = n21332 | n22736 ;
  assign n22738 = ( n2978 & n8177 ) | ( n2978 & n21114 ) | ( n8177 & n21114 ) ;
  assign n22739 = n16971 & ~n22738 ;
  assign n22740 = ~n7239 & n22739 ;
  assign n22741 = n22511 ^ n10519 ^ n4465 ;
  assign n22742 = n16962 ^ n4263 ^ 1'b0 ;
  assign n22743 = n6557 ^ n3728 ^ 1'b0 ;
  assign n22744 = n15764 ^ n2100 ^ 1'b0 ;
  assign n22745 = n10571 & ~n10820 ;
  assign n22746 = n4177 & n18821 ;
  assign n22747 = ~n22745 & n22746 ;
  assign n22748 = ~n10981 & n22747 ;
  assign n22749 = n5309 ^ n1843 ^ 1'b0 ;
  assign n22750 = n8387 & n22749 ;
  assign n22751 = ( ~n22744 & n22748 ) | ( ~n22744 & n22750 ) | ( n22748 & n22750 ) ;
  assign n22752 = n5463 & n17296 ;
  assign n22756 = ~n974 & n11850 ;
  assign n22753 = n5822 ^ n1274 ^ 1'b0 ;
  assign n22754 = ~n16128 & n22753 ;
  assign n22755 = ~n8019 & n22754 ;
  assign n22757 = n22756 ^ n22755 ^ 1'b0 ;
  assign n22758 = n18235 ^ n9777 ^ 1'b0 ;
  assign n22759 = ~n7099 & n22758 ;
  assign n22760 = n8117 & n22759 ;
  assign n22761 = n22760 ^ n6247 ^ 1'b0 ;
  assign n22762 = n7883 ^ n1686 ^ 1'b0 ;
  assign n22763 = n3144 | n22762 ;
  assign n22764 = n22763 ^ n4243 ^ 1'b0 ;
  assign n22765 = n7328 & ~n11432 ;
  assign n22766 = ~n22764 & n22765 ;
  assign n22767 = ( ~n8365 & n18262 ) | ( ~n8365 & n22766 ) | ( n18262 & n22766 ) ;
  assign n22768 = ( n2092 & ~n10109 ) | ( n2092 & n11712 ) | ( ~n10109 & n11712 ) ;
  assign n22769 = n20585 ^ n6721 ^ 1'b0 ;
  assign n22770 = n22769 ^ n3580 ^ 1'b0 ;
  assign n22771 = ~n12329 & n20857 ;
  assign n22772 = ~n18526 & n22771 ;
  assign n22773 = ~n14527 & n22772 ;
  assign n22774 = n16932 & ~n22773 ;
  assign n22775 = n6604 ^ n2965 ^ n895 ;
  assign n22776 = n22774 | n22775 ;
  assign n22777 = n10472 ^ n2267 ^ 1'b0 ;
  assign n22778 = n8403 & n15053 ;
  assign n22779 = n4497 & n22778 ;
  assign n22780 = n1426 & ~n22779 ;
  assign n22781 = ~n11889 & n22780 ;
  assign n22782 = n10132 & ~n22781 ;
  assign n22783 = n22782 ^ n2671 ^ 1'b0 ;
  assign n22784 = n834 & n5956 ;
  assign n22785 = ~n17703 & n22784 ;
  assign n22786 = n8149 & ~n22785 ;
  assign n22787 = n8942 ^ n5529 ^ 1'b0 ;
  assign n22788 = ~n8512 & n22787 ;
  assign n22789 = ( n6405 & n10934 ) | ( n6405 & n22788 ) | ( n10934 & n22788 ) ;
  assign n22790 = ( ~n8738 & n11266 ) | ( ~n8738 & n22789 ) | ( n11266 & n22789 ) ;
  assign n22791 = n7724 ^ n6803 ^ n6564 ;
  assign n22792 = n18387 ^ n16114 ^ 1'b0 ;
  assign n22793 = n4725 ^ n2627 ^ 1'b0 ;
  assign n22794 = n9971 | n22793 ;
  assign n22795 = n14819 ^ n12816 ^ 1'b0 ;
  assign n22796 = n1196 & ~n22795 ;
  assign n22797 = n22796 ^ n19057 ^ 1'b0 ;
  assign n22798 = n22794 | n22797 ;
  assign n22799 = n12813 ^ n3265 ^ 1'b0 ;
  assign n22800 = n12539 | n22799 ;
  assign n22801 = n14917 & ~n22800 ;
  assign n22802 = ~n1381 & n1870 ;
  assign n22803 = n22802 ^ n20340 ^ n1887 ;
  assign n22804 = n3797 ^ n3416 ^ 1'b0 ;
  assign n22805 = n9408 | n12710 ;
  assign n22806 = n2516 | n22805 ;
  assign n22807 = ( n5512 & n6012 ) | ( n5512 & n6862 ) | ( n6012 & n6862 ) ;
  assign n22808 = ( n22804 & n22806 ) | ( n22804 & ~n22807 ) | ( n22806 & ~n22807 ) ;
  assign n22809 = ~n12988 & n19458 ;
  assign n22810 = n2703 & ~n14228 ;
  assign n22811 = n22810 ^ n12168 ^ 1'b0 ;
  assign n22812 = n19158 ^ n160 ^ 1'b0 ;
  assign n22813 = n22811 & n22812 ;
  assign n22814 = n2350 & n18605 ;
  assign n22815 = n22814 ^ n4106 ^ 1'b0 ;
  assign n22816 = n8972 ^ n6083 ^ 1'b0 ;
  assign n22817 = ( n8578 & n17348 ) | ( n8578 & ~n17477 ) | ( n17348 & ~n17477 ) ;
  assign n22818 = n2608 ^ n768 ^ 1'b0 ;
  assign n22819 = n2168 & n10132 ;
  assign n22820 = ~n9962 & n22819 ;
  assign n22821 = n17131 | n22820 ;
  assign n22822 = n6020 & ~n22821 ;
  assign n22823 = n21196 ^ n6344 ^ n3448 ;
  assign n22824 = n22823 ^ n10127 ^ 1'b0 ;
  assign n22825 = n9989 ^ n6375 ^ 1'b0 ;
  assign n22826 = n22825 ^ n8205 ^ 1'b0 ;
  assign n22827 = n6354 & ~n22826 ;
  assign n22828 = ( n357 & ~n2344 ) | ( n357 & n3479 ) | ( ~n2344 & n3479 ) ;
  assign n22829 = n18550 ^ n649 ^ n314 ;
  assign n22830 = n19060 ^ n15982 ^ 1'b0 ;
  assign n22831 = n8049 ^ n7384 ^ 1'b0 ;
  assign n22832 = ( n16672 & n18267 ) | ( n16672 & ~n22831 ) | ( n18267 & ~n22831 ) ;
  assign n22833 = n4668 & ~n22832 ;
  assign n22834 = n6920 ^ n1013 ^ 1'b0 ;
  assign n22835 = ~n20746 & n22834 ;
  assign n22836 = n1900 & n13586 ;
  assign n22837 = n21024 & n22836 ;
  assign n22838 = n18757 ^ n17388 ^ n5897 ;
  assign n22839 = n22838 ^ n17861 ^ 1'b0 ;
  assign n22841 = n2286 & ~n6594 ;
  assign n22842 = n8482 & n22841 ;
  assign n22840 = n20697 | n20704 ;
  assign n22843 = n22842 ^ n22840 ^ n7313 ;
  assign n22845 = ~n743 & n12336 ;
  assign n22846 = n22845 ^ n1627 ^ 1'b0 ;
  assign n22844 = n10681 | n15564 ;
  assign n22847 = n22846 ^ n22844 ^ n14185 ;
  assign n22848 = ( n5760 & ~n6122 ) | ( n5760 & n14664 ) | ( ~n6122 & n14664 ) ;
  assign n22849 = ( n8414 & ~n21053 ) | ( n8414 & n22848 ) | ( ~n21053 & n22848 ) ;
  assign n22850 = n7966 ^ n4445 ^ 1'b0 ;
  assign n22851 = n22850 ^ n6580 ^ 1'b0 ;
  assign n22852 = ( n5728 & ~n16139 ) | ( n5728 & n22851 ) | ( ~n16139 & n22851 ) ;
  assign n22853 = n12593 ^ n1517 ^ 1'b0 ;
  assign n22854 = n15675 ^ n2329 ^ n2248 ;
  assign n22855 = n2239 & n22854 ;
  assign n22856 = ~n22853 & n22855 ;
  assign n22857 = n9883 ^ n1217 ^ 1'b0 ;
  assign n22858 = n16773 ^ n13685 ^ 1'b0 ;
  assign n22859 = n4265 & ~n22858 ;
  assign n22860 = ~n506 & n22859 ;
  assign n22861 = n3727 & n22860 ;
  assign n22862 = n2958 ^ n1056 ^ 1'b0 ;
  assign n22863 = n3063 | n22862 ;
  assign n22864 = n15937 | n22863 ;
  assign n22865 = n9547 ^ x40 ^ 1'b0 ;
  assign n22866 = n6155 | n22865 ;
  assign n22867 = n22864 | n22866 ;
  assign n22868 = ~n9723 & n22867 ;
  assign n22869 = n22868 ^ n1586 ^ 1'b0 ;
  assign n22870 = n14432 ^ n11712 ^ n8941 ;
  assign n22871 = ( ~n5397 & n12503 ) | ( ~n5397 & n22870 ) | ( n12503 & n22870 ) ;
  assign n22872 = ~n239 & n20491 ;
  assign n22873 = n11061 ^ n5020 ^ 1'b0 ;
  assign n22874 = ~n22872 & n22873 ;
  assign n22875 = ( ~n11632 & n16091 ) | ( ~n11632 & n20759 ) | ( n16091 & n20759 ) ;
  assign n22876 = n5098 & n8005 ;
  assign n22877 = n19625 & n22876 ;
  assign n22878 = n2044 & ~n22877 ;
  assign n22879 = n22878 ^ n9423 ^ 1'b0 ;
  assign n22880 = n22879 ^ n8076 ^ 1'b0 ;
  assign n22881 = n19194 ^ n17867 ^ 1'b0 ;
  assign n22882 = ~n11981 & n22881 ;
  assign n22883 = n5263 ^ n4726 ^ 1'b0 ;
  assign n22884 = n22663 ^ n20147 ^ 1'b0 ;
  assign n22885 = n1244 & ~n15176 ;
  assign n22886 = n22885 ^ n10474 ^ 1'b0 ;
  assign n22887 = n4837 ^ x30 ^ 1'b0 ;
  assign n22888 = n22886 & n22887 ;
  assign n22889 = n22888 ^ n17471 ^ n426 ;
  assign n22890 = n8028 ^ n6182 ^ 1'b0 ;
  assign n22891 = x16 & ~n22890 ;
  assign n22892 = ( n1277 & n16919 ) | ( n1277 & n22891 ) | ( n16919 & n22891 ) ;
  assign n22894 = ~n10092 & n21935 ;
  assign n22895 = ~n9369 & n22894 ;
  assign n22893 = n1327 & n17388 ;
  assign n22896 = n22895 ^ n22893 ^ 1'b0 ;
  assign n22897 = n16301 & n19143 ;
  assign n22898 = n4415 & ~n13443 ;
  assign n22899 = ~n16046 & n22898 ;
  assign n22900 = ~n9520 & n22899 ;
  assign n22902 = ~n256 & n525 ;
  assign n22903 = n22902 ^ n228 ^ 1'b0 ;
  assign n22901 = n9242 ^ n4416 ^ 1'b0 ;
  assign n22904 = n22903 ^ n22901 ^ n21040 ;
  assign n22905 = n9065 ^ n4464 ^ 1'b0 ;
  assign n22906 = ( n1314 & n7838 ) | ( n1314 & ~n20847 ) | ( n7838 & ~n20847 ) ;
  assign n22907 = n6604 | n9263 ;
  assign n22908 = ( ~n676 & n2097 ) | ( ~n676 & n9106 ) | ( n2097 & n9106 ) ;
  assign n22909 = n22908 ^ n14190 ^ n9669 ;
  assign n22910 = n22293 ^ n2798 ^ 1'b0 ;
  assign n22911 = n10552 & ~n10558 ;
  assign n22912 = n22911 ^ n14292 ^ 1'b0 ;
  assign n22913 = n16668 ^ n7103 ^ 1'b0 ;
  assign n22914 = ~x3 & n862 ;
  assign n22915 = ( n15610 & ~n16718 ) | ( n15610 & n22914 ) | ( ~n16718 & n22914 ) ;
  assign n22916 = n17842 ^ n7639 ^ 1'b0 ;
  assign n22917 = n17851 ^ n6672 ^ n5215 ;
  assign n22918 = n22917 ^ n6184 ^ n5567 ;
  assign n22919 = n6655 & ~n8461 ;
  assign n22920 = n22919 ^ n19408 ^ n8641 ;
  assign n22921 = n15879 ^ n4841 ^ 1'b0 ;
  assign n22922 = n22921 ^ n15431 ^ n1690 ;
  assign n22923 = ( n6248 & n14745 ) | ( n6248 & ~n22922 ) | ( n14745 & ~n22922 ) ;
  assign n22924 = n4727 ^ n3707 ^ 1'b0 ;
  assign n22925 = ~n5840 & n22924 ;
  assign n22926 = n3373 & n22925 ;
  assign n22927 = n22926 ^ n11493 ^ 1'b0 ;
  assign n22928 = n8606 & ~n22927 ;
  assign n22929 = n22928 ^ n796 ^ 1'b0 ;
  assign n22930 = ( n5149 & n9223 ) | ( n5149 & ~n22383 ) | ( n9223 & ~n22383 ) ;
  assign n22931 = n4155 & ~n22930 ;
  assign n22932 = n22931 ^ n8934 ^ 1'b0 ;
  assign n22933 = n1089 & n4448 ;
  assign n22934 = n22933 ^ n13993 ^ 1'b0 ;
  assign n22935 = ~n3757 & n14512 ;
  assign n22936 = n16007 & n22935 ;
  assign n22937 = ~n2713 & n14053 ;
  assign n22938 = n11335 ^ n7183 ^ 1'b0 ;
  assign n22939 = n22938 ^ n4010 ^ 1'b0 ;
  assign n22940 = n3626 ^ n1889 ^ 1'b0 ;
  assign n22941 = n6492 & ~n22940 ;
  assign n22942 = n16549 ^ n13977 ^ 1'b0 ;
  assign n22943 = n17702 ^ n4129 ^ 1'b0 ;
  assign n22944 = ~n20045 & n22943 ;
  assign n22945 = n22944 ^ n18108 ^ n13637 ;
  assign n22946 = n21709 ^ n9365 ^ n3246 ;
  assign n22947 = ( n636 & n22945 ) | ( n636 & n22946 ) | ( n22945 & n22946 ) ;
  assign n22948 = n19032 ^ n14944 ^ 1'b0 ;
  assign n22949 = n10986 ^ n739 ^ 1'b0 ;
  assign n22950 = n7198 & n22949 ;
  assign n22951 = ~n2006 & n11748 ;
  assign n22952 = n3382 & n22951 ;
  assign n22953 = n17091 & ~n22952 ;
  assign n22954 = n4550 & n22953 ;
  assign n22955 = n2297 | n9034 ;
  assign n22956 = n22955 ^ n3749 ^ 1'b0 ;
  assign n22957 = ( n428 & ~n2473 ) | ( n428 & n19106 ) | ( ~n2473 & n19106 ) ;
  assign n22958 = x59 & n15820 ;
  assign n22959 = n5913 & n22958 ;
  assign n22960 = ( n9193 & ~n21110 ) | ( n9193 & n22959 ) | ( ~n21110 & n22959 ) ;
  assign n22961 = ( ~n4376 & n21069 ) | ( ~n4376 & n22960 ) | ( n21069 & n22960 ) ;
  assign n22962 = ( n12150 & ~n12337 ) | ( n12150 & n22961 ) | ( ~n12337 & n22961 ) ;
  assign n22963 = ( n4699 & n4760 ) | ( n4699 & n14066 ) | ( n4760 & n14066 ) ;
  assign n22964 = ( n3377 & ~n14777 ) | ( n3377 & n16514 ) | ( ~n14777 & n16514 ) ;
  assign n22965 = n6102 | n11984 ;
  assign n22966 = n22965 ^ n11339 ^ 1'b0 ;
  assign n22967 = x91 & n4859 ;
  assign n22968 = n7894 & n22967 ;
  assign n22969 = n22968 ^ n9483 ^ n6619 ;
  assign n22970 = n4207 & ~n6385 ;
  assign n22971 = n3700 & n22970 ;
  assign n22972 = n20884 & ~n22971 ;
  assign n22973 = n22972 ^ n21452 ^ 1'b0 ;
  assign n22974 = n2030 & ~n8187 ;
  assign n22975 = n9960 & n22974 ;
  assign n22976 = n22975 ^ n20504 ^ n16407 ;
  assign n22977 = ( n22969 & n22973 ) | ( n22969 & n22976 ) | ( n22973 & n22976 ) ;
  assign n22978 = ( n11220 & ~n16885 ) | ( n11220 & n22977 ) | ( ~n16885 & n22977 ) ;
  assign n22979 = ~n2237 & n10398 ;
  assign n22980 = n11708 & ~n22979 ;
  assign n22981 = n22978 & n22980 ;
  assign n22982 = x47 & n5465 ;
  assign n22983 = ( x1 & n8660 ) | ( x1 & n22982 ) | ( n8660 & n22982 ) ;
  assign n22984 = n14076 & n16321 ;
  assign n22985 = ~n22983 & n22984 ;
  assign n22986 = n20484 ^ n2931 ^ n436 ;
  assign n22987 = n15580 ^ n7110 ^ 1'b0 ;
  assign n22988 = n11087 & n20575 ;
  assign n22989 = n22988 ^ n19485 ^ n7174 ;
  assign n22990 = n2353 & n7913 ;
  assign n22991 = n6736 ^ n1204 ^ 1'b0 ;
  assign n22992 = n2894 ^ n2513 ^ 1'b0 ;
  assign n22993 = n22991 | n22992 ;
  assign n22994 = ~n4391 & n12345 ;
  assign n22995 = n9286 & n9931 ;
  assign n22996 = n22995 ^ n3360 ^ 1'b0 ;
  assign n22997 = n22994 & n22996 ;
  assign n22998 = n9507 ^ n4892 ^ 1'b0 ;
  assign n22999 = n589 & ~n22998 ;
  assign n23000 = n22999 ^ n9808 ^ 1'b0 ;
  assign n23001 = n182 | n7334 ;
  assign n23002 = n5799 | n7314 ;
  assign n23003 = n8949 | n23002 ;
  assign n23004 = ( ~n6751 & n6926 ) | ( ~n6751 & n23003 ) | ( n6926 & n23003 ) ;
  assign n23005 = n23004 ^ n1402 ^ 1'b0 ;
  assign n23006 = n23001 & ~n23005 ;
  assign n23007 = n23006 ^ n4921 ^ 1'b0 ;
  assign n23009 = n5022 & ~n11789 ;
  assign n23010 = n8981 & n23009 ;
  assign n23008 = n19455 ^ n8429 ^ 1'b0 ;
  assign n23011 = n23010 ^ n23008 ^ 1'b0 ;
  assign n23012 = n11386 & n23011 ;
  assign n23013 = ( n334 & n5502 ) | ( n334 & ~n23012 ) | ( n5502 & ~n23012 ) ;
  assign n23014 = ~n12616 & n17975 ;
  assign n23015 = n7700 ^ n520 ^ 1'b0 ;
  assign n23016 = n9777 ^ n5227 ^ 1'b0 ;
  assign n23017 = n13333 & ~n23016 ;
  assign n23018 = n23015 & n23017 ;
  assign n23019 = n23018 ^ n9565 ^ 1'b0 ;
  assign n23020 = n22602 ^ n11663 ^ 1'b0 ;
  assign n23021 = ~n8984 & n23020 ;
  assign n23022 = ~n7303 & n22119 ;
  assign n23023 = n22995 & n23022 ;
  assign n23024 = n11949 ^ n2432 ^ 1'b0 ;
  assign n23025 = n23024 ^ n13903 ^ 1'b0 ;
  assign n23026 = n8505 ^ n3033 ^ n1583 ;
  assign n23027 = n15319 ^ n13577 ^ 1'b0 ;
  assign n23028 = n11589 ^ n2227 ^ 1'b0 ;
  assign n23029 = n23028 ^ n10554 ^ n9958 ;
  assign n23030 = n4139 & n23029 ;
  assign n23031 = ( n5614 & ~n14368 ) | ( n5614 & n23030 ) | ( ~n14368 & n23030 ) ;
  assign n23032 = n17734 ^ n7448 ^ n2796 ;
  assign n23033 = n23032 ^ n5640 ^ 1'b0 ;
  assign n23034 = n9511 | n23033 ;
  assign n23035 = n23034 ^ n15533 ^ 1'b0 ;
  assign n23036 = n10917 & ~n23035 ;
  assign n23037 = ( n10777 & n17257 ) | ( n10777 & ~n23036 ) | ( n17257 & ~n23036 ) ;
  assign n23038 = n23037 ^ n19476 ^ x15 ;
  assign n23039 = ( n10920 & ~n10980 ) | ( n10920 & n12089 ) | ( ~n10980 & n12089 ) ;
  assign n23040 = n7513 | n23039 ;
  assign n23041 = n2686 & ~n20538 ;
  assign n23042 = n6600 & n23041 ;
  assign n23043 = n11009 & ~n15990 ;
  assign n23044 = n23043 ^ n5697 ^ 1'b0 ;
  assign n23045 = ( n714 & n7813 ) | ( n714 & ~n23044 ) | ( n7813 & ~n23044 ) ;
  assign n23046 = n1918 | n3557 ;
  assign n23047 = n23046 ^ n4710 ^ 1'b0 ;
  assign n23048 = ( n4888 & n9777 ) | ( n4888 & n10990 ) | ( n9777 & n10990 ) ;
  assign n23049 = ~n12485 & n18486 ;
  assign n23050 = n7513 & n8973 ;
  assign n23051 = n23050 ^ n5080 ^ 1'b0 ;
  assign n23052 = n1751 | n17178 ;
  assign n23053 = ~n8220 & n11023 ;
  assign n23054 = n23053 ^ n10270 ^ 1'b0 ;
  assign n23055 = n23054 ^ n8375 ^ 1'b0 ;
  assign n23056 = ( ~n523 & n13607 ) | ( ~n523 & n23055 ) | ( n13607 & n23055 ) ;
  assign n23057 = n10615 & n15724 ;
  assign n23058 = ~n6895 & n7207 ;
  assign n23059 = n23058 ^ n5944 ^ 1'b0 ;
  assign n23060 = n23059 ^ n19895 ^ n3444 ;
  assign n23061 = ( ~n1909 & n23057 ) | ( ~n1909 & n23060 ) | ( n23057 & n23060 ) ;
  assign n23062 = ( n302 & n11293 ) | ( n302 & ~n12597 ) | ( n11293 & ~n12597 ) ;
  assign n23065 = ( n7496 & ~n7743 ) | ( n7496 & n13296 ) | ( ~n7743 & n13296 ) ;
  assign n23063 = n4691 ^ n2252 ^ 1'b0 ;
  assign n23064 = n6732 | n23063 ;
  assign n23066 = n23065 ^ n23064 ^ 1'b0 ;
  assign n23067 = n5843 & n15589 ;
  assign n23068 = n9770 ^ n4741 ^ 1'b0 ;
  assign n23069 = n23068 ^ n11361 ^ n5601 ;
  assign n23071 = n13747 ^ n656 ^ 1'b0 ;
  assign n23070 = n17692 ^ n16555 ^ n13478 ;
  assign n23072 = n23071 ^ n23070 ^ 1'b0 ;
  assign n23073 = n9296 | n20444 ;
  assign n23074 = n3847 ^ n204 ^ 1'b0 ;
  assign n23075 = n18968 | n23074 ;
  assign n23078 = ( x55 & n14787 ) | ( x55 & n17708 ) | ( n14787 & n17708 ) ;
  assign n23076 = ( ~n1761 & n2498 ) | ( ~n1761 & n21614 ) | ( n2498 & n21614 ) ;
  assign n23077 = n7984 | n23076 ;
  assign n23079 = n23078 ^ n23077 ^ 1'b0 ;
  assign n23080 = ~n6336 & n17572 ;
  assign n23081 = n18022 ^ n3792 ^ n1947 ;
  assign n23082 = ~n7909 & n23081 ;
  assign n23083 = n14949 ^ n5188 ^ 1'b0 ;
  assign n23084 = n8610 | n23083 ;
  assign n23085 = n12166 ^ n9661 ^ n2945 ;
  assign n23086 = ( n7913 & n23084 ) | ( n7913 & n23085 ) | ( n23084 & n23085 ) ;
  assign n23087 = n10341 & n21063 ;
  assign n23088 = n23087 ^ n19129 ^ 1'b0 ;
  assign n23089 = ( n4401 & n5431 ) | ( n4401 & n16019 ) | ( n5431 & n16019 ) ;
  assign n23090 = n9931 & n23089 ;
  assign n23091 = n3121 & ~n23090 ;
  assign n23092 = ( ~n6909 & n7649 ) | ( ~n6909 & n21453 ) | ( n7649 & n21453 ) ;
  assign n23093 = n19443 ^ n17738 ^ n1864 ;
  assign n23094 = ~n915 & n11022 ;
  assign n23095 = n23094 ^ n11241 ^ 1'b0 ;
  assign n23096 = n13330 & ~n17879 ;
  assign n23097 = n16197 & n23096 ;
  assign n23098 = n13864 ^ n8475 ^ n1821 ;
  assign n23099 = ( n21110 & n21914 ) | ( n21110 & n23098 ) | ( n21914 & n23098 ) ;
  assign n23100 = ( ~n2535 & n19841 ) | ( ~n2535 & n23099 ) | ( n19841 & n23099 ) ;
  assign n23101 = ~n2020 & n6420 ;
  assign n23102 = n23101 ^ n19058 ^ 1'b0 ;
  assign n23103 = n11032 & n22803 ;
  assign n23104 = ( n4354 & n7238 ) | ( n4354 & ~n10704 ) | ( n7238 & ~n10704 ) ;
  assign n23105 = n2209 & ~n23104 ;
  assign n23106 = n2059 & n23105 ;
  assign n23107 = n13317 & ~n23106 ;
  assign n23108 = n10792 & n23107 ;
  assign n23109 = n6813 & ~n15666 ;
  assign n23110 = ~n4396 & n23109 ;
  assign n23111 = n15806 ^ n14100 ^ 1'b0 ;
  assign n23112 = n14374 ^ n5245 ^ 1'b0 ;
  assign n23113 = n1364 & ~n23112 ;
  assign n23114 = ( n895 & ~n1822 ) | ( n895 & n17242 ) | ( ~n1822 & n17242 ) ;
  assign n23115 = n19873 & ~n22433 ;
  assign n23116 = n23114 & n23115 ;
  assign n23117 = ( ~n6364 & n7224 ) | ( ~n6364 & n19287 ) | ( n7224 & n19287 ) ;
  assign n23118 = ~n23116 & n23117 ;
  assign n23119 = ( ~n237 & n1124 ) | ( ~n237 & n5023 ) | ( n1124 & n5023 ) ;
  assign n23120 = n4021 & n23119 ;
  assign n23121 = ( ~n2971 & n14522 ) | ( ~n2971 & n23120 ) | ( n14522 & n23120 ) ;
  assign n23122 = ( n1076 & n9731 ) | ( n1076 & n11470 ) | ( n9731 & n11470 ) ;
  assign n23123 = n23122 ^ n14723 ^ n9159 ;
  assign n23124 = ( n7929 & ~n10426 ) | ( n7929 & n23123 ) | ( ~n10426 & n23123 ) ;
  assign n23125 = ~n7719 & n11987 ;
  assign n23126 = n6344 & n23125 ;
  assign n23127 = n14463 ^ n1538 ^ n187 ;
  assign n23128 = n2162 & n23127 ;
  assign n23129 = n17601 & n19172 ;
  assign n23130 = ( ~n9591 & n14084 ) | ( ~n9591 & n19821 ) | ( n14084 & n19821 ) ;
  assign n23135 = n1170 & ~n1493 ;
  assign n23134 = ( n1579 & n3877 ) | ( n1579 & n4650 ) | ( n3877 & n4650 ) ;
  assign n23136 = n23135 ^ n23134 ^ 1'b0 ;
  assign n23137 = n23136 ^ n10297 ^ 1'b0 ;
  assign n23138 = ~n6040 & n10735 ;
  assign n23139 = n2697 | n23138 ;
  assign n23140 = n23139 ^ n13118 ^ 1'b0 ;
  assign n23141 = n23137 | n23140 ;
  assign n23133 = n21621 ^ n7189 ^ 1'b0 ;
  assign n23131 = ~n7898 & n21183 ;
  assign n23132 = n23131 ^ n6665 ^ 1'b0 ;
  assign n23142 = n23141 ^ n23133 ^ n23132 ;
  assign n23143 = n21784 ^ n12447 ^ n213 ;
  assign n23144 = n9134 & ~n23010 ;
  assign n23145 = n23144 ^ n22850 ^ n7060 ;
  assign n23146 = n5154 & n13025 ;
  assign n23147 = n13472 & n23146 ;
  assign n23148 = n4843 ^ n1482 ^ 1'b0 ;
  assign n23149 = n866 | n23148 ;
  assign n23150 = n5949 & n23149 ;
  assign n23151 = n22650 ^ n13178 ^ 1'b0 ;
  assign n23152 = n12515 ^ n10722 ^ n9327 ;
  assign n23153 = ~n1387 & n2124 ;
  assign n23154 = n23153 ^ n15191 ^ n12691 ;
  assign n23155 = ~n23034 & n23154 ;
  assign n23156 = ( n5842 & n9324 ) | ( n5842 & n11894 ) | ( n9324 & n11894 ) ;
  assign n23157 = n15468 & n18438 ;
  assign n23158 = n23157 ^ n14279 ^ n10819 ;
  assign n23159 = ~n927 & n14621 ;
  assign n23160 = n23159 ^ n11276 ^ 1'b0 ;
  assign n23161 = n16748 & ~n23160 ;
  assign n23162 = n12316 ^ n11487 ^ n11246 ;
  assign n23163 = n1205 & n23162 ;
  assign n23164 = n15289 ^ n2769 ^ 1'b0 ;
  assign n23165 = ( n136 & n2419 ) | ( n136 & ~n2666 ) | ( n2419 & ~n2666 ) ;
  assign n23166 = n14589 & ~n23165 ;
  assign n23169 = n6908 ^ n2187 ^ n1062 ;
  assign n23167 = n5263 ^ n934 ^ 1'b0 ;
  assign n23168 = n3862 | n23167 ;
  assign n23170 = n23169 ^ n23168 ^ n1608 ;
  assign n23171 = n23170 ^ n1349 ^ n538 ;
  assign n23172 = n22642 ^ n12463 ^ 1'b0 ;
  assign n23173 = n6835 & ~n18044 ;
  assign n23174 = n23173 ^ n3596 ^ 1'b0 ;
  assign n23175 = ( n4602 & ~n22265 ) | ( n4602 & n23174 ) | ( ~n22265 & n23174 ) ;
  assign n23177 = ( n4629 & n5318 ) | ( n4629 & ~n19461 ) | ( n5318 & ~n19461 ) ;
  assign n23178 = n23177 ^ n13496 ^ n11195 ;
  assign n23176 = n13890 & ~n15908 ;
  assign n23179 = n23178 ^ n23176 ^ 1'b0 ;
  assign n23180 = n7887 ^ n2434 ^ 1'b0 ;
  assign n23181 = n2521 & ~n23180 ;
  assign n23183 = n15549 ^ n9120 ^ n4038 ;
  assign n23182 = n15565 ^ n14252 ^ 1'b0 ;
  assign n23184 = n23183 ^ n23182 ^ n6481 ;
  assign n23185 = ( ~n10946 & n11612 ) | ( ~n10946 & n23184 ) | ( n11612 & n23184 ) ;
  assign n23186 = n23185 ^ n11932 ^ 1'b0 ;
  assign n23187 = n5434 | n23186 ;
  assign n23188 = n11510 ^ n5805 ^ n3715 ;
  assign n23189 = n23188 ^ n4378 ^ 1'b0 ;
  assign n23190 = n11040 ^ n5367 ^ n4351 ;
  assign n23191 = n18849 ^ n10674 ^ n834 ;
  assign n23192 = n9205 ^ n8596 ^ 1'b0 ;
  assign n23193 = ~n2478 & n23192 ;
  assign n23194 = n23193 ^ n14245 ^ 1'b0 ;
  assign n23195 = n19524 & ~n23194 ;
  assign n23196 = x108 & ~n2129 ;
  assign n23197 = ( n12456 & ~n12576 ) | ( n12456 & n14839 ) | ( ~n12576 & n14839 ) ;
  assign n23198 = n6191 | n11999 ;
  assign n23199 = n23197 & ~n23198 ;
  assign n23201 = n12322 ^ n3031 ^ 1'b0 ;
  assign n23200 = n16065 ^ n10640 ^ n5336 ;
  assign n23202 = n23201 ^ n23200 ^ n10677 ;
  assign n23203 = n7816 & ~n18451 ;
  assign n23204 = n8992 & n23203 ;
  assign n23205 = n8372 & ~n8469 ;
  assign n23206 = n17278 & n23205 ;
  assign n23208 = ( n1710 & ~n2499 ) | ( n1710 & n6838 ) | ( ~n2499 & n6838 ) ;
  assign n23209 = n6172 & n23208 ;
  assign n23207 = n6977 & n16063 ;
  assign n23210 = n23209 ^ n23207 ^ 1'b0 ;
  assign n23211 = ( n3148 & n9819 ) | ( n3148 & n17070 ) | ( n9819 & n17070 ) ;
  assign n23212 = ( n11135 & n22152 ) | ( n11135 & n23211 ) | ( n22152 & n23211 ) ;
  assign n23214 = n4331 & ~n5561 ;
  assign n23215 = ~n157 & n23214 ;
  assign n23216 = n22618 ^ n9582 ^ 1'b0 ;
  assign n23217 = ~n23215 & n23216 ;
  assign n23213 = n5491 & ~n16948 ;
  assign n23218 = n23217 ^ n23213 ^ 1'b0 ;
  assign n23219 = n2745 ^ n1499 ^ 1'b0 ;
  assign n23220 = n3192 & ~n23219 ;
  assign n23221 = n7946 & ~n10118 ;
  assign n23222 = n11178 ^ n8868 ^ 1'b0 ;
  assign n23223 = n23222 ^ n1814 ^ 1'b0 ;
  assign n23224 = n23223 ^ n12128 ^ n4335 ;
  assign n23225 = n6312 ^ n2848 ^ 1'b0 ;
  assign n23226 = n14961 ^ n5371 ^ 1'b0 ;
  assign n23227 = n17653 ^ n2065 ^ 1'b0 ;
  assign n23228 = n3052 & n23227 ;
  assign n23229 = ( n6180 & n23226 ) | ( n6180 & n23228 ) | ( n23226 & n23228 ) ;
  assign n23230 = n12795 & ~n16968 ;
  assign n23231 = n826 & n23230 ;
  assign n23232 = n982 & ~n5170 ;
  assign n23233 = n23232 ^ n16875 ^ n12295 ;
  assign n23234 = n6192 ^ n2835 ^ n2354 ;
  assign n23235 = ( ~n3971 & n9016 ) | ( ~n3971 & n23234 ) | ( n9016 & n23234 ) ;
  assign n23236 = n19579 ^ n3780 ^ n2407 ;
  assign n23237 = ( ~n1363 & n6704 ) | ( ~n1363 & n20604 ) | ( n6704 & n20604 ) ;
  assign n23238 = n4215 ^ n4002 ^ n2495 ;
  assign n23239 = ( n2098 & n3358 ) | ( n2098 & n10926 ) | ( n3358 & n10926 ) ;
  assign n23240 = ( n2981 & ~n23238 ) | ( n2981 & n23239 ) | ( ~n23238 & n23239 ) ;
  assign n23241 = ( ~n17485 & n23237 ) | ( ~n17485 & n23240 ) | ( n23237 & n23240 ) ;
  assign n23242 = n7965 & n11500 ;
  assign n23243 = ~n5545 & n23242 ;
  assign n23244 = x51 & ~n22862 ;
  assign n23245 = n23243 & n23244 ;
  assign n23246 = ~n19950 & n22258 ;
  assign n23247 = n9167 & ~n23246 ;
  assign n23248 = n6417 | n20370 ;
  assign n23249 = n4605 | n14874 ;
  assign n23250 = n2965 & ~n23249 ;
  assign n23251 = n9698 ^ n3925 ^ n3777 ;
  assign n23252 = n1159 | n5121 ;
  assign n23253 = n23251 & ~n23252 ;
  assign n23254 = n16600 | n23253 ;
  assign n23256 = n2320 ^ n325 ^ 1'b0 ;
  assign n23257 = n23256 ^ n20353 ^ n12425 ;
  assign n23258 = n887 & n23257 ;
  assign n23255 = n15107 ^ n11408 ^ n977 ;
  assign n23259 = n23258 ^ n23255 ^ n1583 ;
  assign n23260 = n15756 ^ n8029 ^ n5153 ;
  assign n23261 = n23260 ^ n12225 ^ n7661 ;
  assign n23262 = n23261 ^ n19278 ^ n6579 ;
  assign n23263 = n23200 ^ n12828 ^ 1'b0 ;
  assign n23264 = n20801 & n23263 ;
  assign n23265 = ~n7727 & n23264 ;
  assign n23266 = n16615 & n19033 ;
  assign n23267 = ~n11286 & n23266 ;
  assign n23268 = n11068 & ~n16606 ;
  assign n23269 = n20178 | n23268 ;
  assign n23270 = n23269 ^ n5779 ^ 1'b0 ;
  assign n23271 = n5875 & n22221 ;
  assign n23272 = n23271 ^ n2660 ^ 1'b0 ;
  assign n23273 = n14156 | n23272 ;
  assign n23274 = n13049 | n23273 ;
  assign n23275 = ~n4188 & n8312 ;
  assign n23276 = n17997 ^ n5414 ^ n5022 ;
  assign n23277 = ~n23275 & n23276 ;
  assign n23278 = n2793 | n2977 ;
  assign n23285 = n8632 ^ n5635 ^ 1'b0 ;
  assign n23286 = ~n3900 & n23285 ;
  assign n23279 = n7339 ^ n1207 ^ n1076 ;
  assign n23280 = ( n7339 & ~n8003 ) | ( n7339 & n23279 ) | ( ~n8003 & n23279 ) ;
  assign n23281 = n23280 ^ n14651 ^ n7829 ;
  assign n23282 = n23281 ^ n22250 ^ n6100 ;
  assign n23283 = n23282 ^ n13434 ^ n2743 ;
  assign n23284 = n16741 | n23283 ;
  assign n23287 = n23286 ^ n23284 ^ n1799 ;
  assign n23288 = ~n1915 & n11124 ;
  assign n23289 = n23288 ^ n1308 ^ 1'b0 ;
  assign n23290 = n9601 & ~n23289 ;
  assign n23291 = n23290 ^ n7127 ^ 1'b0 ;
  assign n23292 = n2919 & n11894 ;
  assign n23293 = ~n10165 & n23292 ;
  assign n23294 = n13452 ^ n11988 ^ 1'b0 ;
  assign n23295 = ~n23293 & n23294 ;
  assign n23296 = n3756 & n23295 ;
  assign n23297 = n19346 ^ n2998 ^ 1'b0 ;
  assign n23298 = n9955 ^ n9383 ^ n360 ;
  assign n23299 = n23004 ^ n2600 ^ 1'b0 ;
  assign n23300 = ( n1240 & n5360 ) | ( n1240 & ~n15416 ) | ( n5360 & ~n15416 ) ;
  assign n23304 = n4742 ^ n4635 ^ n2286 ;
  assign n23305 = n23304 ^ n763 ^ 1'b0 ;
  assign n23306 = n1379 & n23305 ;
  assign n23301 = n9039 ^ n5690 ^ n4849 ;
  assign n23302 = n13667 | n23301 ;
  assign n23303 = n23302 ^ n9256 ^ 1'b0 ;
  assign n23307 = n23306 ^ n23303 ^ n2967 ;
  assign n23308 = n22155 | n23307 ;
  assign n23309 = ( n7783 & n14745 ) | ( n7783 & ~n21080 ) | ( n14745 & ~n21080 ) ;
  assign n23310 = n23309 ^ n16040 ^ 1'b0 ;
  assign n23312 = n3374 & ~n5915 ;
  assign n23313 = n1939 & n23312 ;
  assign n23311 = ~n3970 & n4621 ;
  assign n23314 = n23313 ^ n23311 ^ 1'b0 ;
  assign n23315 = n2692 ^ n2122 ^ n1902 ;
  assign n23316 = ( n890 & n13988 ) | ( n890 & n23315 ) | ( n13988 & n23315 ) ;
  assign n23317 = ~n1676 & n4020 ;
  assign n23318 = n23316 & n23317 ;
  assign n23319 = ( ~n7028 & n8648 ) | ( ~n7028 & n22345 ) | ( n8648 & n22345 ) ;
  assign n23320 = n19636 ^ n9984 ^ n5586 ;
  assign n23322 = n14908 ^ n9129 ^ 1'b0 ;
  assign n23323 = ~n17376 & n23322 ;
  assign n23321 = n8810 & n10011 ;
  assign n23324 = n23323 ^ n23321 ^ 1'b0 ;
  assign n23325 = n13238 ^ n8576 ^ 1'b0 ;
  assign n23326 = ~n23324 & n23325 ;
  assign n23327 = n11115 ^ n6922 ^ 1'b0 ;
  assign n23328 = n3008 & n23327 ;
  assign n23329 = n7216 ^ n541 ^ 1'b0 ;
  assign n23330 = n11819 & n23329 ;
  assign n23331 = x106 & n5935 ;
  assign n23332 = n23331 ^ n20857 ^ 1'b0 ;
  assign n23333 = n23330 & n23332 ;
  assign n23334 = n15999 ^ n13424 ^ n4135 ;
  assign n23335 = n14944 ^ n9829 ^ n2455 ;
  assign n23336 = n16570 ^ n11820 ^ n631 ;
  assign n23337 = ( n1890 & n22978 ) | ( n1890 & n23336 ) | ( n22978 & n23336 ) ;
  assign n23338 = n3007 ^ n2811 ^ 1'b0 ;
  assign n23339 = ( n9341 & ~n14460 ) | ( n9341 & n23338 ) | ( ~n14460 & n23338 ) ;
  assign n23340 = n6408 & n23339 ;
  assign n23341 = n8894 | n20795 ;
  assign n23342 = n20122 ^ n15792 ^ 1'b0 ;
  assign n23343 = ~n21491 & n23342 ;
  assign n23344 = n3774 ^ n2466 ^ 1'b0 ;
  assign n23345 = n154 | n23344 ;
  assign n23346 = n1833 & ~n23345 ;
  assign n23347 = n10519 ^ n6780 ^ 1'b0 ;
  assign n23348 = n19064 ^ n2598 ^ 1'b0 ;
  assign n23349 = n20611 & ~n23348 ;
  assign n23350 = n3132 ^ n2178 ^ n2025 ;
  assign n23351 = ( ~n1492 & n16717 ) | ( ~n1492 & n23350 ) | ( n16717 & n23350 ) ;
  assign n23352 = n5776 & n20488 ;
  assign n23353 = ( n23349 & ~n23351 ) | ( n23349 & n23352 ) | ( ~n23351 & n23352 ) ;
  assign n23354 = n6557 ^ n1146 ^ 1'b0 ;
  assign n23355 = ~n5562 & n21360 ;
  assign n23356 = n1409 & n10236 ;
  assign n23357 = ~n9830 & n23356 ;
  assign n23358 = n4118 & ~n16772 ;
  assign n23359 = n23357 & n23358 ;
  assign n23360 = n20418 ^ n20046 ^ n17073 ;
  assign n23361 = n12965 ^ n12071 ^ n7796 ;
  assign n23362 = n8066 & ~n9045 ;
  assign n23363 = n8936 | n12954 ;
  assign n23364 = n23363 ^ n9087 ^ n8572 ;
  assign n23365 = n820 ^ n495 ^ 1'b0 ;
  assign n23366 = n9357 & n23365 ;
  assign n23367 = n17396 ^ n2897 ^ 1'b0 ;
  assign n23368 = n10767 & ~n23367 ;
  assign n23369 = n8972 ^ n7520 ^ n5513 ;
  assign n23370 = n4839 & ~n21017 ;
  assign n23371 = n17446 ^ n14558 ^ 1'b0 ;
  assign n23372 = n23371 ^ n12736 ^ 1'b0 ;
  assign n23373 = ~n3517 & n6599 ;
  assign n23374 = ~n6599 & n23373 ;
  assign n23375 = n1404 & ~n23374 ;
  assign n23376 = n4800 & n23375 ;
  assign n23377 = n9069 ^ n1859 ^ 1'b0 ;
  assign n23378 = n23376 | n23377 ;
  assign n23379 = n23378 ^ n22462 ^ 1'b0 ;
  assign n23380 = n6607 & ~n22596 ;
  assign n23381 = ~n7358 & n23380 ;
  assign n23382 = n23381 ^ n16182 ^ 1'b0 ;
  assign n23383 = ( ~n9958 & n11093 ) | ( ~n9958 & n14081 ) | ( n11093 & n14081 ) ;
  assign n23384 = n9135 & n9453 ;
  assign n23385 = n23383 & n23384 ;
  assign n23386 = ~n5076 & n12827 ;
  assign n23387 = ( ~n7373 & n19348 ) | ( ~n7373 & n23386 ) | ( n19348 & n23386 ) ;
  assign n23388 = ( n12829 & ~n13451 ) | ( n12829 & n23387 ) | ( ~n13451 & n23387 ) ;
  assign n23389 = n4802 & n7243 ;
  assign n23390 = n6316 & ~n23389 ;
  assign n23391 = n23390 ^ n12062 ^ n7089 ;
  assign n23392 = n23391 ^ n16351 ^ 1'b0 ;
  assign n23393 = n3791 | n15003 ;
  assign n23394 = ( n1692 & n20009 ) | ( n1692 & n23393 ) | ( n20009 & n23393 ) ;
  assign n23395 = n6378 | n22254 ;
  assign n23396 = n23394 | n23395 ;
  assign n23397 = n23396 ^ n9312 ^ n8512 ;
  assign n23398 = n7303 | n10703 ;
  assign n23399 = n11401 & ~n23398 ;
  assign n23400 = ( ~n9338 & n21274 ) | ( ~n9338 & n23399 ) | ( n21274 & n23399 ) ;
  assign n23401 = x107 & n2859 ;
  assign n23402 = n925 & ~n23401 ;
  assign n23403 = n10368 ^ n7075 ^ 1'b0 ;
  assign n23404 = n3455 & n6214 ;
  assign n23405 = ( ~n3152 & n6570 ) | ( ~n3152 & n12289 ) | ( n6570 & n12289 ) ;
  assign n23406 = ( n16566 & n20687 ) | ( n16566 & n23405 ) | ( n20687 & n23405 ) ;
  assign n23407 = ( n7323 & n12736 ) | ( n7323 & ~n21382 ) | ( n12736 & ~n21382 ) ;
  assign n23408 = n23407 ^ x42 ^ 1'b0 ;
  assign n23409 = n13220 ^ n1150 ^ 1'b0 ;
  assign n23410 = n2693 & n23409 ;
  assign n23411 = n4750 & n23410 ;
  assign n23412 = n23411 ^ n915 ^ 1'b0 ;
  assign n23413 = x96 & n4093 ;
  assign n23414 = n23413 ^ n14376 ^ n12313 ;
  assign n23415 = n17312 & n23414 ;
  assign n23416 = n6167 & ~n23415 ;
  assign n23417 = n3750 & ~n12589 ;
  assign n23418 = n23417 ^ n9708 ^ 1'b0 ;
  assign n23419 = ~n8276 & n23418 ;
  assign n23420 = n2641 & ~n4383 ;
  assign n23421 = n23420 ^ n6210 ^ 1'b0 ;
  assign n23424 = n4029 ^ n1550 ^ 1'b0 ;
  assign n23425 = n9007 | n23424 ;
  assign n23426 = n2282 | n23425 ;
  assign n23422 = n16560 ^ n5815 ^ n4400 ;
  assign n23423 = ~n16571 & n23422 ;
  assign n23427 = n23426 ^ n23423 ^ 1'b0 ;
  assign n23428 = n2838 | n5780 ;
  assign n23431 = n9693 ^ n4482 ^ n747 ;
  assign n23429 = n15917 ^ n5351 ^ 1'b0 ;
  assign n23430 = n14563 & ~n23429 ;
  assign n23432 = n23431 ^ n23430 ^ 1'b0 ;
  assign n23434 = ( n2541 & n4873 ) | ( n2541 & n12143 ) | ( n4873 & n12143 ) ;
  assign n23435 = n23434 ^ n18619 ^ 1'b0 ;
  assign n23433 = n13948 & ~n15729 ;
  assign n23436 = n23435 ^ n23433 ^ 1'b0 ;
  assign n23437 = ( ~n2204 & n13916 ) | ( ~n2204 & n23436 ) | ( n13916 & n23436 ) ;
  assign n23438 = n17415 | n18879 ;
  assign n23439 = ~n1219 & n2682 ;
  assign n23440 = n4230 | n6415 ;
  assign n23441 = n7257 | n23440 ;
  assign n23442 = n23439 & n23441 ;
  assign n23443 = n23442 ^ n22246 ^ 1'b0 ;
  assign n23444 = n6624 ^ n3497 ^ 1'b0 ;
  assign n23445 = n7490 | n23444 ;
  assign n23446 = ~n14497 & n23445 ;
  assign n23452 = n5578 ^ n4854 ^ 1'b0 ;
  assign n23450 = n18511 ^ n3853 ^ 1'b0 ;
  assign n23447 = n1226 & n2607 ;
  assign n23448 = n23447 ^ n3485 ^ 1'b0 ;
  assign n23449 = n13462 & ~n23448 ;
  assign n23451 = n23450 ^ n23449 ^ 1'b0 ;
  assign n23453 = n23452 ^ n23451 ^ n21766 ;
  assign n23454 = ( ~n1067 & n1107 ) | ( ~n1067 & n18451 ) | ( n1107 & n18451 ) ;
  assign n23455 = n20670 ^ n12465 ^ n1849 ;
  assign n23456 = n23455 ^ n13858 ^ n11748 ;
  assign n23457 = n10538 ^ n9394 ^ n7959 ;
  assign n23458 = n19804 ^ n11714 ^ 1'b0 ;
  assign n23459 = ~n7911 & n23458 ;
  assign n23460 = n13095 ^ n3287 ^ 1'b0 ;
  assign n23461 = ( ~n4706 & n4967 ) | ( ~n4706 & n11223 ) | ( n4967 & n11223 ) ;
  assign n23462 = n23461 ^ n5170 ^ n4341 ;
  assign n23463 = ~n7913 & n17280 ;
  assign n23464 = n5268 & ~n23463 ;
  assign n23465 = ~x108 & n23464 ;
  assign n23467 = n2077 & n3149 ;
  assign n23466 = n259 | n4062 ;
  assign n23468 = n23467 ^ n23466 ^ 1'b0 ;
  assign n23469 = n22697 ^ n4890 ^ 1'b0 ;
  assign n23470 = n23468 & n23469 ;
  assign n23471 = ~n15927 & n17384 ;
  assign n23472 = ~n8909 & n23471 ;
  assign n23473 = n2192 | n6452 ;
  assign n23474 = n4154 | n7369 ;
  assign n23475 = n23473 & ~n23474 ;
  assign n23476 = n23475 ^ n874 ^ 1'b0 ;
  assign n23477 = ~n3947 & n23476 ;
  assign n23478 = n23477 ^ n16114 ^ 1'b0 ;
  assign n23479 = n18943 | n23478 ;
  assign n23480 = n4580 | n7593 ;
  assign n23481 = n7622 | n23480 ;
  assign n23482 = n17652 | n23481 ;
  assign n23483 = n2205 & ~n23482 ;
  assign n23484 = n23483 ^ n3924 ^ 1'b0 ;
  assign n23485 = ~n20809 & n23484 ;
  assign n23486 = n14213 | n15875 ;
  assign n23487 = n23486 ^ n8468 ^ n1481 ;
  assign n23488 = n1798 & ~n2597 ;
  assign n23489 = n7832 | n10863 ;
  assign n23490 = n8862 ^ n6274 ^ 1'b0 ;
  assign n23491 = n1819 | n19777 ;
  assign n23492 = n23490 & ~n23491 ;
  assign n23493 = n14826 & ~n18902 ;
  assign n23494 = ~n16915 & n23493 ;
  assign n23495 = n6328 ^ n3644 ^ n2265 ;
  assign n23496 = ~n2535 & n23495 ;
  assign n23497 = n23496 ^ n21382 ^ 1'b0 ;
  assign n23498 = ( ~n3171 & n3179 ) | ( ~n3171 & n18024 ) | ( n3179 & n18024 ) ;
  assign n23499 = ( n2072 & n6268 ) | ( n2072 & n12112 ) | ( n6268 & n12112 ) ;
  assign n23500 = n2107 | n3144 ;
  assign n23501 = n23499 | n23500 ;
  assign n23502 = n23501 ^ n10876 ^ n10258 ;
  assign n23504 = n2311 & n2793 ;
  assign n23503 = n8960 ^ n5749 ^ n2356 ;
  assign n23505 = n23504 ^ n23503 ^ n6109 ;
  assign n23506 = ( n2416 & ~n12080 ) | ( n2416 & n18723 ) | ( ~n12080 & n18723 ) ;
  assign n23507 = n23506 ^ n21202 ^ n9849 ;
  assign n23508 = n4714 | n8348 ;
  assign n23509 = n23507 | n23508 ;
  assign n23510 = n7417 ^ n4247 ^ n3326 ;
  assign n23511 = n23510 ^ n22945 ^ 1'b0 ;
  assign n23512 = n8740 | n20263 ;
  assign n23513 = ( n5826 & n14835 ) | ( n5826 & n23452 ) | ( n14835 & n23452 ) ;
  assign n23514 = n23513 ^ n4227 ^ 1'b0 ;
  assign n23515 = n23514 ^ n20924 ^ n1003 ;
  assign n23516 = n3610 | n22476 ;
  assign n23517 = n2537 | n23516 ;
  assign n23518 = ( ~n9506 & n11470 ) | ( ~n9506 & n23517 ) | ( n11470 & n23517 ) ;
  assign n23519 = ( n3488 & n9001 ) | ( n3488 & n11208 ) | ( n9001 & n11208 ) ;
  assign n23520 = ( n266 & ~n6859 ) | ( n266 & n23519 ) | ( ~n6859 & n23519 ) ;
  assign n23521 = ( n3858 & ~n5023 ) | ( n3858 & n23520 ) | ( ~n5023 & n23520 ) ;
  assign n23522 = ( ~n3741 & n14700 ) | ( ~n3741 & n15795 ) | ( n14700 & n15795 ) ;
  assign n23523 = ( n3542 & ~n15021 ) | ( n3542 & n23522 ) | ( ~n15021 & n23522 ) ;
  assign n23526 = ( n1827 & ~n4098 ) | ( n1827 & n7734 ) | ( ~n4098 & n7734 ) ;
  assign n23524 = n1236 ^ n773 ^ 1'b0 ;
  assign n23525 = n1499 & n23524 ;
  assign n23527 = n23526 ^ n23525 ^ 1'b0 ;
  assign n23528 = n11021 | n23527 ;
  assign n23529 = n23528 ^ n3096 ^ 1'b0 ;
  assign n23530 = n23523 & ~n23529 ;
  assign n23531 = n16813 ^ n16021 ^ n3787 ;
  assign n23532 = n23531 ^ n11227 ^ 1'b0 ;
  assign n23533 = n23261 | n23532 ;
  assign n23534 = n23533 ^ n17884 ^ n259 ;
  assign n23535 = n20988 & n23534 ;
  assign n23538 = ~n3838 & n5209 ;
  assign n23536 = ~n1406 & n7652 ;
  assign n23537 = n12450 & n23536 ;
  assign n23539 = n23538 ^ n23537 ^ n2923 ;
  assign n23540 = n7379 | n23539 ;
  assign n23541 = n23540 ^ n5588 ^ 1'b0 ;
  assign n23542 = n23541 ^ n12258 ^ 1'b0 ;
  assign n23543 = ( ~n2200 & n2522 ) | ( ~n2200 & n14548 ) | ( n2522 & n14548 ) ;
  assign n23544 = n3393 ^ n2132 ^ 1'b0 ;
  assign n23545 = n20579 & ~n23544 ;
  assign n23546 = n16566 ^ n1716 ^ 1'b0 ;
  assign n23547 = ~n23127 & n23546 ;
  assign n23548 = n4661 ^ n3650 ^ 1'b0 ;
  assign n23549 = ~n2121 & n23548 ;
  assign n23550 = ( n10313 & ~n19917 ) | ( n10313 & n23549 ) | ( ~n19917 & n23549 ) ;
  assign n23551 = n2077 & n23550 ;
  assign n23554 = n4289 ^ n2298 ^ 1'b0 ;
  assign n23555 = n6690 ^ n6295 ^ n560 ;
  assign n23556 = ( n2207 & n14582 ) | ( n2207 & ~n23555 ) | ( n14582 & ~n23555 ) ;
  assign n23557 = ( ~n1111 & n23554 ) | ( ~n1111 & n23556 ) | ( n23554 & n23556 ) ;
  assign n23558 = n23557 ^ n6683 ^ 1'b0 ;
  assign n23559 = ~n5291 & n23558 ;
  assign n23552 = ~n1652 & n11775 ;
  assign n23553 = n23552 ^ n17864 ^ 1'b0 ;
  assign n23560 = n23559 ^ n23553 ^ n20480 ;
  assign n23561 = ( n2199 & ~n6931 ) | ( n2199 & n14788 ) | ( ~n6931 & n14788 ) ;
  assign n23562 = n547 | n7685 ;
  assign n23563 = n9674 & ~n23562 ;
  assign n23564 = n23563 ^ n20057 ^ n5537 ;
  assign n23565 = n2112 & ~n2634 ;
  assign n23566 = ( ~n984 & n8155 ) | ( ~n984 & n23565 ) | ( n8155 & n23565 ) ;
  assign n23567 = n9021 | n17112 ;
  assign n23568 = n23566 & ~n23567 ;
  assign n23569 = n23568 ^ n11665 ^ n4923 ;
  assign n23570 = n7350 & ~n12936 ;
  assign n23571 = n14997 ^ n11445 ^ 1'b0 ;
  assign n23572 = n2271 & n9441 ;
  assign n23573 = n23571 & n23572 ;
  assign n23574 = n15268 ^ n6847 ^ n662 ;
  assign n23577 = n22074 ^ n20712 ^ n10816 ;
  assign n23575 = n7794 | n20009 ;
  assign n23576 = n23575 ^ n927 ^ 1'b0 ;
  assign n23578 = n23577 ^ n23576 ^ n15191 ;
  assign n23579 = n22407 & ~n23350 ;
  assign n23580 = ~n4396 & n10977 ;
  assign n23581 = n11518 ^ n10280 ^ 1'b0 ;
  assign n23582 = n20962 ^ n8408 ^ 1'b0 ;
  assign n23583 = n3797 & ~n23582 ;
  assign n23584 = n23583 ^ n3120 ^ 1'b0 ;
  assign n23585 = ~n4414 & n5328 ;
  assign n23586 = ( ~n3086 & n3234 ) | ( ~n3086 & n23585 ) | ( n3234 & n23585 ) ;
  assign n23587 = n4038 & ~n23586 ;
  assign n23588 = n23587 ^ n3073 ^ 1'b0 ;
  assign n23590 = n19154 ^ n13002 ^ n5990 ;
  assign n23591 = ( ~n6642 & n14282 ) | ( ~n6642 & n23590 ) | ( n14282 & n23590 ) ;
  assign n23589 = n4736 & n10152 ;
  assign n23592 = n23591 ^ n23589 ^ 1'b0 ;
  assign n23593 = n12276 ^ n10626 ^ n5169 ;
  assign n23594 = ( n870 & n21210 ) | ( n870 & n23222 ) | ( n21210 & n23222 ) ;
  assign n23595 = n3556 & n11628 ;
  assign n23596 = ( n20841 & n23594 ) | ( n20841 & n23595 ) | ( n23594 & n23595 ) ;
  assign n23597 = ( ~n5755 & n5907 ) | ( ~n5755 & n7650 ) | ( n5907 & n7650 ) ;
  assign n23598 = ( n3468 & n8844 ) | ( n3468 & ~n16139 ) | ( n8844 & ~n16139 ) ;
  assign n23599 = ( ~n641 & n7613 ) | ( ~n641 & n9664 ) | ( n7613 & n9664 ) ;
  assign n23600 = n8062 & ~n23599 ;
  assign n23601 = n23598 & n23600 ;
  assign n23602 = n2874 | n7178 ;
  assign n23603 = n12792 ^ n4884 ^ 1'b0 ;
  assign n23604 = n6956 | n23603 ;
  assign n23605 = n15220 | n23604 ;
  assign n23606 = n1065 & n6694 ;
  assign n23607 = n12730 ^ n11458 ^ n1448 ;
  assign n23608 = ( ~n2419 & n4466 ) | ( ~n2419 & n13038 ) | ( n4466 & n13038 ) ;
  assign n23609 = n23607 & n23608 ;
  assign n23610 = ( n308 & n14569 ) | ( n308 & n22250 ) | ( n14569 & n22250 ) ;
  assign n23611 = ( n5238 & ~n23609 ) | ( n5238 & n23610 ) | ( ~n23609 & n23610 ) ;
  assign n23612 = ( ~n12132 & n16838 ) | ( ~n12132 & n17989 ) | ( n16838 & n17989 ) ;
  assign n23613 = n20444 ^ n5566 ^ 1'b0 ;
  assign n23614 = n7311 | n23613 ;
  assign n23615 = ( n4287 & n8313 ) | ( n4287 & ~n11209 ) | ( n8313 & ~n11209 ) ;
  assign n23616 = n21524 | n23615 ;
  assign n23617 = n2436 & ~n23616 ;
  assign n23618 = ~n9309 & n15770 ;
  assign n23619 = n9556 & ~n16923 ;
  assign n23620 = n16923 & n23619 ;
  assign n23621 = n22971 | n23620 ;
  assign n23622 = n22971 & ~n23621 ;
  assign n23623 = ( n11049 & n21263 ) | ( n11049 & n23622 ) | ( n21263 & n23622 ) ;
  assign n23624 = n14448 | n18660 ;
  assign n23625 = n8055 ^ n1007 ^ 1'b0 ;
  assign n23626 = n1863 | n16149 ;
  assign n23627 = n23626 ^ n3341 ^ 1'b0 ;
  assign n23628 = n23090 ^ n2231 ^ 1'b0 ;
  assign n23629 = ~n6107 & n23628 ;
  assign n23631 = n10172 ^ n2504 ^ 1'b0 ;
  assign n23632 = n14599 ^ n6666 ^ 1'b0 ;
  assign n23633 = n23631 & ~n23632 ;
  assign n23634 = ( n10180 & ~n20788 ) | ( n10180 & n23633 ) | ( ~n20788 & n23633 ) ;
  assign n23630 = n4116 | n6967 ;
  assign n23635 = n23634 ^ n23630 ^ 1'b0 ;
  assign n23636 = n18525 ^ n12140 ^ 1'b0 ;
  assign n23637 = x53 & ~n19742 ;
  assign n23638 = n23637 ^ n18770 ^ n1116 ;
  assign n23639 = ( n12585 & n20374 ) | ( n12585 & n23638 ) | ( n20374 & n23638 ) ;
  assign n23640 = ( n4327 & n6083 ) | ( n4327 & ~n17124 ) | ( n6083 & ~n17124 ) ;
  assign n23643 = n20612 ^ n4583 ^ n2364 ;
  assign n23644 = n8729 & n23643 ;
  assign n23645 = n4701 & n23644 ;
  assign n23652 = n3696 | n16136 ;
  assign n23647 = n13477 ^ n5080 ^ n4080 ;
  assign n23648 = n6746 | n23647 ;
  assign n23649 = ~n1902 & n2607 ;
  assign n23650 = n23648 & n23649 ;
  assign n23651 = n9617 | n23650 ;
  assign n23653 = n23652 ^ n23651 ^ 1'b0 ;
  assign n23646 = n4475 & n6768 ;
  assign n23654 = n23653 ^ n23646 ^ 1'b0 ;
  assign n23655 = ( n11615 & n23645 ) | ( n11615 & n23654 ) | ( n23645 & n23654 ) ;
  assign n23641 = ~n8690 & n8890 ;
  assign n23642 = ( n4239 & n19080 ) | ( n4239 & n23641 ) | ( n19080 & n23641 ) ;
  assign n23656 = n23655 ^ n23642 ^ n10551 ;
  assign n23657 = n4198 | n19165 ;
  assign n23658 = ~n9032 & n21704 ;
  assign n23659 = n9511 & n23658 ;
  assign n23660 = n16358 & n21148 ;
  assign n23661 = ~n10121 & n23660 ;
  assign n23662 = n18447 | n21792 ;
  assign n23663 = n1798 & n21376 ;
  assign n23664 = n23663 ^ n15072 ^ 1'b0 ;
  assign n23665 = ( ~x60 & x67 ) | ( ~x60 & n10445 ) | ( x67 & n10445 ) ;
  assign n23666 = n18200 ^ n6547 ^ n3923 ;
  assign n23667 = ( ~n1240 & n11847 ) | ( ~n1240 & n23289 ) | ( n11847 & n23289 ) ;
  assign n23668 = ~n1530 & n3570 ;
  assign n23669 = n23668 ^ n20048 ^ 1'b0 ;
  assign n23672 = n9942 ^ n4834 ^ n4493 ;
  assign n23670 = ~n3004 & n9546 ;
  assign n23671 = n13632 & n23670 ;
  assign n23673 = n23672 ^ n23671 ^ n22971 ;
  assign n23674 = n23673 ^ n13381 ^ n13166 ;
  assign n23675 = n15328 & n20509 ;
  assign n23676 = n23675 ^ n18834 ^ 1'b0 ;
  assign n23677 = n20015 ^ n16168 ^ 1'b0 ;
  assign n23678 = n22476 | n23677 ;
  assign n23679 = n3286 & ~n23678 ;
  assign n23680 = n10824 ^ n4792 ^ 1'b0 ;
  assign n23681 = n18029 & n23680 ;
  assign n23682 = n23681 ^ n12958 ^ 1'b0 ;
  assign n23683 = ( x98 & n3266 ) | ( x98 & ~n10114 ) | ( n3266 & ~n10114 ) ;
  assign n23684 = ( n10239 & n15018 ) | ( n10239 & ~n23683 ) | ( n15018 & ~n23683 ) ;
  assign n23685 = n11361 ^ n7749 ^ 1'b0 ;
  assign n23686 = n8090 & n23685 ;
  assign n23687 = n23684 & ~n23686 ;
  assign n23688 = n9398 ^ n7866 ^ n3731 ;
  assign n23689 = ( n3229 & ~n5172 ) | ( n3229 & n5575 ) | ( ~n5172 & n5575 ) ;
  assign n23690 = n21509 & ~n23689 ;
  assign n23691 = n15366 ^ n6161 ^ 1'b0 ;
  assign n23692 = n5235 & ~n23691 ;
  assign n23693 = ~n4484 & n8734 ;
  assign n23694 = ~n20335 & n23693 ;
  assign n23695 = ~n11689 & n23694 ;
  assign n23696 = n19197 & ~n23695 ;
  assign n23697 = n9193 | n18281 ;
  assign n23698 = n21319 ^ n20994 ^ 1'b0 ;
  assign n23699 = n20168 ^ n6596 ^ 1'b0 ;
  assign n23700 = n19825 ^ n6760 ^ 1'b0 ;
  assign n23701 = n4300 & ~n23700 ;
  assign n23702 = n4322 | n15496 ;
  assign n23703 = n20348 & ~n23702 ;
  assign n23704 = n23703 ^ n7675 ^ 1'b0 ;
  assign n23705 = n927 | n16376 ;
  assign n23706 = n23705 ^ n8329 ^ n4367 ;
  assign n23707 = n15237 & ~n23706 ;
  assign n23708 = n15053 & ~n23707 ;
  assign n23709 = n23708 ^ n4847 ^ 1'b0 ;
  assign n23710 = n7952 & ~n12297 ;
  assign n23711 = n18406 ^ n13924 ^ 1'b0 ;
  assign n23712 = n13096 ^ n6835 ^ n239 ;
  assign n23715 = n14908 ^ n3741 ^ 1'b0 ;
  assign n23713 = ~n4320 & n13663 ;
  assign n23714 = n6657 & n23713 ;
  assign n23716 = n23715 ^ n23714 ^ n3551 ;
  assign n23717 = n23716 ^ n10076 ^ n3948 ;
  assign n23718 = n20262 ^ n12511 ^ n6847 ;
  assign n23719 = n23718 ^ n13159 ^ n531 ;
  assign n23720 = ( ~n188 & n274 ) | ( ~n188 & n23719 ) | ( n274 & n23719 ) ;
  assign n23721 = ( ~n2463 & n4061 ) | ( ~n2463 & n5818 ) | ( n4061 & n5818 ) ;
  assign n23722 = n23721 ^ n13974 ^ 1'b0 ;
  assign n23723 = n23722 ^ n18133 ^ n12578 ;
  assign n23724 = n1128 & ~n5835 ;
  assign n23725 = n15719 | n23724 ;
  assign n23731 = ( n1057 & ~n1621 ) | ( n1057 & n6609 ) | ( ~n1621 & n6609 ) ;
  assign n23730 = n17664 | n22877 ;
  assign n23732 = n23731 ^ n23730 ^ 1'b0 ;
  assign n23726 = ( n2206 & ~n3463 ) | ( n2206 & n10434 ) | ( ~n3463 & n10434 ) ;
  assign n23727 = n969 & n23726 ;
  assign n23728 = ~n13965 & n23727 ;
  assign n23729 = n20556 & ~n23728 ;
  assign n23733 = n23732 ^ n23729 ^ n3185 ;
  assign n23734 = n14861 ^ n4696 ^ 1'b0 ;
  assign n23735 = n13176 ^ n7521 ^ n1649 ;
  assign n23736 = n23735 ^ n23104 ^ n5433 ;
  assign n23737 = ( n11588 & n23734 ) | ( n11588 & n23736 ) | ( n23734 & n23736 ) ;
  assign n23738 = ( n4118 & n5127 ) | ( n4118 & ~n7489 ) | ( n5127 & ~n7489 ) ;
  assign n23739 = ( n6628 & ~n12734 ) | ( n6628 & n22214 ) | ( ~n12734 & n22214 ) ;
  assign n23740 = ( n2805 & n4385 ) | ( n2805 & ~n23739 ) | ( n4385 & ~n23739 ) ;
  assign n23741 = n19594 ^ n5880 ^ 1'b0 ;
  assign n23742 = ( n1422 & n5827 ) | ( n1422 & n23741 ) | ( n5827 & n23741 ) ;
  assign n23743 = n3848 & n4257 ;
  assign n23744 = n6958 & n23743 ;
  assign n23745 = n13269 ^ n8117 ^ 1'b0 ;
  assign n23746 = n21399 & ~n23745 ;
  assign n23747 = ( ~n20410 & n23744 ) | ( ~n20410 & n23746 ) | ( n23744 & n23746 ) ;
  assign n23748 = n2960 & n12375 ;
  assign n23749 = n4986 & ~n23748 ;
  assign n23750 = n23749 ^ n10704 ^ 1'b0 ;
  assign n23751 = n22818 ^ n13109 ^ 1'b0 ;
  assign n23752 = n23344 | n23751 ;
  assign n23753 = n5427 | n21553 ;
  assign n23754 = n6950 ^ x44 ^ 1'b0 ;
  assign n23755 = x49 & ~n903 ;
  assign n23756 = ~n23754 & n23755 ;
  assign n23757 = ( n548 & ~n4953 ) | ( n548 & n5596 ) | ( ~n4953 & n5596 ) ;
  assign n23758 = n10152 ^ n388 ^ 1'b0 ;
  assign n23759 = n2324 & ~n23758 ;
  assign n23760 = ~n23757 & n23759 ;
  assign n23764 = n6123 & n6809 ;
  assign n23761 = n14691 ^ n14402 ^ 1'b0 ;
  assign n23762 = n11379 ^ n5025 ^ 1'b0 ;
  assign n23763 = ~n23761 & n23762 ;
  assign n23765 = n23764 ^ n23763 ^ 1'b0 ;
  assign n23766 = n16431 ^ n13931 ^ 1'b0 ;
  assign n23773 = n16605 & n19076 ;
  assign n23767 = n3867 | n4405 ;
  assign n23768 = n3212 & ~n23767 ;
  assign n23769 = n5021 & ~n23768 ;
  assign n23770 = n13893 & ~n20169 ;
  assign n23771 = n23770 ^ n3116 ^ 1'b0 ;
  assign n23772 = n23769 | n23771 ;
  assign n23774 = n23773 ^ n23772 ^ n12347 ;
  assign n23775 = n831 & n11790 ;
  assign n23776 = n8878 ^ n5784 ^ n2286 ;
  assign n23777 = n23776 ^ n16141 ^ 1'b0 ;
  assign n23778 = ~n2730 & n3007 ;
  assign n23779 = n23778 ^ n1949 ^ 1'b0 ;
  assign n23780 = n23779 ^ n9637 ^ 1'b0 ;
  assign n23781 = n23777 & n23780 ;
  assign n23782 = n1443 & n23781 ;
  assign n23783 = n13067 ^ n9611 ^ 1'b0 ;
  assign n23784 = n13936 & n19408 ;
  assign n23785 = n14743 ^ n3133 ^ n2711 ;
  assign n23786 = ( ~n318 & n17943 ) | ( ~n318 & n23785 ) | ( n17943 & n23785 ) ;
  assign n23787 = n23786 ^ n4092 ^ 1'b0 ;
  assign n23788 = n9041 & ~n23787 ;
  assign n23789 = n6417 ^ n1287 ^ 1'b0 ;
  assign n23790 = n16071 ^ n3780 ^ 1'b0 ;
  assign n23791 = ~n8745 & n10016 ;
  assign n23792 = ( n6038 & n8340 ) | ( n6038 & ~n18354 ) | ( n8340 & ~n18354 ) ;
  assign n23793 = n11544 ^ n6769 ^ 1'b0 ;
  assign n23794 = n6446 & n23793 ;
  assign n23795 = ( n23177 & n23792 ) | ( n23177 & n23794 ) | ( n23792 & n23794 ) ;
  assign n23796 = n19656 ^ n12030 ^ 1'b0 ;
  assign n23799 = n588 & ~n1827 ;
  assign n23800 = n23799 ^ n4993 ^ 1'b0 ;
  assign n23797 = ~n1914 & n23333 ;
  assign n23798 = n23797 ^ n3911 ^ 1'b0 ;
  assign n23801 = n23800 ^ n23798 ^ n13700 ;
  assign n23802 = n15428 ^ n3259 ^ 1'b0 ;
  assign n23803 = n2156 & ~n23802 ;
  assign n23804 = n8910 ^ n2036 ^ 1'b0 ;
  assign n23805 = n20190 & n23804 ;
  assign n23806 = ~n10640 & n16681 ;
  assign n23807 = n17524 ^ n6311 ^ 1'b0 ;
  assign n23808 = n23806 & ~n23807 ;
  assign n23810 = ( n2956 & n16045 ) | ( n2956 & n17294 ) | ( n16045 & n17294 ) ;
  assign n23809 = ( ~n6178 & n7144 ) | ( ~n6178 & n15325 ) | ( n7144 & n15325 ) ;
  assign n23811 = n23810 ^ n23809 ^ 1'b0 ;
  assign n23812 = n16554 ^ n10374 ^ n763 ;
  assign n23813 = ( ~n4864 & n5355 ) | ( ~n4864 & n10735 ) | ( n5355 & n10735 ) ;
  assign n23814 = n21826 | n23378 ;
  assign n23815 = n2655 & n19598 ;
  assign n23816 = n23815 ^ n3792 ^ 1'b0 ;
  assign n23818 = n21062 ^ n16382 ^ n10990 ;
  assign n23817 = n19609 | n21575 ;
  assign n23819 = n23818 ^ n23817 ^ 1'b0 ;
  assign n23820 = ( n3162 & n5718 ) | ( n3162 & ~n17631 ) | ( n5718 & ~n17631 ) ;
  assign n23821 = n11788 & n13120 ;
  assign n23822 = n23821 ^ n10001 ^ 1'b0 ;
  assign n23823 = n12096 & n23822 ;
  assign n23824 = n23820 | n23823 ;
  assign n23825 = n19252 ^ n1212 ^ 1'b0 ;
  assign n23826 = ~n23824 & n23825 ;
  assign n23827 = ( n6714 & n12376 ) | ( n6714 & n21614 ) | ( n12376 & n21614 ) ;
  assign n23828 = n14282 ^ n5839 ^ 1'b0 ;
  assign n23829 = n23827 & n23828 ;
  assign n23830 = n10720 & n23829 ;
  assign n23831 = n11030 & n16411 ;
  assign n23832 = n11082 ^ n9784 ^ n8719 ;
  assign n23833 = n893 & n23832 ;
  assign n23834 = n3468 | n14654 ;
  assign n23835 = n23834 ^ n15346 ^ 1'b0 ;
  assign n23836 = n23835 ^ n16372 ^ 1'b0 ;
  assign n23837 = ( n1622 & n23833 ) | ( n1622 & ~n23836 ) | ( n23833 & ~n23836 ) ;
  assign n23838 = n9512 ^ n5432 ^ 1'b0 ;
  assign n23839 = n19684 & n23838 ;
  assign n23840 = ~n8572 & n23839 ;
  assign n23841 = ( n21771 & n23837 ) | ( n21771 & ~n23840 ) | ( n23837 & ~n23840 ) ;
  assign n23842 = n8344 | n11573 ;
  assign n23843 = n14266 ^ n9106 ^ n2311 ;
  assign n23844 = n6399 | n23843 ;
  assign n23845 = n21266 | n23844 ;
  assign n23846 = n6235 | n12952 ;
  assign n23847 = n10475 ^ x7 ^ 1'b0 ;
  assign n23848 = ( n8547 & n21374 ) | ( n8547 & n23847 ) | ( n21374 & n23847 ) ;
  assign n23849 = n14213 ^ n7434 ^ 1'b0 ;
  assign n23850 = ~n10270 & n13302 ;
  assign n23851 = n23850 ^ n6128 ^ 1'b0 ;
  assign n23852 = n23851 ^ n23836 ^ n12790 ;
  assign n23853 = n8575 ^ n3121 ^ 1'b0 ;
  assign n23854 = n22938 & n23853 ;
  assign n23855 = n23854 ^ n11503 ^ 1'b0 ;
  assign n23856 = x37 & n23855 ;
  assign n23857 = n23856 ^ n22447 ^ n6586 ;
  assign n23858 = n2015 & ~n14728 ;
  assign n23859 = n23858 ^ n5148 ^ 1'b0 ;
  assign n23860 = n3813 & n23859 ;
  assign n23861 = n6041 & n23860 ;
  assign n23864 = ( n6804 & n8951 ) | ( n6804 & ~n22024 ) | ( n8951 & ~n22024 ) ;
  assign n23862 = n7412 ^ n5657 ^ n1663 ;
  assign n23863 = ~n16944 & n23862 ;
  assign n23865 = n23864 ^ n23863 ^ 1'b0 ;
  assign n23866 = n23865 ^ n8065 ^ n1361 ;
  assign n23867 = n7498 ^ n796 ^ 1'b0 ;
  assign n23868 = n22224 ^ n20380 ^ n17897 ;
  assign n23869 = ( n6605 & ~n10945 ) | ( n6605 & n15145 ) | ( ~n10945 & n15145 ) ;
  assign n23870 = n21691 ^ n2738 ^ 1'b0 ;
  assign n23871 = ( n6697 & n23869 ) | ( n6697 & n23870 ) | ( n23869 & n23870 ) ;
  assign n23872 = n23871 ^ n2199 ^ 1'b0 ;
  assign n23873 = n11062 & n14422 ;
  assign n23874 = n16737 | n23873 ;
  assign n23875 = n23872 | n23874 ;
  assign n23876 = n23875 ^ n15579 ^ 1'b0 ;
  assign n23877 = ( n5672 & n11445 ) | ( n5672 & n12945 ) | ( n11445 & n12945 ) ;
  assign n23878 = n23877 ^ n6946 ^ 1'b0 ;
  assign n23879 = n3515 & ~n23878 ;
  assign n23880 = ~n6715 & n10197 ;
  assign n23881 = n20200 & n23880 ;
  assign n23882 = ( n2371 & n7954 ) | ( n2371 & ~n9245 ) | ( n7954 & ~n9245 ) ;
  assign n23883 = n2408 & n23882 ;
  assign n23884 = n23883 ^ n4354 ^ 1'b0 ;
  assign n23888 = ( n636 & n2860 ) | ( n636 & n9472 ) | ( n2860 & n9472 ) ;
  assign n23885 = ( n9996 & n15079 ) | ( n9996 & n19729 ) | ( n15079 & n19729 ) ;
  assign n23886 = n4752 & ~n23885 ;
  assign n23887 = ~n12397 & n23886 ;
  assign n23889 = n23888 ^ n23887 ^ 1'b0 ;
  assign n23890 = n11223 ^ n8469 ^ 1'b0 ;
  assign n23891 = n15770 & ~n23890 ;
  assign n23892 = n21620 | n23253 ;
  assign n23893 = n23892 ^ n10846 ^ 1'b0 ;
  assign n23894 = n12223 ^ n516 ^ 1'b0 ;
  assign n23895 = n5392 ^ n666 ^ n529 ;
  assign n23896 = n4691 & ~n23895 ;
  assign n23897 = ( n4438 & n23894 ) | ( n4438 & n23896 ) | ( n23894 & n23896 ) ;
  assign n23898 = n19026 ^ n16291 ^ 1'b0 ;
  assign n23899 = n23729 ^ n23338 ^ n5034 ;
  assign n23900 = n10626 ^ n8310 ^ n7244 ;
  assign n23901 = n22210 ^ n13319 ^ n8920 ;
  assign n23902 = ( n577 & n4371 ) | ( n577 & n17686 ) | ( n4371 & n17686 ) ;
  assign n23903 = n15270 | n19139 ;
  assign n23904 = n5118 | n23903 ;
  assign n23905 = ( ~n18961 & n23902 ) | ( ~n18961 & n23904 ) | ( n23902 & n23904 ) ;
  assign n23906 = ~n17629 & n23905 ;
  assign n23907 = n14249 | n15877 ;
  assign n23908 = n23907 ^ n17526 ^ 1'b0 ;
  assign n23909 = n8702 | n11106 ;
  assign n23910 = n15996 & n18887 ;
  assign n23911 = n2081 & n3254 ;
  assign n23912 = n23911 ^ n7800 ^ 1'b0 ;
  assign n23913 = n22235 ^ n9569 ^ n5474 ;
  assign n23916 = ~n2390 & n18254 ;
  assign n23917 = n182 & n23916 ;
  assign n23914 = ( n335 & n588 ) | ( n335 & n3030 ) | ( n588 & n3030 ) ;
  assign n23915 = n23914 ^ n8913 ^ 1'b0 ;
  assign n23918 = n23917 ^ n23915 ^ 1'b0 ;
  assign n23919 = n6547 & ~n22409 ;
  assign n23920 = n2568 & ~n3840 ;
  assign n23921 = n23920 ^ n3716 ^ 1'b0 ;
  assign n23922 = n11825 & n14084 ;
  assign n23923 = ~n3556 & n23922 ;
  assign n23924 = ~n4838 & n6046 ;
  assign n23925 = ~n18355 & n23924 ;
  assign n23926 = n16531 ^ n1323 ^ 1'b0 ;
  assign n23927 = n21263 & n23926 ;
  assign n23928 = n9079 ^ n5377 ^ n2770 ;
  assign n23929 = ( n4166 & n19824 ) | ( n4166 & ~n23928 ) | ( n19824 & ~n23928 ) ;
  assign n23930 = n10440 & ~n17182 ;
  assign n23931 = n12395 | n16024 ;
  assign n23932 = n23931 ^ n16838 ^ n14914 ;
  assign n23933 = ( n11885 & ~n12793 ) | ( n11885 & n23932 ) | ( ~n12793 & n23932 ) ;
  assign n23934 = ( ~n4243 & n20759 ) | ( ~n4243 & n23933 ) | ( n20759 & n23933 ) ;
  assign n23936 = n6921 & n12287 ;
  assign n23937 = n23936 ^ n16029 ^ n2711 ;
  assign n23938 = n23937 ^ n8407 ^ n2162 ;
  assign n23939 = n8267 | n23938 ;
  assign n23940 = n8408 | n23939 ;
  assign n23935 = n695 & ~n5353 ;
  assign n23941 = n23940 ^ n23935 ^ n14095 ;
  assign n23942 = ~n19338 & n23450 ;
  assign n23943 = n23942 ^ n10626 ^ 1'b0 ;
  assign n23944 = n18963 ^ n1218 ^ 1'b0 ;
  assign n23945 = ~n14482 & n23944 ;
  assign n23946 = n16389 & n19322 ;
  assign n23947 = n17266 ^ n7125 ^ 1'b0 ;
  assign n23948 = n22872 ^ n4036 ^ n3813 ;
  assign n23949 = ( n3355 & ~n4438 ) | ( n3355 & n23948 ) | ( ~n4438 & n23948 ) ;
  assign n23950 = n19018 ^ x50 ^ 1'b0 ;
  assign n23951 = n20349 ^ n4066 ^ n3974 ;
  assign n23952 = ( n519 & n9526 ) | ( n519 & ~n19764 ) | ( n9526 & ~n19764 ) ;
  assign n23953 = n23586 | n23952 ;
  assign n23954 = ( ~n2239 & n7833 ) | ( ~n2239 & n9828 ) | ( n7833 & n9828 ) ;
  assign n23955 = n9526 | n23954 ;
  assign n23956 = n1217 | n23955 ;
  assign n23957 = n23956 ^ n19271 ^ 1'b0 ;
  assign n23958 = n3364 | n4230 ;
  assign n23959 = ~n9018 & n12915 ;
  assign n23960 = n23958 & n23959 ;
  assign n23962 = n8126 ^ n5533 ^ 1'b0 ;
  assign n23963 = n10219 & ~n23962 ;
  assign n23961 = ~n5142 & n12116 ;
  assign n23964 = n23963 ^ n23961 ^ 1'b0 ;
  assign n23966 = ~n6918 & n9110 ;
  assign n23965 = n3366 & n20382 ;
  assign n23967 = n23966 ^ n23965 ^ 1'b0 ;
  assign n23968 = n7852 & ~n13727 ;
  assign n23974 = n2375 & ~n6036 ;
  assign n23975 = n23974 ^ n2466 ^ 1'b0 ;
  assign n23969 = n21829 ^ n11976 ^ 1'b0 ;
  assign n23970 = n696 | n23969 ;
  assign n23971 = ( ~n6368 & n7501 ) | ( ~n6368 & n23970 ) | ( n7501 & n23970 ) ;
  assign n23972 = n7756 ^ n912 ^ 1'b0 ;
  assign n23973 = ~n23971 & n23972 ;
  assign n23976 = n23975 ^ n23973 ^ n3347 ;
  assign n23977 = n19956 ^ n2735 ^ 1'b0 ;
  assign n23978 = ~n10934 & n23977 ;
  assign n23979 = ~n4657 & n16190 ;
  assign n23980 = n23979 ^ n15829 ^ n8205 ;
  assign n23981 = n5414 & n16132 ;
  assign n23982 = n23981 ^ n2522 ^ 1'b0 ;
  assign n23983 = ~n14874 & n23982 ;
  assign n23984 = ~n9837 & n23983 ;
  assign n23985 = n21441 ^ n4061 ^ 1'b0 ;
  assign n23987 = n6676 ^ n4077 ^ 1'b0 ;
  assign n23988 = n2699 & ~n23987 ;
  assign n23989 = n3124 & n23988 ;
  assign n23990 = ~n19474 & n23989 ;
  assign n23986 = n1456 & ~n2751 ;
  assign n23991 = n23990 ^ n23986 ^ 1'b0 ;
  assign n23992 = n12330 ^ n11469 ^ n1411 ;
  assign n23993 = n5511 ^ n4379 ^ n851 ;
  assign n23994 = n23993 ^ n21034 ^ 1'b0 ;
  assign n23995 = n14137 & n23994 ;
  assign n23996 = ~n6093 & n23995 ;
  assign n23997 = n23996 ^ n7242 ^ 1'b0 ;
  assign n23998 = ( n17900 & ~n23004 ) | ( n17900 & n23997 ) | ( ~n23004 & n23997 ) ;
  assign n23999 = n14177 ^ n11519 ^ 1'b0 ;
  assign n24000 = n22729 ^ n4689 ^ 1'b0 ;
  assign n24001 = n11758 & n24000 ;
  assign n24002 = n24001 ^ n11374 ^ n3715 ;
  assign n24003 = ( n796 & ~n23999 ) | ( n796 & n24002 ) | ( ~n23999 & n24002 ) ;
  assign n24006 = ( n1275 & n17419 ) | ( n1275 & n20491 ) | ( n17419 & n20491 ) ;
  assign n24004 = n8899 ^ n3001 ^ 1'b0 ;
  assign n24005 = n24004 ^ n23024 ^ n5788 ;
  assign n24007 = n24006 ^ n24005 ^ 1'b0 ;
  assign n24009 = n3808 ^ n2813 ^ n1918 ;
  assign n24008 = n167 & ~n5132 ;
  assign n24010 = n24009 ^ n24008 ^ 1'b0 ;
  assign n24011 = n1364 ^ x56 ^ 1'b0 ;
  assign n24012 = ~n24010 & n24011 ;
  assign n24013 = n6605 & n24012 ;
  assign n24014 = ( n3921 & n10754 ) | ( n3921 & n12473 ) | ( n10754 & n12473 ) ;
  assign n24015 = n1771 & n24014 ;
  assign n24016 = ~n13663 & n24015 ;
  assign n24017 = n13557 & ~n24016 ;
  assign n24018 = n13713 & n24017 ;
  assign n24019 = n8592 ^ n3533 ^ 1'b0 ;
  assign n24020 = ( n9835 & ~n18961 ) | ( n9835 & n24019 ) | ( ~n18961 & n24019 ) ;
  assign n24021 = n2730 & n24020 ;
  assign n24022 = n24021 ^ n12727 ^ 1'b0 ;
  assign n24023 = n18470 & ~n24022 ;
  assign n24024 = n6159 & n18755 ;
  assign n24025 = n10007 ^ n4361 ^ 1'b0 ;
  assign n24026 = n24024 & n24025 ;
  assign n24027 = ~n8187 & n10718 ;
  assign n24028 = ~n13871 & n24027 ;
  assign n24029 = ( n354 & ~n2557 ) | ( n354 & n13489 ) | ( ~n2557 & n13489 ) ;
  assign n24030 = n24029 ^ n8528 ^ 1'b0 ;
  assign n24031 = n1757 & ~n3686 ;
  assign n24032 = n6493 & n24031 ;
  assign n24033 = ( n11962 & n16168 ) | ( n11962 & n24032 ) | ( n16168 & n24032 ) ;
  assign n24034 = ( n613 & n2363 ) | ( n613 & ~n8851 ) | ( n2363 & ~n8851 ) ;
  assign n24046 = n7051 & n11118 ;
  assign n24047 = n17992 & n24046 ;
  assign n24035 = n10053 ^ n8777 ^ 1'b0 ;
  assign n24036 = n1762 & n24035 ;
  assign n24037 = ~n3426 & n8324 ;
  assign n24038 = n1691 & ~n24037 ;
  assign n24039 = n24038 ^ n1023 ^ 1'b0 ;
  assign n24040 = n4227 & ~n7551 ;
  assign n24041 = n3382 & n24040 ;
  assign n24042 = ( ~n2768 & n4878 ) | ( ~n2768 & n10463 ) | ( n4878 & n10463 ) ;
  assign n24043 = ( n10382 & n24041 ) | ( n10382 & ~n24042 ) | ( n24041 & ~n24042 ) ;
  assign n24044 = ( n4100 & n14368 ) | ( n4100 & n24043 ) | ( n14368 & n24043 ) ;
  assign n24045 = ( n24036 & n24039 ) | ( n24036 & ~n24044 ) | ( n24039 & ~n24044 ) ;
  assign n24048 = n24047 ^ n24045 ^ n11083 ;
  assign n24049 = n22449 ^ n2108 ^ 1'b0 ;
  assign n24050 = n12036 | n24049 ;
  assign n24051 = ~n11212 & n23441 ;
  assign n24053 = n6281 ^ n6075 ^ 1'b0 ;
  assign n24054 = n9850 & ~n24053 ;
  assign n24052 = n672 & n11331 ;
  assign n24055 = n24054 ^ n24052 ^ 1'b0 ;
  assign n24056 = n2139 ^ n1382 ^ n141 ;
  assign n24057 = n12872 ^ n5692 ^ n983 ;
  assign n24058 = n24056 & n24057 ;
  assign n24059 = ( n3011 & ~n7579 ) | ( n3011 & n24058 ) | ( ~n7579 & n24058 ) ;
  assign n24060 = ( n452 & n9937 ) | ( n452 & n24059 ) | ( n9937 & n24059 ) ;
  assign n24061 = n11546 ^ n318 ^ 1'b0 ;
  assign n24062 = n21590 & n21595 ;
  assign n24063 = ~n24061 & n24062 ;
  assign n24064 = n22624 ^ n13956 ^ 1'b0 ;
  assign n24065 = ~n1230 & n4227 ;
  assign n24066 = n24065 ^ n16431 ^ 1'b0 ;
  assign n24067 = n15443 ^ n8685 ^ 1'b0 ;
  assign n24068 = n19532 ^ n4044 ^ 1'b0 ;
  assign n24069 = ~n12633 & n24068 ;
  assign n24070 = ( n2975 & ~n16364 ) | ( n2975 & n24069 ) | ( ~n16364 & n24069 ) ;
  assign n24071 = n7753 & n10592 ;
  assign n24072 = ~n4294 & n8632 ;
  assign n24073 = n24072 ^ n18812 ^ 1'b0 ;
  assign n24074 = n24071 | n24073 ;
  assign n24075 = n24074 ^ n3303 ^ n635 ;
  assign n24076 = n11483 ^ n2544 ^ n1687 ;
  assign n24077 = n4240 | n17848 ;
  assign n24078 = n13945 & ~n24077 ;
  assign n24079 = n24078 ^ n9349 ^ 1'b0 ;
  assign n24080 = ~n19996 & n24079 ;
  assign n24081 = n737 & n20130 ;
  assign n24082 = n23757 ^ n8350 ^ 1'b0 ;
  assign n24083 = n16192 ^ n7714 ^ n1853 ;
  assign n24084 = ~n14787 & n24083 ;
  assign n24085 = n12716 ^ n4388 ^ n1199 ;
  assign n24086 = n24085 ^ n10693 ^ n7814 ;
  assign n24087 = ( ~n9938 & n12663 ) | ( ~n9938 & n20349 ) | ( n12663 & n20349 ) ;
  assign n24088 = ~n13033 & n23455 ;
  assign n24089 = n4385 | n10314 ;
  assign n24090 = n24089 ^ n16470 ^ 1'b0 ;
  assign n24091 = ~n22144 & n24090 ;
  assign n24092 = n24091 ^ n2142 ^ 1'b0 ;
  assign n24093 = n4109 ^ n296 ^ 1'b0 ;
  assign n24094 = n1274 | n24093 ;
  assign n24095 = n16852 & n24094 ;
  assign n24096 = n18861 ^ n1058 ^ 1'b0 ;
  assign n24097 = ~n19101 & n24096 ;
  assign n24098 = n12440 ^ n11009 ^ n8298 ;
  assign n24099 = n24098 ^ n3439 ^ 1'b0 ;
  assign n24100 = n2915 | n11656 ;
  assign n24101 = n24100 ^ n22976 ^ 1'b0 ;
  assign n24102 = n15741 ^ n6206 ^ n5776 ;
  assign n24103 = ~n953 & n4756 ;
  assign n24104 = n24103 ^ n5650 ^ 1'b0 ;
  assign n24105 = ( ~n11164 & n11393 ) | ( ~n11164 & n24104 ) | ( n11393 & n24104 ) ;
  assign n24106 = ( ~n21818 & n24102 ) | ( ~n21818 & n24105 ) | ( n24102 & n24105 ) ;
  assign n24107 = n24101 | n24106 ;
  assign n24108 = n3985 ^ n3049 ^ n2466 ;
  assign n24109 = n9563 & ~n24108 ;
  assign n24110 = n11031 ^ n6833 ^ n5953 ;
  assign n24111 = n24110 ^ n11008 ^ n1792 ;
  assign n24112 = n1776 | n7937 ;
  assign n24113 = x12 | n24112 ;
  assign n24114 = n19129 ^ n7726 ^ 1'b0 ;
  assign n24115 = n23049 & ~n23739 ;
  assign n24116 = n24115 ^ n13219 ^ 1'b0 ;
  assign n24119 = n7753 | n13841 ;
  assign n24117 = n7074 & n12971 ;
  assign n24118 = n24117 ^ n15808 ^ 1'b0 ;
  assign n24120 = n24119 ^ n24118 ^ n22183 ;
  assign n24121 = x28 & ~n17510 ;
  assign n24122 = ~n3148 & n24121 ;
  assign n24123 = n24122 ^ n9192 ^ n3831 ;
  assign n24124 = n14225 ^ n7565 ^ n3965 ;
  assign n24125 = n22697 ^ n6669 ^ 1'b0 ;
  assign n24126 = n21072 ^ n16586 ^ 1'b0 ;
  assign n24127 = n17828 & ~n24126 ;
  assign n24128 = ~n4984 & n15163 ;
  assign n24129 = n7413 & n24128 ;
  assign n24130 = n10273 ^ n9520 ^ 1'b0 ;
  assign n24131 = n7104 | n11483 ;
  assign n24132 = n24131 ^ n10368 ^ 1'b0 ;
  assign n24133 = n14055 & n19881 ;
  assign n24134 = n21524 ^ n6403 ^ n5721 ;
  assign n24135 = n24134 ^ n6585 ^ 1'b0 ;
  assign n24136 = n24135 ^ n17471 ^ 1'b0 ;
  assign n24137 = n23200 ^ n16979 ^ n9906 ;
  assign n24142 = n6420 ^ n6072 ^ n5070 ;
  assign n24138 = n1776 | n4614 ;
  assign n24139 = n24138 ^ n13447 ^ 1'b0 ;
  assign n24140 = n24139 ^ n11614 ^ 1'b0 ;
  assign n24141 = ~n23857 & n24140 ;
  assign n24143 = n24142 ^ n24141 ^ 1'b0 ;
  assign n24144 = n24143 ^ n11437 ^ n2257 ;
  assign n24145 = ~n4625 & n13796 ;
  assign n24146 = n24145 ^ n3285 ^ 1'b0 ;
  assign n24147 = ( x59 & n4960 ) | ( x59 & ~n8406 ) | ( n4960 & ~n8406 ) ;
  assign n24148 = n7419 ^ n2486 ^ 1'b0 ;
  assign n24149 = n24147 & ~n24148 ;
  assign n24150 = n16321 ^ n915 ^ 1'b0 ;
  assign n24151 = ( n1905 & n18190 ) | ( n1905 & ~n24150 ) | ( n18190 & ~n24150 ) ;
  assign n24155 = n21828 ^ n13434 ^ n1433 ;
  assign n24153 = ( ~n1830 & n12634 ) | ( ~n1830 & n13368 ) | ( n12634 & n13368 ) ;
  assign n24154 = n24153 ^ n20009 ^ 1'b0 ;
  assign n24152 = n12844 ^ n4629 ^ 1'b0 ;
  assign n24156 = n24155 ^ n24154 ^ n24152 ;
  assign n24157 = n7586 ^ n1840 ^ 1'b0 ;
  assign n24158 = n24157 ^ n12157 ^ n8227 ;
  assign n24159 = ( n5759 & n13462 ) | ( n5759 & ~n24158 ) | ( n13462 & ~n24158 ) ;
  assign n24160 = n9846 ^ n1182 ^ 1'b0 ;
  assign n24161 = n1870 ^ n883 ^ 1'b0 ;
  assign n24162 = n24161 ^ n641 ^ 1'b0 ;
  assign n24163 = ~n1943 & n24162 ;
  assign n24164 = ( n719 & n16584 ) | ( n719 & n17287 ) | ( n16584 & n17287 ) ;
  assign n24165 = ( n18659 & ~n24163 ) | ( n18659 & n24164 ) | ( ~n24163 & n24164 ) ;
  assign n24166 = n19554 & ~n24165 ;
  assign n24167 = ~n20367 & n24166 ;
  assign n24168 = n24167 ^ n12913 ^ 1'b0 ;
  assign n24169 = n24168 ^ n4982 ^ 1'b0 ;
  assign n24170 = n15274 ^ n1710 ^ 1'b0 ;
  assign n24171 = n19138 ^ n2036 ^ n1415 ;
  assign n24174 = ( n4526 & n13244 ) | ( n4526 & ~n15650 ) | ( n13244 & ~n15650 ) ;
  assign n24172 = ~n10582 & n19300 ;
  assign n24173 = ~n992 & n24172 ;
  assign n24175 = n24174 ^ n24173 ^ n20015 ;
  assign n24176 = ~n8789 & n20616 ;
  assign n24177 = n22590 ^ n15355 ^ 1'b0 ;
  assign n24178 = n5702 & n24177 ;
  assign n24179 = n10982 ^ n7119 ^ 1'b0 ;
  assign n24180 = n685 | n11736 ;
  assign n24181 = n24179 | n24180 ;
  assign n24182 = n15862 ^ n7655 ^ n3237 ;
  assign n24183 = ( n11437 & n22391 ) | ( n11437 & n24182 ) | ( n22391 & n24182 ) ;
  assign n24184 = n9627 ^ n7118 ^ 1'b0 ;
  assign n24188 = n6215 & n12376 ;
  assign n24189 = ~n11008 & n24188 ;
  assign n24186 = n18472 ^ n2705 ^ 1'b0 ;
  assign n24185 = n15922 & n20576 ;
  assign n24187 = n24186 ^ n24185 ^ 1'b0 ;
  assign n24190 = n24189 ^ n24187 ^ n2292 ;
  assign n24191 = n14954 ^ n4140 ^ n4129 ;
  assign n24192 = n3407 & ~n5471 ;
  assign n24193 = n24192 ^ n5523 ^ 1'b0 ;
  assign n24197 = n5942 ^ n328 ^ 1'b0 ;
  assign n24198 = n1777 & n24197 ;
  assign n24199 = n24198 ^ n6261 ^ 1'b0 ;
  assign n24196 = n917 & n1739 ;
  assign n24200 = n24199 ^ n24196 ^ 1'b0 ;
  assign n24194 = n3118 & ~n3701 ;
  assign n24195 = ~n3648 & n24194 ;
  assign n24201 = n24200 ^ n24195 ^ 1'b0 ;
  assign n24202 = n7006 & ~n15946 ;
  assign n24203 = n24202 ^ n146 ^ 1'b0 ;
  assign n24204 = n24203 ^ n22365 ^ n9427 ;
  assign n24205 = n24204 ^ n3444 ^ 1'b0 ;
  assign n24206 = ~n6100 & n15808 ;
  assign n24207 = n13798 & n24206 ;
  assign n24208 = ~n925 & n4819 ;
  assign n24209 = n458 | n20994 ;
  assign n24210 = n24209 ^ n1758 ^ 1'b0 ;
  assign n24211 = n24210 ^ n19063 ^ 1'b0 ;
  assign n24212 = n12535 | n24211 ;
  assign n24213 = ( n3136 & n12836 ) | ( n3136 & n19730 ) | ( n12836 & n19730 ) ;
  assign n24214 = ( n1553 & ~n18596 ) | ( n1553 & n24186 ) | ( ~n18596 & n24186 ) ;
  assign n24215 = n5527 & ~n24214 ;
  assign n24216 = n24215 ^ n22424 ^ n21830 ;
  assign n24217 = n14827 ^ n12346 ^ n9962 ;
  assign n24218 = ( n8921 & ~n22404 ) | ( n8921 & n24217 ) | ( ~n22404 & n24217 ) ;
  assign n24219 = n24218 ^ n11805 ^ 1'b0 ;
  assign n24220 = ( ~n1561 & n5833 ) | ( ~n1561 & n12099 ) | ( n5833 & n12099 ) ;
  assign n24221 = n24220 ^ n17260 ^ n15035 ;
  assign n24222 = ( ~n10860 & n11253 ) | ( ~n10860 & n24221 ) | ( n11253 & n24221 ) ;
  assign n24223 = n23160 ^ n21667 ^ n19358 ;
  assign n24224 = ( n3840 & n24101 ) | ( n3840 & n24223 ) | ( n24101 & n24223 ) ;
  assign n24225 = n5823 | n7094 ;
  assign n24226 = n5630 | n24225 ;
  assign n24227 = n7174 | n24226 ;
  assign n24228 = n7747 & n24227 ;
  assign n24229 = n3684 | n24228 ;
  assign n24230 = ( n6295 & ~n6890 ) | ( n6295 & n18879 ) | ( ~n6890 & n18879 ) ;
  assign n24231 = ~n5798 & n24230 ;
  assign n24232 = n4184 | n9529 ;
  assign n24233 = n6495 | n15886 ;
  assign n24234 = ( n9761 & n12289 ) | ( n9761 & n24233 ) | ( n12289 & n24233 ) ;
  assign n24235 = n14700 ^ n2151 ^ 1'b0 ;
  assign n24236 = n4347 | n24235 ;
  assign n24237 = n24236 ^ n14716 ^ n1901 ;
  assign n24238 = n10955 ^ n6953 ^ x83 ;
  assign n24239 = n964 & n24238 ;
  assign n24240 = n5077 | n24239 ;
  assign n24241 = n17796 | n24240 ;
  assign n24242 = n24241 ^ n9673 ^ 1'b0 ;
  assign n24248 = n22154 ^ n17664 ^ n16574 ;
  assign n24249 = n24248 ^ n22988 ^ 1'b0 ;
  assign n24250 = n13340 & n24249 ;
  assign n24244 = n10683 | n15046 ;
  assign n24245 = n24244 ^ n11741 ^ 1'b0 ;
  assign n24243 = n4579 & ~n21643 ;
  assign n24246 = n24245 ^ n24243 ^ 1'b0 ;
  assign n24247 = n23195 & n24246 ;
  assign n24251 = n24250 ^ n24247 ^ 1'b0 ;
  assign n24252 = n17822 ^ n13957 ^ n2871 ;
  assign n24253 = ( n804 & n806 ) | ( n804 & ~n6327 ) | ( n806 & ~n6327 ) ;
  assign n24254 = n24253 ^ n21924 ^ n2072 ;
  assign n24255 = n2348 & n24254 ;
  assign n24256 = n209 & n1772 ;
  assign n24257 = n8992 & n24256 ;
  assign n24258 = ( n3100 & n23230 ) | ( n3100 & ~n24257 ) | ( n23230 & ~n24257 ) ;
  assign n24259 = n24258 ^ n8926 ^ n7462 ;
  assign n24260 = ( n6388 & ~n12036 ) | ( n6388 & n14833 ) | ( ~n12036 & n14833 ) ;
  assign n24261 = n9899 ^ n7520 ^ n1801 ;
  assign n24262 = n3942 & n24261 ;
  assign n24263 = ~n6884 & n24262 ;
  assign n24264 = n482 ^ n305 ^ 1'b0 ;
  assign n24265 = n16038 & n24264 ;
  assign n24266 = n6841 & ~n14954 ;
  assign n24267 = ~n17466 & n24266 ;
  assign n24268 = ~n17250 & n24267 ;
  assign n24271 = ( ~n11539 & n12874 ) | ( ~n11539 & n14518 ) | ( n12874 & n14518 ) ;
  assign n24270 = ~n4080 & n19803 ;
  assign n24272 = n24271 ^ n24270 ^ 1'b0 ;
  assign n24269 = n4263 | n11044 ;
  assign n24273 = n24272 ^ n24269 ^ 1'b0 ;
  assign n24274 = ( n1802 & n3429 ) | ( n1802 & ~n15840 ) | ( n3429 & ~n15840 ) ;
  assign n24275 = ~n10066 & n24274 ;
  assign n24277 = n7734 & n17734 ;
  assign n24278 = ~n12825 & n24277 ;
  assign n24276 = n7082 ^ n6491 ^ 1'b0 ;
  assign n24279 = n24278 ^ n24276 ^ 1'b0 ;
  assign n24280 = ~n9125 & n21364 ;
  assign n24281 = n22818 ^ x36 ^ 1'b0 ;
  assign n24282 = n23456 ^ n18722 ^ 1'b0 ;
  assign n24283 = n24281 | n24282 ;
  assign n24284 = ~n1466 & n18645 ;
  assign n24285 = n2006 | n11568 ;
  assign n24286 = ( n1125 & ~n1443 ) | ( n1125 & n2244 ) | ( ~n1443 & n2244 ) ;
  assign n24289 = n4118 & n17290 ;
  assign n24290 = n24289 ^ n7986 ^ 1'b0 ;
  assign n24288 = n3544 & n13977 ;
  assign n24287 = n16858 ^ x4 ^ 1'b0 ;
  assign n24291 = n24290 ^ n24288 ^ n24287 ;
  assign n24292 = n2671 & ~n22586 ;
  assign n24293 = n24292 ^ n10079 ^ 1'b0 ;
  assign n24294 = n6124 & n24293 ;
  assign n24295 = n24294 ^ n22476 ^ 1'b0 ;
  assign n24296 = n18092 ^ n4597 ^ 1'b0 ;
  assign n24297 = n9314 & ~n24296 ;
  assign n24298 = n24297 ^ n14928 ^ 1'b0 ;
  assign n24299 = n9471 & n20683 ;
  assign n24300 = n4406 & ~n10288 ;
  assign n24301 = n24300 ^ n4174 ^ 1'b0 ;
  assign n24302 = ~n933 & n5730 ;
  assign n24303 = ~n10285 & n24302 ;
  assign n24304 = ( n4858 & ~n13047 ) | ( n4858 & n16199 ) | ( ~n13047 & n16199 ) ;
  assign n24305 = n13628 | n20582 ;
  assign n24306 = n8311 ^ n2706 ^ n1934 ;
  assign n24307 = n21494 ^ n1205 ^ 1'b0 ;
  assign n24308 = n13398 | n24307 ;
  assign n24309 = n8928 ^ n6962 ^ n5322 ;
  assign n24310 = n10002 ^ n5088 ^ 1'b0 ;
  assign n24311 = ~n24309 & n24310 ;
  assign n24312 = ( n24306 & ~n24308 ) | ( n24306 & n24311 ) | ( ~n24308 & n24311 ) ;
  assign n24313 = ~n2154 & n18131 ;
  assign n24315 = ~n4087 & n20957 ;
  assign n24316 = n24315 ^ n1252 ^ 1'b0 ;
  assign n24314 = n20607 ^ n2175 ^ 1'b0 ;
  assign n24317 = n24316 ^ n24314 ^ n22172 ;
  assign n24318 = n16447 ^ n11535 ^ n707 ;
  assign n24319 = n24318 ^ n21115 ^ 1'b0 ;
  assign n24320 = n1289 | n4980 ;
  assign n24321 = ( n1496 & n12269 ) | ( n1496 & n15458 ) | ( n12269 & n15458 ) ;
  assign n24322 = n2638 & ~n24321 ;
  assign n24323 = ~n6515 & n24322 ;
  assign n24324 = n4243 | n19426 ;
  assign n24325 = n11319 | n17010 ;
  assign n24326 = n24325 ^ n144 ^ 1'b0 ;
  assign n24327 = n8093 & ~n16387 ;
  assign n24328 = n3502 & n24327 ;
  assign n24329 = ( n10469 & ~n15804 ) | ( n10469 & n24328 ) | ( ~n15804 & n24328 ) ;
  assign n24330 = ( n4432 & ~n4436 ) | ( n4432 & n5249 ) | ( ~n4436 & n5249 ) ;
  assign n24331 = n24330 ^ n23180 ^ 1'b0 ;
  assign n24332 = n14691 | n17758 ;
  assign n24334 = n15371 ^ n15193 ^ 1'b0 ;
  assign n24333 = n12018 | n13595 ;
  assign n24335 = n24334 ^ n24333 ^ 1'b0 ;
  assign n24336 = n3633 & ~n7096 ;
  assign n24337 = n982 | n7711 ;
  assign n24338 = n24337 ^ n14644 ^ 1'b0 ;
  assign n24339 = n15526 ^ n1345 ^ 1'b0 ;
  assign n24340 = ( n6293 & n10730 ) | ( n6293 & ~n24339 ) | ( n10730 & ~n24339 ) ;
  assign n24341 = n24340 ^ n15076 ^ 1'b0 ;
  assign n24342 = n11733 & n24341 ;
  assign n24343 = n871 | n11261 ;
  assign n24344 = ~n3752 & n14814 ;
  assign n24345 = n7516 & n24344 ;
  assign n24346 = n3626 & ~n14012 ;
  assign n24347 = n171 & n24346 ;
  assign n24348 = ~n10238 & n24347 ;
  assign n24349 = n24345 & ~n24348 ;
  assign n24352 = n1962 & n5546 ;
  assign n24350 = ~n10855 & n12759 ;
  assign n24351 = n24350 ^ n15881 ^ 1'b0 ;
  assign n24353 = n24352 ^ n24351 ^ n22703 ;
  assign n24354 = n5210 ^ n2419 ^ 1'b0 ;
  assign n24355 = n18022 & ~n24354 ;
  assign n24356 = ( n8793 & n13285 ) | ( n8793 & ~n14801 ) | ( n13285 & ~n14801 ) ;
  assign n24357 = n18906 ^ n7900 ^ 1'b0 ;
  assign n24358 = ~n2703 & n11879 ;
  assign n24359 = x2 & n3629 ;
  assign n24360 = n24359 ^ n1212 ^ 1'b0 ;
  assign n24361 = n4125 ^ n3632 ^ 1'b0 ;
  assign n24362 = n24360 & n24361 ;
  assign n24363 = n5219 | n16738 ;
  assign n24364 = n17179 ^ n16091 ^ n12543 ;
  assign n24365 = n4823 ^ n4061 ^ n2502 ;
  assign n24366 = n24365 ^ n22623 ^ n11159 ;
  assign n24367 = ~n3858 & n22458 ;
  assign n24369 = n2520 ^ n1092 ^ 1'b0 ;
  assign n24370 = n19342 & n24369 ;
  assign n24368 = ~n916 & n9350 ;
  assign n24371 = n24370 ^ n24368 ^ 1'b0 ;
  assign n24372 = ~n14643 & n17093 ;
  assign n24378 = n7994 ^ n889 ^ 1'b0 ;
  assign n24374 = ( n8019 & n8133 ) | ( n8019 & n10451 ) | ( n8133 & n10451 ) ;
  assign n24373 = n3505 & ~n9398 ;
  assign n24375 = n24374 ^ n24373 ^ 1'b0 ;
  assign n24376 = n24375 ^ n12336 ^ n953 ;
  assign n24377 = n24376 ^ n8640 ^ 1'b0 ;
  assign n24379 = n24378 ^ n24377 ^ n23835 ;
  assign n24380 = ~n6385 & n24379 ;
  assign n24385 = n19031 ^ n10593 ^ 1'b0 ;
  assign n24381 = n2878 ^ n1839 ^ 1'b0 ;
  assign n24382 = n24381 ^ n10231 ^ 1'b0 ;
  assign n24383 = n1783 | n24382 ;
  assign n24384 = n24383 ^ n4859 ^ 1'b0 ;
  assign n24386 = n24385 ^ n24384 ^ n23786 ;
  assign n24387 = ( n2284 & ~n13878 ) | ( n2284 & n23840 ) | ( ~n13878 & n23840 ) ;
  assign n24388 = n16162 ^ n13684 ^ 1'b0 ;
  assign n24389 = n4348 & n24388 ;
  assign n24390 = ~n2670 & n24389 ;
  assign n24391 = n24390 ^ n10229 ^ 1'b0 ;
  assign n24392 = n24391 ^ n22952 ^ n17516 ;
  assign n24393 = n12407 ^ n8408 ^ 1'b0 ;
  assign n24394 = n12218 | n24393 ;
  assign n24395 = n16072 ^ n14140 ^ n10200 ;
  assign n24396 = n16412 & ~n24395 ;
  assign n24397 = n10324 | n24396 ;
  assign n24398 = n12150 ^ n10213 ^ n1280 ;
  assign n24399 = n1493 | n24398 ;
  assign n24400 = n24399 ^ n15295 ^ 1'b0 ;
  assign n24401 = ( n10529 & n16630 ) | ( n10529 & n20766 ) | ( n16630 & n20766 ) ;
  assign n24402 = ( ~n10668 & n15661 ) | ( ~n10668 & n16467 ) | ( n15661 & n16467 ) ;
  assign n24403 = n10787 & n24402 ;
  assign n24404 = ( n465 & n1209 ) | ( n465 & n17570 ) | ( n1209 & n17570 ) ;
  assign n24405 = ~n22600 & n24404 ;
  assign n24406 = ( n8593 & n24403 ) | ( n8593 & n24405 ) | ( n24403 & n24405 ) ;
  assign n24407 = n9378 & n16827 ;
  assign n24409 = n7720 ^ n3221 ^ n1521 ;
  assign n24410 = ( ~n6281 & n12510 ) | ( ~n6281 & n24409 ) | ( n12510 & n24409 ) ;
  assign n24408 = n725 | n8183 ;
  assign n24411 = n24410 ^ n24408 ^ n1318 ;
  assign n24412 = ( ~n3616 & n5766 ) | ( ~n3616 & n13713 ) | ( n5766 & n13713 ) ;
  assign n24413 = n3499 | n24412 ;
  assign n24414 = n24413 ^ n1006 ^ 1'b0 ;
  assign n24415 = n16023 ^ n15786 ^ n997 ;
  assign n24416 = n24415 ^ n5322 ^ 1'b0 ;
  assign n24417 = n24416 ^ n21875 ^ n21226 ;
  assign n24418 = n21625 ^ n15589 ^ 1'b0 ;
  assign n24419 = ~n24417 & n24418 ;
  assign n24420 = n4034 & n22449 ;
  assign n24421 = n12550 & n24420 ;
  assign n24422 = ~n8154 & n11243 ;
  assign n24423 = x93 & ~n3746 ;
  assign n24424 = n24423 ^ n11701 ^ 1'b0 ;
  assign n24425 = n24422 | n24424 ;
  assign n24426 = n13953 & ~n14582 ;
  assign n24427 = n24426 ^ n19017 ^ 1'b0 ;
  assign n24428 = ( n6578 & n22252 ) | ( n6578 & ~n23757 ) | ( n22252 & ~n23757 ) ;
  assign n24429 = n19068 | n24428 ;
  assign n24430 = n18724 & ~n24429 ;
  assign n24431 = n17814 ^ n4222 ^ n3340 ;
  assign n24432 = n23988 ^ n1523 ^ 1'b0 ;
  assign n24433 = ~n2931 & n3829 ;
  assign n24434 = n24433 ^ n14098 ^ n1609 ;
  assign n24435 = n8344 ^ n3757 ^ 1'b0 ;
  assign n24436 = n10869 ^ n6420 ^ 1'b0 ;
  assign n24437 = n10329 | n24436 ;
  assign n24438 = ( n3416 & n9460 ) | ( n3416 & ~n20497 ) | ( n9460 & ~n20497 ) ;
  assign n24439 = n20603 ^ n19902 ^ 1'b0 ;
  assign n24440 = n24438 & ~n24439 ;
  assign n24441 = n19962 ^ n15654 ^ n2889 ;
  assign n24443 = n7913 & n23208 ;
  assign n24442 = n12973 ^ n6500 ^ 1'b0 ;
  assign n24444 = n24443 ^ n24442 ^ n14902 ;
  assign n24445 = n9155 ^ n8963 ^ 1'b0 ;
  assign n24446 = n5420 | n24445 ;
  assign n24447 = n21001 | n24446 ;
  assign n24448 = n2971 & ~n24447 ;
  assign n24449 = x52 & ~n12627 ;
  assign n24450 = n24449 ^ n10857 ^ 1'b0 ;
  assign n24451 = ( n158 & n16475 ) | ( n158 & n24450 ) | ( n16475 & n24450 ) ;
  assign n24452 = n24102 ^ n15888 ^ 1'b0 ;
  assign n24453 = n13894 ^ n2370 ^ 1'b0 ;
  assign n24454 = ~n24452 & n24453 ;
  assign n24455 = ~n8359 & n10176 ;
  assign n24456 = n24455 ^ n7284 ^ 1'b0 ;
  assign n24457 = n11022 & n22022 ;
  assign n24458 = n24457 ^ n12225 ^ 1'b0 ;
  assign n24459 = n8721 ^ n8308 ^ 1'b0 ;
  assign n24460 = ( n1620 & ~n12406 ) | ( n1620 & n16266 ) | ( ~n12406 & n16266 ) ;
  assign n24461 = ~n17617 & n24460 ;
  assign n24462 = ( n2929 & ~n20435 ) | ( n2929 & n24461 ) | ( ~n20435 & n24461 ) ;
  assign n24463 = n9159 ^ n4013 ^ n3775 ;
  assign n24464 = ( ~n1959 & n6895 ) | ( ~n1959 & n17627 ) | ( n6895 & n17627 ) ;
  assign n24465 = n24464 ^ n1632 ^ 1'b0 ;
  assign n24466 = ~n5305 & n11027 ;
  assign n24467 = n24090 ^ n10624 ^ n5186 ;
  assign n24468 = n24467 ^ n13368 ^ n1562 ;
  assign n24469 = ( n12932 & n19311 ) | ( n12932 & n24468 ) | ( n19311 & n24468 ) ;
  assign n24470 = n13119 ^ n3838 ^ 1'b0 ;
  assign n24471 = ~n20716 & n24470 ;
  assign n24472 = n15735 & n24471 ;
  assign n24473 = n18655 ^ n1110 ^ 1'b0 ;
  assign n24474 = n24473 ^ n14790 ^ n12735 ;
  assign n24475 = n11565 ^ n2371 ^ 1'b0 ;
  assign n24476 = n24474 | n24475 ;
  assign n24482 = ( n1760 & ~n11890 ) | ( n1760 & n20744 ) | ( ~n11890 & n20744 ) ;
  assign n24477 = n7112 ^ n3958 ^ 1'b0 ;
  assign n24478 = n5890 & n24477 ;
  assign n24479 = ~n12150 & n24478 ;
  assign n24480 = n14539 & n24479 ;
  assign n24481 = n24480 ^ n22613 ^ 1'b0 ;
  assign n24483 = n24482 ^ n24481 ^ n20275 ;
  assign n24484 = n24483 ^ n4148 ^ 1'b0 ;
  assign n24485 = n9937 & ~n24484 ;
  assign n24486 = n9069 ^ n2737 ^ 1'b0 ;
  assign n24487 = ~n10428 & n24486 ;
  assign n24488 = n3925 & n6909 ;
  assign n24489 = n24488 ^ n10120 ^ 1'b0 ;
  assign n24490 = ~n2337 & n24489 ;
  assign n24491 = ~x110 & n24490 ;
  assign n24492 = ( n1314 & n9661 ) | ( n1314 & n24491 ) | ( n9661 & n24491 ) ;
  assign n24493 = ( n1485 & n6145 ) | ( n1485 & ~n6148 ) | ( n6145 & ~n6148 ) ;
  assign n24494 = ( n8391 & n18883 ) | ( n8391 & ~n24493 ) | ( n18883 & ~n24493 ) ;
  assign n24495 = n10980 ^ n10581 ^ 1'b0 ;
  assign n24496 = ( n5805 & n6485 ) | ( n5805 & ~n16344 ) | ( n6485 & ~n16344 ) ;
  assign n24497 = ~n610 & n16963 ;
  assign n24498 = n24497 ^ n23955 ^ 1'b0 ;
  assign n24499 = ( n3095 & ~n4543 ) | ( n3095 & n13393 ) | ( ~n4543 & n13393 ) ;
  assign n24500 = n5121 ^ n708 ^ 1'b0 ;
  assign n24501 = n9177 | n24500 ;
  assign n24502 = n24499 & ~n24501 ;
  assign n24503 = n22898 ^ n18041 ^ 1'b0 ;
  assign n24504 = n18057 ^ n4557 ^ n1915 ;
  assign n24505 = ( ~n11489 & n14455 ) | ( ~n11489 & n19129 ) | ( n14455 & n19129 ) ;
  assign n24506 = ~n21470 & n24505 ;
  assign n24507 = n20054 ^ n2844 ^ 1'b0 ;
  assign n24508 = n20043 ^ n4082 ^ 1'b0 ;
  assign n24509 = n21729 & n24508 ;
  assign n24510 = n24507 & n24509 ;
  assign n24518 = n3441 ^ x12 ^ 1'b0 ;
  assign n24519 = ~n9245 & n24518 ;
  assign n24511 = n12254 | n14804 ;
  assign n24512 = n18846 | n24511 ;
  assign n24513 = n24512 ^ n7532 ^ x127 ;
  assign n24514 = ~n2243 & n24513 ;
  assign n24515 = n9860 & ~n24514 ;
  assign n24516 = n24515 ^ n23134 ^ 1'b0 ;
  assign n24517 = n4851 | n24516 ;
  assign n24520 = n24519 ^ n24517 ^ 1'b0 ;
  assign n24521 = n3553 & n3606 ;
  assign n24522 = n24521 ^ n6827 ^ 1'b0 ;
  assign n24523 = n6821 ^ n4376 ^ 1'b0 ;
  assign n24524 = n5509 & n24523 ;
  assign n24525 = n24524 ^ n6340 ^ 1'b0 ;
  assign n24526 = ( ~n10120 & n24522 ) | ( ~n10120 & n24525 ) | ( n24522 & n24525 ) ;
  assign n24528 = n5687 & n11961 ;
  assign n24527 = n3668 & ~n4594 ;
  assign n24529 = n24528 ^ n24527 ^ 1'b0 ;
  assign n24530 = n24529 ^ n16698 ^ 1'b0 ;
  assign n24533 = n12344 ^ n2668 ^ 1'b0 ;
  assign n24531 = n22759 ^ n22476 ^ n8429 ;
  assign n24532 = n10141 & ~n24531 ;
  assign n24534 = n24533 ^ n24532 ^ n3485 ;
  assign n24535 = n5837 ^ n1901 ^ 1'b0 ;
  assign n24536 = n1065 & ~n24535 ;
  assign n24537 = n24536 ^ n3391 ^ 1'b0 ;
  assign n24538 = n5900 | n24537 ;
  assign n24539 = n15187 ^ n6669 ^ 1'b0 ;
  assign n24540 = ( n4861 & ~n16929 ) | ( n4861 & n24539 ) | ( ~n16929 & n24539 ) ;
  assign n24541 = n24540 ^ n3429 ^ 1'b0 ;
  assign n24542 = ~n3514 & n24541 ;
  assign n24543 = n8578 & ~n20392 ;
  assign n24544 = n24543 ^ n6330 ^ 1'b0 ;
  assign n24545 = n8198 | n11193 ;
  assign n24546 = n24545 ^ n4960 ^ 1'b0 ;
  assign n24547 = n8117 ^ n3467 ^ 1'b0 ;
  assign n24548 = n24546 | n24547 ;
  assign n24549 = n24548 ^ n15927 ^ 1'b0 ;
  assign n24550 = ~n19208 & n24549 ;
  assign n24551 = n15629 ^ n7763 ^ 1'b0 ;
  assign n24552 = n10699 | n24551 ;
  assign n24553 = n4336 | n20119 ;
  assign n24554 = n4296 & ~n10582 ;
  assign n24555 = ~n24553 & n24554 ;
  assign n24556 = ( n1276 & ~n5857 ) | ( n1276 & n24555 ) | ( ~n5857 & n24555 ) ;
  assign n24557 = n24556 ^ n15632 ^ 1'b0 ;
  assign n24558 = n23781 & ~n24557 ;
  assign n24559 = ( n441 & n4137 ) | ( n441 & n15219 ) | ( n4137 & n15219 ) ;
  assign n24560 = ( n1451 & n9327 ) | ( n1451 & n22903 ) | ( n9327 & n22903 ) ;
  assign n24561 = ( n8791 & ~n17744 ) | ( n8791 & n24560 ) | ( ~n17744 & n24560 ) ;
  assign n24563 = n7705 | n23728 ;
  assign n24564 = n24563 ^ n18363 ^ 1'b0 ;
  assign n24562 = ~n6140 & n11119 ;
  assign n24565 = n24564 ^ n24562 ^ 1'b0 ;
  assign n24566 = n15650 ^ n5886 ^ 1'b0 ;
  assign n24567 = n24566 ^ n6418 ^ 1'b0 ;
  assign n24568 = ~n5914 & n24567 ;
  assign n24569 = n8301 & ~n15674 ;
  assign n24570 = ~n15306 & n24569 ;
  assign n24571 = ( n393 & n1050 ) | ( n393 & n11566 ) | ( n1050 & n11566 ) ;
  assign n24572 = n24571 ^ n7874 ^ n3971 ;
  assign n24573 = n7647 & ~n12376 ;
  assign n24574 = n24573 ^ n8765 ^ n431 ;
  assign n24575 = ( ~n10411 & n10866 ) | ( ~n10411 & n12329 ) | ( n10866 & n12329 ) ;
  assign n24576 = n24575 ^ n14455 ^ n12913 ;
  assign n24577 = n24576 ^ n7738 ^ 1'b0 ;
  assign n24581 = n10874 ^ n9726 ^ n6910 ;
  assign n24578 = n7903 ^ n3131 ^ 1'b0 ;
  assign n24579 = n22726 & ~n24578 ;
  assign n24580 = ( n8394 & ~n10547 ) | ( n8394 & n24579 ) | ( ~n10547 & n24579 ) ;
  assign n24582 = n24581 ^ n24580 ^ 1'b0 ;
  assign n24583 = n3892 & n11753 ;
  assign n24584 = n4822 & n24583 ;
  assign n24585 = n16313 ^ n1566 ^ 1'b0 ;
  assign n24586 = ( n5349 & n9628 ) | ( n5349 & n24585 ) | ( n9628 & n24585 ) ;
  assign n24587 = ~n800 & n3494 ;
  assign n24588 = n24586 & n24587 ;
  assign n24589 = ( x53 & n7148 ) | ( x53 & n23832 ) | ( n7148 & n23832 ) ;
  assign n24590 = ( n1864 & ~n6353 ) | ( n1864 & n24589 ) | ( ~n6353 & n24589 ) ;
  assign n24591 = ( ~n1017 & n3110 ) | ( ~n1017 & n7679 ) | ( n3110 & n7679 ) ;
  assign n24594 = ( n8164 & n13296 ) | ( n8164 & ~n15662 ) | ( n13296 & ~n15662 ) ;
  assign n24592 = ~n8845 & n10777 ;
  assign n24593 = n24592 ^ n8691 ^ 1'b0 ;
  assign n24595 = n24594 ^ n24593 ^ 1'b0 ;
  assign n24596 = ~n2545 & n9142 ;
  assign n24597 = n13109 | n18336 ;
  assign n24598 = n24597 ^ n6048 ^ 1'b0 ;
  assign n24599 = n8705 ^ n3415 ^ 1'b0 ;
  assign n24600 = ~n8256 & n12540 ;
  assign n24601 = ~n5136 & n24600 ;
  assign n24602 = n8199 | n21085 ;
  assign n24603 = n17572 ^ n16256 ^ n13445 ;
  assign n24604 = ( x113 & n2934 ) | ( x113 & n10258 ) | ( n2934 & n10258 ) ;
  assign n24605 = n19284 ^ n11841 ^ n4735 ;
  assign n24606 = n24605 ^ n12662 ^ 1'b0 ;
  assign n24607 = n24446 ^ n24002 ^ n9931 ;
  assign n24614 = n13369 & ~n20132 ;
  assign n24615 = ~n3084 & n24614 ;
  assign n24608 = n5428 & n9303 ;
  assign n24609 = n24608 ^ n1920 ^ 1'b0 ;
  assign n24610 = n8343 ^ n6140 ^ 1'b0 ;
  assign n24611 = ~n5071 & n24610 ;
  assign n24612 = ~n3633 & n24611 ;
  assign n24613 = n24609 & n24612 ;
  assign n24616 = n24615 ^ n24613 ^ 1'b0 ;
  assign n24617 = n10587 & ~n24616 ;
  assign n24618 = ( n11978 & n15492 ) | ( n11978 & n24617 ) | ( n15492 & n24617 ) ;
  assign n24619 = ( n1842 & ~n7122 ) | ( n1842 & n24455 ) | ( ~n7122 & n24455 ) ;
  assign n24620 = n18435 ^ n2834 ^ 1'b0 ;
  assign n24621 = ( n19615 & n19924 ) | ( n19615 & n24620 ) | ( n19924 & n24620 ) ;
  assign n24622 = n24621 ^ n12995 ^ 1'b0 ;
  assign n24623 = n7315 ^ n5727 ^ 1'b0 ;
  assign n24624 = n7415 | n24623 ;
  assign n24625 = ( n969 & n10413 ) | ( n969 & ~n14697 ) | ( n10413 & ~n14697 ) ;
  assign n24626 = ~n12908 & n24625 ;
  assign n24627 = n24626 ^ n16787 ^ 1'b0 ;
  assign n24628 = n5354 | n12869 ;
  assign n24629 = n24628 ^ n24447 ^ 1'b0 ;
  assign n24630 = n11415 & ~n21309 ;
  assign n24631 = ( n7863 & n10950 ) | ( n7863 & n11155 ) | ( n10950 & n11155 ) ;
  assign n24632 = n1400 | n18070 ;
  assign n24633 = n24632 ^ n8853 ^ 1'b0 ;
  assign n24634 = ( n4435 & n15723 ) | ( n4435 & ~n24633 ) | ( n15723 & ~n24633 ) ;
  assign n24635 = n6555 ^ n4885 ^ n1690 ;
  assign n24636 = ( n1691 & n24634 ) | ( n1691 & ~n24635 ) | ( n24634 & ~n24635 ) ;
  assign n24637 = n11614 | n17000 ;
  assign n24638 = n24637 ^ n7175 ^ 1'b0 ;
  assign n24639 = ( n8133 & n18670 ) | ( n8133 & n24638 ) | ( n18670 & n24638 ) ;
  assign n24640 = ( n10047 & n12710 ) | ( n10047 & n16698 ) | ( n12710 & n16698 ) ;
  assign n24641 = n9443 ^ n5017 ^ 1'b0 ;
  assign n24642 = ~n7110 & n24641 ;
  assign n24643 = n24642 ^ n3351 ^ n3118 ;
  assign n24644 = n24643 ^ n3037 ^ 1'b0 ;
  assign n24645 = ( n18500 & n24640 ) | ( n18500 & n24644 ) | ( n24640 & n24644 ) ;
  assign n24646 = n8255 ^ n7053 ^ n5340 ;
  assign n24647 = ( n260 & ~n7249 ) | ( n260 & n21504 ) | ( ~n7249 & n21504 ) ;
  assign n24648 = ( n4169 & n24646 ) | ( n4169 & n24647 ) | ( n24646 & n24647 ) ;
  assign n24649 = n14952 ^ n13213 ^ 1'b0 ;
  assign n24650 = ~n1451 & n24649 ;
  assign n24651 = n1426 | n20116 ;
  assign n24652 = n23551 ^ n12932 ^ 1'b0 ;
  assign n24653 = ~n13448 & n24652 ;
  assign n24654 = n10989 | n16214 ;
  assign n24655 = n24654 ^ n6932 ^ n732 ;
  assign n24656 = n24655 ^ n5079 ^ 1'b0 ;
  assign n24657 = n6731 ^ n4594 ^ 1'b0 ;
  assign n24658 = n13774 ^ n5827 ^ n1176 ;
  assign n24661 = ( ~n2344 & n11462 ) | ( ~n2344 & n12500 ) | ( n11462 & n12500 ) ;
  assign n24660 = ( n1732 & n2833 ) | ( n1732 & n8087 ) | ( n2833 & n8087 ) ;
  assign n24659 = n1973 & ~n10643 ;
  assign n24662 = n24661 ^ n24660 ^ n24659 ;
  assign n24663 = ( ~n5398 & n9581 ) | ( ~n5398 & n24662 ) | ( n9581 & n24662 ) ;
  assign n24664 = n23634 ^ n2344 ^ 1'b0 ;
  assign n24665 = n22634 ^ n14755 ^ 1'b0 ;
  assign n24666 = n3896 | n22274 ;
  assign n24667 = ( n495 & n9670 ) | ( n495 & ~n19425 ) | ( n9670 & ~n19425 ) ;
  assign n24668 = n6223 ^ n4686 ^ 1'b0 ;
  assign n24669 = n8676 | n24668 ;
  assign n24670 = n7314 | n24669 ;
  assign n24671 = n11691 ^ n8391 ^ n791 ;
  assign n24672 = n24671 ^ n7284 ^ n6485 ;
  assign n24673 = n432 & ~n3988 ;
  assign n24674 = n13865 | n24673 ;
  assign n24675 = n22167 ^ n13888 ^ n4322 ;
  assign n24676 = n18071 & ~n24675 ;
  assign n24677 = ~n4510 & n24676 ;
  assign n24680 = ( ~n505 & n829 ) | ( ~n505 & n4618 ) | ( n829 & n4618 ) ;
  assign n24678 = ~n6919 & n9269 ;
  assign n24679 = n24678 ^ n1004 ^ 1'b0 ;
  assign n24681 = n24680 ^ n24679 ^ n10197 ;
  assign n24682 = n10238 | n24681 ;
  assign n24683 = n16183 | n24682 ;
  assign n24685 = ~n5127 & n15191 ;
  assign n24686 = n24685 ^ n19175 ^ 1'b0 ;
  assign n24684 = ~n7404 & n23588 ;
  assign n24687 = n24686 ^ n24684 ^ 1'b0 ;
  assign n24688 = ( ~n1100 & n3599 ) | ( ~n1100 & n6797 ) | ( n3599 & n6797 ) ;
  assign n24689 = n5331 & ~n24688 ;
  assign n24690 = n24689 ^ n5171 ^ 1'b0 ;
  assign n24691 = ( ~n16931 & n17135 ) | ( ~n16931 & n24690 ) | ( n17135 & n24690 ) ;
  assign n24692 = n21161 ^ n11859 ^ 1'b0 ;
  assign n24693 = n2868 & n15580 ;
  assign n24694 = n23870 ^ n20797 ^ 1'b0 ;
  assign n24695 = ( n19879 & n22144 ) | ( n19879 & ~n24694 ) | ( n22144 & ~n24694 ) ;
  assign n24696 = ~n8350 & n10359 ;
  assign n24697 = n24696 ^ n9803 ^ n4457 ;
  assign n24698 = n20004 ^ n773 ^ 1'b0 ;
  assign n24699 = n8259 ^ n1666 ^ 1'b0 ;
  assign n24700 = n24699 ^ n20244 ^ n14354 ;
  assign n24701 = n12603 & n24700 ;
  assign n24702 = n24701 ^ n12372 ^ 1'b0 ;
  assign n24703 = ~n3701 & n15056 ;
  assign n24704 = n17290 & ~n23037 ;
  assign n24705 = n24704 ^ n22239 ^ 1'b0 ;
  assign n24706 = n23504 ^ n7830 ^ 1'b0 ;
  assign n24707 = n3179 | n9069 ;
  assign n24708 = n24707 ^ n15846 ^ 1'b0 ;
  assign n24709 = n24708 ^ n9611 ^ n1789 ;
  assign n24710 = ( n17745 & ~n19430 ) | ( n17745 & n23275 ) | ( ~n19430 & n23275 ) ;
  assign n24711 = ~n325 & n7734 ;
  assign n24712 = n24711 ^ n18644 ^ 1'b0 ;
  assign n24713 = n24712 ^ n3330 ^ 1'b0 ;
  assign n24714 = n12285 ^ n3355 ^ 1'b0 ;
  assign n24715 = n24714 ^ n23152 ^ 1'b0 ;
  assign n24716 = n19435 & n24715 ;
  assign n24717 = n3008 & n18380 ;
  assign n24718 = ~n24716 & n24717 ;
  assign n24719 = n5403 & ~n23258 ;
  assign n24720 = n4615 & ~n6497 ;
  assign n24721 = n15878 & n24720 ;
  assign n24722 = n24721 ^ n8243 ^ 1'b0 ;
  assign n24723 = n10162 ^ n851 ^ 1'b0 ;
  assign n24724 = n4579 & n24723 ;
  assign n24725 = n24724 ^ n1938 ^ 1'b0 ;
  assign n24726 = n265 | n24725 ;
  assign n24727 = n24726 ^ n3232 ^ n1964 ;
  assign n24728 = ( n11931 & n24722 ) | ( n11931 & n24727 ) | ( n24722 & n24727 ) ;
  assign n24729 = n985 | n20045 ;
  assign n24730 = n24729 ^ n10785 ^ n2550 ;
  assign n24731 = n23484 ^ n2342 ^ n347 ;
  assign n24732 = n24731 ^ n5442 ^ 1'b0 ;
  assign n24733 = n12257 & n24732 ;
  assign n24734 = ~n2793 & n20342 ;
  assign n24735 = n24734 ^ n4445 ^ 1'b0 ;
  assign n24736 = n5922 & n11342 ;
  assign n24737 = n17109 ^ n6624 ^ 1'b0 ;
  assign n24738 = ( n14088 & n22137 ) | ( n14088 & n24737 ) | ( n22137 & n24737 ) ;
  assign n24739 = n15826 ^ n7698 ^ n2665 ;
  assign n24740 = n24739 ^ n9246 ^ 1'b0 ;
  assign n24741 = n23238 ^ n18712 ^ 1'b0 ;
  assign n24742 = n14685 & ~n22326 ;
  assign n24743 = n14171 & n24742 ;
  assign n24744 = n24743 ^ n9691 ^ 1'b0 ;
  assign n24745 = ( n8949 & ~n10105 ) | ( n8949 & n16287 ) | ( ~n10105 & n16287 ) ;
  assign n24746 = n4465 & n24745 ;
  assign n24747 = ( n980 & ~n8412 ) | ( n980 & n16158 ) | ( ~n8412 & n16158 ) ;
  assign n24748 = n24747 ^ n7555 ^ 1'b0 ;
  assign n24749 = n2657 ^ n182 ^ 1'b0 ;
  assign n24750 = n8243 | n24749 ;
  assign n24751 = n24750 ^ n3643 ^ n2413 ;
  assign n24752 = n24751 ^ n16638 ^ 1'b0 ;
  assign n24753 = n18640 & n24752 ;
  assign n24754 = n6901 ^ n3148 ^ 1'b0 ;
  assign n24755 = ~n1007 & n24754 ;
  assign n24756 = n22537 ^ n14521 ^ 1'b0 ;
  assign n24757 = n16983 & n24756 ;
  assign n24758 = ( n9198 & n24755 ) | ( n9198 & ~n24757 ) | ( n24755 & ~n24757 ) ;
  assign n24759 = n15574 ^ n4509 ^ n3007 ;
  assign n24760 = ( ~n1379 & n23223 ) | ( ~n1379 & n24759 ) | ( n23223 & n24759 ) ;
  assign n24761 = ~n10995 & n15194 ;
  assign n24762 = n1800 & n22216 ;
  assign n24763 = ~n15239 & n24762 ;
  assign n24764 = n24763 ^ n9855 ^ 1'b0 ;
  assign n24765 = ( n5697 & n24761 ) | ( n5697 & ~n24764 ) | ( n24761 & ~n24764 ) ;
  assign n24766 = n13788 ^ n6546 ^ 1'b0 ;
  assign n24767 = n134 | n24586 ;
  assign n24768 = n24767 ^ n12301 ^ 1'b0 ;
  assign n24769 = n6891 & ~n11967 ;
  assign n24770 = ( n10357 & n16840 ) | ( n10357 & n24769 ) | ( n16840 & n24769 ) ;
  assign n24771 = ( n1628 & n2082 ) | ( n1628 & n8265 ) | ( n2082 & n8265 ) ;
  assign n24772 = ( n13713 & n20352 ) | ( n13713 & n23729 ) | ( n20352 & n23729 ) ;
  assign n24773 = n10581 ^ n8891 ^ n6456 ;
  assign n24774 = n7729 & ~n9581 ;
  assign n24775 = n24774 ^ n15604 ^ 1'b0 ;
  assign n24776 = ~n14902 & n24775 ;
  assign n24777 = n23967 ^ n18073 ^ 1'b0 ;
  assign n24778 = n19848 & n24777 ;
  assign n24779 = n22170 ^ n9439 ^ 1'b0 ;
  assign n24780 = n7900 ^ n3542 ^ 1'b0 ;
  assign n24781 = ~n5154 & n24780 ;
  assign n24782 = n18496 & n24781 ;
  assign n24783 = n19507 ^ n7622 ^ 1'b0 ;
  assign n24784 = n5810 | n24783 ;
  assign n24786 = x127 & ~n8621 ;
  assign n24787 = n1910 & n24786 ;
  assign n24785 = n11022 & ~n17730 ;
  assign n24788 = n24787 ^ n24785 ^ 1'b0 ;
  assign n24789 = n15330 ^ n1481 ^ 1'b0 ;
  assign n24790 = n6159 & n16062 ;
  assign n24791 = ~n24789 & n24790 ;
  assign n24792 = n3799 | n4726 ;
  assign n24793 = n9368 & ~n24792 ;
  assign n24794 = n24793 ^ n24696 ^ n19702 ;
  assign n24795 = n22449 ^ n17197 ^ n14313 ;
  assign n24796 = n13567 ^ n12730 ^ 1'b0 ;
  assign n24797 = n8606 & n24796 ;
  assign n24798 = ( ~n5730 & n11570 ) | ( ~n5730 & n24797 ) | ( n11570 & n24797 ) ;
  assign n24799 = n16099 ^ n12867 ^ 1'b0 ;
  assign n24800 = n2871 & ~n24799 ;
  assign n24801 = n14089 ^ n9548 ^ 1'b0 ;
  assign n24802 = n1346 & ~n24801 ;
  assign n24803 = n1291 & n5652 ;
  assign n24804 = n7714 & ~n24803 ;
  assign n24805 = n24804 ^ n2301 ^ 1'b0 ;
  assign n24806 = ~n11513 & n16684 ;
  assign n24807 = ( n1040 & ~n4286 ) | ( n1040 & n14905 ) | ( ~n4286 & n14905 ) ;
  assign n24808 = n10141 & n10816 ;
  assign n24809 = n21179 & n24808 ;
  assign n24810 = n24809 ^ n8309 ^ 1'b0 ;
  assign n24811 = ~n12323 & n24810 ;
  assign n24812 = n24807 & ~n24811 ;
  assign n24814 = ~n1611 & n3896 ;
  assign n24813 = n19823 ^ n6333 ^ 1'b0 ;
  assign n24815 = n24814 ^ n24813 ^ n5120 ;
  assign n24817 = n7940 ^ n6196 ^ n1986 ;
  assign n24818 = n24817 ^ n23718 ^ n9598 ;
  assign n24816 = ~n2822 & n18662 ;
  assign n24819 = n24818 ^ n24816 ^ 1'b0 ;
  assign n24820 = n24819 ^ n3548 ^ 1'b0 ;
  assign n24821 = n8193 | n24820 ;
  assign n24822 = n15176 ^ n1306 ^ 1'b0 ;
  assign n24823 = n24822 ^ n11211 ^ n5473 ;
  assign n24824 = ~n5935 & n7534 ;
  assign n24825 = n24823 & n24824 ;
  assign n24826 = ~n4014 & n20981 ;
  assign n24827 = ( n1455 & ~n9984 ) | ( n1455 & n24826 ) | ( ~n9984 & n24826 ) ;
  assign n24828 = n20667 ^ n13938 ^ 1'b0 ;
  assign n24829 = n24828 ^ n20350 ^ n17906 ;
  assign n24830 = n17944 ^ n5876 ^ 1'b0 ;
  assign n24831 = n24830 ^ n12336 ^ n8452 ;
  assign n24832 = n17108 ^ n13288 ^ 1'b0 ;
  assign n24833 = n10084 & n14648 ;
  assign n24834 = n9466 & n10285 ;
  assign n24835 = n8116 & n22148 ;
  assign n24836 = ~n22287 & n24835 ;
  assign n24837 = n21580 & ~n24229 ;
  assign n24838 = n24837 ^ n14141 ^ 1'b0 ;
  assign n24839 = ~n214 & n16637 ;
  assign n24842 = n1820 | n3499 ;
  assign n24843 = n6856 | n24842 ;
  assign n24840 = ~n10750 & n20268 ;
  assign n24841 = n24840 ^ n14578 ^ 1'b0 ;
  assign n24844 = n24843 ^ n24841 ^ n20912 ;
  assign n24845 = ( n20066 & n24839 ) | ( n20066 & n24844 ) | ( n24839 & n24844 ) ;
  assign n24846 = n18779 ^ n13181 ^ n12881 ;
  assign n24847 = n19939 ^ n13873 ^ 1'b0 ;
  assign n24848 = n8528 & ~n24847 ;
  assign n24849 = ( ~n15118 & n16973 ) | ( ~n15118 & n24848 ) | ( n16973 & n24848 ) ;
  assign n24850 = ( n1501 & ~n2114 ) | ( n1501 & n5853 ) | ( ~n2114 & n5853 ) ;
  assign n24851 = ~n5440 & n24850 ;
  assign n24853 = n6358 ^ n2023 ^ 1'b0 ;
  assign n24852 = n11537 | n18771 ;
  assign n24854 = n24853 ^ n24852 ^ 1'b0 ;
  assign n24855 = n22141 ^ n4908 ^ 1'b0 ;
  assign n24856 = n9620 ^ x9 ^ 1'b0 ;
  assign n24857 = n1185 & ~n2424 ;
  assign n24858 = n23792 & n23872 ;
  assign n24859 = n18244 ^ n3238 ^ 1'b0 ;
  assign n24860 = n18527 & ~n24859 ;
  assign n24861 = ( ~n4150 & n10922 ) | ( ~n4150 & n11253 ) | ( n10922 & n11253 ) ;
  assign n24862 = n6975 ^ n6751 ^ n6300 ;
  assign n24863 = n2543 & ~n4623 ;
  assign n24864 = n24863 ^ n5159 ^ n4986 ;
  assign n24865 = n24864 ^ n21481 ^ 1'b0 ;
  assign n24866 = n24865 ^ n14887 ^ n6135 ;
  assign n24867 = ( n24861 & n24862 ) | ( n24861 & ~n24866 ) | ( n24862 & ~n24866 ) ;
  assign n24868 = n16051 ^ n11964 ^ n5390 ;
  assign n24869 = n5535 & ~n12576 ;
  assign n24870 = n24869 ^ n16776 ^ 1'b0 ;
  assign n24871 = n24868 & ~n24870 ;
  assign n24872 = ( n7704 & ~n20855 ) | ( n7704 & n24871 ) | ( ~n20855 & n24871 ) ;
  assign n24873 = n2426 & n7239 ;
  assign n24874 = n20663 & ~n24873 ;
  assign n24875 = n24874 ^ n15632 ^ 1'b0 ;
  assign n24876 = n8005 ^ n2240 ^ 1'b0 ;
  assign n24877 = n370 & n24876 ;
  assign n24878 = n11082 & ~n11948 ;
  assign n24879 = n14019 ^ n1484 ^ 1'b0 ;
  assign n24880 = n9445 & n24879 ;
  assign n24881 = n6591 ^ n539 ^ 1'b0 ;
  assign n24882 = ( n5627 & n8869 ) | ( n5627 & ~n24881 ) | ( n8869 & ~n24881 ) ;
  assign n24883 = n17912 ^ n3108 ^ n2145 ;
  assign n24884 = n23754 ^ n11785 ^ 1'b0 ;
  assign n24885 = n19653 ^ n9919 ^ n5570 ;
  assign n24886 = n24884 & ~n24885 ;
  assign n24891 = n439 | n1219 ;
  assign n24892 = n24891 ^ n5365 ^ 1'b0 ;
  assign n24893 = ( n1646 & n3900 ) | ( n1646 & n24892 ) | ( n3900 & n24892 ) ;
  assign n24894 = n24893 ^ n9425 ^ n6023 ;
  assign n24887 = ~n11660 & n13017 ;
  assign n24888 = n24887 ^ n11368 ^ n8908 ;
  assign n24889 = ( n10057 & ~n15673 ) | ( n10057 & n24888 ) | ( ~n15673 & n24888 ) ;
  assign n24890 = n4544 & ~n24889 ;
  assign n24895 = n24894 ^ n24890 ^ 1'b0 ;
  assign n24896 = n6169 | n8436 ;
  assign n24898 = n6420 & n18222 ;
  assign n24897 = n3325 & n10831 ;
  assign n24899 = n24898 ^ n24897 ^ n10300 ;
  assign n24900 = n15986 ^ n9483 ^ n1801 ;
  assign n24901 = ( ~n4488 & n18476 ) | ( ~n4488 & n24694 ) | ( n18476 & n24694 ) ;
  assign n24902 = n9699 ^ n7077 ^ 1'b0 ;
  assign n24903 = n2964 | n24902 ;
  assign n24904 = ( ~n1240 & n19638 ) | ( ~n1240 & n24903 ) | ( n19638 & n24903 ) ;
  assign n24905 = n16693 ^ n7477 ^ n4344 ;
  assign n24906 = n24905 ^ n5273 ^ 1'b0 ;
  assign n24907 = n10203 | n17131 ;
  assign n24908 = n24907 ^ n18307 ^ 1'b0 ;
  assign n24909 = n16199 ^ n14030 ^ 1'b0 ;
  assign n24910 = n4952 | n24909 ;
  assign n24911 = n24144 & ~n24910 ;
  assign n24912 = n24911 ^ n2179 ^ 1'b0 ;
  assign n24913 = n1019 & ~n12942 ;
  assign n24914 = n24913 ^ n3258 ^ 1'b0 ;
  assign n24915 = n13805 ^ n1820 ^ 1'b0 ;
  assign n24916 = n24914 & n24915 ;
  assign n24917 = n9180 ^ n4329 ^ 1'b0 ;
  assign n24918 = n13231 ^ n4297 ^ 1'b0 ;
  assign n24919 = n19008 | n24918 ;
  assign n24920 = n24047 ^ n19691 ^ n1198 ;
  assign n24921 = ( n2420 & ~n6146 ) | ( n2420 & n19476 ) | ( ~n6146 & n19476 ) ;
  assign n24922 = ( ~n2059 & n4424 ) | ( ~n2059 & n4804 ) | ( n4424 & n4804 ) ;
  assign n24923 = n24922 ^ n1819 ^ 1'b0 ;
  assign n24924 = ( n6559 & ~n23280 ) | ( n6559 & n24923 ) | ( ~n23280 & n24923 ) ;
  assign n24926 = n6500 & ~n14633 ;
  assign n24927 = n24926 ^ n16042 ^ 1'b0 ;
  assign n24925 = n1266 ^ n186 ^ 1'b0 ;
  assign n24928 = n24927 ^ n24925 ^ n7536 ;
  assign n24929 = n2911 | n5137 ;
  assign n24930 = ~n15216 & n24929 ;
  assign n24931 = n21691 ^ n15947 ^ n5835 ;
  assign n24932 = n6144 & ~n24931 ;
  assign n24933 = ~n24930 & n24932 ;
  assign n24934 = n6451 & ~n10825 ;
  assign n24935 = n15650 & ~n16932 ;
  assign n24936 = n24935 ^ n20484 ^ 1'b0 ;
  assign n24937 = ( n3742 & n3777 ) | ( n3742 & ~n14422 ) | ( n3777 & ~n14422 ) ;
  assign n24938 = n7798 | n24937 ;
  assign n24939 = ~n1553 & n8289 ;
  assign n24940 = n18187 ^ n4042 ^ n1462 ;
  assign n24941 = n4943 & ~n7205 ;
  assign n24942 = n2869 & n24941 ;
  assign n24943 = n24942 ^ n2836 ^ 1'b0 ;
  assign n24944 = n11268 ^ n774 ^ 1'b0 ;
  assign n24945 = n2165 & n24944 ;
  assign n24946 = n1591 & ~n24566 ;
  assign n24947 = n24946 ^ n20354 ^ 1'b0 ;
  assign n24948 = n6894 & ~n24947 ;
  assign n24949 = n24948 ^ n10600 ^ 1'b0 ;
  assign n24950 = n1032 & ~n1388 ;
  assign n24951 = ~n3195 & n8379 ;
  assign n24952 = n11868 ^ n2559 ^ 1'b0 ;
  assign n24953 = ( n8394 & n13168 ) | ( n8394 & ~n24952 ) | ( n13168 & ~n24952 ) ;
  assign n24954 = n5064 & n8899 ;
  assign n24958 = n11010 ^ x32 ^ 1'b0 ;
  assign n24957 = n4039 & ~n7931 ;
  assign n24959 = n24958 ^ n24957 ^ 1'b0 ;
  assign n24955 = ( n5900 & ~n14368 ) | ( n5900 & n17586 ) | ( ~n14368 & n17586 ) ;
  assign n24956 = n24955 ^ n20714 ^ n12855 ;
  assign n24960 = n24959 ^ n24956 ^ n1022 ;
  assign n24961 = n22817 ^ n14482 ^ 1'b0 ;
  assign n24962 = n8591 | n18549 ;
  assign n24963 = n18597 ^ n13234 ^ 1'b0 ;
  assign n24964 = n16342 & n24963 ;
  assign n24968 = n13207 ^ n4081 ^ 1'b0 ;
  assign n24969 = ( ~n2606 & n4783 ) | ( ~n2606 & n24968 ) | ( n4783 & n24968 ) ;
  assign n24965 = n7947 & n22199 ;
  assign n24966 = ~n501 & n24965 ;
  assign n24967 = n1128 | n24966 ;
  assign n24970 = n24969 ^ n24967 ^ 1'b0 ;
  assign n24971 = n18375 ^ n18139 ^ n12339 ;
  assign n24972 = n24971 ^ n23137 ^ n17967 ;
  assign n24973 = ~n6143 & n6625 ;
  assign n24974 = n24973 ^ n23144 ^ n19032 ;
  assign n24975 = n2969 | n10182 ;
  assign n24976 = n3340 | n4588 ;
  assign n24977 = n994 & ~n24976 ;
  assign n24978 = n3153 & ~n11234 ;
  assign n24979 = ~n9685 & n24973 ;
  assign n24980 = n8394 & n24979 ;
  assign n24981 = n4092 & ~n24980 ;
  assign n24982 = n24978 & n24981 ;
  assign n24983 = n4719 & n19666 ;
  assign n24984 = n24983 ^ n5336 ^ 1'b0 ;
  assign n24985 = ( n2224 & n3144 ) | ( n2224 & ~n20267 ) | ( n3144 & ~n20267 ) ;
  assign n24986 = n6515 & ~n18549 ;
  assign n24987 = ~n24985 & n24986 ;
  assign n24988 = n3097 & n13562 ;
  assign n24989 = n24988 ^ n14474 ^ 1'b0 ;
  assign n24990 = n19131 | n24989 ;
  assign n24991 = ( n2242 & n19532 ) | ( n2242 & ~n24990 ) | ( n19532 & ~n24990 ) ;
  assign n24992 = ( n10103 & ~n13661 ) | ( n10103 & n17438 ) | ( ~n13661 & n17438 ) ;
  assign n24993 = n2212 & n17987 ;
  assign n24994 = n24993 ^ n6113 ^ 1'b0 ;
  assign n24995 = ( n752 & n5186 ) | ( n752 & n24994 ) | ( n5186 & n24994 ) ;
  assign n24996 = n306 & n16340 ;
  assign n24997 = n3684 & n24996 ;
  assign n24998 = n13933 ^ n13493 ^ 1'b0 ;
  assign n24999 = ~n6703 & n8757 ;
  assign n25000 = n24998 & n24999 ;
  assign n25001 = n7478 ^ n4503 ^ 1'b0 ;
  assign n25002 = n2671 & ~n25001 ;
  assign n25003 = n10209 | n25002 ;
  assign n25004 = n6417 | n8827 ;
  assign n25005 = n25004 ^ n20601 ^ 1'b0 ;
  assign n25009 = n4772 & ~n8475 ;
  assign n25010 = n25009 ^ n23280 ^ n7248 ;
  assign n25006 = n9283 | n22862 ;
  assign n25007 = n470 | n25006 ;
  assign n25008 = n25007 ^ n6706 ^ 1'b0 ;
  assign n25011 = n25010 ^ n25008 ^ n20470 ;
  assign n25012 = ( n4712 & n12938 ) | ( n4712 & n25011 ) | ( n12938 & n25011 ) ;
  assign n25013 = n16387 ^ n13368 ^ n3943 ;
  assign n25014 = n21609 ^ n18941 ^ 1'b0 ;
  assign n25015 = n4093 & ~n17380 ;
  assign n25016 = n3926 & n5630 ;
  assign n25017 = n25016 ^ n3436 ^ 1'b0 ;
  assign n25018 = n25017 ^ n9848 ^ n4859 ;
  assign n25019 = n3234 | n21251 ;
  assign n25020 = n25018 & ~n25019 ;
  assign n25021 = n5214 | n7684 ;
  assign n25022 = n23761 & ~n25021 ;
  assign n25023 = n25022 ^ n1105 ^ 1'b0 ;
  assign n25024 = n4907 ^ n3790 ^ x7 ;
  assign n25025 = n13264 | n25024 ;
  assign n25026 = n25025 ^ n2090 ^ 1'b0 ;
  assign n25027 = ~n25023 & n25026 ;
  assign n25028 = n6068 & ~n22072 ;
  assign n25029 = ( n12820 & n25027 ) | ( n12820 & n25028 ) | ( n25027 & n25028 ) ;
  assign n25030 = ~n1258 & n15840 ;
  assign n25031 = n25030 ^ n14577 ^ 1'b0 ;
  assign n25032 = ( ~n6823 & n22976 ) | ( ~n6823 & n25031 ) | ( n22976 & n25031 ) ;
  assign n25033 = n23405 ^ n18022 ^ 1'b0 ;
  assign n25034 = ~n5266 & n8964 ;
  assign n25036 = n8505 ^ n204 ^ 1'b0 ;
  assign n25035 = n357 | n12593 ;
  assign n25037 = n25036 ^ n25035 ^ 1'b0 ;
  assign n25038 = n18786 ^ n14756 ^ n1198 ;
  assign n25040 = n8541 | n18475 ;
  assign n25041 = n25040 ^ n13061 ^ 1'b0 ;
  assign n25039 = n6370 ^ n5234 ^ 1'b0 ;
  assign n25042 = n25041 ^ n25039 ^ 1'b0 ;
  assign n25043 = ( n2494 & n5751 ) | ( n2494 & ~n7560 ) | ( n5751 & ~n7560 ) ;
  assign n25044 = n24533 & ~n25043 ;
  assign n25047 = n11921 ^ n3688 ^ 1'b0 ;
  assign n25045 = n2053 & ~n4550 ;
  assign n25046 = ~n906 & n25045 ;
  assign n25048 = n25047 ^ n25046 ^ n555 ;
  assign n25049 = ~n19842 & n25048 ;
  assign n25050 = n7700 & n16173 ;
  assign n25051 = ~n11620 & n25050 ;
  assign n25054 = n10764 ^ n6206 ^ n4733 ;
  assign n25052 = n11108 & ~n21367 ;
  assign n25053 = n25052 ^ n8946 ^ 1'b0 ;
  assign n25055 = n25054 ^ n25053 ^ n2491 ;
  assign n25056 = n14026 & ~n25055 ;
  assign n25057 = ( n2222 & n3101 ) | ( n2222 & ~n8116 ) | ( n3101 & ~n8116 ) ;
  assign n25058 = n25057 ^ n16004 ^ 1'b0 ;
  assign n25059 = n11202 & ~n24170 ;
  assign n25060 = n25059 ^ n6092 ^ 1'b0 ;
  assign n25064 = n2116 | n2246 ;
  assign n25061 = n24539 ^ n6775 ^ x108 ;
  assign n25062 = ~n9245 & n13410 ;
  assign n25063 = ~n25061 & n25062 ;
  assign n25065 = n25064 ^ n25063 ^ n11314 ;
  assign n25066 = n1864 | n4946 ;
  assign n25067 = n25066 ^ n6469 ^ 1'b0 ;
  assign n25069 = n594 & ~n2316 ;
  assign n25070 = n25069 ^ n18381 ^ 1'b0 ;
  assign n25068 = n22406 ^ n5863 ^ n583 ;
  assign n25071 = n25070 ^ n25068 ^ n747 ;
  assign n25072 = n25067 | n25071 ;
  assign n25073 = n6522 | n13804 ;
  assign n25074 = n808 | n25073 ;
  assign n25075 = n24294 & ~n25074 ;
  assign n25076 = ( ~n783 & n1625 ) | ( ~n783 & n5259 ) | ( n1625 & n5259 ) ;
  assign n25077 = n7240 ^ n4305 ^ 1'b0 ;
  assign n25078 = n25076 & ~n25077 ;
  assign n25079 = ( n15893 & n22564 ) | ( n15893 & n25078 ) | ( n22564 & n25078 ) ;
  assign n25080 = n5006 | n18438 ;
  assign n25081 = n25080 ^ n8162 ^ 1'b0 ;
  assign n25082 = n9565 & ~n25081 ;
  assign n25083 = n5521 & ~n9298 ;
  assign n25086 = n13185 ^ n7141 ^ n6175 ;
  assign n25084 = n15739 ^ n7957 ^ 1'b0 ;
  assign n25085 = ~n15023 & n25084 ;
  assign n25087 = n25086 ^ n25085 ^ 1'b0 ;
  assign n25088 = n25087 ^ n21568 ^ 1'b0 ;
  assign n25090 = n10259 ^ n4114 ^ n3485 ;
  assign n25089 = n2996 | n8297 ;
  assign n25091 = n25090 ^ n25089 ^ 1'b0 ;
  assign n25092 = ~n19020 & n25091 ;
  assign n25093 = n8619 ^ n7024 ^ 1'b0 ;
  assign n25094 = n7726 | n25093 ;
  assign n25095 = n19687 ^ n18093 ^ n16135 ;
  assign n25096 = n24681 ^ n24612 ^ n11160 ;
  assign n25097 = n1430 & ~n14083 ;
  assign n25098 = n23434 & n25097 ;
  assign n25099 = n25098 ^ n10803 ^ n498 ;
  assign n25100 = n21930 ^ n20253 ^ n17750 ;
  assign n25101 = n5492 | n18776 ;
  assign n25102 = n25101 ^ n14402 ^ 1'b0 ;
  assign n25103 = n18838 ^ n11814 ^ n5929 ;
  assign n25104 = ( n1287 & n13177 ) | ( n1287 & ~n19430 ) | ( n13177 & ~n19430 ) ;
  assign n25105 = n25104 ^ n8124 ^ 1'b0 ;
  assign n25106 = n25103 & ~n25105 ;
  assign n25107 = ~n2899 & n11253 ;
  assign n25108 = n25107 ^ n20402 ^ 1'b0 ;
  assign n25109 = ~n4285 & n19714 ;
  assign n25110 = n21424 ^ n16840 ^ n7239 ;
  assign n25111 = n1116 & n4917 ;
  assign n25112 = n540 | n23655 ;
  assign n25113 = n6791 & ~n17162 ;
  assign n25114 = n25113 ^ n6256 ^ 1'b0 ;
  assign n25115 = n4948 | n17451 ;
  assign n25116 = n1837 | n25115 ;
  assign n25119 = n4049 | n5919 ;
  assign n25120 = n25119 ^ n17418 ^ 1'b0 ;
  assign n25117 = ( ~n8058 & n10997 ) | ( ~n8058 & n21010 ) | ( n10997 & n21010 ) ;
  assign n25118 = n11102 | n25117 ;
  assign n25121 = n25120 ^ n25118 ^ 1'b0 ;
  assign n25122 = n17277 ^ n11447 ^ 1'b0 ;
  assign n25123 = n13211 & ~n25122 ;
  assign n25124 = ( n10364 & n10773 ) | ( n10364 & ~n25123 ) | ( n10773 & ~n25123 ) ;
  assign n25131 = n6059 ^ n2191 ^ 1'b0 ;
  assign n25132 = n8748 & n25131 ;
  assign n25129 = n8432 ^ n5850 ^ 1'b0 ;
  assign n25125 = n3672 & n8812 ;
  assign n25126 = n5395 & n13674 ;
  assign n25127 = n25125 & n25126 ;
  assign n25128 = ( n6439 & n9728 ) | ( n6439 & n25127 ) | ( n9728 & n25127 ) ;
  assign n25130 = n25129 ^ n25128 ^ n3565 ;
  assign n25133 = n25132 ^ n25130 ^ n1586 ;
  assign n25134 = n10184 & n13299 ;
  assign n25135 = n25134 ^ n18483 ^ n12514 ;
  assign n25136 = n11260 ^ n826 ^ 1'b0 ;
  assign n25137 = n3045 & n6938 ;
  assign n25138 = n25137 ^ n8142 ^ 1'b0 ;
  assign n25139 = n18316 ^ n14011 ^ 1'b0 ;
  assign n25140 = ~n19248 & n25139 ;
  assign n25141 = n16201 ^ n7042 ^ 1'b0 ;
  assign n25142 = n15045 ^ n12290 ^ n6187 ;
  assign n25143 = ~n2204 & n21685 ;
  assign n25144 = n25143 ^ n10318 ^ 1'b0 ;
  assign n25145 = ~n18659 & n25144 ;
  assign n25146 = ~n19471 & n25145 ;
  assign n25147 = ~n5088 & n6881 ;
  assign n25148 = n12921 | n25147 ;
  assign n25149 = n25146 & ~n25148 ;
  assign n25150 = ~n1201 & n1880 ;
  assign n25151 = n25150 ^ n19705 ^ n8046 ;
  assign n25152 = n20718 | n25151 ;
  assign n25153 = x97 & ~n3858 ;
  assign n25154 = n25153 ^ n14868 ^ 1'b0 ;
  assign n25155 = n1404 & ~n5850 ;
  assign n25156 = n7413 & n25155 ;
  assign n25157 = n16394 ^ n13381 ^ 1'b0 ;
  assign n25158 = n767 & ~n8227 ;
  assign n25159 = n12417 | n25158 ;
  assign n25160 = n9866 ^ n2896 ^ 1'b0 ;
  assign n25161 = n15155 & n18537 ;
  assign n25162 = ~n11885 & n25161 ;
  assign n25163 = n6858 ^ n547 ^ 1'b0 ;
  assign n25164 = n6498 & n25163 ;
  assign n25165 = n14799 ^ n8630 ^ 1'b0 ;
  assign n25166 = n25164 & n25165 ;
  assign n25167 = n2453 & n3822 ;
  assign n25168 = n25167 ^ n8215 ^ 1'b0 ;
  assign n25169 = ( n23501 & ~n24376 ) | ( n23501 & n25168 ) | ( ~n24376 & n25168 ) ;
  assign n25170 = n25169 ^ n24507 ^ n9087 ;
  assign n25171 = ~n11217 & n15836 ;
  assign n25172 = n25171 ^ n10481 ^ n7623 ;
  assign n25173 = n8237 ^ n4760 ^ 1'b0 ;
  assign n25174 = n605 & ~n25173 ;
  assign n25175 = n14619 ^ n13566 ^ n2200 ;
  assign n25176 = ~n25174 & n25175 ;
  assign n25177 = n19012 ^ n6493 ^ n1007 ;
  assign n25178 = ( n7365 & n22450 ) | ( n7365 & n25177 ) | ( n22450 & n25177 ) ;
  assign n25179 = n25178 ^ n22512 ^ n11727 ;
  assign n25180 = ~n10590 & n25179 ;
  assign n25181 = n3570 & n8152 ;
  assign n25182 = ( n2629 & n10688 ) | ( n2629 & ~n25181 ) | ( n10688 & ~n25181 ) ;
  assign n25183 = n25182 ^ n23856 ^ n20344 ;
  assign n25184 = ( n8495 & ~n12730 ) | ( n8495 & n25183 ) | ( ~n12730 & n25183 ) ;
  assign n25185 = n15331 & ~n21330 ;
  assign n25186 = n25185 ^ n10716 ^ 1'b0 ;
  assign n25187 = n23504 ^ n21732 ^ n12033 ;
  assign n25188 = n24166 ^ n21744 ^ 1'b0 ;
  assign n25189 = ~n25187 & n25188 ;
  assign n25190 = n8452 & ~n14013 ;
  assign n25191 = ~n985 & n25190 ;
  assign n25192 = n25191 ^ n12183 ^ n3991 ;
  assign n25193 = n12699 ^ n2878 ^ 1'b0 ;
  assign n25194 = n3255 | n25193 ;
  assign n25195 = n25194 ^ n3790 ^ 1'b0 ;
  assign n25196 = ~n25192 & n25195 ;
  assign n25197 = n18616 ^ n5368 ^ 1'b0 ;
  assign n25198 = n9458 ^ n307 ^ 1'b0 ;
  assign n25199 = x37 & ~n25198 ;
  assign n25200 = n25199 ^ n13726 ^ n4386 ;
  assign n25201 = ( n1891 & n14448 ) | ( n1891 & ~n20101 ) | ( n14448 & ~n20101 ) ;
  assign n25202 = n11601 ^ n2762 ^ 1'b0 ;
  assign n25203 = n854 | n8038 ;
  assign n25204 = n16867 ^ n5172 ^ 1'b0 ;
  assign n25205 = ~n4944 & n5255 ;
  assign n25206 = n3955 & n25205 ;
  assign n25207 = n23764 | n25206 ;
  assign n25208 = ( n866 & ~n22359 ) | ( n866 & n23135 ) | ( ~n22359 & n23135 ) ;
  assign n25209 = n11692 ^ n9028 ^ 1'b0 ;
  assign n25210 = n18394 ^ n270 ^ 1'b0 ;
  assign n25211 = ( x22 & n1318 ) | ( x22 & ~n25210 ) | ( n1318 & ~n25210 ) ;
  assign n25216 = n11628 & n20357 ;
  assign n25212 = n1666 & ~n1863 ;
  assign n25213 = n25212 ^ n6446 ^ n432 ;
  assign n25214 = ( ~n6168 & n10158 ) | ( ~n6168 & n25213 ) | ( n10158 & n25213 ) ;
  assign n25215 = ( n3062 & n12291 ) | ( n3062 & ~n25214 ) | ( n12291 & ~n25214 ) ;
  assign n25217 = n25216 ^ n25215 ^ n24700 ;
  assign n25218 = n25217 ^ n22647 ^ n9710 ;
  assign n25219 = ( n699 & n11893 ) | ( n699 & n18063 ) | ( n11893 & n18063 ) ;
  assign n25220 = ( n10796 & n13106 ) | ( n10796 & n25219 ) | ( n13106 & n25219 ) ;
  assign n25221 = n25071 ^ n4100 ^ n2562 ;
  assign n25222 = n20408 ^ n13614 ^ n7898 ;
  assign n25225 = n6243 ^ n5216 ^ n2536 ;
  assign n25223 = n7230 ^ n2127 ^ 1'b0 ;
  assign n25224 = n3824 & ~n25223 ;
  assign n25226 = n25225 ^ n25224 ^ 1'b0 ;
  assign n25227 = ( n5396 & n17481 ) | ( n5396 & ~n25226 ) | ( n17481 & ~n25226 ) ;
  assign n25228 = n25227 ^ n20475 ^ 1'b0 ;
  assign n25229 = n22160 ^ n17516 ^ 1'b0 ;
  assign n25234 = n4278 & n10846 ;
  assign n25235 = n25234 ^ n21476 ^ 1'b0 ;
  assign n25230 = n7204 ^ x96 ^ 1'b0 ;
  assign n25231 = ~n11183 & n25230 ;
  assign n25232 = n25231 ^ n12447 ^ 1'b0 ;
  assign n25233 = n24029 | n25232 ;
  assign n25236 = n25235 ^ n25233 ^ 1'b0 ;
  assign n25237 = n12721 ^ n4283 ^ 1'b0 ;
  assign n25238 = ~n1612 & n5294 ;
  assign n25239 = ( n7926 & n8114 ) | ( n7926 & n25238 ) | ( n8114 & n25238 ) ;
  assign n25240 = n5969 ^ n2259 ^ n328 ;
  assign n25241 = n25240 ^ n1073 ^ 1'b0 ;
  assign n25242 = ( n1954 & n3304 ) | ( n1954 & n6375 ) | ( n3304 & n6375 ) ;
  assign n25243 = n25242 ^ n6450 ^ 1'b0 ;
  assign n25244 = n19674 & n21483 ;
  assign n25245 = n25244 ^ n19753 ^ 1'b0 ;
  assign n25246 = n18438 ^ n8999 ^ 1'b0 ;
  assign n25247 = n9902 & ~n25246 ;
  assign n25248 = ~n12130 & n23068 ;
  assign n25249 = n9630 & n25248 ;
  assign n25250 = n25249 ^ n21900 ^ 1'b0 ;
  assign n25251 = ( n4679 & n7384 ) | ( n4679 & ~n14952 ) | ( n7384 & ~n14952 ) ;
  assign n25252 = n20305 | n25251 ;
  assign n25253 = n25252 ^ n11505 ^ 1'b0 ;
  assign n25254 = n25250 | n25253 ;
  assign n25255 = n16156 ^ n4299 ^ n2801 ;
  assign n25256 = n1079 | n3074 ;
  assign n25257 = n25255 & ~n25256 ;
  assign n25258 = n25257 ^ n14801 ^ 1'b0 ;
  assign n25259 = ~n25254 & n25258 ;
  assign n25260 = n9226 | n23716 ;
  assign n25271 = n10025 | n20618 ;
  assign n25272 = n15397 | n25271 ;
  assign n25263 = n14297 ^ n3637 ^ n1348 ;
  assign n25264 = n7586 ^ n6109 ^ 1'b0 ;
  assign n25265 = ( n2646 & n4872 ) | ( n2646 & ~n25264 ) | ( n4872 & ~n25264 ) ;
  assign n25266 = n2487 & ~n25265 ;
  assign n25267 = n25266 ^ n14560 ^ 1'b0 ;
  assign n25268 = n25267 ^ n10856 ^ n9373 ;
  assign n25269 = n2242 & n25268 ;
  assign n25270 = n25263 & n25269 ;
  assign n25261 = ( n11717 & n20267 ) | ( n11717 & n24922 ) | ( n20267 & n24922 ) ;
  assign n25262 = n25261 ^ n3301 ^ n365 ;
  assign n25273 = n25272 ^ n25270 ^ n25262 ;
  assign n25274 = ( n12895 & n18689 ) | ( n12895 & ~n23046 ) | ( n18689 & ~n23046 ) ;
  assign n25278 = n976 | n4283 ;
  assign n25279 = n25278 ^ n2937 ^ 1'b0 ;
  assign n25280 = n6581 & ~n25279 ;
  assign n25275 = n8208 & ~n12713 ;
  assign n25276 = ~n9002 & n25275 ;
  assign n25277 = ~n4129 & n25276 ;
  assign n25281 = n25280 ^ n25277 ^ 1'b0 ;
  assign n25285 = n5415 ^ n5021 ^ 1'b0 ;
  assign n25286 = n5878 | n25285 ;
  assign n25287 = n7976 | n25286 ;
  assign n25288 = n25287 ^ n14432 ^ 1'b0 ;
  assign n25289 = n21583 ^ n13550 ^ n7914 ;
  assign n25290 = n25289 ^ n19576 ^ 1'b0 ;
  assign n25291 = n25288 & n25290 ;
  assign n25282 = n7585 & n13624 ;
  assign n25283 = ~n10706 & n25282 ;
  assign n25284 = n11318 & ~n25283 ;
  assign n25292 = n25291 ^ n25284 ^ 1'b0 ;
  assign n25293 = n18483 & ~n24318 ;
  assign n25294 = n11661 ^ n10634 ^ 1'b0 ;
  assign n25295 = n25293 & ~n25294 ;
  assign n25296 = ( n361 & ~n3185 ) | ( n361 & n8514 ) | ( ~n3185 & n8514 ) ;
  assign n25297 = n3943 & ~n12770 ;
  assign n25298 = n25296 & n25297 ;
  assign n25299 = n12713 ^ n9887 ^ 1'b0 ;
  assign n25300 = n21170 & n25299 ;
  assign n25301 = n25300 ^ n18056 ^ n2801 ;
  assign n25302 = n3756 ^ n848 ^ n636 ;
  assign n25303 = n22285 ^ n13888 ^ 1'b0 ;
  assign n25304 = n25303 ^ n18888 ^ n6803 ;
  assign n25305 = ( n14391 & n20152 ) | ( n14391 & ~n25304 ) | ( n20152 & ~n25304 ) ;
  assign n25306 = ( n2242 & n4433 ) | ( n2242 & n6604 ) | ( n4433 & n6604 ) ;
  assign n25307 = ( n13088 & n14564 ) | ( n13088 & ~n25306 ) | ( n14564 & ~n25306 ) ;
  assign n25308 = ~n5873 & n10828 ;
  assign n25309 = ~n7539 & n25308 ;
  assign n25310 = ~n1363 & n9565 ;
  assign n25311 = n25309 & n25310 ;
  assign n25312 = ( ~n3844 & n6644 ) | ( ~n3844 & n8645 ) | ( n6644 & n8645 ) ;
  assign n25313 = n15155 & ~n21524 ;
  assign n25314 = n25312 & n25313 ;
  assign n25315 = n12316 ^ n7216 ^ 1'b0 ;
  assign n25316 = n22664 & ~n25315 ;
  assign n25317 = n17911 & n18285 ;
  assign n25318 = n25317 ^ n13455 ^ 1'b0 ;
  assign n25319 = n3118 & n3719 ;
  assign n25320 = n3229 & n25319 ;
  assign n25321 = n25320 ^ n227 ^ 1'b0 ;
  assign n25322 = n8944 ^ n1972 ^ 1'b0 ;
  assign n25323 = ~n15564 & n25322 ;
  assign n25324 = n15986 ^ n12199 ^ n6858 ;
  assign n25325 = n3501 & ~n8653 ;
  assign n25326 = n25325 ^ n10162 ^ 1'b0 ;
  assign n25327 = n9875 & n25326 ;
  assign n25328 = ( n7845 & n13177 ) | ( n7845 & ~n16108 ) | ( n13177 & ~n16108 ) ;
  assign n25329 = ~n18771 & n25328 ;
  assign n25330 = ~n16753 & n25329 ;
  assign n25331 = n9587 & n11462 ;
  assign n25332 = ~n2281 & n4713 ;
  assign n25333 = n25332 ^ n20053 ^ 1'b0 ;
  assign n25334 = n11007 ^ n8297 ^ n3483 ;
  assign n25335 = ( ~n1418 & n5234 ) | ( ~n1418 & n11319 ) | ( n5234 & n11319 ) ;
  assign n25336 = n25335 ^ n18315 ^ 1'b0 ;
  assign n25337 = ~n2869 & n25336 ;
  assign n25338 = n25337 ^ n14742 ^ 1'b0 ;
  assign n25339 = n25338 ^ n6363 ^ 1'b0 ;
  assign n25340 = ( n565 & ~n5059 ) | ( n565 & n25339 ) | ( ~n5059 & n25339 ) ;
  assign n25341 = ( n7649 & ~n13829 ) | ( n7649 & n22999 ) | ( ~n13829 & n22999 ) ;
  assign n25342 = n4015 & ~n19873 ;
  assign n25343 = n13095 | n21176 ;
  assign n25344 = n14009 | n25343 ;
  assign n25345 = n7056 & n25344 ;
  assign n25346 = ~n6656 & n25345 ;
  assign n25347 = n25346 ^ n17886 ^ n11489 ;
  assign n25348 = n8501 & ~n25347 ;
  assign n25349 = n25348 ^ n15736 ^ 1'b0 ;
  assign n25350 = n2676 & ~n7784 ;
  assign n25351 = n25350 ^ n794 ^ 1'b0 ;
  assign n25352 = n21072 ^ n13502 ^ 1'b0 ;
  assign n25353 = ( n2592 & n10449 ) | ( n2592 & n17197 ) | ( n10449 & n17197 ) ;
  assign n25354 = n8651 | n14680 ;
  assign n25355 = ( ~n2649 & n3844 ) | ( ~n2649 & n25354 ) | ( n3844 & n25354 ) ;
  assign n25356 = n10410 ^ n9041 ^ 1'b0 ;
  assign n25357 = n25356 ^ n11222 ^ n2760 ;
  assign n25358 = ( n226 & n13612 ) | ( n226 & n17778 ) | ( n13612 & n17778 ) ;
  assign n25359 = ( n17957 & ~n19931 ) | ( n17957 & n23436 ) | ( ~n19931 & n23436 ) ;
  assign n25360 = ~n7404 & n17073 ;
  assign n25361 = n7261 & n25360 ;
  assign n25363 = n2146 & ~n7419 ;
  assign n25364 = n25363 ^ n23867 ^ 1'b0 ;
  assign n25362 = n2596 & ~n20273 ;
  assign n25365 = n25364 ^ n25362 ^ 1'b0 ;
  assign n25368 = x113 & ~n13522 ;
  assign n25366 = n3056 ^ n598 ^ 1'b0 ;
  assign n25367 = n25366 ^ n14157 ^ n10613 ;
  assign n25369 = n25368 ^ n25367 ^ n15639 ;
  assign n25370 = n7827 ^ n3988 ^ 1'b0 ;
  assign n25371 = ( ~n3598 & n18349 ) | ( ~n3598 & n24903 ) | ( n18349 & n24903 ) ;
  assign n25372 = ( n1759 & n7234 ) | ( n1759 & n11868 ) | ( n7234 & n11868 ) ;
  assign n25373 = n15149 ^ n592 ^ 1'b0 ;
  assign n25374 = n25372 & ~n25373 ;
  assign n25377 = ( ~n10407 & n19187 ) | ( ~n10407 & n23895 ) | ( n19187 & n23895 ) ;
  assign n25375 = n9561 & ~n13405 ;
  assign n25376 = n14629 | n25375 ;
  assign n25378 = n25377 ^ n25376 ^ 1'b0 ;
  assign n25381 = n11522 ^ n11331 ^ 1'b0 ;
  assign n25379 = n4598 ^ n357 ^ 1'b0 ;
  assign n25380 = n7468 & ~n25379 ;
  assign n25382 = n25381 ^ n25380 ^ 1'b0 ;
  assign n25383 = n14176 ^ n11816 ^ n5891 ;
  assign n25384 = n25383 ^ n18901 ^ n942 ;
  assign n25386 = ~n565 & n4415 ;
  assign n25387 = n9158 & n25386 ;
  assign n25388 = ( x40 & n21817 ) | ( x40 & n25387 ) | ( n21817 & n25387 ) ;
  assign n25385 = ~n5173 & n11191 ;
  assign n25389 = n25388 ^ n25385 ^ n20377 ;
  assign n25390 = ( n6144 & n7661 ) | ( n6144 & ~n14041 ) | ( n7661 & ~n14041 ) ;
  assign n25391 = n3672 | n14416 ;
  assign n25392 = n464 | n25391 ;
  assign n25393 = n3946 & ~n25392 ;
  assign n25394 = ( n3791 & n22434 ) | ( n3791 & n25393 ) | ( n22434 & n25393 ) ;
  assign n25395 = ~n2363 & n8529 ;
  assign n25396 = n9645 ^ n2746 ^ 1'b0 ;
  assign n25397 = ~n7781 & n25396 ;
  assign n25398 = ~n10079 & n25397 ;
  assign n25399 = n7807 ^ n4367 ^ 1'b0 ;
  assign n25400 = ~n25398 & n25399 ;
  assign n25401 = ( n533 & ~n3271 ) | ( n533 & n25400 ) | ( ~n3271 & n25400 ) ;
  assign n25402 = n7215 & n25401 ;
  assign n25403 = n25402 ^ n15201 ^ 1'b0 ;
  assign n25404 = n11592 ^ n5169 ^ 1'b0 ;
  assign n25405 = n23524 ^ n5094 ^ 1'b0 ;
  assign n25406 = ~n24593 & n25405 ;
  assign n25407 = n1343 & n5270 ;
  assign n25408 = n2355 | n3074 ;
  assign n25409 = ( ~n7016 & n25407 ) | ( ~n7016 & n25408 ) | ( n25407 & n25408 ) ;
  assign n25410 = ( n4699 & n10440 ) | ( n4699 & ~n16833 ) | ( n10440 & ~n16833 ) ;
  assign n25411 = n15788 ^ n6236 ^ 1'b0 ;
  assign n25412 = n13708 ^ n3959 ^ 1'b0 ;
  assign n25413 = ~n25411 & n25412 ;
  assign n25414 = n5437 | n9106 ;
  assign n25415 = n9566 | n25414 ;
  assign n25416 = ( ~n16557 & n21727 ) | ( ~n16557 & n25415 ) | ( n21727 & n25415 ) ;
  assign n25417 = n18062 ^ n4219 ^ 1'b0 ;
  assign n25418 = n25416 & ~n25417 ;
  assign n25419 = ( n14068 & ~n14904 ) | ( n14068 & n20220 ) | ( ~n14904 & n20220 ) ;
  assign n25420 = n7236 ^ n3403 ^ 1'b0 ;
  assign n25421 = ( ~n4710 & n16989 ) | ( ~n4710 & n25420 ) | ( n16989 & n25420 ) ;
  assign n25422 = n25421 ^ n14069 ^ 1'b0 ;
  assign n25423 = n17598 ^ n5121 ^ 1'b0 ;
  assign n25424 = ( n652 & n15112 ) | ( n652 & n25423 ) | ( n15112 & n25423 ) ;
  assign n25425 = n22903 ^ n9942 ^ 1'b0 ;
  assign n25426 = n8038 | n20629 ;
  assign n25427 = n23648 ^ n3343 ^ n742 ;
  assign n25428 = n25427 ^ n20188 ^ 1'b0 ;
  assign n25429 = n25426 | n25428 ;
  assign n25430 = n17508 ^ n14639 ^ n5428 ;
  assign n25431 = n7591 ^ n7319 ^ 1'b0 ;
  assign n25432 = n23635 & n25431 ;
  assign n25433 = n1811 & ~n10657 ;
  assign n25434 = ~n2701 & n25433 ;
  assign n25435 = n4999 ^ n4302 ^ 1'b0 ;
  assign n25436 = n25435 ^ n15918 ^ 1'b0 ;
  assign n25437 = n20957 ^ n7195 ^ 1'b0 ;
  assign n25438 = n6697 ^ n1813 ^ 1'b0 ;
  assign n25439 = n25438 ^ n19977 ^ n4349 ;
  assign n25440 = n20547 ^ n17941 ^ 1'b0 ;
  assign n25441 = n1129 | n9370 ;
  assign n25442 = n3334 | n11665 ;
  assign n25443 = n25441 | n25442 ;
  assign n25444 = ( ~n3405 & n7622 ) | ( ~n3405 & n23032 ) | ( n7622 & n23032 ) ;
  assign n25445 = ~n6043 & n25444 ;
  assign n25446 = n1809 & n25445 ;
  assign n25447 = n17578 ^ n7067 ^ 1'b0 ;
  assign n25448 = ( n21676 & n23180 ) | ( n21676 & ~n25447 ) | ( n23180 & ~n25447 ) ;
  assign n25449 = ( ~n1306 & n17127 ) | ( ~n1306 & n25448 ) | ( n17127 & n25448 ) ;
  assign n25450 = n9160 ^ n8336 ^ 1'b0 ;
  assign n25451 = n3619 & ~n4594 ;
  assign n25452 = n8592 ^ n5156 ^ 1'b0 ;
  assign n25453 = ( n933 & ~n8058 ) | ( n933 & n25452 ) | ( ~n8058 & n25452 ) ;
  assign n25454 = ( n880 & n5068 ) | ( n880 & ~n25453 ) | ( n5068 & ~n25453 ) ;
  assign n25455 = n7913 & n17989 ;
  assign n25456 = n7521 | n15290 ;
  assign n25457 = n4156 & n25456 ;
  assign n25458 = n5411 ^ n2871 ^ 1'b0 ;
  assign n25459 = n14051 & ~n25458 ;
  assign n25460 = n11140 & ~n12339 ;
  assign n25461 = n5270 & n25460 ;
  assign n25462 = n25461 ^ n11937 ^ n3171 ;
  assign n25463 = n12514 | n19814 ;
  assign n25464 = n25463 ^ n11131 ^ 1'b0 ;
  assign n25465 = ( n19866 & n20283 ) | ( n19866 & ~n25464 ) | ( n20283 & ~n25464 ) ;
  assign n25466 = n6824 | n7931 ;
  assign n25467 = n10454 ^ n2994 ^ n409 ;
  assign n25471 = n7092 ^ n4505 ^ 1'b0 ;
  assign n25472 = n21221 & n25471 ;
  assign n25468 = n3980 | n11451 ;
  assign n25469 = n25468 ^ n13083 ^ 1'b0 ;
  assign n25470 = n1760 | n25469 ;
  assign n25473 = n25472 ^ n25470 ^ 1'b0 ;
  assign n25474 = n16606 ^ n13666 ^ n9620 ;
  assign n25475 = n25473 & ~n25474 ;
  assign n25476 = n5091 ^ n4397 ^ 1'b0 ;
  assign n25477 = n13945 ^ n3619 ^ 1'b0 ;
  assign n25478 = n3777 & n25477 ;
  assign n25479 = n19753 ^ n9941 ^ 1'b0 ;
  assign n25480 = n12966 & ~n25479 ;
  assign n25481 = n18387 ^ n17020 ^ x16 ;
  assign n25482 = ( ~n24887 & n25480 ) | ( ~n24887 & n25481 ) | ( n25480 & n25481 ) ;
  assign n25485 = n5492 ^ n5131 ^ n4446 ;
  assign n25486 = n25485 ^ n9546 ^ 1'b0 ;
  assign n25487 = n3614 | n25486 ;
  assign n25488 = n3015 & ~n8637 ;
  assign n25489 = n25488 ^ n15475 ^ 1'b0 ;
  assign n25490 = n25487 | n25489 ;
  assign n25484 = n13458 ^ n9841 ^ n2285 ;
  assign n25483 = n3111 & ~n18207 ;
  assign n25491 = n25490 ^ n25484 ^ n25483 ;
  assign n25492 = n8591 ^ n7035 ^ 1'b0 ;
  assign n25493 = n12306 ^ n5045 ^ 1'b0 ;
  assign n25494 = n7539 & ~n25493 ;
  assign n25495 = n25494 ^ n22208 ^ 1'b0 ;
  assign n25496 = ( n14915 & n25492 ) | ( n14915 & ~n25495 ) | ( n25492 & ~n25495 ) ;
  assign n25497 = n11270 | n17729 ;
  assign n25498 = ( n4888 & n5154 ) | ( n4888 & ~n7882 ) | ( n5154 & ~n7882 ) ;
  assign n25499 = ( n1656 & ~n6361 ) | ( n1656 & n25498 ) | ( ~n6361 & n25498 ) ;
  assign n25500 = n10114 & ~n16921 ;
  assign n25501 = n25500 ^ n5041 ^ 1'b0 ;
  assign n25504 = ~n11661 & n12792 ;
  assign n25502 = n19594 & ~n21224 ;
  assign n25503 = n23142 | n25502 ;
  assign n25505 = n25504 ^ n25503 ^ 1'b0 ;
  assign n25506 = n12827 | n16519 ;
  assign n25507 = ( ~n13740 & n15757 ) | ( ~n13740 & n19443 ) | ( n15757 & n19443 ) ;
  assign n25508 = ( ~n1277 & n4657 ) | ( ~n1277 & n25507 ) | ( n4657 & n25507 ) ;
  assign n25509 = ( n4451 & n13413 ) | ( n4451 & n17758 ) | ( n13413 & n17758 ) ;
  assign n25510 = n15297 & ~n17200 ;
  assign n25511 = n25510 ^ n806 ^ 1'b0 ;
  assign n25512 = ( n1867 & ~n7028 ) | ( n1867 & n17406 ) | ( ~n7028 & n17406 ) ;
  assign n25513 = n16699 ^ n1601 ^ 1'b0 ;
  assign n25514 = n8360 & n19642 ;
  assign n25515 = n25514 ^ n12563 ^ 1'b0 ;
  assign n25519 = n11019 ^ n4238 ^ 1'b0 ;
  assign n25520 = n25164 & ~n25519 ;
  assign n25521 = ( ~n15523 & n15647 ) | ( ~n15523 & n25520 ) | ( n15647 & n25520 ) ;
  assign n25517 = n7183 & n9675 ;
  assign n25518 = n2074 | n25517 ;
  assign n25516 = n4351 & n7959 ;
  assign n25522 = n25521 ^ n25518 ^ n25516 ;
  assign n25523 = ( n3782 & n8943 ) | ( n3782 & ~n9708 ) | ( n8943 & ~n9708 ) ;
  assign n25524 = n20322 ^ n12431 ^ 1'b0 ;
  assign n25525 = n15735 | n24910 ;
  assign n25526 = n7752 & ~n25525 ;
  assign n25527 = n22769 ^ n2908 ^ 1'b0 ;
  assign n25528 = n24405 | n25527 ;
  assign n25529 = ( n10182 & n25526 ) | ( n10182 & n25528 ) | ( n25526 & n25528 ) ;
  assign n25530 = n6358 & ~n6517 ;
  assign n25531 = n6551 & n25530 ;
  assign n25532 = n20795 ^ n10393 ^ 1'b0 ;
  assign n25533 = n25531 | n25532 ;
  assign n25534 = n786 & ~n2962 ;
  assign n25535 = n12929 & ~n25534 ;
  assign n25536 = n5885 & ~n25535 ;
  assign n25537 = n945 | n24037 ;
  assign n25538 = n25537 ^ n3346 ^ 1'b0 ;
  assign n25539 = n25536 & n25538 ;
  assign n25540 = n1529 | n9362 ;
  assign n25541 = n1899 | n25540 ;
  assign n25542 = n866 & ~n1792 ;
  assign n25543 = n14597 & n25542 ;
  assign n25544 = ( ~n3286 & n17406 ) | ( ~n3286 & n25543 ) | ( n17406 & n25543 ) ;
  assign n25545 = ( n4310 & ~n4624 ) | ( n4310 & n6672 ) | ( ~n4624 & n6672 ) ;
  assign n25546 = n25545 ^ n13802 ^ n2671 ;
  assign n25547 = ( n2652 & n8158 ) | ( n2652 & ~n25546 ) | ( n8158 & ~n25546 ) ;
  assign n25548 = n11082 ^ n3611 ^ 1'b0 ;
  assign n25549 = n18905 ^ n14420 ^ 1'b0 ;
  assign n25550 = n11247 ^ n6013 ^ 1'b0 ;
  assign n25551 = n20054 | n25550 ;
  assign n25552 = ( n474 & ~n20235 ) | ( n474 & n25551 ) | ( ~n20235 & n25551 ) ;
  assign n25553 = ( n14867 & ~n25423 ) | ( n14867 & n25552 ) | ( ~n25423 & n25552 ) ;
  assign n25554 = ~n3035 & n3407 ;
  assign n25555 = n25554 ^ n354 ^ 1'b0 ;
  assign n25556 = n7719 ^ n6572 ^ n1517 ;
  assign n25557 = ( ~n6732 & n9721 ) | ( ~n6732 & n25556 ) | ( n9721 & n25556 ) ;
  assign n25558 = n20059 ^ n18405 ^ n15490 ;
  assign n25559 = ~n25557 & n25558 ;
  assign n25561 = n4545 ^ n1262 ^ n477 ;
  assign n25562 = ( n2296 & ~n6277 ) | ( n2296 & n25561 ) | ( ~n6277 & n25561 ) ;
  assign n25560 = n9472 ^ n5151 ^ n4534 ;
  assign n25563 = n25562 ^ n25560 ^ n7220 ;
  assign n25564 = n1267 | n25563 ;
  assign n25565 = n15151 & ~n25564 ;
  assign n25566 = n5405 & ~n10391 ;
  assign n25567 = n2472 & ~n15036 ;
  assign n25568 = n17918 ^ n15863 ^ n10469 ;
  assign n25569 = n25568 ^ n3050 ^ n1540 ;
  assign n25570 = ( n11213 & n14799 ) | ( n11213 & ~n25526 ) | ( n14799 & ~n25526 ) ;
  assign n25571 = n10318 ^ n8298 ^ n6066 ;
  assign n25572 = n12996 ^ n4964 ^ 1'b0 ;
  assign n25573 = ~n1780 & n4044 ;
  assign n25574 = n1289 & ~n11134 ;
  assign n25575 = ~n25573 & n25574 ;
  assign n25576 = n4546 | n13119 ;
  assign n25577 = n25576 ^ n4970 ^ 1'b0 ;
  assign n25578 = ( n6221 & n13999 ) | ( n6221 & n25577 ) | ( n13999 & n25577 ) ;
  assign n25579 = n21252 & n25578 ;
  assign n25580 = n25579 ^ n9464 ^ 1'b0 ;
  assign n25581 = n7261 ^ n4644 ^ 1'b0 ;
  assign n25582 = n20231 ^ n7809 ^ 1'b0 ;
  assign n25583 = n3209 & ~n9488 ;
  assign n25584 = n25583 ^ n23425 ^ n10193 ;
  assign n25585 = n17298 ^ n2947 ^ 1'b0 ;
  assign n25586 = ~n6059 & n25585 ;
  assign n25587 = n25586 ^ n8056 ^ 1'b0 ;
  assign n25588 = n23211 & ~n25587 ;
  assign n25589 = n10203 ^ n8496 ^ n3393 ;
  assign n25590 = n3677 & n8922 ;
  assign n25591 = ~n25589 & n25590 ;
  assign n25593 = n4167 & n17228 ;
  assign n25592 = n2618 & n24156 ;
  assign n25594 = n25593 ^ n25592 ^ 1'b0 ;
  assign n25597 = n21121 ^ n891 ^ 1'b0 ;
  assign n25598 = n6947 & n25597 ;
  assign n25595 = n13724 | n17860 ;
  assign n25596 = n25595 ^ n8324 ^ 1'b0 ;
  assign n25599 = n25598 ^ n25596 ^ n556 ;
  assign n25600 = n25599 ^ n16839 ^ n1279 ;
  assign n25601 = ( n2038 & n2343 ) | ( n2038 & n9158 ) | ( n2343 & n9158 ) ;
  assign n25609 = n19875 ^ n6183 ^ n2272 ;
  assign n25610 = n11310 & n25609 ;
  assign n25611 = n25610 ^ n1111 ^ 1'b0 ;
  assign n25604 = n3471 & n5390 ;
  assign n25605 = n25604 ^ n1628 ^ 1'b0 ;
  assign n25606 = n2011 & n25605 ;
  assign n25607 = n25606 ^ n15383 ^ n13505 ;
  assign n25608 = n7763 & ~n25607 ;
  assign n25612 = n25611 ^ n25608 ^ n7848 ;
  assign n25602 = n3181 ^ n2199 ^ 1'b0 ;
  assign n25603 = ~n9120 & n25602 ;
  assign n25613 = n25612 ^ n25603 ^ 1'b0 ;
  assign n25614 = n25613 ^ n11531 ^ n5766 ;
  assign n25615 = ~n3030 & n4701 ;
  assign n25616 = n15463 ^ n628 ^ 1'b0 ;
  assign n25617 = n14664 & n25616 ;
  assign n25618 = n4740 & ~n25617 ;
  assign n25619 = ~n19430 & n25618 ;
  assign n25620 = n8606 & ~n16150 ;
  assign n25621 = n9713 & n25620 ;
  assign n25622 = n25621 ^ n5112 ^ 1'b0 ;
  assign n25623 = ~n1149 & n25622 ;
  assign n25625 = n1887 & n5902 ;
  assign n25624 = x66 & ~n19097 ;
  assign n25626 = n25625 ^ n25624 ^ 1'b0 ;
  assign n25627 = ( n15154 & n15478 ) | ( n15154 & n23037 ) | ( n15478 & n23037 ) ;
  assign n25628 = n1342 | n5414 ;
  assign n25629 = ~n2332 & n25628 ;
  assign n25630 = ~n8499 & n9581 ;
  assign n25631 = n25630 ^ n20767 ^ 1'b0 ;
  assign n25632 = n14157 ^ n9324 ^ n1309 ;
  assign n25633 = n25632 ^ n754 ^ x21 ;
  assign n25634 = ( n2723 & n2773 ) | ( n2723 & n7299 ) | ( n2773 & n7299 ) ;
  assign n25635 = n25634 ^ x18 ^ 1'b0 ;
  assign n25636 = ~n15353 & n25635 ;
  assign n25637 = n15129 ^ x79 ^ 1'b0 ;
  assign n25638 = n25636 & ~n25637 ;
  assign n25639 = n19780 & n25638 ;
  assign n25640 = ~n6422 & n25639 ;
  assign n25642 = n4141 & n25043 ;
  assign n25643 = n25642 ^ n3098 ^ 1'b0 ;
  assign n25641 = n7620 & n22303 ;
  assign n25644 = n25643 ^ n25641 ^ 1'b0 ;
  assign n25646 = n10183 ^ n5745 ^ n3847 ;
  assign n25645 = n5940 ^ n3703 ^ n736 ;
  assign n25647 = n25646 ^ n25645 ^ 1'b0 ;
  assign n25648 = n17635 | n25647 ;
  assign n25649 = ~n21152 & n25648 ;
  assign n25650 = ( n8601 & ~n24019 ) | ( n8601 & n25649 ) | ( ~n24019 & n25649 ) ;
  assign n25651 = n25650 ^ n5263 ^ 1'b0 ;
  assign n25652 = n6617 & n25651 ;
  assign n25653 = n2876 & ~n19664 ;
  assign n25654 = n2949 & ~n9274 ;
  assign n25655 = n25654 ^ n1869 ^ 1'b0 ;
  assign n25656 = ( ~n1590 & n7778 ) | ( ~n1590 & n15418 ) | ( n7778 & n15418 ) ;
  assign n25657 = ( n473 & n19149 ) | ( n473 & n21822 ) | ( n19149 & n21822 ) ;
  assign n25658 = ( ~n1776 & n5929 ) | ( ~n1776 & n23116 ) | ( n5929 & n23116 ) ;
  assign n25660 = n5786 ^ n2197 ^ 1'b0 ;
  assign n25659 = ( n1253 & n4051 ) | ( n1253 & ~n4745 ) | ( n4051 & ~n4745 ) ;
  assign n25661 = n25660 ^ n25659 ^ n23966 ;
  assign n25662 = n8343 ^ n346 ^ 1'b0 ;
  assign n25663 = n25661 & n25662 ;
  assign n25664 = n14617 ^ n9715 ^ n3715 ;
  assign n25665 = ~n13522 & n25664 ;
  assign n25666 = n17668 | n25665 ;
  assign n25667 = n25666 ^ n10202 ^ 1'b0 ;
  assign n25668 = ~n6503 & n7797 ;
  assign n25669 = n13267 ^ n9913 ^ 1'b0 ;
  assign n25670 = n6493 & n25669 ;
  assign n25671 = n25670 ^ n16368 ^ 1'b0 ;
  assign n25672 = n25668 | n25671 ;
  assign n25673 = ~n17330 & n19089 ;
  assign n25674 = n3861 & n25673 ;
  assign n25675 = n19594 ^ n10935 ^ 1'b0 ;
  assign n25676 = n17482 & n25675 ;
  assign n25677 = n25676 ^ n14867 ^ 1'b0 ;
  assign n25678 = n19148 & n25677 ;
  assign n25679 = n826 | n4710 ;
  assign n25680 = n4239 | n25679 ;
  assign n25681 = ( ~n4414 & n6324 ) | ( ~n4414 & n25680 ) | ( n6324 & n25680 ) ;
  assign n25682 = ( ~n1718 & n10564 ) | ( ~n1718 & n25681 ) | ( n10564 & n25681 ) ;
  assign n25683 = n3121 | n20244 ;
  assign n25684 = n2751 & ~n3220 ;
  assign n25685 = n25684 ^ n6038 ^ 1'b0 ;
  assign n25686 = n25685 ^ n2610 ^ 1'b0 ;
  assign n25687 = n10058 & ~n23117 ;
  assign n25688 = n24387 ^ n11933 ^ 1'b0 ;
  assign n25689 = n5702 & n25688 ;
  assign n25690 = n5041 ^ n940 ^ 1'b0 ;
  assign n25691 = n6297 & n10581 ;
  assign n25692 = n2670 & n25691 ;
  assign n25693 = n25692 ^ n10412 ^ 1'b0 ;
  assign n25694 = n19084 ^ n7459 ^ 1'b0 ;
  assign n25695 = n25694 ^ n24009 ^ n19031 ;
  assign n25697 = ~n2515 & n12916 ;
  assign n25698 = ~n13927 & n25697 ;
  assign n25696 = ( n5712 & n14271 ) | ( n5712 & ~n23017 ) | ( n14271 & ~n23017 ) ;
  assign n25699 = n25698 ^ n25696 ^ n25366 ;
  assign n25701 = n20247 ^ n8018 ^ n304 ;
  assign n25702 = ( x92 & n9803 ) | ( x92 & ~n25701 ) | ( n9803 & ~n25701 ) ;
  assign n25700 = n2115 & n22811 ;
  assign n25703 = n25702 ^ n25700 ^ n2347 ;
  assign n25704 = ( n2389 & n4661 ) | ( n2389 & ~n7361 ) | ( n4661 & ~n7361 ) ;
  assign n25705 = n25704 ^ n12376 ^ 1'b0 ;
  assign n25706 = ~n10663 & n25705 ;
  assign n25707 = n12091 & n12823 ;
  assign n25708 = ~n24467 & n25707 ;
  assign n25709 = n25708 ^ n3542 ^ 1'b0 ;
  assign n25710 = x79 & ~n25709 ;
  assign n25711 = n15746 ^ n15302 ^ 1'b0 ;
  assign n25712 = n25711 ^ n20194 ^ n9901 ;
  assign n25713 = n22222 ^ n6072 ^ n1154 ;
  assign n25715 = n23599 ^ n12919 ^ n374 ;
  assign n25714 = n2734 & n4323 ;
  assign n25716 = n25715 ^ n25714 ^ 1'b0 ;
  assign n25717 = n15256 ^ n11747 ^ n406 ;
  assign n25718 = n25716 & n25717 ;
  assign n25719 = ( ~n5442 & n15783 ) | ( ~n5442 & n22560 ) | ( n15783 & n22560 ) ;
  assign n25720 = ~n15667 & n20536 ;
  assign n25721 = ~n485 & n15536 ;
  assign n25722 = ~n1324 & n5903 ;
  assign n25723 = ( n7070 & n11047 ) | ( n7070 & n21780 ) | ( n11047 & n21780 ) ;
  assign n25724 = n7476 ^ n139 ^ 1'b0 ;
  assign n25725 = ~n224 & n25724 ;
  assign n25726 = n7040 & n10300 ;
  assign n25727 = ~n434 & n12138 ;
  assign n25728 = n25727 ^ n7108 ^ 1'b0 ;
  assign n25729 = ( n21344 & n25726 ) | ( n21344 & ~n25728 ) | ( n25726 & ~n25728 ) ;
  assign n25730 = ~n25725 & n25729 ;
  assign n25731 = n25010 ^ n17836 ^ 1'b0 ;
  assign n25732 = n4942 & n9218 ;
  assign n25733 = ~n15727 & n25732 ;
  assign n25734 = ~n20604 & n25733 ;
  assign n25735 = n7788 & ~n9002 ;
  assign n25736 = n25735 ^ n208 ^ 1'b0 ;
  assign n25737 = ~n23928 & n25736 ;
  assign n25738 = n9691 & n25737 ;
  assign n25739 = n2593 & n25738 ;
  assign n25740 = n9203 | n13574 ;
  assign n25741 = n14746 & ~n25740 ;
  assign n25742 = n16778 ^ n5556 ^ x71 ;
  assign n25743 = n14745 ^ n7449 ^ 1'b0 ;
  assign n25744 = ( n7547 & ~n25742 ) | ( n7547 & n25743 ) | ( ~n25742 & n25743 ) ;
  assign n25745 = ( n296 & n10219 ) | ( n296 & n17729 ) | ( n10219 & n17729 ) ;
  assign n25746 = n5381 | n25745 ;
  assign n25747 = n25744 | n25746 ;
  assign n25748 = n11769 ^ n7852 ^ 1'b0 ;
  assign n25749 = n14767 & n25748 ;
  assign n25750 = ( n9299 & n16940 ) | ( n9299 & ~n25749 ) | ( n16940 & ~n25749 ) ;
  assign n25751 = ( ~n1686 & n7814 ) | ( ~n1686 & n8199 ) | ( n7814 & n8199 ) ;
  assign n25752 = n25751 ^ n3965 ^ 1'b0 ;
  assign n25753 = n3465 & n7062 ;
  assign n25754 = n25753 ^ n21329 ^ n11730 ;
  assign n25755 = n25754 ^ n13914 ^ n1962 ;
  assign n25756 = n17823 | n25755 ;
  assign n25758 = n18369 ^ n6139 ^ n3175 ;
  assign n25757 = n1561 & ~n5729 ;
  assign n25759 = n25758 ^ n25757 ^ n22470 ;
  assign n25760 = n13997 ^ n13152 ^ x25 ;
  assign n25761 = n1819 | n25760 ;
  assign n25762 = n11049 ^ n5969 ^ n295 ;
  assign n25763 = n15888 & ~n25762 ;
  assign n25764 = n25763 ^ n9777 ^ 1'b0 ;
  assign n25765 = ~n2053 & n11437 ;
  assign n25766 = n25765 ^ n11629 ^ 1'b0 ;
  assign n25767 = n16716 & ~n25766 ;
  assign n25768 = n13973 ^ n8661 ^ n5880 ;
  assign n25769 = n2535 | n25768 ;
  assign n25770 = n23421 & n25769 ;
  assign n25771 = n3049 & n14455 ;
  assign n25772 = n1510 & n25771 ;
  assign n25773 = n10330 | n25772 ;
  assign n25774 = n25773 ^ n12606 ^ 1'b0 ;
  assign n25775 = ( n5493 & n19744 ) | ( n5493 & ~n24889 ) | ( n19744 & ~n24889 ) ;
  assign n25776 = n8669 ^ n7457 ^ n979 ;
  assign n25777 = ( n3625 & n4138 ) | ( n3625 & ~n25776 ) | ( n4138 & ~n25776 ) ;
  assign n25778 = n4744 ^ n4432 ^ 1'b0 ;
  assign n25779 = n8964 | n25778 ;
  assign n25780 = n25779 ^ n23859 ^ n7300 ;
  assign n25781 = n5578 & ~n8245 ;
  assign n25783 = n19524 ^ n5941 ^ n3411 ;
  assign n25782 = n6063 ^ n4663 ^ n4022 ;
  assign n25784 = n25783 ^ n25782 ^ n18670 ;
  assign n25785 = ( n4419 & ~n7113 ) | ( n4419 & n9307 ) | ( ~n7113 & n9307 ) ;
  assign n25786 = ~n543 & n25785 ;
  assign n25787 = n11616 & n25786 ;
  assign n25788 = n22963 | n25787 ;
  assign n25789 = n10295 & ~n25788 ;
  assign n25790 = n9603 ^ n7006 ^ n4723 ;
  assign n25791 = n24978 ^ n11283 ^ 1'b0 ;
  assign n25792 = n25790 | n25791 ;
  assign n25793 = x102 & n14061 ;
  assign n25794 = n25793 ^ n7192 ^ 1'b0 ;
  assign n25795 = ( ~n12102 & n16577 ) | ( ~n12102 & n25794 ) | ( n16577 & n25794 ) ;
  assign n25796 = ( ~n7296 & n10642 ) | ( ~n7296 & n25117 ) | ( n10642 & n25117 ) ;
  assign n25797 = n25795 & ~n25796 ;
  assign n25798 = n25797 ^ n22188 ^ 1'b0 ;
  assign n25799 = n4516 ^ n695 ^ 1'b0 ;
  assign n25800 = n15659 | n25799 ;
  assign n25801 = n23389 ^ n2277 ^ x80 ;
  assign n25802 = n21038 & ~n24446 ;
  assign n25803 = n25802 ^ n230 ^ 1'b0 ;
  assign n25804 = n14221 ^ n3757 ^ 1'b0 ;
  assign n25809 = ( n2279 & n2984 ) | ( n2279 & n10346 ) | ( n2984 & n10346 ) ;
  assign n25805 = n11967 ^ n1585 ^ 1'b0 ;
  assign n25806 = n7430 | n25805 ;
  assign n25807 = ( ~n7732 & n12679 ) | ( ~n7732 & n25806 ) | ( n12679 & n25806 ) ;
  assign n25808 = n2386 | n25807 ;
  assign n25810 = n25809 ^ n25808 ^ 1'b0 ;
  assign n25811 = ( ~n2272 & n25804 ) | ( ~n2272 & n25810 ) | ( n25804 & n25810 ) ;
  assign n25812 = n9932 & n13455 ;
  assign n25813 = ~n23178 & n25812 ;
  assign n25814 = ~n18919 & n25813 ;
  assign n25815 = n16302 & ~n19474 ;
  assign n25816 = n1591 | n25815 ;
  assign n25817 = n19162 & ~n25816 ;
  assign n25818 = n6148 | n25817 ;
  assign n25819 = n25818 ^ n13869 ^ 1'b0 ;
  assign n25820 = n14903 ^ n14092 ^ 1'b0 ;
  assign n25821 = n3883 | n25820 ;
  assign n25822 = n12887 ^ n7727 ^ 1'b0 ;
  assign n25823 = n2876 & n25822 ;
  assign n25824 = n767 | n25782 ;
  assign n25825 = n25420 ^ n24182 ^ n19387 ;
  assign n25826 = n1171 | n18254 ;
  assign n25827 = ( n4718 & n17528 ) | ( n4718 & ~n25826 ) | ( n17528 & ~n25826 ) ;
  assign n25828 = n25827 ^ n5145 ^ 1'b0 ;
  assign n25829 = n19966 ^ n16620 ^ n3312 ;
  assign n25830 = ~n15690 & n17371 ;
  assign n25831 = ( n1131 & ~n18222 ) | ( n1131 & n25830 ) | ( ~n18222 & n25830 ) ;
  assign n25832 = n9478 | n25255 ;
  assign n25833 = n3819 & ~n25832 ;
  assign n25834 = n18769 ^ n4093 ^ 1'b0 ;
  assign n25835 = ~n25833 & n25834 ;
  assign n25836 = n16149 ^ n6066 ^ n3218 ;
  assign n25837 = n21059 & n25836 ;
  assign n25838 = ~n25835 & n25837 ;
  assign n25839 = ~n22848 & n24485 ;
  assign n25840 = n25839 ^ n20948 ^ 1'b0 ;
  assign n25841 = n12270 ^ n5182 ^ 1'b0 ;
  assign n25842 = n12710 ^ n5915 ^ n365 ;
  assign n25843 = n7492 & n25070 ;
  assign n25848 = n11310 ^ n10954 ^ 1'b0 ;
  assign n25846 = ( n776 & ~n5134 ) | ( n776 & n5519 ) | ( ~n5134 & n5519 ) ;
  assign n25844 = n8032 ^ n5654 ^ n1527 ;
  assign n25845 = ~n4741 & n25844 ;
  assign n25847 = n25846 ^ n25845 ^ 1'b0 ;
  assign n25849 = n25848 ^ n25847 ^ n5622 ;
  assign n25850 = n25210 ^ n17277 ^ n9547 ;
  assign n25851 = ~n19052 & n24085 ;
  assign n25852 = ( n5392 & n18841 ) | ( n5392 & n25851 ) | ( n18841 & n25851 ) ;
  assign n25853 = n21830 ^ n7555 ^ 1'b0 ;
  assign n25858 = n14289 ^ n2217 ^ 1'b0 ;
  assign n25859 = n2029 & ~n25858 ;
  assign n25860 = n5862 | n7030 ;
  assign n25861 = ( ~n454 & n25859 ) | ( ~n454 & n25860 ) | ( n25859 & n25860 ) ;
  assign n25854 = n13816 ^ n637 ^ 1'b0 ;
  assign n25855 = n11770 | n25854 ;
  assign n25856 = n25855 ^ n3024 ^ 1'b0 ;
  assign n25857 = ~n18880 & n25856 ;
  assign n25862 = n25861 ^ n25857 ^ 1'b0 ;
  assign n25863 = ~n2013 & n15397 ;
  assign n25864 = n25863 ^ n2832 ^ 1'b0 ;
  assign n25865 = n25864 ^ n1678 ^ 1'b0 ;
  assign n25866 = n327 | n5526 ;
  assign n25867 = n16647 & ~n25866 ;
  assign n25868 = n24507 ^ n11835 ^ n5888 ;
  assign n25869 = n3169 | n16750 ;
  assign n25870 = n14204 | n25869 ;
  assign n25871 = ( ~n6155 & n18649 ) | ( ~n6155 & n25870 ) | ( n18649 & n25870 ) ;
  assign n25872 = ( n144 & n159 ) | ( n144 & n783 ) | ( n159 & n783 ) ;
  assign n25873 = n25872 ^ n6119 ^ n2269 ;
  assign n25874 = n8888 | n25873 ;
  assign n25875 = ( ~n2824 & n4757 ) | ( ~n2824 & n7110 ) | ( n4757 & n7110 ) ;
  assign n25876 = n25875 ^ n15589 ^ 1'b0 ;
  assign n25877 = ~n23568 & n25876 ;
  assign n25878 = n2522 & ~n5265 ;
  assign n25879 = n16162 & n16929 ;
  assign n25880 = ~n10531 & n21994 ;
  assign n25881 = n25880 ^ n13511 ^ n930 ;
  assign n25882 = n5421 | n12139 ;
  assign n25883 = n1407 & ~n8331 ;
  assign n25884 = ~n25882 & n25883 ;
  assign n25885 = n25884 ^ n15754 ^ n9717 ;
  assign n25886 = n25242 ^ n827 ^ 1'b0 ;
  assign n25887 = n2039 & n25886 ;
  assign n25888 = ~n415 & n25887 ;
  assign n25889 = n2305 ^ n2162 ^ 1'b0 ;
  assign n25890 = n2827 & ~n25889 ;
  assign n25891 = n23182 & n25890 ;
  assign n25892 = n5159 ^ n1689 ^ 1'b0 ;
  assign n25893 = n10047 & ~n14902 ;
  assign n25894 = ~n4390 & n25893 ;
  assign n25895 = n25894 ^ n15040 ^ n8117 ;
  assign n25896 = ( n9613 & n25892 ) | ( n9613 & n25895 ) | ( n25892 & n25895 ) ;
  assign n25897 = n16746 ^ n6506 ^ n6002 ;
  assign n25898 = n5421 & n17120 ;
  assign n25899 = n10380 ^ n6439 ^ 1'b0 ;
  assign n25902 = n6202 ^ n3748 ^ 1'b0 ;
  assign n25903 = n1467 | n25902 ;
  assign n25900 = n10872 ^ n4474 ^ n3086 ;
  assign n25901 = n18653 & n25900 ;
  assign n25904 = n25903 ^ n25901 ^ 1'b0 ;
  assign n25905 = n6931 & n21179 ;
  assign n25906 = n25905 ^ n4716 ^ 1'b0 ;
  assign n25907 = ~n13009 & n25906 ;
  assign n25908 = n1150 & ~n10049 ;
  assign n25909 = n25908 ^ n16203 ^ n14773 ;
  assign n25910 = n7816 & ~n25909 ;
  assign n25911 = n5476 & n25910 ;
  assign n25912 = n3965 & ~n6793 ;
  assign n25913 = n25912 ^ n10439 ^ 1'b0 ;
  assign n25917 = n6382 ^ n3030 ^ 1'b0 ;
  assign n25914 = ( n2031 & n5718 ) | ( n2031 & ~n15405 ) | ( n5718 & ~n15405 ) ;
  assign n25915 = n5937 & ~n12463 ;
  assign n25916 = ~n25914 & n25915 ;
  assign n25918 = n25917 ^ n25916 ^ n6590 ;
  assign n25919 = n6668 ^ n6123 ^ 1'b0 ;
  assign n25920 = ~n5991 & n15343 ;
  assign n25921 = n15619 & n25920 ;
  assign n25922 = n25921 ^ n11679 ^ n11365 ;
  assign n25923 = ( n6332 & n8268 ) | ( n6332 & ~n11312 ) | ( n8268 & ~n11312 ) ;
  assign n25925 = n3198 & ~n8835 ;
  assign n25924 = n4927 | n15619 ;
  assign n25926 = n25925 ^ n25924 ^ 1'b0 ;
  assign n25927 = n4220 | n7768 ;
  assign n25928 = n21480 & ~n25927 ;
  assign n25929 = n12450 ^ n7605 ^ 1'b0 ;
  assign n25930 = n4012 | n8820 ;
  assign n25931 = n25930 ^ n12514 ^ 1'b0 ;
  assign n25933 = n13255 | n13696 ;
  assign n25932 = n2569 & n5657 ;
  assign n25934 = n25933 ^ n25932 ^ 1'b0 ;
  assign n25935 = ( n4792 & ~n22804 ) | ( n4792 & n25934 ) | ( ~n22804 & n25934 ) ;
  assign n25936 = ~n885 & n14221 ;
  assign n25937 = n3131 | n25936 ;
  assign n25938 = n11696 & ~n25937 ;
  assign n25939 = n25938 ^ n14216 ^ 1'b0 ;
  assign n25940 = n196 | n5909 ;
  assign n25941 = n25289 ^ n7232 ^ 1'b0 ;
  assign n25942 = ( n16563 & n25940 ) | ( n16563 & n25941 ) | ( n25940 & n25941 ) ;
  assign n25943 = ( n153 & ~n5304 ) | ( n153 & n13989 ) | ( ~n5304 & n13989 ) ;
  assign n25944 = n25943 ^ n12787 ^ 1'b0 ;
  assign n25945 = ~n9344 & n17686 ;
  assign n25946 = n19061 & n25945 ;
  assign n25947 = ~n3322 & n3457 ;
  assign n25948 = n25947 ^ n10722 ^ 1'b0 ;
  assign n25949 = n5808 | n17949 ;
  assign n25950 = n25948 | n25949 ;
  assign n25952 = n6040 ^ n3346 ^ n1874 ;
  assign n25953 = n17916 & n25952 ;
  assign n25951 = n1525 & n21224 ;
  assign n25954 = n25953 ^ n25951 ^ 1'b0 ;
  assign n25955 = ( n8930 & n11027 ) | ( n8930 & ~n23499 ) | ( n11027 & ~n23499 ) ;
  assign n25956 = n25955 ^ n13461 ^ n3390 ;
  assign n25957 = ( ~n7432 & n8414 ) | ( ~n7432 & n12363 ) | ( n8414 & n12363 ) ;
  assign n25958 = ( ~n2609 & n3287 ) | ( ~n2609 & n13814 ) | ( n3287 & n13814 ) ;
  assign n25959 = n25958 ^ n17342 ^ 1'b0 ;
  assign n25960 = n11346 ^ n4680 ^ 1'b0 ;
  assign n25961 = n7124 | n25960 ;
  assign n25962 = ~n4810 & n5765 ;
  assign n25963 = n25962 ^ n13370 ^ 1'b0 ;
  assign n25964 = n9109 & n25963 ;
  assign n25965 = n25964 ^ n21447 ^ 1'b0 ;
  assign n25966 = ( n3468 & n3775 ) | ( n3468 & ~n25965 ) | ( n3775 & ~n25965 ) ;
  assign n25967 = n23580 | n25966 ;
  assign n25968 = n25967 ^ n4878 ^ 1'b0 ;
  assign n25969 = n14716 ^ n14300 ^ 1'b0 ;
  assign n25970 = n23051 ^ n1278 ^ 1'b0 ;
  assign n25971 = n9076 & n25970 ;
  assign n25972 = n893 ^ n846 ^ 1'b0 ;
  assign n25973 = n17852 & n25972 ;
  assign n25974 = ( ~x63 & n17617 ) | ( ~x63 & n21110 ) | ( n17617 & n21110 ) ;
  assign n25975 = ( n7487 & n16404 ) | ( n7487 & n16648 ) | ( n16404 & n16648 ) ;
  assign n25976 = n290 & ~n8339 ;
  assign n25977 = n25976 ^ n21424 ^ 1'b0 ;
  assign n25981 = ( n878 & ~n1666 ) | ( n878 & n16750 ) | ( ~n1666 & n16750 ) ;
  assign n25982 = n25981 ^ n25859 ^ n21887 ;
  assign n25983 = n24423 ^ n15627 ^ 1'b0 ;
  assign n25984 = ~n25982 & n25983 ;
  assign n25978 = n5476 | n13862 ;
  assign n25979 = n25978 ^ n3030 ^ 1'b0 ;
  assign n25980 = n12869 | n25979 ;
  assign n25985 = n25984 ^ n25980 ^ 1'b0 ;
  assign n25986 = ( n8030 & n10219 ) | ( n8030 & ~n25985 ) | ( n10219 & ~n25985 ) ;
  assign n25987 = ( ~n2813 & n6946 ) | ( ~n2813 & n16258 ) | ( n6946 & n16258 ) ;
  assign n25988 = ( n1108 & ~n8883 ) | ( n1108 & n25987 ) | ( ~n8883 & n25987 ) ;
  assign n25989 = n25988 ^ n12631 ^ n2197 ;
  assign n25990 = ( n6802 & n19097 ) | ( n6802 & n20318 ) | ( n19097 & n20318 ) ;
  assign n25991 = ~n5759 & n12889 ;
  assign n25992 = n7844 & n25991 ;
  assign n25993 = n23611 & ~n25992 ;
  assign n25994 = n25990 & n25993 ;
  assign n25995 = n19944 ^ n14369 ^ 1'b0 ;
  assign n25996 = ( ~n20476 & n22908 ) | ( ~n20476 & n23954 ) | ( n22908 & n23954 ) ;
  assign n25997 = n18016 ^ n17570 ^ 1'b0 ;
  assign n25998 = n632 | n15802 ;
  assign n25999 = ( n4530 & n8988 ) | ( n4530 & ~n9842 ) | ( n8988 & ~n9842 ) ;
  assign n26000 = n4864 & ~n10494 ;
  assign n26001 = n26000 ^ n7752 ^ 1'b0 ;
  assign n26002 = ~n3694 & n4232 ;
  assign n26003 = n26002 ^ n9860 ^ 1'b0 ;
  assign n26004 = n24669 ^ n6072 ^ 1'b0 ;
  assign n26005 = ~n13140 & n26004 ;
  assign n26007 = ~n1365 & n2787 ;
  assign n26006 = n2829 & n10652 ;
  assign n26008 = n26007 ^ n26006 ^ 1'b0 ;
  assign n26009 = n9544 ^ n1693 ^ 1'b0 ;
  assign n26010 = n2742 | n19075 ;
  assign n26011 = n26010 ^ n19002 ^ 1'b0 ;
  assign n26012 = n10537 ^ n8823 ^ 1'b0 ;
  assign n26013 = n838 & n26012 ;
  assign n26014 = n26013 ^ n11135 ^ 1'b0 ;
  assign n26015 = x94 & ~n26014 ;
  assign n26016 = ( n5321 & n6065 ) | ( n5321 & ~n7409 ) | ( n6065 & ~n7409 ) ;
  assign n26017 = n26016 ^ n12563 ^ 1'b0 ;
  assign n26018 = n17483 | n26017 ;
  assign n26019 = n6921 & n9536 ;
  assign n26020 = n26019 ^ n1555 ^ 1'b0 ;
  assign n26021 = ( n9838 & n26018 ) | ( n9838 & n26020 ) | ( n26018 & n26020 ) ;
  assign n26022 = ~n6489 & n12416 ;
  assign n26023 = n4021 & n26022 ;
  assign n26024 = ( n22422 & n22794 ) | ( n22422 & ~n26023 ) | ( n22794 & ~n26023 ) ;
  assign n26025 = n6483 & n6668 ;
  assign n26026 = ( ~n2315 & n3121 ) | ( ~n2315 & n22345 ) | ( n3121 & n22345 ) ;
  assign n26027 = n26026 ^ n12164 ^ 1'b0 ;
  assign n26028 = n26025 | n26027 ;
  assign n26029 = n12025 | n26028 ;
  assign n26030 = n26029 ^ n17929 ^ 1'b0 ;
  assign n26031 = n4624 & ~n14852 ;
  assign n26032 = n4129 & n20177 ;
  assign n26033 = n26032 ^ n24555 ^ 1'b0 ;
  assign n26034 = n3874 ^ n1671 ^ 1'b0 ;
  assign n26035 = n4221 ^ n1189 ^ 1'b0 ;
  assign n26036 = n11918 ^ n7910 ^ 1'b0 ;
  assign n26037 = n4850 & ~n26036 ;
  assign n26038 = ( ~n425 & n557 ) | ( ~n425 & n26037 ) | ( n557 & n26037 ) ;
  assign n26039 = n19472 ^ n18219 ^ n16991 ;
  assign n26040 = n26039 ^ x65 ^ 1'b0 ;
  assign n26043 = n8272 ^ n7614 ^ 1'b0 ;
  assign n26041 = n3028 & n5008 ;
  assign n26042 = ~n2416 & n26041 ;
  assign n26044 = n26043 ^ n26042 ^ n9967 ;
  assign n26045 = ~n8076 & n14438 ;
  assign n26046 = n26045 ^ n17811 ^ 1'b0 ;
  assign n26047 = ~n13350 & n22719 ;
  assign n26048 = n8697 & n26047 ;
  assign n26049 = n26048 ^ n20543 ^ n2104 ;
  assign n26050 = n24724 & n26049 ;
  assign n26051 = n19940 & n26050 ;
  assign n26057 = n10780 | n21152 ;
  assign n26058 = n19468 & ~n26057 ;
  assign n26055 = n551 & n6147 ;
  assign n26056 = n26055 ^ n10629 ^ 1'b0 ;
  assign n26052 = n23413 ^ n3010 ^ n1242 ;
  assign n26053 = n26052 ^ n17411 ^ x47 ;
  assign n26054 = n26053 ^ n2093 ^ n1100 ;
  assign n26059 = n26058 ^ n26056 ^ n26054 ;
  assign n26060 = n20221 & ~n26059 ;
  assign n26061 = n14891 & n26060 ;
  assign n26062 = n16757 & ~n26061 ;
  assign n26063 = n2887 & n3386 ;
  assign n26064 = n26063 ^ n10360 ^ 1'b0 ;
  assign n26065 = ( n9108 & n15144 ) | ( n9108 & ~n16306 ) | ( n15144 & ~n16306 ) ;
  assign n26066 = n7421 ^ n4275 ^ 1'b0 ;
  assign n26067 = n26066 ^ n23557 ^ n2829 ;
  assign n26068 = n26067 ^ n9279 ^ n1437 ;
  assign n26069 = ( n1798 & n9607 ) | ( n1798 & ~n13030 ) | ( n9607 & ~n13030 ) ;
  assign n26070 = n26069 ^ n22562 ^ n13168 ;
  assign n26071 = n5302 & n21203 ;
  assign n26072 = ~n12624 & n19397 ;
  assign n26073 = ( n3325 & n26071 ) | ( n3325 & n26072 ) | ( n26071 & n26072 ) ;
  assign n26074 = n6274 ^ n1986 ^ 1'b0 ;
  assign n26075 = n12335 ^ n7725 ^ n6204 ;
  assign n26076 = n22960 | n26075 ;
  assign n26077 = n1368 | n8789 ;
  assign n26078 = n26077 ^ n23448 ^ 1'b0 ;
  assign n26079 = ( n8757 & n10417 ) | ( n8757 & ~n10963 ) | ( n10417 & ~n10963 ) ;
  assign n26080 = ~n5004 & n26079 ;
  assign n26081 = n4990 & n26080 ;
  assign n26082 = n13882 ^ x77 ^ 1'b0 ;
  assign n26083 = n16982 & n26082 ;
  assign n26084 = n8156 ^ n3633 ^ 1'b0 ;
  assign n26085 = n26083 | n26084 ;
  assign n26086 = n3206 ^ n357 ^ 1'b0 ;
  assign n26087 = ( n8424 & ~n20611 ) | ( n8424 & n26086 ) | ( ~n20611 & n26086 ) ;
  assign n26088 = n26087 ^ n25181 ^ n2011 ;
  assign n26089 = n21397 ^ n15373 ^ n4719 ;
  assign n26090 = ( n3139 & n13222 ) | ( n3139 & n23871 ) | ( n13222 & n23871 ) ;
  assign n26091 = n16772 ^ n13672 ^ n4818 ;
  assign n26092 = n26091 ^ n23390 ^ n8079 ;
  assign n26093 = n19113 ^ n12414 ^ n4632 ;
  assign n26094 = n17012 ^ n15196 ^ n611 ;
  assign n26095 = ~n18030 & n26094 ;
  assign n26096 = n11763 & ~n26095 ;
  assign n26097 = n26096 ^ n11452 ^ 1'b0 ;
  assign n26098 = n1882 | n26097 ;
  assign n26099 = n10156 & n18864 ;
  assign n26100 = ( n6298 & n18766 ) | ( n6298 & ~n26094 ) | ( n18766 & ~n26094 ) ;
  assign n26101 = n19615 ^ n9615 ^ 1'b0 ;
  assign n26102 = ( n380 & n7168 ) | ( n380 & ~n19208 ) | ( n7168 & ~n19208 ) ;
  assign n26103 = n6657 ^ n3724 ^ 1'b0 ;
  assign n26104 = ~n23686 & n26103 ;
  assign n26105 = n26102 & n26104 ;
  assign n26106 = ( n344 & ~n19757 ) | ( n344 & n21620 ) | ( ~n19757 & n21620 ) ;
  assign n26107 = n2366 & n9837 ;
  assign n26108 = n12763 & ~n26107 ;
  assign n26109 = ( n3373 & n7211 ) | ( n3373 & ~n24581 ) | ( n7211 & ~n24581 ) ;
  assign n26110 = ~n4018 & n13482 ;
  assign n26111 = n26109 & n26110 ;
  assign n26112 = n1244 & ~n13698 ;
  assign n26113 = n18635 & n20499 ;
  assign n26114 = n6607 | n7208 ;
  assign n26115 = ( n2121 & n2530 ) | ( n2121 & ~n25856 ) | ( n2530 & ~n25856 ) ;
  assign n26116 = n3283 ^ n3200 ^ 1'b0 ;
  assign n26117 = n26116 ^ n4890 ^ 1'b0 ;
  assign n26118 = ( n12790 & ~n21221 ) | ( n12790 & n26117 ) | ( ~n21221 & n26117 ) ;
  assign n26123 = ( n8661 & ~n18225 ) | ( n8661 & n20733 ) | ( ~n18225 & n20733 ) ;
  assign n26122 = ( n6823 & n7115 ) | ( n6823 & ~n13752 ) | ( n7115 & ~n13752 ) ;
  assign n26119 = ~n4567 & n9295 ;
  assign n26120 = n26119 ^ n1691 ^ 1'b0 ;
  assign n26121 = ( n12123 & n17629 ) | ( n12123 & n26120 ) | ( n17629 & n26120 ) ;
  assign n26124 = n26123 ^ n26122 ^ n26121 ;
  assign n26125 = ( n4593 & n15632 ) | ( n4593 & n26124 ) | ( n15632 & n26124 ) ;
  assign n26126 = n11905 ^ n8530 ^ n1123 ;
  assign n26127 = n6222 & n18595 ;
  assign n26129 = n7913 & n7914 ;
  assign n26130 = n26129 ^ n8723 ^ 1'b0 ;
  assign n26131 = n5402 | n26130 ;
  assign n26128 = n574 & n5971 ;
  assign n26132 = n26131 ^ n26128 ^ 1'b0 ;
  assign n26135 = n3433 & n4290 ;
  assign n26133 = n4070 & n10149 ;
  assign n26134 = n26133 ^ n1546 ^ n1084 ;
  assign n26136 = n26135 ^ n26134 ^ n2960 ;
  assign n26137 = ( n7233 & n13145 ) | ( n7233 & n22850 ) | ( n13145 & n22850 ) ;
  assign n26138 = n5593 | n26137 ;
  assign n26139 = ( n6486 & n19978 ) | ( n6486 & n25557 ) | ( n19978 & n25557 ) ;
  assign n26140 = n1786 & n26139 ;
  assign n26141 = n13893 & n16168 ;
  assign n26142 = n12782 & n26141 ;
  assign n26143 = n13854 | n23990 ;
  assign n26144 = n26143 ^ n9694 ^ 1'b0 ;
  assign n26145 = ( n12470 & n14672 ) | ( n12470 & n19490 ) | ( n14672 & n19490 ) ;
  assign n26146 = n26145 ^ n17992 ^ n206 ;
  assign n26147 = n5665 & n26146 ;
  assign n26148 = n4477 ^ n4137 ^ 1'b0 ;
  assign n26149 = ( n13353 & n14086 ) | ( n13353 & n26148 ) | ( n14086 & n26148 ) ;
  assign n26150 = n26149 ^ n19271 ^ n15354 ;
  assign n26151 = n6692 & n11025 ;
  assign n26152 = n20490 ^ n8117 ^ n8074 ;
  assign n26153 = n26152 ^ n7816 ^ 1'b0 ;
  assign n26154 = n2894 | n13432 ;
  assign n26155 = n8113 | n26154 ;
  assign n26156 = n26155 ^ n6260 ^ 1'b0 ;
  assign n26157 = n23879 & n26156 ;
  assign n26158 = n7817 | n13498 ;
  assign n26159 = n26158 ^ n7456 ^ 1'b0 ;
  assign n26160 = n554 | n5370 ;
  assign n26161 = n26160 ^ n5513 ^ 1'b0 ;
  assign n26162 = n17304 & n26161 ;
  assign n26163 = n10904 & ~n12645 ;
  assign n26164 = n4476 & n26163 ;
  assign n26165 = ( n3419 & n7806 ) | ( n3419 & ~n12892 ) | ( n7806 & ~n12892 ) ;
  assign n26166 = n21710 ^ n17876 ^ n6310 ;
  assign n26167 = n2343 & ~n5779 ;
  assign n26168 = n26167 ^ n3398 ^ 1'b0 ;
  assign n26169 = n26166 & ~n26168 ;
  assign n26170 = ( n3032 & n26165 ) | ( n3032 & n26169 ) | ( n26165 & n26169 ) ;
  assign n26171 = n7843 ^ n4289 ^ 1'b0 ;
  assign n26173 = n1887 & ~n12910 ;
  assign n26172 = n12248 & ~n13434 ;
  assign n26174 = n26173 ^ n26172 ^ 1'b0 ;
  assign n26175 = n26174 ^ n22968 ^ n19115 ;
  assign n26176 = ( ~n1431 & n22930 ) | ( ~n1431 & n26175 ) | ( n22930 & n26175 ) ;
  assign n26177 = n19132 ^ n17339 ^ 1'b0 ;
  assign n26179 = n6250 ^ n2934 ^ 1'b0 ;
  assign n26180 = ~n4263 & n26179 ;
  assign n26178 = n6564 ^ n1551 ^ n436 ;
  assign n26181 = n26180 ^ n26178 ^ 1'b0 ;
  assign n26182 = ~n10433 & n22908 ;
  assign n26183 = n9216 & n26182 ;
  assign n26184 = n23097 | n26183 ;
  assign n26185 = n12039 | n26184 ;
  assign n26186 = n15617 ^ n11229 ^ n6079 ;
  assign n26187 = n16165 | n26186 ;
  assign n26188 = n13696 ^ n3481 ^ n708 ;
  assign n26189 = n1235 | n4492 ;
  assign n26190 = n25507 ^ n7644 ^ 1'b0 ;
  assign n26191 = n22634 ^ n16109 ^ n12484 ;
  assign n26192 = n26191 ^ n535 ^ 1'b0 ;
  assign n26193 = n5836 & n14002 ;
  assign n26194 = n26192 & n26193 ;
  assign n26195 = n6975 & ~n7175 ;
  assign n26196 = n14401 ^ n4910 ^ 1'b0 ;
  assign n26197 = ( n5040 & n10276 ) | ( n5040 & n26196 ) | ( n10276 & n26196 ) ;
  assign n26198 = n12208 ^ n9675 ^ 1'b0 ;
  assign n26199 = ~n5328 & n26198 ;
  assign n26200 = n26199 ^ n16684 ^ 1'b0 ;
  assign n26201 = ( ~n13319 & n23528 ) | ( ~n13319 & n26200 ) | ( n23528 & n26200 ) ;
  assign n26202 = n742 & ~n19860 ;
  assign n26203 = n21078 ^ n1077 ^ 1'b0 ;
  assign n26204 = n1343 & ~n26203 ;
  assign n26205 = n2922 & n26204 ;
  assign n26206 = n3519 & ~n3988 ;
  assign n26207 = n26206 ^ n10315 ^ 1'b0 ;
  assign n26208 = n12923 | n14407 ;
  assign n26209 = n26208 ^ n6059 ^ 1'b0 ;
  assign n26210 = n204 & ~n8159 ;
  assign n26211 = n7937 & n26210 ;
  assign n26212 = ( ~n4091 & n9855 ) | ( ~n4091 & n26211 ) | ( n9855 & n26211 ) ;
  assign n26213 = n6787 & n19202 ;
  assign n26214 = n26213 ^ n233 ^ 1'b0 ;
  assign n26215 = ( ~n10916 & n12560 ) | ( ~n10916 & n26214 ) | ( n12560 & n26214 ) ;
  assign n26216 = n13158 ^ n1761 ^ 1'b0 ;
  assign n26217 = n26216 ^ n9059 ^ n8791 ;
  assign n26218 = n4525 | n26217 ;
  assign n26219 = ( n2792 & ~n8909 ) | ( n2792 & n26218 ) | ( ~n8909 & n26218 ) ;
  assign n26220 = ( n3027 & n7627 ) | ( n3027 & ~n17504 ) | ( n7627 & ~n17504 ) ;
  assign n26222 = ( n5996 & n6891 ) | ( n5996 & ~n10846 ) | ( n6891 & ~n10846 ) ;
  assign n26221 = n11964 ^ n8468 ^ n7149 ;
  assign n26223 = n26222 ^ n26221 ^ n16013 ;
  assign n26224 = n25908 ^ n11337 ^ 1'b0 ;
  assign n26225 = n26223 & n26224 ;
  assign n26226 = n21349 | n21500 ;
  assign n26227 = n5582 & n21368 ;
  assign n26228 = n26227 ^ n24059 ^ 1'b0 ;
  assign n26229 = n4315 | n11770 ;
  assign n26230 = n17420 | n17802 ;
  assign n26231 = n9347 | n26230 ;
  assign n26232 = ~x122 & n13629 ;
  assign n26233 = ~n259 & n3033 ;
  assign n26234 = n19248 & n26233 ;
  assign n26235 = n19063 & ~n26234 ;
  assign n26236 = n10831 & ~n19684 ;
  assign n26237 = n26236 ^ n9263 ^ 1'b0 ;
  assign n26238 = n15110 & n26237 ;
  assign n26239 = ( ~n7188 & n11373 ) | ( ~n7188 & n26238 ) | ( n11373 & n26238 ) ;
  assign n26240 = n19998 ^ n5800 ^ n2209 ;
  assign n26241 = ( n15042 & n20582 ) | ( n15042 & n26240 ) | ( n20582 & n26240 ) ;
  assign n26242 = n26241 ^ n8641 ^ 1'b0 ;
  assign n26243 = n3195 ^ n1250 ^ 1'b0 ;
  assign n26244 = n11566 & n26243 ;
  assign n26245 = n26244 ^ n18670 ^ n14164 ;
  assign n26246 = ~n11260 & n17419 ;
  assign n26247 = n23081 ^ n16029 ^ n5129 ;
  assign n26248 = ~n13074 & n26247 ;
  assign n26249 = n3124 & ~n3790 ;
  assign n26250 = n26249 ^ n5266 ^ 1'b0 ;
  assign n26251 = n1399 | n1480 ;
  assign n26252 = n18982 ^ n16673 ^ 1'b0 ;
  assign n26253 = n26252 ^ n20548 ^ n11894 ;
  assign n26254 = n15036 ^ n12500 ^ 1'b0 ;
  assign n26255 = n13515 ^ n5997 ^ n5885 ;
  assign n26256 = n26255 ^ n14684 ^ 1'b0 ;
  assign n26257 = n23643 ^ n22207 ^ n6999 ;
  assign n26259 = n19444 ^ n1193 ^ x64 ;
  assign n26258 = ~n16780 & n22386 ;
  assign n26260 = n26259 ^ n26258 ^ 1'b0 ;
  assign n26261 = ~n12936 & n15294 ;
  assign n26262 = n26261 ^ n7998 ^ 1'b0 ;
  assign n26263 = n2253 | n9734 ;
  assign n26264 = n26263 ^ n9082 ^ 1'b0 ;
  assign n26265 = n23350 ^ n460 ^ 1'b0 ;
  assign n26266 = n577 | n26265 ;
  assign n26267 = n26266 ^ n24237 ^ 1'b0 ;
  assign n26268 = n26267 ^ n21887 ^ 1'b0 ;
  assign n26269 = n5683 & n8744 ;
  assign n26270 = n26269 ^ n1534 ^ 1'b0 ;
  assign n26271 = ~x113 & n1642 ;
  assign n26272 = n26271 ^ n20005 ^ n6425 ;
  assign n26273 = ( n10149 & n10771 ) | ( n10149 & ~n14071 ) | ( n10771 & ~n14071 ) ;
  assign n26274 = n11621 ^ n5498 ^ 1'b0 ;
  assign n26275 = n22115 & ~n26274 ;
  assign n26276 = n26275 ^ n25906 ^ 1'b0 ;
  assign n26277 = n15709 & n21872 ;
  assign n26278 = n26277 ^ n5133 ^ 1'b0 ;
  assign n26279 = n26278 ^ n16446 ^ 1'b0 ;
  assign n26280 = n6486 & n26279 ;
  assign n26281 = n10051 ^ n3984 ^ 1'b0 ;
  assign n26282 = ( n4252 & ~n26280 ) | ( n4252 & n26281 ) | ( ~n26280 & n26281 ) ;
  assign n26284 = n13920 ^ n9925 ^ 1'b0 ;
  assign n26285 = n16502 & n26284 ;
  assign n26286 = n17942 & n26285 ;
  assign n26283 = n7494 & n8829 ;
  assign n26287 = n26286 ^ n26283 ^ 1'b0 ;
  assign n26288 = ( n2702 & ~n6967 ) | ( n2702 & n9060 ) | ( ~n6967 & n9060 ) ;
  assign n26289 = n26288 ^ n13670 ^ 1'b0 ;
  assign n26290 = ~n8412 & n26289 ;
  assign n26291 = n26290 ^ n9335 ^ 1'b0 ;
  assign n26292 = n10125 & ~n13118 ;
  assign n26293 = n26292 ^ n5068 ^ 1'b0 ;
  assign n26294 = n19977 ^ n8342 ^ 1'b0 ;
  assign n26295 = n26293 & n26294 ;
  assign n26296 = n14906 | n18978 ;
  assign n26297 = n26023 ^ n13097 ^ 1'b0 ;
  assign n26298 = n1893 & n26297 ;
  assign n26299 = ~n23999 & n26298 ;
  assign n26300 = n7676 ^ n6170 ^ n3964 ;
  assign n26301 = n24714 & n26300 ;
  assign n26302 = n26301 ^ n20994 ^ 1'b0 ;
  assign n26303 = n4703 ^ n1754 ^ 1'b0 ;
  assign n26304 = n2381 | n26303 ;
  assign n26305 = n9593 & ~n26304 ;
  assign n26306 = n26305 ^ n11618 ^ 1'b0 ;
  assign n26307 = n26306 ^ n19490 ^ n3374 ;
  assign n26308 = n3704 ^ n1686 ^ 1'b0 ;
  assign n26309 = n26308 ^ n18834 ^ n16733 ;
  assign n26310 = n16735 ^ n3902 ^ n2744 ;
  assign n26311 = n6207 | n13104 ;
  assign n26312 = n819 | n26311 ;
  assign n26313 = n12250 ^ n7806 ^ n4489 ;
  assign n26314 = n26313 ^ n17677 ^ 1'b0 ;
  assign n26315 = n26314 ^ n18079 ^ 1'b0 ;
  assign n26316 = n26312 & n26315 ;
  assign n26317 = ~n19018 & n26316 ;
  assign n26318 = ~n2165 & n18701 ;
  assign n26319 = n7339 ^ n2325 ^ n1519 ;
  assign n26320 = x127 | n11622 ;
  assign n26321 = n11466 ^ n11053 ^ n10837 ;
  assign n26322 = ( n5578 & ~n26320 ) | ( n5578 & n26321 ) | ( ~n26320 & n26321 ) ;
  assign n26323 = n14717 ^ n13330 ^ 1'b0 ;
  assign n26324 = ( n26319 & n26322 ) | ( n26319 & ~n26323 ) | ( n26322 & ~n26323 ) ;
  assign n26325 = n19405 | n21723 ;
  assign n26326 = n26325 ^ n4973 ^ 1'b0 ;
  assign n26327 = n26324 | n26326 ;
  assign n26328 = n13708 ^ n6172 ^ 1'b0 ;
  assign n26329 = n14526 & n26328 ;
  assign n26330 = n2420 & ~n11659 ;
  assign n26331 = n26330 ^ n25210 ^ n3166 ;
  assign n26332 = n4109 & n26331 ;
  assign n26333 = n20915 & n26332 ;
  assign n26334 = n24381 ^ n12345 ^ n2849 ;
  assign n26335 = ~n10056 & n26334 ;
  assign n26336 = n14522 & ~n20374 ;
  assign n26337 = n12864 ^ n4086 ^ 1'b0 ;
  assign n26339 = n14749 | n26056 ;
  assign n26338 = n833 & ~n1456 ;
  assign n26340 = n26339 ^ n26338 ^ n13587 ;
  assign n26341 = n10038 & ~n15971 ;
  assign n26342 = n10751 ^ n1864 ^ n1173 ;
  assign n26343 = n16773 ^ n2655 ^ n2458 ;
  assign n26344 = n23124 | n26343 ;
  assign n26345 = n26342 & ~n26344 ;
  assign n26347 = ( ~n1009 & n3235 ) | ( ~n1009 & n10196 ) | ( n3235 & n10196 ) ;
  assign n26346 = ~n7752 & n16699 ;
  assign n26348 = n26347 ^ n26346 ^ 1'b0 ;
  assign n26349 = n1032 & n7475 ;
  assign n26350 = n26349 ^ n23607 ^ 1'b0 ;
  assign n26351 = n9746 & n19490 ;
  assign n26352 = n827 | n10961 ;
  assign n26353 = n599 | n13939 ;
  assign n26354 = n4087 | n13900 ;
  assign n26355 = n1032 | n26354 ;
  assign n26356 = ( ~n251 & n575 ) | ( ~n251 & n4722 ) | ( n575 & n4722 ) ;
  assign n26357 = n2550 & ~n18373 ;
  assign n26358 = ~n26356 & n26357 ;
  assign n26359 = ~n3682 & n11215 ;
  assign n26360 = n1718 & n26359 ;
  assign n26361 = n1858 | n10839 ;
  assign n26362 = ( ~n3790 & n4354 ) | ( ~n3790 & n13088 ) | ( n4354 & n13088 ) ;
  assign n26363 = ( ~n3046 & n23672 ) | ( ~n3046 & n26362 ) | ( n23672 & n26362 ) ;
  assign n26364 = ( ~n14751 & n14968 ) | ( ~n14751 & n17744 ) | ( n14968 & n17744 ) ;
  assign n26365 = n2694 | n12631 ;
  assign n26366 = n26365 ^ n8721 ^ n5171 ;
  assign n26368 = n10186 ^ n2286 ^ 1'b0 ;
  assign n26369 = ~n10000 & n26368 ;
  assign n26367 = ~n5479 & n23338 ;
  assign n26370 = n26369 ^ n26367 ^ n14554 ;
  assign n26371 = n8052 ^ n5079 ^ 1'b0 ;
  assign n26372 = n8508 | n26371 ;
  assign n26373 = n2042 | n26372 ;
  assign n26374 = n3432 | n26373 ;
  assign n26375 = n26016 ^ n24201 ^ 1'b0 ;
  assign n26376 = ~n23932 & n26375 ;
  assign n26377 = n23555 ^ n20094 ^ n9664 ;
  assign n26378 = ~n9007 & n11448 ;
  assign n26379 = n26377 & n26378 ;
  assign n26380 = n10998 | n17350 ;
  assign n26381 = n26380 ^ n3447 ^ 1'b0 ;
  assign n26382 = n9398 ^ n341 ^ 1'b0 ;
  assign n26383 = n9614 & ~n15305 ;
  assign n26384 = n26382 & n26383 ;
  assign n26385 = n26384 ^ n25064 ^ n2285 ;
  assign n26386 = n6799 | n19329 ;
  assign n26387 = n2296 | n3070 ;
  assign n26388 = n26387 ^ n3874 ^ 1'b0 ;
  assign n26389 = ( n24292 & n26386 ) | ( n24292 & ~n26388 ) | ( n26386 & ~n26388 ) ;
  assign n26390 = n16162 ^ n10465 ^ n2911 ;
  assign n26391 = n26390 ^ n4628 ^ 1'b0 ;
  assign n26392 = n10330 | n26391 ;
  assign n26393 = ~n9580 & n26392 ;
  assign n26394 = ( n2900 & n18583 ) | ( n2900 & ~n21611 ) | ( n18583 & ~n21611 ) ;
  assign n26395 = n20472 ^ n6583 ^ 1'b0 ;
  assign n26397 = n8373 ^ n7152 ^ n1527 ;
  assign n26396 = n1328 & ~n12923 ;
  assign n26398 = n26397 ^ n26396 ^ 1'b0 ;
  assign n26399 = n15119 & ~n17800 ;
  assign n26400 = n13413 ^ n10314 ^ 1'b0 ;
  assign n26401 = ~n188 & n26400 ;
  assign n26402 = n15837 & n23372 ;
  assign n26403 = n26402 ^ n4436 ^ 1'b0 ;
  assign n26404 = ( n7602 & n12763 ) | ( n7602 & n21794 ) | ( n12763 & n21794 ) ;
  assign n26405 = n5036 & n7177 ;
  assign n26406 = ( ~n3118 & n10562 ) | ( ~n3118 & n26405 ) | ( n10562 & n26405 ) ;
  assign n26407 = n6114 & ~n11937 ;
  assign n26408 = n26407 ^ n16362 ^ n5506 ;
  assign n26409 = n26408 ^ n1934 ^ 1'b0 ;
  assign n26410 = n19723 | n26120 ;
  assign n26411 = n20181 ^ n3625 ^ 1'b0 ;
  assign n26412 = n23726 & ~n26411 ;
  assign n26413 = n5870 | n7770 ;
  assign n26414 = ( n10018 & n23905 ) | ( n10018 & n26413 ) | ( n23905 & n26413 ) ;
  assign n26415 = n6916 ^ n2455 ^ 1'b0 ;
  assign n26416 = n7088 & ~n26415 ;
  assign n26417 = n26416 ^ n23165 ^ n4162 ;
  assign n26418 = n26417 ^ n16600 ^ 1'b0 ;
  assign n26419 = n26414 & ~n26418 ;
  assign n26420 = ~n9091 & n11053 ;
  assign n26421 = n9324 & n26420 ;
  assign n26422 = ~n1994 & n18154 ;
  assign n26423 = n17590 | n20076 ;
  assign n26424 = n26423 ^ n15381 ^ 1'b0 ;
  assign n26425 = n13863 ^ n9556 ^ 1'b0 ;
  assign n26426 = n9024 & ~n26425 ;
  assign n26427 = n14324 & n19925 ;
  assign n26428 = n26427 ^ n14097 ^ n10231 ;
  assign n26431 = n3919 ^ n1475 ^ n1055 ;
  assign n26432 = ~n7132 & n26431 ;
  assign n26433 = n1723 & n26432 ;
  assign n26429 = n13026 & ~n18608 ;
  assign n26430 = n7384 & n26429 ;
  assign n26434 = n26433 ^ n26430 ^ n6027 ;
  assign n26435 = n26434 ^ n20046 ^ n12798 ;
  assign n26436 = n19366 ^ n16362 ^ n2100 ;
  assign n26437 = n6624 & n26436 ;
  assign n26438 = n26437 ^ n7450 ^ 1'b0 ;
  assign n26439 = ( n1043 & n8323 ) | ( n1043 & ~n26438 ) | ( n8323 & ~n26438 ) ;
  assign n26440 = n17912 ^ n16350 ^ n15126 ;
  assign n26441 = ( ~n2095 & n2455 ) | ( ~n2095 & n6572 ) | ( n2455 & n6572 ) ;
  assign n26442 = n6128 | n20144 ;
  assign n26443 = n16697 | n26442 ;
  assign n26444 = n13204 ^ n10824 ^ 1'b0 ;
  assign n26445 = n26443 & ~n26444 ;
  assign n26446 = n17434 ^ n12437 ^ 1'b0 ;
  assign n26447 = n7636 & n26446 ;
  assign n26448 = n14353 & n26447 ;
  assign n26449 = n5554 ^ n5503 ^ 1'b0 ;
  assign n26450 = n19049 ^ n6985 ^ 1'b0 ;
  assign n26451 = n2794 & n26450 ;
  assign n26452 = n6134 ^ n2136 ^ 1'b0 ;
  assign n26453 = n26452 ^ n3836 ^ n2124 ;
  assign n26454 = ~n3215 & n26453 ;
  assign n26455 = n26454 ^ n2361 ^ 1'b0 ;
  assign n26456 = ~n6781 & n26455 ;
  assign n26457 = n7951 ^ n505 ^ 1'b0 ;
  assign n26458 = ~n26456 & n26457 ;
  assign n26461 = n16171 ^ n7863 ^ 1'b0 ;
  assign n26459 = n5347 & n5848 ;
  assign n26460 = n16208 & n26459 ;
  assign n26462 = n26461 ^ n26460 ^ n7509 ;
  assign n26463 = n141 & n2802 ;
  assign n26464 = ~n9585 & n26463 ;
  assign n26465 = ~n9145 & n26464 ;
  assign n26466 = ~n10105 & n14776 ;
  assign n26467 = ( ~n6169 & n18181 ) | ( ~n6169 & n26466 ) | ( n18181 & n26466 ) ;
  assign n26468 = n7436 & n7948 ;
  assign n26469 = n19704 & n25383 ;
  assign n26475 = n12911 & n16657 ;
  assign n26476 = n10596 & n26475 ;
  assign n26472 = n15430 ^ n2442 ^ x90 ;
  assign n26473 = n26472 ^ n5776 ^ n1409 ;
  assign n26470 = ~n2858 & n7376 ;
  assign n26471 = ~n18057 & n26470 ;
  assign n26474 = n26473 ^ n26471 ^ n3790 ;
  assign n26477 = n26476 ^ n26474 ^ n8883 ;
  assign n26478 = n17367 ^ n5730 ^ n1632 ;
  assign n26479 = n4181 & n12938 ;
  assign n26480 = n3879 & n26479 ;
  assign n26481 = n7806 ^ n5260 ^ 1'b0 ;
  assign n26482 = ~n1372 & n26481 ;
  assign n26483 = n26482 ^ n13091 ^ n8944 ;
  assign n26484 = ( n11519 & ~n26480 ) | ( n11519 & n26483 ) | ( ~n26480 & n26483 ) ;
  assign n26485 = n3235 ^ n1080 ^ 1'b0 ;
  assign n26486 = n12524 & ~n26485 ;
  assign n26487 = n20043 ^ n1256 ^ 1'b0 ;
  assign n26489 = n18363 ^ n4847 ^ 1'b0 ;
  assign n26490 = n9378 & ~n26489 ;
  assign n26488 = n7853 | n18364 ;
  assign n26491 = n26490 ^ n26488 ^ 1'b0 ;
  assign n26492 = n9841 | n25807 ;
  assign n26493 = n3619 ^ x127 ^ 1'b0 ;
  assign n26494 = n26493 ^ n16477 ^ n3271 ;
  assign n26495 = ~n5727 & n6455 ;
  assign n26496 = n22650 & n26495 ;
  assign n26497 = n18696 | n26496 ;
  assign n26501 = n7741 ^ n5233 ^ 1'b0 ;
  assign n26499 = n2178 ^ x56 ^ 1'b0 ;
  assign n26500 = ( n9748 & n11848 ) | ( n9748 & n26499 ) | ( n11848 & n26499 ) ;
  assign n26498 = ~n22305 & n23101 ;
  assign n26502 = n26501 ^ n26500 ^ n26498 ;
  assign n26503 = n12395 ^ n3889 ^ 1'b0 ;
  assign n26504 = n12530 & n26503 ;
  assign n26505 = n24005 & n26504 ;
  assign n26506 = n9770 & n23948 ;
  assign n26507 = ~n3788 & n26506 ;
  assign n26508 = ~n508 & n26507 ;
  assign n26509 = ( ~n2326 & n7717 ) | ( ~n2326 & n15408 ) | ( n7717 & n15408 ) ;
  assign n26510 = n4818 & n19590 ;
  assign n26511 = n1068 & n4000 ;
  assign n26512 = n26511 ^ n5780 ^ 1'b0 ;
  assign n26513 = n26510 & n26512 ;
  assign n26514 = n26513 ^ n16962 ^ n9043 ;
  assign n26515 = n16114 ^ n1880 ^ 1'b0 ;
  assign n26516 = n13232 ^ n10710 ^ 1'b0 ;
  assign n26517 = n4006 | n26516 ;
  assign n26518 = ( n20444 & n26515 ) | ( n20444 & ~n26517 ) | ( n26515 & ~n26517 ) ;
  assign n26519 = n16698 ^ n9817 ^ n6071 ;
  assign n26520 = n23145 ^ n656 ^ 1'b0 ;
  assign n26521 = ~n11533 & n26520 ;
  assign n26525 = ( n4928 & n5880 ) | ( n4928 & ~n13737 ) | ( n5880 & ~n13737 ) ;
  assign n26523 = n8970 & ~n12185 ;
  assign n26524 = n26523 ^ n1615 ^ 1'b0 ;
  assign n26522 = ( n1710 & n11601 ) | ( n1710 & ~n19886 ) | ( n11601 & ~n19886 ) ;
  assign n26526 = n26525 ^ n26524 ^ n26522 ;
  assign n26527 = n12234 ^ n829 ^ 1'b0 ;
  assign n26528 = n13849 & ~n26527 ;
  assign n26529 = n26528 ^ n5434 ^ 1'b0 ;
  assign n26530 = n20986 | n26529 ;
  assign n26531 = n466 & ~n10187 ;
  assign n26532 = n26531 ^ n25181 ^ 1'b0 ;
  assign n26533 = ( n1137 & n15191 ) | ( n1137 & ~n26532 ) | ( n15191 & ~n26532 ) ;
  assign n26534 = n16607 ^ n13314 ^ 1'b0 ;
  assign n26535 = ( ~n16077 & n19837 ) | ( ~n16077 & n26534 ) | ( n19837 & n26534 ) ;
  assign n26536 = n7902 ^ n2189 ^ 1'b0 ;
  assign n26537 = n13127 & n20234 ;
  assign n26538 = ( n652 & ~n3354 ) | ( n652 & n4256 ) | ( ~n3354 & n4256 ) ;
  assign n26539 = ( n2511 & n22328 ) | ( n2511 & ~n26538 ) | ( n22328 & ~n26538 ) ;
  assign n26540 = ( n26536 & n26537 ) | ( n26536 & n26539 ) | ( n26537 & n26539 ) ;
  assign n26541 = n4402 & ~n9268 ;
  assign n26542 = n26541 ^ n8273 ^ 1'b0 ;
  assign n26543 = n4401 ^ n4140 ^ n669 ;
  assign n26544 = n26543 ^ n23405 ^ n4212 ;
  assign n26545 = n4277 & ~n13810 ;
  assign n26546 = ~n26544 & n26545 ;
  assign n26547 = n17471 & n26072 ;
  assign n26548 = n26547 ^ n3718 ^ 1'b0 ;
  assign n26549 = n23832 ^ n9245 ^ 1'b0 ;
  assign n26550 = ( n15752 & n23238 ) | ( n15752 & ~n26549 ) | ( n23238 & ~n26549 ) ;
  assign n26551 = n4445 & n14175 ;
  assign n26552 = ~n13865 & n26551 ;
  assign n26553 = n26552 ^ n21063 ^ n7507 ;
  assign n26554 = n6364 & n23119 ;
  assign n26555 = ( n2845 & n19589 ) | ( n2845 & n26554 ) | ( n19589 & n26554 ) ;
  assign n26556 = ~n8570 & n10180 ;
  assign n26557 = ~n15992 & n26556 ;
  assign n26558 = n23201 ^ n2624 ^ 1'b0 ;
  assign n26559 = ~n14150 & n26558 ;
  assign n26560 = ( n17447 & n26557 ) | ( n17447 & n26559 ) | ( n26557 & n26559 ) ;
  assign n26562 = n11487 & ~n19842 ;
  assign n26561 = n8820 ^ n5514 ^ n776 ;
  assign n26563 = n26562 ^ n26561 ^ n2081 ;
  assign n26564 = n11404 ^ n5395 ^ 1'b0 ;
  assign n26565 = ( n1372 & n5679 ) | ( n1372 & n17434 ) | ( n5679 & n17434 ) ;
  assign n26566 = n26565 ^ n3527 ^ 1'b0 ;
  assign n26567 = n26564 & n26566 ;
  assign n26568 = n21189 ^ n2244 ^ 1'b0 ;
  assign n26569 = n26567 & ~n26568 ;
  assign n26570 = n10531 ^ n1435 ^ 1'b0 ;
  assign n26571 = n1204 & n20490 ;
  assign n26572 = n26571 ^ n25257 ^ n22733 ;
  assign n26573 = n2043 & ~n14846 ;
  assign n26574 = n7913 ^ n406 ^ 1'b0 ;
  assign n26575 = ~n26573 & n26574 ;
  assign n26576 = ( n656 & ~n16214 ) | ( n656 & n18087 ) | ( ~n16214 & n18087 ) ;
  assign n26577 = n26576 ^ n12332 ^ n6786 ;
  assign n26578 = n8288 ^ n2301 ^ n1621 ;
  assign n26579 = n26578 ^ n7845 ^ 1'b0 ;
  assign n26580 = ( ~n7740 & n9391 ) | ( ~n7740 & n26579 ) | ( n9391 & n26579 ) ;
  assign n26581 = ~n3633 & n11710 ;
  assign n26582 = ~n15035 & n26581 ;
  assign n26583 = ( ~n5068 & n8368 ) | ( ~n5068 & n22537 ) | ( n8368 & n22537 ) ;
  assign n26584 = ( n16711 & n18408 ) | ( n16711 & ~n26583 ) | ( n18408 & ~n26583 ) ;
  assign n26585 = n15608 ^ n15533 ^ n4493 ;
  assign n26586 = n17625 & n26585 ;
  assign n26587 = n26584 & n26586 ;
  assign n26588 = n19738 ^ n16302 ^ 1'b0 ;
  assign n26589 = n26588 ^ n2965 ^ 1'b0 ;
  assign n26590 = n14560 ^ n1676 ^ 1'b0 ;
  assign n26591 = n17178 & ~n26590 ;
  assign n26592 = n7990 & ~n8802 ;
  assign n26593 = n15173 & n20373 ;
  assign n26594 = n26593 ^ n8269 ^ 1'b0 ;
  assign n26595 = n26592 & ~n26594 ;
  assign n26596 = n19132 ^ n7898 ^ 1'b0 ;
  assign n26597 = n9515 ^ n8782 ^ n8099 ;
  assign n26599 = ~n6042 & n11716 ;
  assign n26600 = ~n11787 & n26599 ;
  assign n26598 = n17775 ^ n8793 ^ 1'b0 ;
  assign n26601 = n26600 ^ n26598 ^ n1089 ;
  assign n26602 = ( ~n8178 & n10259 ) | ( ~n8178 & n23867 ) | ( n10259 & n23867 ) ;
  assign n26603 = ( n3383 & n20876 ) | ( n3383 & ~n22807 ) | ( n20876 & ~n22807 ) ;
  assign n26604 = n12388 ^ n486 ^ n256 ;
  assign n26605 = n26604 ^ n18303 ^ 1'b0 ;
  assign n26606 = ~n18846 & n26605 ;
  assign n26607 = n26606 ^ n23820 ^ 1'b0 ;
  assign n26608 = n21627 ^ n982 ^ 1'b0 ;
  assign n26609 = n21376 & n26608 ;
  assign n26610 = n9067 ^ n5797 ^ 1'b0 ;
  assign n26611 = n11957 & n26610 ;
  assign n26612 = n26611 ^ n4783 ^ 1'b0 ;
  assign n26613 = n20144 | n26612 ;
  assign n26614 = n13489 ^ n7382 ^ n3371 ;
  assign n26615 = n15070 & n26614 ;
  assign n26616 = n26615 ^ n11496 ^ 1'b0 ;
  assign n26617 = n25645 ^ n1586 ^ 1'b0 ;
  assign n26618 = n308 | n17151 ;
  assign n26619 = n26618 ^ n2336 ^ 1'b0 ;
  assign n26620 = n10219 & n19762 ;
  assign n26621 = n26620 ^ n18023 ^ 1'b0 ;
  assign n26622 = n14048 & n23195 ;
  assign n26623 = n21620 & n26622 ;
  assign n26624 = n9163 & ~n22517 ;
  assign n26625 = n12749 ^ n9455 ^ 1'b0 ;
  assign n26627 = n11524 ^ n7175 ^ 1'b0 ;
  assign n26628 = n26319 | n26627 ;
  assign n26629 = ( n3782 & n11187 ) | ( n3782 & ~n26628 ) | ( n11187 & ~n26628 ) ;
  assign n26626 = n19948 | n22877 ;
  assign n26630 = n26629 ^ n26626 ^ 1'b0 ;
  assign n26631 = n14619 ^ n14564 ^ n5631 ;
  assign n26632 = n26631 ^ n22324 ^ 1'b0 ;
  assign n26633 = ( ~n8746 & n12236 ) | ( ~n8746 & n18688 ) | ( n12236 & n18688 ) ;
  assign n26634 = ( n3498 & ~n10206 ) | ( n3498 & n22706 ) | ( ~n10206 & n22706 ) ;
  assign n26635 = n18834 ^ n7832 ^ n2108 ;
  assign n26636 = ( n1051 & n22200 ) | ( n1051 & n26635 ) | ( n22200 & n26635 ) ;
  assign n26637 = n25048 & n26636 ;
  assign n26641 = n9101 ^ n6694 ^ n2472 ;
  assign n26638 = n26452 ^ n6999 ^ n6124 ;
  assign n26639 = n26638 ^ n2316 ^ 1'b0 ;
  assign n26640 = n2272 | n26639 ;
  assign n26642 = n26641 ^ n26640 ^ 1'b0 ;
  assign n26644 = n1678 & n11386 ;
  assign n26645 = ~n9257 & n26644 ;
  assign n26643 = ~n5088 & n13234 ;
  assign n26646 = n26645 ^ n26643 ^ 1'b0 ;
  assign n26647 = n4048 & ~n8675 ;
  assign n26648 = n16711 ^ n2192 ^ 1'b0 ;
  assign n26649 = n3473 & ~n26648 ;
  assign n26650 = ( n18117 & n26647 ) | ( n18117 & n26649 ) | ( n26647 & n26649 ) ;
  assign n26651 = ( n3756 & ~n25306 ) | ( n3756 & n26650 ) | ( ~n25306 & n26650 ) ;
  assign n26652 = n12724 ^ x76 ^ 1'b0 ;
  assign n26653 = n26652 ^ n25648 ^ n2762 ;
  assign n26654 = n25869 ^ n23209 ^ 1'b0 ;
  assign n26655 = n1934 & n6016 ;
  assign n26656 = n26655 ^ n8838 ^ 1'b0 ;
  assign n26657 = n4462 | n10984 ;
  assign n26658 = n26657 ^ n2608 ^ 1'b0 ;
  assign n26659 = n646 & ~n3110 ;
  assign n26660 = n24006 ^ n9142 ^ n3885 ;
  assign n26661 = n22813 & ~n26660 ;
  assign n26662 = ( ~x37 & n9766 ) | ( ~x37 & n11849 ) | ( n9766 & n11849 ) ;
  assign n26663 = ( n1776 & ~n3817 ) | ( n1776 & n9613 ) | ( ~n3817 & n9613 ) ;
  assign n26664 = n8426 ^ n4446 ^ n3389 ;
  assign n26665 = n26664 ^ n3645 ^ n269 ;
  assign n26666 = n24898 ^ n5513 ^ 1'b0 ;
  assign n26667 = n26666 ^ n8688 ^ n6637 ;
  assign n26668 = n26667 ^ n14300 ^ n6816 ;
  assign n26669 = n11626 ^ n7710 ^ n2891 ;
  assign n26670 = n18821 ^ n2430 ^ 1'b0 ;
  assign n26671 = n24409 & n26670 ;
  assign n26672 = n3909 & n9565 ;
  assign n26673 = n26672 ^ n10957 ^ n5791 ;
  assign n26674 = n21471 ^ n7613 ^ n557 ;
  assign n26675 = ~n3696 & n9643 ;
  assign n26676 = n6966 | n26675 ;
  assign n26677 = n26135 & ~n26676 ;
  assign n26678 = n21963 ^ n16418 ^ 1'b0 ;
  assign n26679 = x14 & ~n26678 ;
  assign n26680 = n883 & ~n8873 ;
  assign n26681 = n26680 ^ n5542 ^ 1'b0 ;
  assign n26682 = n6488 & n26300 ;
  assign n26683 = n26681 & n26682 ;
  assign n26684 = n8525 & ~n14301 ;
  assign n26685 = n26684 ^ n6016 ^ 1'b0 ;
  assign n26686 = n26685 ^ n24828 ^ n11431 ;
  assign n26687 = ( n3965 & ~n17148 ) | ( n3965 & n23869 ) | ( ~n17148 & n23869 ) ;
  assign n26688 = n20720 ^ n17528 ^ n2359 ;
  assign n26689 = n25569 ^ n7300 ^ 1'b0 ;
  assign n26691 = ( x95 & ~n1780 ) | ( x95 & n5798 ) | ( ~n1780 & n5798 ) ;
  assign n26692 = n26691 ^ n7985 ^ n6199 ;
  assign n26693 = n173 & ~n26692 ;
  assign n26694 = n23873 & n26693 ;
  assign n26690 = ~n1441 & n20220 ;
  assign n26695 = n26694 ^ n26690 ^ 1'b0 ;
  assign n26696 = n3105 & n7232 ;
  assign n26697 = n26696 ^ n3824 ^ 1'b0 ;
  assign n26698 = x61 & n18860 ;
  assign n26699 = n26698 ^ n7611 ^ 1'b0 ;
  assign n26700 = n18235 & n26699 ;
  assign n26701 = n26700 ^ n18753 ^ 1'b0 ;
  assign n26702 = n243 | n2305 ;
  assign n26703 = n9617 & ~n26702 ;
  assign n26704 = x83 & ~n16445 ;
  assign n26705 = n21414 ^ n3807 ^ n1813 ;
  assign n26706 = n26705 ^ n2038 ^ 1'b0 ;
  assign n26707 = n26706 ^ n16127 ^ n10019 ;
  assign n26708 = n14883 ^ n7608 ^ 1'b0 ;
  assign n26709 = n269 & ~n26708 ;
  assign n26710 = n2762 & n26709 ;
  assign n26711 = ~n3606 & n26710 ;
  assign n26712 = n11162 | n26152 ;
  assign n26713 = n26712 ^ n2614 ^ 1'b0 ;
  assign n26714 = n1371 ^ n406 ^ 1'b0 ;
  assign n26715 = ~n5631 & n26714 ;
  assign n26716 = n20424 ^ n897 ^ 1'b0 ;
  assign n26717 = n19636 & n26716 ;
  assign n26718 = ( n938 & ~n4584 ) | ( n938 & n8685 ) | ( ~n4584 & n8685 ) ;
  assign n26723 = n12698 ^ n7639 ^ n4436 ;
  assign n26720 = n4658 & n7112 ;
  assign n26721 = n26720 ^ n808 ^ 1'b0 ;
  assign n26722 = ~n1732 & n26721 ;
  assign n26724 = n26723 ^ n26722 ^ 1'b0 ;
  assign n26719 = n22006 ^ n16709 ^ n4092 ;
  assign n26725 = n26724 ^ n26719 ^ n16629 ;
  assign n26728 = ~n5839 & n19642 ;
  assign n26726 = n14203 ^ n12511 ^ 1'b0 ;
  assign n26727 = ~n13416 & n26726 ;
  assign n26729 = n26728 ^ n26727 ^ n6391 ;
  assign n26730 = n4075 & ~n16766 ;
  assign n26731 = n26730 ^ n15392 ^ 1'b0 ;
  assign n26732 = n5887 | n18451 ;
  assign n26733 = n26732 ^ n8220 ^ 1'b0 ;
  assign n26734 = n15833 ^ n2901 ^ 1'b0 ;
  assign n26736 = n1622 & ~n3186 ;
  assign n26737 = n26736 ^ n8683 ^ 1'b0 ;
  assign n26735 = ( n627 & n7429 ) | ( n627 & n13956 ) | ( n7429 & n13956 ) ;
  assign n26738 = n26737 ^ n26735 ^ n144 ;
  assign n26739 = n4775 | n10989 ;
  assign n26740 = ( n12250 & ~n22529 ) | ( n12250 & n26739 ) | ( ~n22529 & n26739 ) ;
  assign n26741 = n8993 & ~n14310 ;
  assign n26742 = n17601 ^ n7971 ^ 1'b0 ;
  assign n26743 = n2744 & n26742 ;
  assign n26744 = ( n10105 & n25815 ) | ( n10105 & n26743 ) | ( n25815 & n26743 ) ;
  assign n26745 = n7098 | n11777 ;
  assign n26746 = ~n24888 & n26745 ;
  assign n26747 = ~n8704 & n26746 ;
  assign n26748 = n14228 ^ n1754 ^ 1'b0 ;
  assign n26749 = n2839 & ~n26748 ;
  assign n26750 = n3086 & ~n4380 ;
  assign n26751 = n26750 ^ n24422 ^ 1'b0 ;
  assign n26752 = n6702 | n8446 ;
  assign n26753 = n26751 | n26752 ;
  assign n26755 = ~n236 & n527 ;
  assign n26756 = n26755 ^ n806 ^ 1'b0 ;
  assign n26757 = n10024 & ~n26756 ;
  assign n26754 = n23993 ^ n8329 ^ 1'b0 ;
  assign n26758 = n26757 ^ n26754 ^ 1'b0 ;
  assign n26759 = n26758 ^ n8541 ^ 1'b0 ;
  assign n26760 = n22803 & ~n26628 ;
  assign n26761 = n20603 & n26760 ;
  assign n26762 = n7926 & n22646 ;
  assign n26763 = ~n23139 & n26762 ;
  assign n26764 = n26763 ^ n4832 ^ 1'b0 ;
  assign n26765 = ( n5647 & n15996 ) | ( n5647 & n26764 ) | ( n15996 & n26764 ) ;
  assign n26766 = ( n3749 & n9942 ) | ( n3749 & ~n20428 ) | ( n9942 & ~n20428 ) ;
  assign n26767 = n19884 ^ n9544 ^ n7436 ;
  assign n26768 = n4497 | n21277 ;
  assign n26769 = ( n9327 & ~n14252 ) | ( n9327 & n20729 ) | ( ~n14252 & n20729 ) ;
  assign n26770 = ( n11021 & n26768 ) | ( n11021 & ~n26769 ) | ( n26768 & ~n26769 ) ;
  assign n26771 = n19160 & n21599 ;
  assign n26772 = n10400 & n26771 ;
  assign n26773 = n14505 | n26772 ;
  assign n26774 = x110 | n26773 ;
  assign n26776 = n6002 ^ n1089 ^ 1'b0 ;
  assign n26777 = n4726 | n17228 ;
  assign n26778 = n13060 | n26777 ;
  assign n26779 = n26776 & n26778 ;
  assign n26780 = n26779 ^ n6074 ^ 1'b0 ;
  assign n26775 = ~n1090 & n12543 ;
  assign n26781 = n26780 ^ n26775 ^ 1'b0 ;
  assign n26782 = n2227 | n25388 ;
  assign n26783 = n13333 ^ n4848 ^ 1'b0 ;
  assign n26784 = n26782 & n26783 ;
  assign n26786 = ~n7853 & n12895 ;
  assign n26785 = ( n6406 & ~n7242 ) | ( n6406 & n7921 ) | ( ~n7242 & n7921 ) ;
  assign n26787 = n26786 ^ n26785 ^ 1'b0 ;
  assign n26788 = n8479 ^ n8469 ^ 1'b0 ;
  assign n26789 = n26787 & n26788 ;
  assign n26790 = ( n165 & n3791 ) | ( n165 & ~n12550 ) | ( n3791 & ~n12550 ) ;
  assign n26791 = ( ~n3055 & n4091 ) | ( ~n3055 & n26790 ) | ( n4091 & n26790 ) ;
  assign n26792 = ~n7528 & n15126 ;
  assign n26793 = n17221 & n25386 ;
  assign n26794 = n26793 ^ n18915 ^ 1'b0 ;
  assign n26795 = ~n24174 & n26794 ;
  assign n26796 = n10866 & n26795 ;
  assign n26797 = n26796 ^ n25938 ^ n1934 ;
  assign n26798 = n13814 | n22420 ;
  assign n26799 = n2200 ^ n911 ^ 1'b0 ;
  assign n26800 = n3271 | n26799 ;
  assign n26801 = ~n2615 & n20957 ;
  assign n26802 = n26800 & n26801 ;
  assign n26803 = n449 & n25606 ;
  assign n26804 = ~n11406 & n26803 ;
  assign n26805 = n20444 ^ n18371 ^ 1'b0 ;
  assign n26806 = n21199 ^ n14919 ^ 1'b0 ;
  assign n26807 = n26805 & ~n26806 ;
  assign n26808 = ~n7772 & n8361 ;
  assign n26809 = n26808 ^ n2267 ^ 1'b0 ;
  assign n26810 = n9544 ^ n5965 ^ 1'b0 ;
  assign n26811 = n26809 & n26810 ;
  assign n26812 = n3260 & n14622 ;
  assign n26813 = n26812 ^ n11530 ^ 1'b0 ;
  assign n26814 = ( n5792 & ~n24968 ) | ( n5792 & n25698 ) | ( ~n24968 & n25698 ) ;
  assign n26815 = n1002 | n26814 ;
  assign n26816 = ~n22081 & n26815 ;
  assign n26819 = n17861 ^ n11518 ^ 1'b0 ;
  assign n26817 = n10261 ^ n5328 ^ 1'b0 ;
  assign n26818 = n2253 | n26817 ;
  assign n26820 = n26819 ^ n26818 ^ n11381 ;
  assign n26821 = n11656 ^ n1683 ^ n598 ;
  assign n26822 = n26821 ^ n6845 ^ n2621 ;
  assign n26823 = ~n11512 & n12994 ;
  assign n26824 = n4644 & n26823 ;
  assign n26825 = n3587 | n26824 ;
  assign n26826 = n11522 | n26825 ;
  assign n26827 = n1083 & ~n1504 ;
  assign n26828 = n8987 & n26827 ;
  assign n26829 = n10989 & ~n26828 ;
  assign n26830 = x114 & n26829 ;
  assign n26831 = n26830 ^ n15546 ^ 1'b0 ;
  assign n26832 = n6067 & ~n10474 ;
  assign n26833 = n26832 ^ n7254 ^ 1'b0 ;
  assign n26834 = n23689 | n26833 ;
  assign n26835 = x39 & n9740 ;
  assign n26836 = n26835 ^ n5127 ^ 1'b0 ;
  assign n26837 = n5297 & ~n13654 ;
  assign n26838 = n26836 | n26837 ;
  assign n26839 = n22054 | n26838 ;
  assign n26840 = n26839 ^ n10351 ^ 1'b0 ;
  assign n26841 = n26503 ^ n12842 ^ 1'b0 ;
  assign n26842 = n23323 ^ n16175 ^ n4821 ;
  assign n26843 = ( ~n144 & n3781 ) | ( ~n144 & n6344 ) | ( n3781 & n6344 ) ;
  assign n26844 = ( n14252 & ~n17941 ) | ( n14252 & n26843 ) | ( ~n17941 & n26843 ) ;
  assign n26845 = n15719 ^ n9789 ^ 1'b0 ;
  assign n26846 = n8600 & ~n26845 ;
  assign n26847 = n14307 ^ n5265 ^ 1'b0 ;
  assign n26848 = n26846 | n26847 ;
  assign n26849 = n6699 ^ n3679 ^ 1'b0 ;
  assign n26850 = ~n3827 & n26849 ;
  assign n26851 = n21629 ^ n14051 ^ n2057 ;
  assign n26852 = ( n3964 & n23281 ) | ( n3964 & ~n26851 ) | ( n23281 & ~n26851 ) ;
  assign n26855 = n845 | n8222 ;
  assign n26856 = n26855 ^ n2948 ^ 1'b0 ;
  assign n26853 = n15858 ^ n2701 ^ n1110 ;
  assign n26854 = n12678 | n26853 ;
  assign n26857 = n26856 ^ n26854 ^ 1'b0 ;
  assign n26858 = n947 & ~n26857 ;
  assign n26859 = ~n26852 & n26858 ;
  assign n26860 = ( n8972 & n17625 ) | ( n8972 & ~n18001 ) | ( n17625 & ~n18001 ) ;
  assign n26861 = ( n132 & n6143 ) | ( n132 & ~n26860 ) | ( n6143 & ~n26860 ) ;
  assign n26862 = n8038 & n20460 ;
  assign n26863 = ( n17064 & n17843 ) | ( n17064 & ~n26862 ) | ( n17843 & ~n26862 ) ;
  assign n26864 = n24105 ^ n4097 ^ n2423 ;
  assign n26865 = n17030 ^ n16282 ^ 1'b0 ;
  assign n26866 = n9280 | n9440 ;
  assign n26867 = n4535 ^ n3388 ^ 1'b0 ;
  assign n26868 = n333 & ~n11253 ;
  assign n26870 = x37 | n197 ;
  assign n26869 = x120 & ~n12563 ;
  assign n26871 = n26870 ^ n26869 ^ 1'b0 ;
  assign n26872 = n15563 ^ n9541 ^ n5387 ;
  assign n26873 = ( n14605 & n26405 ) | ( n14605 & n26872 ) | ( n26405 & n26872 ) ;
  assign n26875 = n3398 & ~n4564 ;
  assign n26876 = n26875 ^ n7052 ^ 1'b0 ;
  assign n26877 = ~n25255 & n26876 ;
  assign n26874 = n8738 & n14389 ;
  assign n26878 = n26877 ^ n26874 ^ n19575 ;
  assign n26879 = n6276 ^ n5556 ^ n523 ;
  assign n26881 = n8838 ^ n4089 ^ n2883 ;
  assign n26880 = n8943 ^ n6020 ^ 1'b0 ;
  assign n26882 = n26881 ^ n26880 ^ n5364 ;
  assign n26883 = n2634 & n14769 ;
  assign n26884 = n1612 & ~n10076 ;
  assign n26885 = n26884 ^ n5058 ^ 1'b0 ;
  assign n26886 = ~n26883 & n26885 ;
  assign n26887 = n24205 ^ n16410 ^ 1'b0 ;
  assign n26888 = n6811 & ~n26887 ;
  assign n26889 = n1404 & n18161 ;
  assign n26890 = ~n7030 & n13090 ;
  assign n26891 = n13961 ^ n5151 ^ 1'b0 ;
  assign n26892 = n22303 ^ n4673 ^ 1'b0 ;
  assign n26893 = ~n26891 & n26892 ;
  assign n26894 = n7095 ^ n2363 ^ 1'b0 ;
  assign n26895 = n16618 & n26894 ;
  assign n26896 = n26895 ^ n12889 ^ n9517 ;
  assign n26897 = n14308 & n19063 ;
  assign n26898 = ( n4609 & ~n9706 ) | ( n4609 & n26897 ) | ( ~n9706 & n26897 ) ;
  assign n26899 = ( ~n1462 & n10202 ) | ( ~n1462 & n26898 ) | ( n10202 & n26898 ) ;
  assign n26900 = ( n4745 & ~n10176 ) | ( n4745 & n23304 ) | ( ~n10176 & n23304 ) ;
  assign n26901 = ~n1354 & n26900 ;
  assign n26902 = ~n16903 & n26901 ;
  assign n26903 = ( n11386 & n21571 ) | ( n11386 & ~n26902 ) | ( n21571 & ~n26902 ) ;
  assign n26904 = n5953 ^ n4847 ^ n4690 ;
  assign n26905 = n21312 ^ n14348 ^ 1'b0 ;
  assign n26906 = n26904 & ~n26905 ;
  assign n26908 = n5984 | n12510 ;
  assign n26909 = n26908 ^ n3782 ^ 1'b0 ;
  assign n26910 = n26909 ^ n21629 ^ n9448 ;
  assign n26907 = ~n4145 & n6674 ;
  assign n26911 = n26910 ^ n26907 ^ 1'b0 ;
  assign n26912 = n16346 & n26911 ;
  assign n26913 = n26912 ^ n19326 ^ 1'b0 ;
  assign n26916 = n5320 | n6976 ;
  assign n26917 = n26916 ^ n3590 ^ 1'b0 ;
  assign n26918 = n26917 ^ n20247 ^ n12699 ;
  assign n26914 = n25981 ^ n22511 ^ n3751 ;
  assign n26915 = ~n12102 & n26914 ;
  assign n26919 = n26918 ^ n26915 ^ 1'b0 ;
  assign n26920 = ~n13199 & n15922 ;
  assign n26921 = ~n7756 & n26920 ;
  assign n26922 = n1067 & n23591 ;
  assign n26923 = n8972 & n26922 ;
  assign n26924 = ( n15984 & n19339 ) | ( n15984 & ~n26923 ) | ( n19339 & ~n26923 ) ;
  assign n26925 = n11404 ^ n4405 ^ 1'b0 ;
  assign n26926 = ( n8225 & ~n22091 ) | ( n8225 & n26925 ) | ( ~n22091 & n26925 ) ;
  assign n26927 = ( n3738 & n6564 ) | ( n3738 & n14509 ) | ( n6564 & n14509 ) ;
  assign n26928 = ( n9324 & n21319 ) | ( n9324 & n26927 ) | ( n21319 & n26927 ) ;
  assign n26929 = n6557 | n13705 ;
  assign n26930 = n4087 & ~n26929 ;
  assign n26931 = n26930 ^ n16053 ^ n15355 ;
  assign n26932 = n9696 | n12054 ;
  assign n26933 = n26932 ^ n7121 ^ 1'b0 ;
  assign n26934 = n26933 ^ n24054 ^ n20247 ;
  assign n26935 = n17252 ^ n5227 ^ 1'b0 ;
  assign n26936 = n4492 | n26935 ;
  assign n26937 = n656 & ~n7600 ;
  assign n26938 = n26056 & n26937 ;
  assign n26939 = n23476 & ~n23595 ;
  assign n26941 = n10801 ^ n1940 ^ n1449 ;
  assign n26942 = x108 & n26941 ;
  assign n26940 = n3177 & n12680 ;
  assign n26943 = n26942 ^ n26940 ^ 1'b0 ;
  assign n26944 = ~n2511 & n4140 ;
  assign n26945 = n7956 & n26944 ;
  assign n26946 = n5580 ^ n1096 ^ 1'b0 ;
  assign n26947 = ( n23686 & n26945 ) | ( n23686 & n26946 ) | ( n26945 & n26946 ) ;
  assign n26948 = n8621 | n18198 ;
  assign n26949 = n15290 | n26948 ;
  assign n26950 = n26949 ^ n934 ^ 1'b0 ;
  assign n26951 = n8253 | n26950 ;
  assign n26952 = n6480 & ~n9008 ;
  assign n26953 = n5522 & n19177 ;
  assign n26954 = ( ~n511 & n26952 ) | ( ~n511 & n26953 ) | ( n26952 & n26953 ) ;
  assign n26955 = ( n8808 & n26951 ) | ( n8808 & n26954 ) | ( n26951 & n26954 ) ;
  assign n26956 = ( n1019 & n16607 ) | ( n1019 & ~n20048 ) | ( n16607 & ~n20048 ) ;
  assign n26957 = n10411 ^ n4414 ^ 1'b0 ;
  assign n26958 = n9350 & n26957 ;
  assign n26959 = ( n4852 & n23643 ) | ( n4852 & ~n26958 ) | ( n23643 & ~n26958 ) ;
  assign n26960 = n3596 & n18951 ;
  assign n26961 = n26960 ^ n22483 ^ n3885 ;
  assign n26962 = n20989 | n21814 ;
  assign n26963 = n24143 ^ n141 ^ 1'b0 ;
  assign n26964 = ( n2857 & n7102 ) | ( n2857 & n8396 ) | ( n7102 & n8396 ) ;
  assign n26965 = ( n681 & n6482 ) | ( n681 & n26964 ) | ( n6482 & n26964 ) ;
  assign n26966 = n934 & n26965 ;
  assign n26967 = n689 & ~n13749 ;
  assign n26968 = n26967 ^ n17884 ^ 1'b0 ;
  assign n26969 = n26968 ^ n24540 ^ 1'b0 ;
  assign n26970 = n8597 & ~n20095 ;
  assign n26971 = ( n13974 & ~n16241 ) | ( n13974 & n22151 ) | ( ~n16241 & n22151 ) ;
  assign n26972 = ( n5238 & ~n18915 ) | ( n5238 & n26971 ) | ( ~n18915 & n26971 ) ;
  assign n26973 = n5674 ^ n2543 ^ 1'b0 ;
  assign n26974 = ( ~n8361 & n12003 ) | ( ~n8361 & n25372 ) | ( n12003 & n25372 ) ;
  assign n26975 = n16997 & n26974 ;
  assign n26976 = n5993 & n26975 ;
  assign n26977 = n6161 ^ n4508 ^ 1'b0 ;
  assign n26978 = ( ~n897 & n4057 ) | ( ~n897 & n7076 ) | ( n4057 & n7076 ) ;
  assign n26979 = n6371 & ~n26978 ;
  assign n26980 = ~n4339 & n26979 ;
  assign n26981 = n8436 | n24313 ;
  assign n26982 = n10495 | n20633 ;
  assign n26983 = n22064 ^ n19780 ^ 1'b0 ;
  assign n26984 = ~n15183 & n24942 ;
  assign n26985 = n24057 & ~n26984 ;
  assign n26986 = ( n6125 & ~n12890 ) | ( n6125 & n26985 ) | ( ~n12890 & n26985 ) ;
  assign n26987 = n12645 ^ n4497 ^ 1'b0 ;
  assign n26988 = n10838 & n26987 ;
  assign n26989 = ( n1385 & n23295 ) | ( n1385 & n26988 ) | ( n23295 & n26988 ) ;
  assign n26990 = n26989 ^ n22832 ^ 1'b0 ;
  assign n26991 = n6797 ^ n5282 ^ 1'b0 ;
  assign n26992 = n25645 ^ n9620 ^ n7725 ;
  assign n26993 = ~n10599 & n26992 ;
  assign n26994 = ( n6386 & n18005 ) | ( n6386 & n20633 ) | ( n18005 & n20633 ) ;
  assign n26995 = n26994 ^ n5345 ^ 1'b0 ;
  assign n26996 = n8584 & n26995 ;
  assign n26997 = x11 & n2894 ;
  assign n26998 = ~n3992 & n8230 ;
  assign n26999 = n26998 ^ n15645 ^ 1'b0 ;
  assign n27000 = ( n4253 & ~n26997 ) | ( n4253 & n26999 ) | ( ~n26997 & n26999 ) ;
  assign n27001 = n10284 & n27000 ;
  assign n27002 = n25534 ^ n25217 ^ n15026 ;
  assign n27003 = n13540 ^ n2665 ^ 1'b0 ;
  assign n27004 = n27002 & n27003 ;
  assign n27005 = ( n2329 & n4800 ) | ( n2329 & n12912 ) | ( n4800 & n12912 ) ;
  assign n27006 = ( n13431 & ~n22305 ) | ( n13431 & n27005 ) | ( ~n22305 & n27005 ) ;
  assign n27007 = n3154 & n3792 ;
  assign n27008 = n17944 & ~n18904 ;
  assign n27009 = n27007 & ~n27008 ;
  assign n27010 = n12490 ^ n11679 ^ n8318 ;
  assign n27011 = n10850 ^ n8643 ^ n1625 ;
  assign n27012 = ( n566 & n11628 ) | ( n566 & ~n27011 ) | ( n11628 & ~n27011 ) ;
  assign n27013 = ~n5115 & n9962 ;
  assign n27014 = n27013 ^ n14035 ^ 1'b0 ;
  assign n27015 = n23074 ^ n15586 ^ 1'b0 ;
  assign n27016 = n3152 & ~n27015 ;
  assign n27017 = n10176 ^ n6780 ^ 1'b0 ;
  assign n27018 = n10036 & ~n27017 ;
  assign n27021 = ~n3468 & n6316 ;
  assign n27019 = n11275 ^ n10388 ^ 1'b0 ;
  assign n27020 = n27019 ^ n13837 ^ 1'b0 ;
  assign n27022 = n27021 ^ n27020 ^ n6534 ;
  assign n27023 = ( ~n9254 & n9921 ) | ( ~n9254 & n15804 ) | ( n9921 & n15804 ) ;
  assign n27024 = n22524 ^ n1032 ^ 1'b0 ;
  assign n27025 = n12356 ^ n11356 ^ n6551 ;
  assign n27026 = n4135 & n13940 ;
  assign n27027 = ~n27025 & n27026 ;
  assign n27028 = ( n10715 & n21540 ) | ( n10715 & n27027 ) | ( n21540 & n27027 ) ;
  assign n27029 = ~n1088 & n9383 ;
  assign n27030 = ~n18511 & n27029 ;
  assign n27031 = n1467 | n11260 ;
  assign n27032 = n6366 & ~n27031 ;
  assign n27033 = n3576 & ~n21748 ;
  assign n27034 = ~n6581 & n27033 ;
  assign n27035 = ( n5753 & ~n6674 ) | ( n5753 & n15936 ) | ( ~n6674 & n15936 ) ;
  assign n27036 = n15816 & n27035 ;
  assign n27038 = n20356 ^ n18756 ^ n4304 ;
  assign n27037 = ( n5262 & n7409 ) | ( n5262 & n21040 ) | ( n7409 & n21040 ) ;
  assign n27039 = n27038 ^ n27037 ^ n8352 ;
  assign n27040 = n6022 & ~n10923 ;
  assign n27041 = n16191 | n27040 ;
  assign n27042 = n27041 ^ n15585 ^ n15079 ;
  assign n27044 = ~n10190 & n11002 ;
  assign n27045 = n25206 & n27044 ;
  assign n27043 = n4874 & ~n15385 ;
  assign n27046 = n27045 ^ n27043 ^ 1'b0 ;
  assign n27047 = n27046 ^ n9714 ^ n1986 ;
  assign n27048 = ( n1435 & n4608 ) | ( n1435 & n19227 ) | ( n4608 & n19227 ) ;
  assign n27049 = ( ~n6436 & n17008 ) | ( ~n6436 & n19028 ) | ( n17008 & n19028 ) ;
  assign n27050 = n2662 | n5728 ;
  assign n27051 = n27050 ^ n12866 ^ 1'b0 ;
  assign n27052 = n983 & n4465 ;
  assign n27053 = ~n25835 & n27052 ;
  assign n27054 = n5218 & ~n14965 ;
  assign n27055 = n27054 ^ n13698 ^ 1'b0 ;
  assign n27056 = n27055 ^ n15912 ^ 1'b0 ;
  assign n27057 = n27053 | n27056 ;
  assign n27058 = n23768 ^ n15075 ^ 1'b0 ;
  assign n27059 = n14912 ^ n3828 ^ 1'b0 ;
  assign n27060 = n9951 ^ n3913 ^ n668 ;
  assign n27061 = ~n12035 & n12404 ;
  assign n27062 = n2110 & n6268 ;
  assign n27063 = n26615 | n27062 ;
  assign n27065 = n3357 ^ n2224 ^ 1'b0 ;
  assign n27066 = ~n12183 & n27065 ;
  assign n27067 = ( n4334 & n7565 ) | ( n4334 & ~n27066 ) | ( n7565 & ~n27066 ) ;
  assign n27068 = n27067 ^ n23718 ^ n12260 ;
  assign n27064 = ~n9971 & n13479 ;
  assign n27069 = n27068 ^ n27064 ^ n11869 ;
  assign n27070 = ~n3488 & n10754 ;
  assign n27071 = n10929 & n27070 ;
  assign n27074 = n12335 ^ n357 ^ 1'b0 ;
  assign n27072 = n16673 ^ n2165 ^ n1862 ;
  assign n27073 = ~n13696 & n27072 ;
  assign n27075 = n27074 ^ n27073 ^ 1'b0 ;
  assign n27076 = ~n6926 & n9806 ;
  assign n27077 = n27076 ^ n3754 ^ 1'b0 ;
  assign n27078 = n21341 ^ n11196 ^ 1'b0 ;
  assign n27079 = ( n7810 & ~n21218 ) | ( n7810 & n26776 ) | ( ~n21218 & n26776 ) ;
  assign n27080 = ~n2631 & n7978 ;
  assign n27081 = n27080 ^ n804 ^ 1'b0 ;
  assign n27082 = ~n24982 & n27081 ;
  assign n27083 = ( n2417 & n21551 ) | ( n2417 & n27082 ) | ( n21551 & n27082 ) ;
  assign n27084 = n15565 ^ n11455 ^ n5635 ;
  assign n27085 = n202 & n27084 ;
  assign n27086 = n27085 ^ n7792 ^ 1'b0 ;
  assign n27087 = ~n13124 & n21611 ;
  assign n27088 = ~n8970 & n27087 ;
  assign n27089 = n1295 & n8955 ;
  assign n27090 = ~n19912 & n27089 ;
  assign n27091 = n13928 ^ n7361 ^ 1'b0 ;
  assign n27092 = n2610 & ~n27091 ;
  assign n27093 = ( n7786 & n11994 ) | ( n7786 & ~n27092 ) | ( n11994 & ~n27092 ) ;
  assign n27094 = n9770 ^ n993 ^ 1'b0 ;
  assign n27095 = n27093 | n27094 ;
  assign n27096 = n16410 ^ n1612 ^ 1'b0 ;
  assign n27097 = ~n27095 & n27096 ;
  assign n27098 = ( ~n3888 & n12864 ) | ( ~n3888 & n21017 ) | ( n12864 & n21017 ) ;
  assign n27099 = n27098 ^ n15236 ^ n5993 ;
  assign n27100 = n10637 ^ n7578 ^ n5417 ;
  assign n27101 = ~n24239 & n25790 ;
  assign n27102 = n17432 & ~n27101 ;
  assign n27103 = n27100 & n27102 ;
  assign n27104 = n24986 ^ n5044 ^ 1'b0 ;
  assign n27105 = n23344 ^ n9368 ^ 1'b0 ;
  assign n27106 = n27105 ^ n13212 ^ 1'b0 ;
  assign n27107 = ~n19825 & n27106 ;
  assign n27108 = n6910 & n27107 ;
  assign n27109 = n7621 ^ n3406 ^ 1'b0 ;
  assign n27112 = n488 & n3001 ;
  assign n27113 = n562 & n27112 ;
  assign n27114 = n16983 | n27113 ;
  assign n27110 = n10755 ^ n8320 ^ 1'b0 ;
  assign n27111 = n9691 | n27110 ;
  assign n27115 = n27114 ^ n27111 ^ n6492 ;
  assign n27117 = n2744 & n12889 ;
  assign n27118 = n5170 & n27117 ;
  assign n27116 = n25074 ^ n14914 ^ n13123 ;
  assign n27119 = n27118 ^ n27116 ^ 1'b0 ;
  assign n27120 = ~n5201 & n27119 ;
  assign n27121 = n27120 ^ n22214 ^ 1'b0 ;
  assign n27122 = n12063 ^ n9273 ^ 1'b0 ;
  assign n27123 = ~n22356 & n27122 ;
  assign n27126 = n20113 ^ n2824 ^ 1'b0 ;
  assign n27124 = x33 & x113 ;
  assign n27125 = n27124 ^ n3836 ^ 1'b0 ;
  assign n27127 = n27126 ^ n27125 ^ n11621 ;
  assign n27128 = n23997 ^ n8512 ^ n337 ;
  assign n27129 = n6059 | n12250 ;
  assign n27130 = n27129 ^ n10886 ^ 1'b0 ;
  assign n27131 = n27130 ^ n20394 ^ n8742 ;
  assign n27132 = n3192 & n11032 ;
  assign n27133 = n16982 & n27132 ;
  assign n27134 = ( ~n2858 & n24161 ) | ( ~n2858 & n24712 ) | ( n24161 & n24712 ) ;
  assign n27135 = ( n1024 & n27133 ) | ( n1024 & ~n27134 ) | ( n27133 & ~n27134 ) ;
  assign n27136 = n7798 & n27135 ;
  assign n27137 = n9104 | n10751 ;
  assign n27138 = ( x48 & n895 ) | ( x48 & n13573 ) | ( n895 & n13573 ) ;
  assign n27139 = n5228 | n27138 ;
  assign n27140 = n2430 & n23200 ;
  assign n27141 = n12427 | n15902 ;
  assign n27142 = n3841 & ~n16987 ;
  assign n27143 = n27142 ^ n5454 ^ 1'b0 ;
  assign n27144 = n21333 & ~n27143 ;
  assign n27145 = n27144 ^ n23650 ^ 1'b0 ;
  assign n27146 = n27145 ^ n11503 ^ n10398 ;
  assign n27147 = n9534 ^ n8532 ^ n3489 ;
  assign n27148 = n27147 ^ n2207 ^ 1'b0 ;
  assign n27149 = n3134 | n7955 ;
  assign n27150 = n27149 ^ n26407 ^ 1'b0 ;
  assign n27151 = n27150 ^ n25502 ^ 1'b0 ;
  assign n27152 = n8922 ^ n8669 ^ 1'b0 ;
  assign n27153 = n9061 | n20608 ;
  assign n27154 = n147 & ~n18061 ;
  assign n27155 = n27154 ^ n9039 ^ 1'b0 ;
  assign n27156 = n4131 | n20048 ;
  assign n27157 = n23506 ^ n13025 ^ 1'b0 ;
  assign n27158 = n6447 ^ n3349 ^ 1'b0 ;
  assign n27159 = n27158 ^ n23113 ^ n17250 ;
  assign n27161 = ~n672 & n5528 ;
  assign n27160 = n10412 ^ n2469 ^ 1'b0 ;
  assign n27162 = n27161 ^ n27160 ^ n6995 ;
  assign n27163 = n7627 | n8010 ;
  assign n27164 = n27162 | n27163 ;
  assign n27165 = ( n12333 & n13625 ) | ( n12333 & n27164 ) | ( n13625 & n27164 ) ;
  assign n27166 = n2639 & n20142 ;
  assign n27167 = n27166 ^ n15632 ^ 1'b0 ;
  assign n27168 = ~n479 & n27167 ;
  assign n27169 = n21560 & n27168 ;
  assign n27170 = n27169 ^ n5247 ^ 1'b0 ;
  assign n27171 = ( n8536 & n13144 ) | ( n8536 & n20322 ) | ( n13144 & n20322 ) ;
  assign n27172 = n7271 ^ n1404 ^ n866 ;
  assign n27173 = n4688 ^ n2331 ^ 1'b0 ;
  assign n27174 = n27172 | n27173 ;
  assign n27175 = n11599 ^ n11469 ^ n6999 ;
  assign n27176 = ( n6966 & n12151 ) | ( n6966 & ~n27175 ) | ( n12151 & ~n27175 ) ;
  assign n27177 = n27176 ^ n6410 ^ 1'b0 ;
  assign n27178 = n6520 | n15700 ;
  assign n27179 = x41 | n27178 ;
  assign n27180 = n2626 ^ n1738 ^ n1339 ;
  assign n27181 = n1646 & n27180 ;
  assign n27182 = n22586 & n27181 ;
  assign n27183 = n27182 ^ n11606 ^ 1'b0 ;
  assign n27184 = n3504 | n11334 ;
  assign n27185 = n2486 & n15387 ;
  assign n27186 = n19249 & n27185 ;
  assign n27187 = n27186 ^ n10770 ^ n6288 ;
  assign n27188 = n13871 ^ n12750 ^ 1'b0 ;
  assign n27189 = n21704 & n27188 ;
  assign n27190 = n27189 ^ n22724 ^ 1'b0 ;
  assign n27191 = ~n3416 & n7188 ;
  assign n27192 = n27191 ^ n15910 ^ n2459 ;
  assign n27193 = n9848 & n17249 ;
  assign n27194 = ( n7503 & n27192 ) | ( n7503 & ~n27193 ) | ( n27192 & ~n27193 ) ;
  assign n27195 = n9944 & n26909 ;
  assign n27196 = ~n21576 & n27195 ;
  assign n27197 = n1760 | n23116 ;
  assign n27198 = n27197 ^ n2421 ^ 1'b0 ;
  assign n27199 = n6480 ^ n1855 ^ 1'b0 ;
  assign n27200 = n27198 & n27199 ;
  assign n27201 = n7669 & ~n18336 ;
  assign n27202 = n27201 ^ n21163 ^ 1'b0 ;
  assign n27203 = n18136 & ~n25275 ;
  assign n27204 = n8392 ^ n2304 ^ 1'b0 ;
  assign n27205 = ( n2592 & n22537 ) | ( n2592 & n27204 ) | ( n22537 & n27204 ) ;
  assign n27206 = ~n2372 & n26699 ;
  assign n27207 = n27206 ^ n2959 ^ 1'b0 ;
  assign n27208 = ( ~n6859 & n7551 ) | ( ~n6859 & n27207 ) | ( n7551 & n27207 ) ;
  assign n27209 = n11229 ^ n2369 ^ 1'b0 ;
  assign n27210 = n14846 & n27209 ;
  assign n27211 = n1205 | n17912 ;
  assign n27212 = n14251 | n27211 ;
  assign n27213 = n23736 ^ n20048 ^ 1'b0 ;
  assign n27214 = n8572 | n27213 ;
  assign n27215 = n689 | n21778 ;
  assign n27216 = n27215 ^ n22999 ^ 1'b0 ;
  assign n27217 = n5362 & ~n11833 ;
  assign n27218 = n27217 ^ n17804 ^ 1'b0 ;
  assign n27219 = ( n4765 & n11587 ) | ( n4765 & n27218 ) | ( n11587 & n27218 ) ;
  assign n27220 = n27219 ^ n18601 ^ n6614 ;
  assign n27224 = n11114 ^ n307 ^ x116 ;
  assign n27221 = ~n1212 & n23684 ;
  assign n27222 = n5351 | n6163 ;
  assign n27223 = n27221 | n27222 ;
  assign n27225 = n27224 ^ n27223 ^ n8564 ;
  assign n27226 = n23756 ^ n18587 ^ 1'b0 ;
  assign n27227 = n18638 & ~n27226 ;
  assign n27228 = ( n13738 & n27225 ) | ( n13738 & ~n27227 ) | ( n27225 & ~n27227 ) ;
  assign n27229 = n22379 ^ n16818 ^ n16183 ;
  assign n27230 = ( n1739 & n17837 ) | ( n1739 & ~n27229 ) | ( n17837 & ~n27229 ) ;
  assign n27236 = n3811 & n5332 ;
  assign n27237 = n27236 ^ n2389 ^ 1'b0 ;
  assign n27238 = n27237 ^ n3162 ^ 1'b0 ;
  assign n27233 = n18441 ^ n16948 ^ 1'b0 ;
  assign n27234 = n3845 & ~n27233 ;
  assign n27235 = ~n7923 & n27234 ;
  assign n27231 = n683 ^ n192 ^ 1'b0 ;
  assign n27232 = ~n14447 & n27231 ;
  assign n27239 = n27238 ^ n27235 ^ n27232 ;
  assign n27240 = ( n248 & ~n6452 ) | ( n248 & n10866 ) | ( ~n6452 & n10866 ) ;
  assign n27241 = n14531 | n22023 ;
  assign n27242 = n27241 ^ n4588 ^ 1'b0 ;
  assign n27243 = ~n3547 & n6838 ;
  assign n27244 = n27243 ^ n7254 ^ 1'b0 ;
  assign n27245 = n27244 ^ n24313 ^ 1'b0 ;
  assign n27246 = n27242 | n27245 ;
  assign n27247 = n19300 ^ n17629 ^ 1'b0 ;
  assign n27248 = ~n5040 & n27247 ;
  assign n27249 = n15355 & n27248 ;
  assign n27250 = n27249 ^ n2010 ^ 1'b0 ;
  assign n27251 = ( n10018 & ~n10934 ) | ( n10018 & n16514 ) | ( ~n10934 & n16514 ) ;
  assign n27252 = n5609 ^ n4765 ^ 1'b0 ;
  assign n27253 = n27251 & n27252 ;
  assign n27254 = n23165 & ~n27253 ;
  assign n27255 = n3223 & ~n6480 ;
  assign n27256 = n1509 | n27255 ;
  assign n27257 = n27256 ^ n1683 ^ 1'b0 ;
  assign n27258 = n1426 & ~n14172 ;
  assign n27259 = n27258 ^ n7033 ^ 1'b0 ;
  assign n27260 = n1083 & n1673 ;
  assign n27261 = n27260 ^ n6394 ^ 1'b0 ;
  assign n27262 = n17974 ^ n10908 ^ n8087 ;
  assign n27263 = ( n4033 & n6413 ) | ( n4033 & ~n11849 ) | ( n6413 & ~n11849 ) ;
  assign n27264 = n11210 & ~n27263 ;
  assign n27265 = n17067 ^ n4949 ^ 1'b0 ;
  assign n27266 = ~n23135 & n27265 ;
  assign n27267 = ( n22960 & ~n24461 ) | ( n22960 & n27266 ) | ( ~n24461 & n27266 ) ;
  assign n27268 = n26724 ^ n6621 ^ 1'b0 ;
  assign n27269 = n4006 | n22510 ;
  assign n27270 = n27269 ^ n13166 ^ 1'b0 ;
  assign n27271 = n7228 ^ n1927 ^ n260 ;
  assign n27272 = ( n3803 & n10049 ) | ( n3803 & n27271 ) | ( n10049 & n27271 ) ;
  assign n27273 = ( n3206 & n27270 ) | ( n3206 & n27272 ) | ( n27270 & n27272 ) ;
  assign n27274 = ( n22426 & n26573 ) | ( n22426 & n27273 ) | ( n26573 & n27273 ) ;
  assign n27275 = n5384 & ~n22433 ;
  assign n27276 = ~n3479 & n4628 ;
  assign n27277 = n27276 ^ n25726 ^ n25655 ;
  assign n27278 = ~n24299 & n27277 ;
  assign n27279 = n3084 ^ n481 ^ 1'b0 ;
  assign n27280 = n8763 ^ n7375 ^ 1'b0 ;
  assign n27281 = n1455 & n6733 ;
  assign n27282 = n9539 ^ n5131 ^ 1'b0 ;
  assign n27283 = n3763 & ~n27282 ;
  assign n27284 = ( n14721 & n27281 ) | ( n14721 & ~n27283 ) | ( n27281 & ~n27283 ) ;
  assign n27285 = n27280 & n27284 ;
  assign n27287 = n13219 ^ n10219 ^ n8156 ;
  assign n27286 = n3715 ^ n3692 ^ 1'b0 ;
  assign n27288 = n27287 ^ n27286 ^ n9607 ;
  assign n27289 = n27288 ^ n13696 ^ n6032 ;
  assign n27290 = n20030 ^ n4060 ^ 1'b0 ;
  assign n27291 = ~n10953 & n14872 ;
  assign n27292 = ~n1653 & n27291 ;
  assign n27293 = ( ~n993 & n27290 ) | ( ~n993 & n27292 ) | ( n27290 & n27292 ) ;
  assign n27294 = ( n2340 & n11815 ) | ( n2340 & n27293 ) | ( n11815 & n27293 ) ;
  assign n27295 = n10883 & n20121 ;
  assign n27296 = n10225 & ~n27281 ;
  assign n27297 = ~n24033 & n27296 ;
  assign n27298 = n11578 ^ n7897 ^ x17 ;
  assign n27299 = n9855 & n27298 ;
  assign n27300 = n27299 ^ n11868 ^ 1'b0 ;
  assign n27301 = n27300 ^ n19033 ^ 1'b0 ;
  assign n27302 = n3496 | n27301 ;
  assign n27303 = n18766 | n18916 ;
  assign n27304 = n27303 ^ n934 ^ 1'b0 ;
  assign n27306 = n4265 & n14350 ;
  assign n27305 = n14474 | n23837 ;
  assign n27307 = n27306 ^ n27305 ^ n15707 ;
  assign n27308 = n14605 ^ n8626 ^ 1'b0 ;
  assign n27309 = n6419 | n12973 ;
  assign n27310 = n15741 | n27309 ;
  assign n27311 = n27310 ^ n19066 ^ 1'b0 ;
  assign n27312 = ( n5109 & n18095 ) | ( n5109 & n21266 ) | ( n18095 & n21266 ) ;
  assign n27313 = n2865 | n14149 ;
  assign n27314 = n2865 & ~n27313 ;
  assign n27315 = n27314 ^ n21240 ^ 1'b0 ;
  assign n27316 = ~n4313 & n27315 ;
  assign n27317 = ~n12517 & n27316 ;
  assign n27318 = n27317 ^ n24922 ^ 1'b0 ;
  assign n27319 = n9842 ^ n976 ^ n523 ;
  assign n27320 = n27319 ^ n10708 ^ 1'b0 ;
  assign n27321 = n19527 | n27320 ;
  assign n27322 = n9440 & ~n9521 ;
  assign n27323 = ~n469 & n27322 ;
  assign n27324 = x125 & ~n22788 ;
  assign n27325 = n27324 ^ n3230 ^ 1'b0 ;
  assign n27326 = n27323 | n27325 ;
  assign n27327 = n7204 | n21439 ;
  assign n27328 = ~n27326 & n27327 ;
  assign n27329 = n27321 & n27328 ;
  assign n27330 = n7384 | n10528 ;
  assign n27331 = n20735 ^ n7143 ^ 1'b0 ;
  assign n27332 = n7375 | n27331 ;
  assign n27333 = n27332 ^ n21547 ^ 1'b0 ;
  assign n27334 = n25453 | n27333 ;
  assign n27335 = n1352 | n2335 ;
  assign n27336 = n27335 ^ n2199 ^ 1'b0 ;
  assign n27337 = n27336 ^ n11931 ^ n2561 ;
  assign n27338 = ~n1250 & n1264 ;
  assign n27339 = ~n368 & n27338 ;
  assign n27340 = n19419 ^ n3105 ^ 1'b0 ;
  assign n27341 = n10785 & n27340 ;
  assign n27342 = ( ~n3965 & n27339 ) | ( ~n3965 & n27341 ) | ( n27339 & n27341 ) ;
  assign n27343 = ( ~n1096 & n17167 ) | ( ~n1096 & n27342 ) | ( n17167 & n27342 ) ;
  assign n27344 = n9594 | n12896 ;
  assign n27345 = n27344 ^ n13673 ^ n1666 ;
  assign n27346 = n27343 & ~n27345 ;
  assign n27347 = ( ~n19444 & n27337 ) | ( ~n19444 & n27346 ) | ( n27337 & n27346 ) ;
  assign n27349 = ~n8043 & n9229 ;
  assign n27348 = n24982 ^ n19935 ^ n4438 ;
  assign n27350 = n27349 ^ n27348 ^ 1'b0 ;
  assign n27351 = ( n5336 & ~n15151 ) | ( n5336 & n26578 ) | ( ~n15151 & n26578 ) ;
  assign n27352 = n27351 ^ n17186 ^ 1'b0 ;
  assign n27353 = n2409 | n14700 ;
  assign n27354 = n27353 ^ n15369 ^ n9364 ;
  assign n27356 = n2732 & ~n10839 ;
  assign n27357 = n27356 ^ n15993 ^ 1'b0 ;
  assign n27355 = n3777 & n4834 ;
  assign n27358 = n27357 ^ n27355 ^ n27162 ;
  assign n27359 = ~n15568 & n27358 ;
  assign n27360 = n597 | n3481 ;
  assign n27361 = ~n4062 & n27360 ;
  assign n27362 = n349 & n27361 ;
  assign n27363 = n10989 & ~n27362 ;
  assign n27364 = n27363 ^ n1543 ^ 1'b0 ;
  assign n27365 = n17846 | n27364 ;
  assign n27366 = n3295 & n14266 ;
  assign n27367 = n19665 ^ n296 ^ 1'b0 ;
  assign n27368 = n20268 ^ n7239 ^ 1'b0 ;
  assign n27369 = n27368 ^ n14691 ^ n5295 ;
  assign n27370 = n987 & n16840 ;
  assign n27371 = n27370 ^ n26472 ^ 1'b0 ;
  assign n27372 = n22854 & ~n27371 ;
  assign n27373 = ~n9725 & n16735 ;
  assign n27374 = ~n16735 & n27373 ;
  assign n27375 = ( n2086 & n4466 ) | ( n2086 & ~n27374 ) | ( n4466 & ~n27374 ) ;
  assign n27376 = ~n8650 & n27375 ;
  assign n27377 = n21062 ^ n13281 ^ 1'b0 ;
  assign n27378 = n4329 & n25157 ;
  assign n27379 = n27378 ^ n4644 ^ 1'b0 ;
  assign n27380 = ( ~n10586 & n12704 ) | ( ~n10586 & n12983 ) | ( n12704 & n12983 ) ;
  assign n27381 = n9931 ^ n7712 ^ 1'b0 ;
  assign n27382 = ~n27380 & n27381 ;
  assign n27383 = ( ~n1022 & n6273 ) | ( ~n1022 & n9272 ) | ( n6273 & n9272 ) ;
  assign n27384 = n15432 ^ n3766 ^ 1'b0 ;
  assign n27385 = n27383 & n27384 ;
  assign n27386 = n9925 & ~n10854 ;
  assign n27387 = n27386 ^ n9047 ^ 1'b0 ;
  assign n27388 = ( n17078 & n21438 ) | ( n17078 & n27387 ) | ( n21438 & n27387 ) ;
  assign n27389 = n8575 & ~n15797 ;
  assign n27390 = n4628 & n27389 ;
  assign n27391 = n27390 ^ n24254 ^ 1'b0 ;
  assign n27392 = n9955 ^ n7026 ^ n5270 ;
  assign n27393 = ( n4165 & ~n12879 ) | ( n4165 & n27392 ) | ( ~n12879 & n27392 ) ;
  assign n27394 = ( n1182 & ~n3340 ) | ( n1182 & n15086 ) | ( ~n3340 & n15086 ) ;
  assign n27395 = n701 & ~n4739 ;
  assign n27396 = ( n13792 & n24014 ) | ( n13792 & n27395 ) | ( n24014 & n27395 ) ;
  assign n27397 = ( n27393 & n27394 ) | ( n27393 & n27396 ) | ( n27394 & n27396 ) ;
  assign n27398 = ( n15940 & ~n16856 ) | ( n15940 & n20352 ) | ( ~n16856 & n20352 ) ;
  assign n27399 = n8017 ^ n3215 ^ 1'b0 ;
  assign n27400 = ( n14829 & n16941 ) | ( n14829 & ~n27399 ) | ( n16941 & ~n27399 ) ;
  assign n27401 = n8593 & n27400 ;
  assign n27402 = ( ~n618 & n3181 ) | ( ~n618 & n15723 ) | ( n3181 & n15723 ) ;
  assign n27403 = n19114 & ~n27402 ;
  assign n27404 = ~n24147 & n27403 ;
  assign n27405 = n3067 & n11229 ;
  assign n27406 = ~n1213 & n15047 ;
  assign n27407 = n8253 ^ n3668 ^ n2350 ;
  assign n27408 = n27407 ^ n901 ^ 1'b0 ;
  assign n27409 = ( ~n18061 & n20965 ) | ( ~n18061 & n21460 ) | ( n20965 & n21460 ) ;
  assign n27410 = ( n1579 & n24405 ) | ( n1579 & n27409 ) | ( n24405 & n27409 ) ;
  assign n27411 = ~x76 & n15985 ;
  assign n27412 = ( ~n4884 & n17034 ) | ( ~n4884 & n27411 ) | ( n17034 & n27411 ) ;
  assign n27413 = n4399 ^ n601 ^ 1'b0 ;
  assign n27414 = ~n25055 & n27413 ;
  assign n27415 = n16931 & n21161 ;
  assign n27416 = n18492 ^ n15221 ^ 1'b0 ;
  assign n27418 = n12198 ^ n2165 ^ n694 ;
  assign n27417 = ~n5057 & n23549 ;
  assign n27419 = n27418 ^ n27417 ^ 1'b0 ;
  assign n27420 = n7227 & n18055 ;
  assign n27421 = n27420 ^ n2593 ^ 1'b0 ;
  assign n27422 = n4808 & ~n7430 ;
  assign n27423 = n10835 ^ n1740 ^ 1'b0 ;
  assign n27424 = n13198 & ~n27423 ;
  assign n27425 = n11769 & n27424 ;
  assign n27426 = n17646 & n27425 ;
  assign n27427 = ( n5076 & n9674 ) | ( n5076 & ~n27426 ) | ( n9674 & ~n27426 ) ;
  assign n27428 = n8721 ^ n8480 ^ 1'b0 ;
  assign n27429 = ~n26338 & n27428 ;
  assign n27430 = n8133 ^ n3854 ^ 1'b0 ;
  assign n27431 = ( ~n2626 & n27429 ) | ( ~n2626 & n27430 ) | ( n27429 & n27430 ) ;
  assign n27433 = ( ~n1162 & n3897 ) | ( ~n1162 & n16509 ) | ( n3897 & n16509 ) ;
  assign n27432 = n15922 ^ n755 ^ 1'b0 ;
  assign n27434 = n27433 ^ n27432 ^ n1326 ;
  assign n27435 = n20797 ^ n13110 ^ 1'b0 ;
  assign n27436 = n4680 | n27435 ;
  assign n27437 = ( ~n3015 & n19322 ) | ( ~n3015 & n27436 ) | ( n19322 & n27436 ) ;
  assign n27438 = n27437 ^ n6129 ^ 1'b0 ;
  assign n27439 = n27438 ^ n23431 ^ 1'b0 ;
  assign n27440 = n2018 & ~n15486 ;
  assign n27441 = n27439 & n27440 ;
  assign n27442 = n1065 & ~n15788 ;
  assign n27443 = n22033 & ~n26405 ;
  assign n27444 = ~n8331 & n24539 ;
  assign n27445 = n9076 ^ n4461 ^ 1'b0 ;
  assign n27446 = ( n3235 & n27444 ) | ( n3235 & n27445 ) | ( n27444 & n27445 ) ;
  assign n27447 = n23933 ^ n18877 ^ n1783 ;
  assign n27448 = ( ~n3837 & n7199 ) | ( ~n3837 & n27447 ) | ( n7199 & n27447 ) ;
  assign n27450 = ( ~n6728 & n24589 ) | ( ~n6728 & n26675 ) | ( n24589 & n26675 ) ;
  assign n27449 = n2736 | n8191 ;
  assign n27451 = n27450 ^ n27449 ^ 1'b0 ;
  assign n27452 = ( ~n2631 & n4754 ) | ( ~n2631 & n27451 ) | ( n4754 & n27451 ) ;
  assign n27453 = n10516 ^ n4819 ^ 1'b0 ;
  assign n27454 = n27453 ^ n6261 ^ 1'b0 ;
  assign n27456 = n9309 | n9552 ;
  assign n27455 = n22664 ^ n12570 ^ n2139 ;
  assign n27457 = n27456 ^ n27455 ^ n12766 ;
  assign n27458 = n3656 & n23539 ;
  assign n27459 = n27458 ^ n21079 ^ 1'b0 ;
  assign n27460 = n27457 | n27459 ;
  assign n27461 = ( n3046 & n6287 ) | ( n3046 & ~n10903 ) | ( n6287 & ~n10903 ) ;
  assign n27462 = n9964 & ~n27461 ;
  assign n27463 = n4758 & ~n9366 ;
  assign n27464 = n15236 & ~n22025 ;
  assign n27465 = n27464 ^ n5753 ^ 1'b0 ;
  assign n27469 = n234 & n3816 ;
  assign n27466 = n908 | n8055 ;
  assign n27467 = n27466 ^ n7551 ^ 1'b0 ;
  assign n27468 = n18537 & ~n27467 ;
  assign n27470 = n27469 ^ n27468 ^ 1'b0 ;
  assign n27471 = n3688 & ~n15696 ;
  assign n27472 = n8583 & n27471 ;
  assign n27473 = n447 & n27472 ;
  assign n27474 = ( n11220 & n12338 ) | ( n11220 & n25507 ) | ( n12338 & n25507 ) ;
  assign n27475 = n23988 ^ n9944 ^ 1'b0 ;
  assign n27476 = ~n22096 & n27475 ;
  assign n27477 = n9151 & n27476 ;
  assign n27478 = n17773 | n21884 ;
  assign n27480 = ~n5512 & n5670 ;
  assign n27479 = n6674 & n15704 ;
  assign n27481 = n27480 ^ n27479 ^ n10453 ;
  assign n27482 = n2261 & ~n15881 ;
  assign n27483 = n3175 | n6370 ;
  assign n27484 = n27483 ^ n3929 ^ 1'b0 ;
  assign n27485 = n23142 & n27484 ;
  assign n27486 = n3301 & ~n6954 ;
  assign n27487 = n7124 & n27486 ;
  assign n27488 = n5831 ^ n3262 ^ 1'b0 ;
  assign n27489 = n23279 & n27488 ;
  assign n27490 = ( n8993 & ~n27487 ) | ( n8993 & n27489 ) | ( ~n27487 & n27489 ) ;
  assign n27491 = n2681 & n27490 ;
  assign n27493 = n9972 ^ n9913 ^ 1'b0 ;
  assign n27492 = n5526 | n9533 ;
  assign n27494 = n27493 ^ n27492 ^ 1'b0 ;
  assign n27495 = n9425 ^ n4432 ^ 1'b0 ;
  assign n27496 = ~n5965 & n27495 ;
  assign n27499 = n759 | n4964 ;
  assign n27500 = n27499 ^ n12140 ^ n7378 ;
  assign n27501 = ( n7531 & n16612 ) | ( n7531 & ~n27500 ) | ( n16612 & ~n27500 ) ;
  assign n27497 = n5149 | n18506 ;
  assign n27498 = n6175 & ~n27497 ;
  assign n27502 = n27501 ^ n27498 ^ n6623 ;
  assign n27505 = n1464 | n10929 ;
  assign n27506 = n27505 ^ n11930 ^ 1'b0 ;
  assign n27507 = n796 & n3848 ;
  assign n27508 = n3221 | n4260 ;
  assign n27509 = ~n27507 & n27508 ;
  assign n27510 = n27506 & n27509 ;
  assign n27503 = n8431 | n19617 ;
  assign n27504 = n27503 ^ n1837 ^ 1'b0 ;
  assign n27511 = n27510 ^ n27504 ^ n16150 ;
  assign n27513 = n13701 | n20716 ;
  assign n27514 = n2481 & ~n27513 ;
  assign n27512 = n22922 ^ n4628 ^ n3376 ;
  assign n27515 = n27514 ^ n27512 ^ 1'b0 ;
  assign n27519 = ~n7244 & n12750 ;
  assign n27517 = n11789 ^ n8990 ^ n6572 ;
  assign n27516 = n9637 & ~n16102 ;
  assign n27518 = n27517 ^ n27516 ^ 1'b0 ;
  assign n27520 = n27519 ^ n27518 ^ n1626 ;
  assign n27521 = n26203 ^ n6748 ^ n3274 ;
  assign n27522 = ~n14447 & n27521 ;
  assign n27523 = n3546 | n13078 ;
  assign n27524 = n27523 ^ n1184 ^ 1'b0 ;
  assign n27525 = n27522 | n27524 ;
  assign n27526 = n22726 ^ n1851 ^ 1'b0 ;
  assign n27527 = n3121 | n27526 ;
  assign n27528 = n26525 & ~n27527 ;
  assign n27529 = n11277 ^ n1845 ^ 1'b0 ;
  assign n27530 = ~n9748 & n11213 ;
  assign n27531 = ~n3619 & n27530 ;
  assign n27532 = n4543 & ~n27531 ;
  assign n27533 = n27532 ^ n1811 ^ 1'b0 ;
  assign n27534 = n19430 ^ n16188 ^ n7469 ;
  assign n27535 = n27534 ^ n24168 ^ 1'b0 ;
  assign n27536 = n11738 ^ n7783 ^ 1'b0 ;
  assign n27537 = ( ~n3640 & n5301 ) | ( ~n3640 & n27536 ) | ( n5301 & n27536 ) ;
  assign n27538 = ~n1063 & n14664 ;
  assign n27539 = n21384 & n27538 ;
  assign n27540 = n27539 ^ n18092 ^ 1'b0 ;
  assign n27541 = n26286 ^ n21625 ^ 1'b0 ;
  assign n27542 = n3290 & n21078 ;
  assign n27543 = n27542 ^ n845 ^ 1'b0 ;
  assign n27544 = ( n5122 & ~n7737 ) | ( n5122 & n27543 ) | ( ~n7737 & n27543 ) ;
  assign n27545 = n26079 ^ n17516 ^ n296 ;
  assign n27546 = ~n4964 & n10162 ;
  assign n27547 = n13810 & n27546 ;
  assign n27548 = n8187 | n27547 ;
  assign n27549 = n27548 ^ n25732 ^ 1'b0 ;
  assign n27550 = n17530 ^ n14594 ^ 1'b0 ;
  assign n27551 = n10584 & n27550 ;
  assign n27552 = n27551 ^ n20056 ^ n5753 ;
  assign n27553 = n2420 & n15287 ;
  assign n27554 = n4239 ^ n1634 ^ x84 ;
  assign n27558 = n9529 | n23084 ;
  assign n27559 = n27558 ^ n5384 ^ 1'b0 ;
  assign n27560 = n27559 ^ n25344 ^ n1053 ;
  assign n27555 = ~n2535 & n8361 ;
  assign n27556 = ~n877 & n27555 ;
  assign n27557 = ( ~n17284 & n21131 ) | ( ~n17284 & n27556 ) | ( n21131 & n27556 ) ;
  assign n27561 = n27560 ^ n27557 ^ n12104 ;
  assign n27562 = n2998 & ~n10373 ;
  assign n27563 = n10265 & n27562 ;
  assign n27564 = ~n16618 & n27563 ;
  assign n27565 = n5189 & ~n26061 ;
  assign n27566 = n7152 ^ n2483 ^ 1'b0 ;
  assign n27567 = n1040 & ~n27566 ;
  assign n27568 = n27567 ^ n18760 ^ 1'b0 ;
  assign n27569 = n10134 | n27568 ;
  assign n27570 = ( n9314 & ~n10372 ) | ( n9314 & n20965 ) | ( ~n10372 & n20965 ) ;
  assign n27571 = ( x27 & n291 ) | ( x27 & ~n15040 ) | ( n291 & ~n15040 ) ;
  assign n27572 = ( n12827 & n15514 ) | ( n12827 & ~n27571 ) | ( n15514 & ~n27571 ) ;
  assign n27573 = n20132 ^ n15022 ^ n13559 ;
  assign n27574 = n23534 ^ n5254 ^ 1'b0 ;
  assign n27575 = n22758 ^ n1338 ^ 1'b0 ;
  assign n27576 = ~n2697 & n27575 ;
  assign n27577 = ( n16576 & ~n27574 ) | ( n16576 & n27576 ) | ( ~n27574 & n27576 ) ;
  assign n27578 = n22347 ^ n2697 ^ 1'b0 ;
  assign n27579 = n6827 ^ n3550 ^ 1'b0 ;
  assign n27580 = n6498 & n27579 ;
  assign n27581 = n3240 & ~n3775 ;
  assign n27582 = n12519 | n27319 ;
  assign n27583 = n27582 ^ n1962 ^ 1'b0 ;
  assign n27584 = n6493 & ~n14812 ;
  assign n27585 = n27584 ^ n9607 ^ 1'b0 ;
  assign n27586 = n5086 | n13576 ;
  assign n27587 = n27586 ^ n13485 ^ 1'b0 ;
  assign n27588 = n26434 ^ n18509 ^ n219 ;
  assign n27589 = ( x120 & n2376 ) | ( x120 & n2508 ) | ( n2376 & n2508 ) ;
  assign n27590 = ( n12853 & ~n14757 ) | ( n12853 & n27589 ) | ( ~n14757 & n27589 ) ;
  assign n27591 = ( n6210 & n16657 ) | ( n6210 & ~n21062 ) | ( n16657 & ~n21062 ) ;
  assign n27592 = ~n14249 & n18842 ;
  assign n27593 = n23794 & n27592 ;
  assign n27594 = ( n2590 & n5068 ) | ( n2590 & ~n27453 ) | ( n5068 & ~n27453 ) ;
  assign n27595 = n27594 ^ n19954 ^ 1'b0 ;
  assign n27596 = n26822 & n27595 ;
  assign n27597 = n17561 & n27596 ;
  assign n27598 = n1816 & n22214 ;
  assign n27599 = ~n23349 & n27598 ;
  assign n27600 = n1911 | n3626 ;
  assign n27601 = n6082 | n27600 ;
  assign n27602 = n2589 & ~n7720 ;
  assign n27603 = ~n14670 & n27602 ;
  assign n27604 = n23238 ^ n8825 ^ n5510 ;
  assign n27607 = ( n328 & n3262 ) | ( n328 & ~n11253 ) | ( n3262 & ~n11253 ) ;
  assign n27605 = ( n2041 & n6214 ) | ( n2041 & ~n12823 ) | ( n6214 & ~n12823 ) ;
  assign n27606 = ( n14407 & n15892 ) | ( n14407 & ~n27605 ) | ( n15892 & ~n27605 ) ;
  assign n27608 = n27607 ^ n27606 ^ n15702 ;
  assign n27609 = n26240 ^ n10616 ^ 1'b0 ;
  assign n27613 = n5110 & ~n15962 ;
  assign n27614 = n27613 ^ n15400 ^ 1'b0 ;
  assign n27610 = ( n4582 & n13834 ) | ( n4582 & ~n16754 ) | ( n13834 & ~n16754 ) ;
  assign n27611 = n12864 & n26949 ;
  assign n27612 = n27610 & n27611 ;
  assign n27615 = n27614 ^ n27612 ^ 1'b0 ;
  assign n27616 = n23063 ^ n898 ^ 1'b0 ;
  assign n27617 = n19562 | n27616 ;
  assign n27618 = n11371 & ~n11471 ;
  assign n27619 = n27618 ^ n22040 ^ 1'b0 ;
  assign n27620 = n10283 ^ n7129 ^ 1'b0 ;
  assign n27621 = n728 & n27620 ;
  assign n27622 = ~n27609 & n27621 ;
  assign n27623 = ~n17537 & n18527 ;
  assign n27624 = n27623 ^ n6059 ^ 1'b0 ;
  assign n27625 = n7940 ^ n3134 ^ 1'b0 ;
  assign n27626 = n7550 | n27625 ;
  assign n27627 = n1839 & ~n27626 ;
  assign n27628 = n27627 ^ n16716 ^ 1'b0 ;
  assign n27629 = n9626 | n27628 ;
  assign n27631 = n12170 ^ n5578 ^ 1'b0 ;
  assign n27632 = n1682 | n27631 ;
  assign n27630 = ( ~n3405 & n13965 ) | ( ~n3405 & n22744 ) | ( n13965 & n22744 ) ;
  assign n27633 = n27632 ^ n27630 ^ 1'b0 ;
  assign n27634 = n27633 ^ n19881 ^ n10342 ;
  assign n27635 = ( n19020 & ~n26133 ) | ( n19020 & n27238 ) | ( ~n26133 & n27238 ) ;
  assign n27636 = n19414 ^ n10656 ^ 1'b0 ;
  assign n27637 = ( ~n19898 & n24423 ) | ( ~n19898 & n27636 ) | ( n24423 & n27636 ) ;
  assign n27638 = n14172 ^ n11908 ^ n2867 ;
  assign n27639 = n4880 ^ n1370 ^ n357 ;
  assign n27640 = n27639 ^ n7263 ^ 1'b0 ;
  assign n27641 = n6617 & ~n27640 ;
  assign n27642 = ( n2252 & n13705 ) | ( n2252 & n27360 ) | ( n13705 & n27360 ) ;
  assign n27643 = n27642 ^ n8808 ^ 1'b0 ;
  assign n27644 = n23304 ^ n4663 ^ 1'b0 ;
  assign n27645 = ~n10876 & n17822 ;
  assign n27646 = n3527 | n12096 ;
  assign n27647 = n1973 ^ n1870 ^ n1387 ;
  assign n27648 = n27647 ^ n2048 ^ 1'b0 ;
  assign n27649 = ~n14619 & n27648 ;
  assign n27650 = ( ~n1229 & n27646 ) | ( ~n1229 & n27649 ) | ( n27646 & n27649 ) ;
  assign n27651 = n19206 ^ n18052 ^ n8469 ;
  assign n27652 = n11521 ^ n1387 ^ 1'b0 ;
  assign n27653 = n27652 ^ n17446 ^ n2876 ;
  assign n27654 = n3749 & n27653 ;
  assign n27655 = n27654 ^ n20015 ^ n11270 ;
  assign n27656 = ( n20625 & n27284 ) | ( n20625 & ~n27655 ) | ( n27284 & ~n27655 ) ;
  assign n27657 = n2879 | n4000 ;
  assign n27658 = n18328 ^ n1406 ^ 1'b0 ;
  assign n27659 = n7411 | n27658 ;
  assign n27661 = n4834 ^ n3590 ^ 1'b0 ;
  assign n27660 = n16407 & ~n25112 ;
  assign n27662 = n27661 ^ n27660 ^ 1'b0 ;
  assign n27663 = n6569 & n13263 ;
  assign n27664 = ~n2798 & n27663 ;
  assign n27665 = n2713 & n6984 ;
  assign n27670 = n6016 & n8079 ;
  assign n27671 = ~n21257 & n27670 ;
  assign n27666 = n2361 & ~n18957 ;
  assign n27667 = n27666 ^ n14627 ^ 1'b0 ;
  assign n27668 = ~n296 & n27667 ;
  assign n27669 = n27668 ^ n216 ^ 1'b0 ;
  assign n27672 = n27671 ^ n27669 ^ n19598 ;
  assign n27673 = n13204 & ~n14155 ;
  assign n27674 = ( n8258 & n11769 ) | ( n8258 & ~n17117 ) | ( n11769 & ~n17117 ) ;
  assign n27675 = n27674 ^ n9460 ^ n3274 ;
  assign n27676 = ( n851 & n14575 ) | ( n851 & ~n27675 ) | ( n14575 & ~n27675 ) ;
  assign n27677 = n22823 ^ n12957 ^ n5535 ;
  assign n27678 = n4699 | n25448 ;
  assign n27680 = n1716 & ~n7635 ;
  assign n27679 = n1189 & ~n9108 ;
  assign n27681 = n27680 ^ n27679 ^ 1'b0 ;
  assign n27683 = n7875 ^ n2423 ^ 1'b0 ;
  assign n27682 = n2110 | n13925 ;
  assign n27684 = n27683 ^ n27682 ^ 1'b0 ;
  assign n27685 = n15595 & ~n25692 ;
  assign n27686 = ~n7883 & n12333 ;
  assign n27687 = n17337 ^ n1024 ^ 1'b0 ;
  assign n27688 = n18682 & ~n27687 ;
  assign n27689 = n25306 | n27688 ;
  assign n27690 = ( n567 & ~n16090 ) | ( n567 & n19870 ) | ( ~n16090 & n19870 ) ;
  assign n27691 = ( n17968 & ~n27606 ) | ( n17968 & n27690 ) | ( ~n27606 & n27690 ) ;
  assign n27692 = n27130 ^ n3737 ^ 1'b0 ;
  assign n27693 = n16638 | n22634 ;
  assign n27694 = n27692 & ~n27693 ;
  assign n27695 = n6714 & ~n25558 ;
  assign n27696 = n27694 & n27695 ;
  assign n27697 = n4100 ^ n2373 ^ 1'b0 ;
  assign n27698 = n5543 | n27697 ;
  assign n27699 = n3347 & n26238 ;
  assign n27700 = n27698 & n27699 ;
  assign n27701 = n8582 ^ n1521 ^ 1'b0 ;
  assign n27702 = n14164 ^ n11258 ^ 1'b0 ;
  assign n27703 = ( n3723 & n23074 ) | ( n3723 & ~n27702 ) | ( n23074 & ~n27702 ) ;
  assign n27704 = n27703 ^ n16136 ^ n7103 ;
  assign n27705 = ~n7152 & n18696 ;
  assign n27706 = ( n4828 & n12449 ) | ( n4828 & n23208 ) | ( n12449 & n23208 ) ;
  assign n27707 = n27706 ^ n2112 ^ n1366 ;
  assign n27708 = n23528 ^ n12849 ^ 1'b0 ;
  assign n27709 = n9782 ^ n6930 ^ 1'b0 ;
  assign n27710 = n16803 & ~n27709 ;
  assign n27711 = n27710 ^ n10591 ^ 1'b0 ;
  assign n27712 = n23055 & n27711 ;
  assign n27715 = ~n11984 & n15113 ;
  assign n27716 = n17009 & n27715 ;
  assign n27713 = n11364 | n17082 ;
  assign n27714 = n3775 & n27713 ;
  assign n27717 = n27716 ^ n27714 ^ 1'b0 ;
  assign n27718 = n266 & ~n10001 ;
  assign n27719 = n27718 ^ n12541 ^ 1'b0 ;
  assign n27720 = n3907 & n27719 ;
  assign n27722 = n23455 ^ n6859 ^ 1'b0 ;
  assign n27721 = n8941 & n17855 ;
  assign n27723 = n27722 ^ n27721 ^ 1'b0 ;
  assign n27725 = ~n11582 & n13479 ;
  assign n27726 = n27725 ^ n360 ^ 1'b0 ;
  assign n27727 = ( n8273 & n22565 ) | ( n8273 & n27726 ) | ( n22565 & n27726 ) ;
  assign n27724 = n315 | n5631 ;
  assign n27728 = n27727 ^ n27724 ^ n25017 ;
  assign n27729 = n10735 ^ n2383 ^ 1'b0 ;
  assign n27730 = ~n6403 & n27729 ;
  assign n27731 = n27730 ^ n25171 ^ 1'b0 ;
  assign n27732 = n15862 ^ n1247 ^ 1'b0 ;
  assign n27733 = n3900 | n16578 ;
  assign n27734 = n27733 ^ n9661 ^ n809 ;
  assign n27735 = n9383 & n22091 ;
  assign n27736 = n27735 ^ n17375 ^ 1'b0 ;
  assign n27737 = n14308 & ~n17947 ;
  assign n27738 = ~n1640 & n27737 ;
  assign n27739 = ~n916 & n14204 ;
  assign n27740 = ( n15893 & n18005 ) | ( n15893 & ~n27739 ) | ( n18005 & ~n27739 ) ;
  assign n27741 = ~n20326 & n27740 ;
  assign n27742 = n27738 & n27741 ;
  assign n27743 = n10854 & n15480 ;
  assign n27744 = ( n4882 & n8493 ) | ( n4882 & ~n9805 ) | ( n8493 & ~n9805 ) ;
  assign n27745 = n23520 ^ n22512 ^ n13399 ;
  assign n27746 = ~n531 & n22056 ;
  assign n27747 = ~n24443 & n27746 ;
  assign n27748 = n27747 ^ n16593 ^ 1'b0 ;
  assign n27749 = n15477 ^ n15126 ^ 1'b0 ;
  assign n27750 = ~n15146 & n26911 ;
  assign n27751 = ( ~n9183 & n16727 ) | ( ~n9183 & n27484 ) | ( n16727 & n27484 ) ;
  assign n27752 = n27751 ^ n8658 ^ 1'b0 ;
  assign n27753 = n23582 | n27752 ;
  assign n27754 = n6527 | n8587 ;
  assign n27755 = n27754 ^ n13381 ^ 1'b0 ;
  assign n27756 = n328 | n3640 ;
  assign n27757 = n8309 | n27756 ;
  assign n27758 = ~n4819 & n27757 ;
  assign n27759 = n24334 ^ n17741 ^ 1'b0 ;
  assign n27760 = n25987 ^ n6055 ^ 1'b0 ;
  assign n27761 = n23847 & ~n27760 ;
  assign n27762 = ~n26941 & n27761 ;
  assign n27763 = ~n17380 & n27762 ;
  assign n27764 = n676 & ~n1086 ;
  assign n27765 = n27764 ^ n5857 ^ 1'b0 ;
  assign n27766 = ( n4179 & ~n15169 ) | ( n4179 & n27765 ) | ( ~n15169 & n27765 ) ;
  assign n27767 = n10341 & n13181 ;
  assign n27768 = n27767 ^ n13574 ^ 1'b0 ;
  assign n27769 = n27766 & ~n27768 ;
  assign n27770 = n2057 & ~n9317 ;
  assign n27771 = n3660 | n27770 ;
  assign n27772 = ( n2381 & n9773 ) | ( n2381 & ~n15757 ) | ( n9773 & ~n15757 ) ;
  assign n27773 = n12800 & ~n27772 ;
  assign n27774 = n8227 & n27773 ;
  assign n27775 = ~n5446 & n13060 ;
  assign n27776 = n27774 & n27775 ;
  assign n27777 = n590 & n17330 ;
  assign n27778 = n24942 ^ n8137 ^ 1'b0 ;
  assign n27779 = ~n8331 & n27778 ;
  assign n27780 = n27779 ^ n22898 ^ n6163 ;
  assign n27781 = ( n7934 & n14489 ) | ( n7934 & n18972 ) | ( n14489 & n18972 ) ;
  assign n27782 = ~n5261 & n26314 ;
  assign n27783 = n27782 ^ n21864 ^ 1'b0 ;
  assign n27784 = ( n13519 & n15408 ) | ( n13519 & ~n27783 ) | ( n15408 & ~n27783 ) ;
  assign n27785 = ( ~n1447 & n6130 ) | ( ~n1447 & n24311 ) | ( n6130 & n24311 ) ;
  assign n27786 = n21590 ^ n10036 ^ n2544 ;
  assign n27787 = n1282 | n3154 ;
  assign n27788 = n11616 & ~n27787 ;
  assign n27789 = n13856 ^ n6440 ^ 1'b0 ;
  assign n27790 = n17248 | n27789 ;
  assign n27791 = n27790 ^ n3071 ^ 1'b0 ;
  assign n27792 = n4765 & ~n9414 ;
  assign n27793 = n17157 & n27792 ;
  assign n27794 = n2140 & ~n27793 ;
  assign n27795 = n21438 & n27794 ;
  assign n27796 = ( n13844 & n26416 ) | ( n13844 & n27795 ) | ( n26416 & n27795 ) ;
  assign n27797 = ~n15387 & n27796 ;
  assign n27798 = n531 | n21251 ;
  assign n27799 = n27798 ^ n3850 ^ n1074 ;
  assign n27800 = n17133 ^ n9617 ^ 1'b0 ;
  assign n27801 = n21207 & ~n22631 ;
  assign n27802 = n7337 ^ n3913 ^ 1'b0 ;
  assign n27803 = n8381 ^ n8230 ^ 1'b0 ;
  assign n27804 = n8106 & ~n18827 ;
  assign n27805 = x81 & n8938 ;
  assign n27806 = n27805 ^ n827 ^ 1'b0 ;
  assign n27807 = n18496 ^ n12212 ^ n1842 ;
  assign n27808 = n12654 & n27807 ;
  assign n27809 = n27808 ^ n3633 ^ 1'b0 ;
  assign n27810 = n9158 & ~n11164 ;
  assign n27811 = ( ~n2277 & n22308 ) | ( ~n2277 & n26198 ) | ( n22308 & n26198 ) ;
  assign n27812 = n266 & n1645 ;
  assign n27813 = n27812 ^ n25738 ^ n24489 ;
  assign n27814 = ( n2289 & ~n3310 ) | ( n2289 & n9935 ) | ( ~n3310 & n9935 ) ;
  assign n27815 = n27814 ^ n17970 ^ n7192 ;
  assign n27816 = n7191 & n23162 ;
  assign n27817 = n11618 & n27816 ;
  assign n27818 = n27817 ^ n15531 ^ n13986 ;
  assign n27819 = n27818 ^ n14461 ^ 1'b0 ;
  assign n27820 = n6109 ^ n349 ^ 1'b0 ;
  assign n27821 = ~n20030 & n27820 ;
  assign n27822 = ( n2209 & ~n6215 ) | ( n2209 & n9675 ) | ( ~n6215 & n9675 ) ;
  assign n27823 = n7291 | n27822 ;
  assign n27824 = n14412 | n27823 ;
  assign n27825 = n27114 ^ n8708 ^ x17 ;
  assign n27826 = n27825 ^ n3754 ^ 1'b0 ;
  assign n27827 = n9556 & ~n27826 ;
  assign n27828 = n5665 & n14116 ;
  assign n27829 = n1720 & n27828 ;
  assign n27830 = ( n3787 & ~n8562 ) | ( n3787 & n23057 ) | ( ~n8562 & n23057 ) ;
  assign n27831 = n27830 ^ n22383 ^ n5730 ;
  assign n27832 = n7968 ^ n4481 ^ 1'b0 ;
  assign n27833 = n11211 ^ n8545 ^ n796 ;
  assign n27834 = ( n17407 & n27832 ) | ( n17407 & ~n27833 ) | ( n27832 & ~n27833 ) ;
  assign n27835 = ( ~n1740 & n11833 ) | ( ~n1740 & n16765 ) | ( n11833 & n16765 ) ;
  assign n27836 = n14618 ^ n4894 ^ 1'b0 ;
  assign n27837 = ( n10609 & n14900 ) | ( n10609 & ~n18542 ) | ( n14900 & ~n18542 ) ;
  assign n27838 = n18250 ^ n14368 ^ 1'b0 ;
  assign n27839 = n9324 | n27838 ;
  assign n27840 = n27839 ^ n20735 ^ n2272 ;
  assign n27841 = n27840 ^ n10510 ^ 1'b0 ;
  assign n27842 = ( ~n1276 & n4380 ) | ( ~n1276 & n7207 ) | ( n4380 & n7207 ) ;
  assign n27843 = n2977 & ~n27842 ;
  assign n27844 = n27843 ^ n21385 ^ 1'b0 ;
  assign n27845 = n23894 ^ n19216 ^ 1'b0 ;
  assign n27846 = n12338 & ~n27845 ;
  assign n27847 = n27846 ^ x21 ^ 1'b0 ;
  assign n27848 = n3091 ^ n2543 ^ n2513 ;
  assign n27849 = n27848 ^ n8565 ^ 1'b0 ;
  assign n27850 = n5068 | n27849 ;
  assign n27851 = n26694 ^ n1068 ^ 1'b0 ;
  assign n27852 = n10304 & n17851 ;
  assign n27853 = n5301 & n27852 ;
  assign n27854 = n27853 ^ n18850 ^ n14418 ;
  assign n27855 = n13957 ^ n2819 ^ 1'b0 ;
  assign n27856 = n27855 ^ n23001 ^ n17553 ;
  assign n27857 = ~n7725 & n17009 ;
  assign n27858 = ( n1518 & n9573 ) | ( n1518 & ~n12633 ) | ( n9573 & ~n12633 ) ;
  assign n27859 = ( ~n16279 & n27857 ) | ( ~n16279 & n27858 ) | ( n27857 & n27858 ) ;
  assign n27860 = ( ~n208 & n2060 ) | ( ~n208 & n9958 ) | ( n2060 & n9958 ) ;
  assign n27861 = n5868 & ~n19097 ;
  assign n27862 = n27861 ^ n1962 ^ 1'b0 ;
  assign n27863 = n4055 ^ n2343 ^ 1'b0 ;
  assign n27864 = ~n2573 & n27863 ;
  assign n27865 = n331 & n10862 ;
  assign n27866 = n20729 ^ n11805 ^ 1'b0 ;
  assign n27867 = n27865 & n27866 ;
  assign n27868 = n1636 | n27429 ;
  assign n27871 = ~n2767 & n10379 ;
  assign n27872 = n10359 & n27871 ;
  assign n27869 = n1376 | n12342 ;
  assign n27870 = n27869 ^ n17006 ^ 1'b0 ;
  assign n27873 = n27872 ^ n27870 ^ n7119 ;
  assign n27874 = n6892 ^ n5453 ^ n3750 ;
  assign n27875 = n21817 ^ n1972 ^ 1'b0 ;
  assign n27876 = ( n9698 & n25558 ) | ( n9698 & n27875 ) | ( n25558 & n27875 ) ;
  assign n27877 = n366 & ~n9364 ;
  assign n27878 = n15317 ^ n14053 ^ n9373 ;
  assign n27879 = n27878 ^ n18215 ^ 1'b0 ;
  assign n27880 = n10660 ^ n2029 ^ 1'b0 ;
  assign n27881 = n9391 & ~n27880 ;
  assign n27882 = n3896 | n9246 ;
  assign n27883 = n25762 ^ n23579 ^ 1'b0 ;
  assign n27884 = n25272 & n27883 ;
  assign n27885 = n2363 & n3625 ;
  assign n27886 = ~n16955 & n27885 ;
  assign n27888 = ( n3149 & ~n15918 ) | ( n3149 & n18030 ) | ( ~n15918 & n18030 ) ;
  assign n27887 = n7100 | n27830 ;
  assign n27889 = n27888 ^ n27887 ^ 1'b0 ;
  assign n27890 = ( ~n4605 & n6191 ) | ( ~n4605 & n27889 ) | ( n6191 & n27889 ) ;
  assign n27891 = ~n16670 & n25716 ;
  assign n27892 = ( x51 & n20484 ) | ( x51 & n23307 ) | ( n20484 & n23307 ) ;
  assign n27893 = n8385 ^ n7984 ^ 1'b0 ;
  assign n27894 = n14965 ^ n11246 ^ n9175 ;
  assign n27895 = n27894 ^ n12652 ^ 1'b0 ;
  assign n27896 = n27893 & ~n27895 ;
  assign n27897 = ~n6173 & n24914 ;
  assign n27898 = ~n2774 & n27897 ;
  assign n27900 = n12125 ^ n6274 ^ 1'b0 ;
  assign n27901 = n4240 | n27900 ;
  assign n27899 = ~n14678 & n16813 ;
  assign n27902 = n27901 ^ n27899 ^ 1'b0 ;
  assign n27903 = n5593 ^ n2329 ^ 1'b0 ;
  assign n27904 = n7611 | n27903 ;
  assign n27905 = n27098 ^ n15976 ^ 1'b0 ;
  assign n27906 = ( n14097 & ~n27607 ) | ( n14097 & n27905 ) | ( ~n27607 & n27905 ) ;
  assign n27909 = ( n5984 & n9951 ) | ( n5984 & ~n12195 ) | ( n9951 & ~n12195 ) ;
  assign n27907 = n1658 & n6629 ;
  assign n27908 = n8832 & n27907 ;
  assign n27910 = n27909 ^ n27908 ^ n22383 ;
  assign n27911 = x67 & n501 ;
  assign n27912 = n12407 & n27911 ;
  assign n27913 = ( n1264 & n25250 ) | ( n1264 & ~n27912 ) | ( n25250 & ~n27912 ) ;
  assign n27914 = ( n5641 & ~n6879 ) | ( n5641 & n9473 ) | ( ~n6879 & n9473 ) ;
  assign n27916 = n6005 ^ n4020 ^ n1493 ;
  assign n27915 = n15118 | n25742 ;
  assign n27917 = n27916 ^ n27915 ^ 1'b0 ;
  assign n27918 = n1653 & n22719 ;
  assign n27919 = ~n27773 & n27918 ;
  assign n27920 = n12185 | n16049 ;
  assign n27921 = n11289 & ~n27920 ;
  assign n27925 = n8554 ^ n5779 ^ n2854 ;
  assign n27926 = n1855 | n27925 ;
  assign n27922 = n23641 | n27683 ;
  assign n27923 = n12233 | n27922 ;
  assign n27924 = n15331 & n27923 ;
  assign n27927 = n27926 ^ n27924 ^ 1'b0 ;
  assign n27928 = n18103 ^ n6754 ^ 1'b0 ;
  assign n27929 = n9714 | n27928 ;
  assign n27930 = ( ~n4254 & n27927 ) | ( ~n4254 & n27929 ) | ( n27927 & n27929 ) ;
  assign n27931 = n14362 ^ n4782 ^ 1'b0 ;
  assign n27932 = ( ~n5570 & n27242 ) | ( ~n5570 & n27931 ) | ( n27242 & n27931 ) ;
  assign n27934 = n5050 & ~n8137 ;
  assign n27933 = ~n5883 & n6186 ;
  assign n27935 = n27934 ^ n27933 ^ n23331 ;
  assign n27936 = ( n5305 & n22216 ) | ( n5305 & n24037 ) | ( n22216 & n24037 ) ;
  assign n27937 = ~n1558 & n27936 ;
  assign n27938 = n14619 & n27937 ;
  assign n27939 = ~n12690 & n27938 ;
  assign n27940 = n8427 ^ n1447 ^ 1'b0 ;
  assign n27941 = n15228 | n27940 ;
  assign n27944 = ( n2056 & n2062 ) | ( n2056 & n3407 ) | ( n2062 & n3407 ) ;
  assign n27942 = ~n12369 & n23137 ;
  assign n27943 = n5490 & ~n27942 ;
  assign n27945 = n27944 ^ n27943 ^ 1'b0 ;
  assign n27947 = n846 & n5202 ;
  assign n27946 = n5915 ^ n786 ^ x105 ;
  assign n27948 = n27947 ^ n27946 ^ n14594 ;
  assign n27949 = n16885 ^ n7174 ^ n5522 ;
  assign n27950 = n27949 ^ n4840 ^ n502 ;
  assign n27956 = n1726 & n13174 ;
  assign n27957 = n4247 & n27956 ;
  assign n27951 = ( n5018 & ~n19753 ) | ( n5018 & n22634 ) | ( ~n19753 & n22634 ) ;
  assign n27952 = n18353 & ~n27951 ;
  assign n27953 = n11062 ^ n9077 ^ n1069 ;
  assign n27954 = n7724 & n27953 ;
  assign n27955 = ( n6699 & ~n27952 ) | ( n6699 & n27954 ) | ( ~n27952 & n27954 ) ;
  assign n27958 = n27957 ^ n27955 ^ n11848 ;
  assign n27962 = ( n2377 & ~n4039 ) | ( n2377 & n6571 ) | ( ~n4039 & n6571 ) ;
  assign n27959 = ( n1443 & ~n3257 ) | ( n1443 & n3293 ) | ( ~n3257 & n3293 ) ;
  assign n27960 = n27959 ^ n23162 ^ x113 ;
  assign n27961 = n11957 & n27960 ;
  assign n27963 = n27962 ^ n27961 ^ 1'b0 ;
  assign n27964 = n4815 ^ n485 ^ 1'b0 ;
  assign n27965 = ( n612 & ~n16641 ) | ( n612 & n27964 ) | ( ~n16641 & n27964 ) ;
  assign n27966 = n25568 | n27115 ;
  assign n27967 = n27965 & ~n27966 ;
  assign n27968 = n9324 ^ n6744 ^ 1'b0 ;
  assign n27969 = n3268 | n5084 ;
  assign n27970 = n5381 & ~n27969 ;
  assign n27971 = n27970 ^ n4511 ^ 1'b0 ;
  assign n27972 = ~n27968 & n27971 ;
  assign n27973 = n5827 ^ n2797 ^ n1132 ;
  assign n27974 = n6402 ^ n5801 ^ n3401 ;
  assign n27975 = n10998 & n16285 ;
  assign n27976 = n27975 ^ n27767 ^ 1'b0 ;
  assign n27977 = ( ~n24985 & n27974 ) | ( ~n24985 & n27976 ) | ( n27974 & n27976 ) ;
  assign n27979 = n5498 & n13984 ;
  assign n27978 = n26211 ^ n11659 ^ n9341 ;
  assign n27980 = n27979 ^ n27978 ^ n4421 ;
  assign n27981 = n1316 & ~n22975 ;
  assign n27982 = n27981 ^ n9152 ^ 1'b0 ;
  assign n27983 = x32 & ~n9926 ;
  assign n27987 = n6421 | n15464 ;
  assign n27988 = n22625 & ~n27987 ;
  assign n27984 = ~n4429 & n14785 ;
  assign n27985 = n4177 & n27984 ;
  assign n27986 = n27985 ^ n17343 ^ 1'b0 ;
  assign n27989 = n27988 ^ n27986 ^ n11799 ;
  assign n27990 = n4477 | n6831 ;
  assign n27991 = n27990 ^ n8558 ^ 1'b0 ;
  assign n27992 = n9993 & n27991 ;
  assign n27993 = n23763 ^ n18951 ^ 1'b0 ;
  assign n27994 = n2433 | n18838 ;
  assign n27995 = n27994 ^ n8630 ^ 1'b0 ;
  assign n27996 = n12252 ^ n9143 ^ n1957 ;
  assign n27997 = n23456 & ~n27996 ;
  assign n27998 = ~n10460 & n27997 ;
  assign n27999 = n10683 ^ n10617 ^ 1'b0 ;
  assign n28000 = ( n11319 & ~n20132 ) | ( n11319 & n21417 ) | ( ~n20132 & n21417 ) ;
  assign n28004 = n9607 & ~n23823 ;
  assign n28005 = n17437 & n28004 ;
  assign n28001 = ~n2910 & n4791 ;
  assign n28002 = ~n21499 & n28001 ;
  assign n28003 = n8432 & ~n28002 ;
  assign n28006 = n28005 ^ n28003 ^ n23556 ;
  assign n28007 = ( n3657 & n13442 ) | ( n3657 & ~n20046 ) | ( n13442 & ~n20046 ) ;
  assign n28008 = ( n13196 & n13281 ) | ( n13196 & n15381 ) | ( n13281 & n15381 ) ;
  assign n28009 = n2839 | n4486 ;
  assign n28010 = ~n1075 & n28009 ;
  assign n28011 = n12849 & n16516 ;
  assign n28012 = n28011 ^ n24446 ^ 1'b0 ;
  assign n28013 = n14726 ^ n4525 ^ 1'b0 ;
  assign n28014 = n372 & ~n1851 ;
  assign n28015 = n10359 & n28014 ;
  assign n28016 = ( ~n1332 & n5569 ) | ( ~n1332 & n21400 ) | ( n5569 & n21400 ) ;
  assign n28020 = n24761 ^ n24507 ^ 1'b0 ;
  assign n28017 = n5002 & n22666 ;
  assign n28018 = n11560 & ~n28017 ;
  assign n28019 = n28018 ^ n1837 ^ 1'b0 ;
  assign n28021 = n28020 ^ n28019 ^ n8577 ;
  assign n28022 = ( n7417 & n15583 ) | ( n7417 & ~n28021 ) | ( n15583 & ~n28021 ) ;
  assign n28023 = n1329 | n11427 ;
  assign n28024 = ( n7244 & ~n23422 ) | ( n7244 & n28023 ) | ( ~n23422 & n28023 ) ;
  assign n28025 = n26206 ^ n8679 ^ n5353 ;
  assign n28026 = n17371 ^ n8795 ^ 1'b0 ;
  assign n28027 = ~n15649 & n28026 ;
  assign n28028 = n28027 ^ n16278 ^ 1'b0 ;
  assign n28029 = ~n2865 & n28028 ;
  assign n28030 = n5267 | n13695 ;
  assign n28031 = n17744 ^ n9373 ^ 1'b0 ;
  assign n28032 = n924 & n28031 ;
  assign n28033 = n18589 ^ n18136 ^ n7886 ;
  assign n28034 = n740 & ~n28033 ;
  assign n28035 = n4292 & n14266 ;
  assign n28036 = n28035 ^ n16987 ^ 1'b0 ;
  assign n28037 = n28036 ^ n20797 ^ 1'b0 ;
  assign n28038 = ~n708 & n21691 ;
  assign n28039 = ~n23209 & n28038 ;
  assign n28040 = n23970 ^ n11433 ^ n9192 ;
  assign n28041 = n17070 | n28040 ;
  assign n28042 = n28039 & ~n28041 ;
  assign n28043 = n7710 ^ x24 ^ 1'b0 ;
  assign n28044 = n5673 & ~n14015 ;
  assign n28045 = ~n28043 & n28044 ;
  assign n28046 = ( n8535 & ~n20610 ) | ( n8535 & n28045 ) | ( ~n20610 & n28045 ) ;
  assign n28047 = n28046 ^ n22379 ^ n20416 ;
  assign n28049 = n3165 ^ n601 ^ 1'b0 ;
  assign n28048 = ( ~n1861 & n21680 ) | ( ~n1861 & n23136 ) | ( n21680 & n23136 ) ;
  assign n28050 = n28049 ^ n28048 ^ n16779 ;
  assign n28051 = n14635 ^ n5902 ^ n3382 ;
  assign n28052 = ( n1154 & ~n3635 ) | ( n1154 & n22546 ) | ( ~n3635 & n22546 ) ;
  assign n28053 = n3238 & n26052 ;
  assign n28054 = n28053 ^ n6975 ^ 1'b0 ;
  assign n28055 = n191 & n28054 ;
  assign n28056 = n28055 ^ n19345 ^ 1'b0 ;
  assign n28057 = ~n28052 & n28056 ;
  assign n28058 = ~n5811 & n14967 ;
  assign n28059 = n3037 | n28058 ;
  assign n28060 = n14827 | n28059 ;
  assign n28061 = ~n17399 & n28060 ;
  assign n28062 = n28061 ^ n2320 ^ 1'b0 ;
  assign n28063 = n6023 ^ n1715 ^ 1'b0 ;
  assign n28064 = n469 & ~n8090 ;
  assign n28065 = n28064 ^ n8364 ^ 1'b0 ;
  assign n28066 = ~n15778 & n19944 ;
  assign n28067 = ~n28065 & n28066 ;
  assign n28068 = ~n4401 & n20259 ;
  assign n28069 = n5905 & n28068 ;
  assign n28070 = ~n4821 & n21018 ;
  assign n28071 = ( n1250 & ~n13714 ) | ( n1250 & n27319 ) | ( ~n13714 & n27319 ) ;
  assign n28072 = n2667 & n4819 ;
  assign n28073 = n28072 ^ n5037 ^ 1'b0 ;
  assign n28074 = ( n471 & ~n10942 ) | ( n471 & n18916 ) | ( ~n10942 & n18916 ) ;
  assign n28075 = n28074 ^ n8183 ^ 1'b0 ;
  assign n28076 = n28073 & n28075 ;
  assign n28077 = n28076 ^ n12457 ^ 1'b0 ;
  assign n28078 = ~n10351 & n14213 ;
  assign n28079 = ~x125 & n28078 ;
  assign n28080 = ~n280 & n13612 ;
  assign n28081 = n28080 ^ n3921 ^ 1'b0 ;
  assign n28082 = n1271 & ~n28081 ;
  assign n28083 = n2442 & n28082 ;
  assign n28084 = n25551 ^ n1542 ^ 1'b0 ;
  assign n28085 = n27300 | n28084 ;
  assign n28086 = n7752 ^ n2573 ^ 1'b0 ;
  assign n28087 = ~n28085 & n28086 ;
  assign n28088 = n437 | n1555 ;
  assign n28089 = n9534 ^ n6277 ^ n4033 ;
  assign n28090 = n2131 | n28089 ;
  assign n28091 = n17662 | n20697 ;
  assign n28092 = n28091 ^ n6215 ^ 1'b0 ;
  assign n28093 = n24274 & n28092 ;
  assign n28094 = n10586 & n19106 ;
  assign n28095 = ( n9024 & n17472 ) | ( n9024 & ~n21226 ) | ( n17472 & ~n21226 ) ;
  assign n28096 = n13938 ^ n13706 ^ n4421 ;
  assign n28097 = ( n4070 & ~n9508 ) | ( n4070 & n14041 ) | ( ~n9508 & n14041 ) ;
  assign n28098 = n10934 | n28097 ;
  assign n28099 = n25070 ^ n18099 ^ n10771 ;
  assign n28100 = n7024 & n28099 ;
  assign n28101 = n5971 & ~n15285 ;
  assign n28102 = n28101 ^ n1980 ^ 1'b0 ;
  assign n28103 = n3074 | n14569 ;
  assign n28104 = n623 & ~n28103 ;
  assign n28105 = n7349 | n7364 ;
  assign n28106 = n3020 & ~n28105 ;
  assign n28107 = ~n4136 & n9963 ;
  assign n28108 = n28107 ^ n11240 ^ n10616 ;
  assign n28109 = n28108 ^ n20186 ^ n15727 ;
  assign n28110 = n8227 | n18222 ;
  assign n28112 = ( n2860 & ~n8250 ) | ( n2860 & n8279 ) | ( ~n8250 & n8279 ) ;
  assign n28111 = n12431 ^ n8316 ^ n3521 ;
  assign n28113 = n28112 ^ n28111 ^ n5307 ;
  assign n28114 = ( ~n544 & n1067 ) | ( ~n544 & n17127 ) | ( n1067 & n17127 ) ;
  assign n28117 = n1234 & n26737 ;
  assign n28118 = ( n9190 & ~n21951 ) | ( n9190 & n28117 ) | ( ~n21951 & n28117 ) ;
  assign n28115 = n8149 & ~n9280 ;
  assign n28116 = n28115 ^ n4254 ^ 1'b0 ;
  assign n28119 = n28118 ^ n28116 ^ n3229 ;
  assign n28121 = n242 & n310 ;
  assign n28122 = n28121 ^ n4637 ^ 1'b0 ;
  assign n28123 = n4804 & ~n26222 ;
  assign n28124 = n28122 & n28123 ;
  assign n28120 = n4409 & n22379 ;
  assign n28125 = n28124 ^ n28120 ^ 1'b0 ;
  assign n28126 = n3311 | n12324 ;
  assign n28127 = n28126 ^ n10629 ^ 1'b0 ;
  assign n28128 = n8284 & n27327 ;
  assign n28129 = n28128 ^ n14009 ^ 1'b0 ;
  assign n28130 = n3836 | n11784 ;
  assign n28131 = n28130 ^ n5044 ^ 1'b0 ;
  assign n28132 = n26829 ^ n6931 ^ 1'b0 ;
  assign n28133 = n28132 ^ x82 ^ 1'b0 ;
  assign n28134 = ( n5229 & ~n24585 ) | ( n5229 & n28133 ) | ( ~n24585 & n28133 ) ;
  assign n28135 = n11552 ^ n4376 ^ 1'b0 ;
  assign n28136 = n12485 ^ n7237 ^ n3688 ;
  assign n28137 = n22800 | n28136 ;
  assign n28138 = ( n15118 & ~n28135 ) | ( n15118 & n28137 ) | ( ~n28135 & n28137 ) ;
  assign n28139 = n13550 & n18245 ;
  assign n28140 = ~n164 & n9582 ;
  assign n28141 = n28139 & n28140 ;
  assign n28142 = n588 & ~n3538 ;
  assign n28143 = n12460 & n28142 ;
  assign n28144 = n1777 & ~n28143 ;
  assign n28145 = ~n28141 & n28144 ;
  assign n28146 = n4377 & n4772 ;
  assign n28147 = ( n3161 & ~n3739 ) | ( n3161 & n28146 ) | ( ~n3739 & n28146 ) ;
  assign n28148 = n5030 ^ n352 ^ 1'b0 ;
  assign n28149 = n8791 & n28148 ;
  assign n28150 = n28149 ^ n26979 ^ n7647 ;
  assign n28152 = n13115 ^ n9373 ^ n1435 ;
  assign n28153 = n28152 ^ n24009 ^ 1'b0 ;
  assign n28151 = n6021 & n11118 ;
  assign n28154 = n28153 ^ n28151 ^ 1'b0 ;
  assign n28155 = n13193 ^ n5639 ^ n3666 ;
  assign n28156 = n28155 ^ n3164 ^ 1'b0 ;
  assign n28157 = n7657 & n28156 ;
  assign n28158 = ( n346 & ~n4701 ) | ( n346 & n24404 ) | ( ~n4701 & n24404 ) ;
  assign n28159 = ( ~n182 & n577 ) | ( ~n182 & n28158 ) | ( n577 & n28158 ) ;
  assign n28160 = n968 | n28159 ;
  assign n28161 = n28160 ^ n6918 ^ 1'b0 ;
  assign n28162 = n28161 ^ n26503 ^ n8997 ;
  assign n28163 = n6614 & ~n20251 ;
  assign n28164 = n26758 & n28163 ;
  assign n28165 = n6462 & ~n10275 ;
  assign n28166 = ~n7625 & n28165 ;
  assign n28167 = n5709 & n16807 ;
  assign n28168 = n28166 & n28167 ;
  assign n28169 = n11242 ^ n1620 ^ 1'b0 ;
  assign n28170 = n14887 ^ n1805 ^ 1'b0 ;
  assign n28171 = ( n12772 & ~n14743 ) | ( n12772 & n19809 ) | ( ~n14743 & n19809 ) ;
  assign n28172 = ( n3175 & ~n6405 ) | ( n3175 & n11253 ) | ( ~n6405 & n11253 ) ;
  assign n28173 = n10980 ^ n7444 ^ 1'b0 ;
  assign n28174 = x124 & ~n28173 ;
  assign n28175 = n4208 ^ n483 ^ 1'b0 ;
  assign n28176 = n28174 & n28175 ;
  assign n28177 = n14723 & n28176 ;
  assign n28178 = ( n3367 & n4512 ) | ( n3367 & ~n20720 ) | ( n4512 & ~n20720 ) ;
  assign n28179 = n329 & n23635 ;
  assign n28180 = ~n16397 & n28179 ;
  assign n28181 = n18999 | n26997 ;
  assign n28182 = n6092 ^ n4142 ^ 1'b0 ;
  assign n28183 = n28182 ^ n26699 ^ n13137 ;
  assign n28184 = ( n10132 & n12096 ) | ( n10132 & ~n28183 ) | ( n12096 & ~n28183 ) ;
  assign n28185 = n28184 ^ n5683 ^ 1'b0 ;
  assign n28186 = n209 & n1922 ;
  assign n28187 = ~n15428 & n28186 ;
  assign n28188 = n28187 ^ n21419 ^ 1'b0 ;
  assign n28189 = ~n5267 & n7979 ;
  assign n28190 = ~n157 & n28189 ;
  assign n28191 = n869 & ~n28190 ;
  assign n28192 = n28191 ^ n7024 ^ 1'b0 ;
  assign n28193 = ~n25487 & n28192 ;
  assign n28194 = n17301 ^ n11364 ^ n1962 ;
  assign n28195 = ( ~x69 & n10214 ) | ( ~x69 & n19944 ) | ( n10214 & n19944 ) ;
  assign n28196 = n26933 ^ n20147 ^ 1'b0 ;
  assign n28197 = n11978 | n28196 ;
  assign n28198 = n12383 & ~n18712 ;
  assign n28199 = n28198 ^ n7081 ^ 1'b0 ;
  assign n28200 = n21161 & ~n28199 ;
  assign n28201 = n28200 ^ n11886 ^ 1'b0 ;
  assign n28205 = n13984 ^ n5403 ^ n749 ;
  assign n28202 = n1466 & n9916 ;
  assign n28203 = ~n10314 & n28202 ;
  assign n28204 = n7124 | n28203 ;
  assign n28206 = n28205 ^ n28204 ^ 1'b0 ;
  assign n28207 = n20738 & n25578 ;
  assign n28208 = n10109 & n28207 ;
  assign n28209 = n5263 ^ n1739 ^ n887 ;
  assign n28210 = ~n3365 & n10136 ;
  assign n28211 = n28209 & n28210 ;
  assign n28216 = n2836 & n3262 ;
  assign n28217 = n28216 ^ x54 ^ 1'b0 ;
  assign n28212 = ( n1399 & n8779 ) | ( n1399 & n10980 ) | ( n8779 & n10980 ) ;
  assign n28213 = n28212 ^ n15201 ^ n9192 ;
  assign n28214 = n10334 ^ n2199 ^ 1'b0 ;
  assign n28215 = ( n13997 & n28213 ) | ( n13997 & ~n28214 ) | ( n28213 & ~n28214 ) ;
  assign n28218 = n28217 ^ n28215 ^ n2921 ;
  assign n28219 = ~n8576 & n14284 ;
  assign n28220 = n28219 ^ n13170 ^ n2459 ;
  assign n28221 = n10092 ^ n5940 ^ n4387 ;
  assign n28222 = ( n2819 & ~n3043 ) | ( n2819 & n9174 ) | ( ~n3043 & n9174 ) ;
  assign n28223 = n3684 | n7104 ;
  assign n28224 = ~n8538 & n28223 ;
  assign n28225 = n574 & n28224 ;
  assign n28226 = n17729 | n18670 ;
  assign n28229 = n2788 & n7129 ;
  assign n28230 = n28229 ^ n3405 ^ 1'b0 ;
  assign n28231 = n28230 ^ n11749 ^ 1'b0 ;
  assign n28232 = n25578 & ~n28231 ;
  assign n28233 = ( n13919 & n20871 ) | ( n13919 & n28232 ) | ( n20871 & n28232 ) ;
  assign n28227 = n7816 | n17575 ;
  assign n28228 = n28227 ^ n11659 ^ n11322 ;
  assign n28234 = n28233 ^ n28228 ^ 1'b0 ;
  assign n28235 = n6870 & n27000 ;
  assign n28236 = n1955 | n28235 ;
  assign n28237 = ~n18451 & n28236 ;
  assign n28238 = n28234 & n28237 ;
  assign n28239 = ( n308 & ~n760 ) | ( n308 & n11739 ) | ( ~n760 & n11739 ) ;
  assign n28240 = n28239 ^ x60 ^ 1'b0 ;
  assign n28241 = n28240 ^ n7998 ^ n5753 ;
  assign n28242 = ~n15228 & n17404 ;
  assign n28243 = n28242 ^ n1266 ^ 1'b0 ;
  assign n28244 = ~n16254 & n28243 ;
  assign n28245 = n8572 ^ n5639 ^ n1135 ;
  assign n28246 = n28245 ^ n25265 ^ n333 ;
  assign n28247 = n1074 & ~n28246 ;
  assign n28248 = x112 & n28247 ;
  assign n28249 = n16180 ^ n6473 ^ n4626 ;
  assign n28250 = ( n21155 & ~n28248 ) | ( n21155 & n28249 ) | ( ~n28248 & n28249 ) ;
  assign n28251 = ( n2272 & ~n6683 ) | ( n2272 & n7979 ) | ( ~n6683 & n7979 ) ;
  assign n28252 = ( n1348 & n3565 ) | ( n1348 & n14333 ) | ( n3565 & n14333 ) ;
  assign n28253 = n28252 ^ n18429 ^ 1'b0 ;
  assign n28254 = ( n28250 & n28251 ) | ( n28250 & ~n28253 ) | ( n28251 & ~n28253 ) ;
  assign n28255 = n17627 ^ n12549 ^ n7624 ;
  assign n28256 = n13726 ^ n13598 ^ 1'b0 ;
  assign n28257 = n28255 & ~n28256 ;
  assign n28258 = ( ~n19934 & n21553 ) | ( ~n19934 & n25129 ) | ( n21553 & n25129 ) ;
  assign n28259 = n28258 ^ n4283 ^ 1'b0 ;
  assign n28260 = n5506 & n9561 ;
  assign n28261 = ~n3935 & n28260 ;
  assign n28262 = n1905 | n19835 ;
  assign n28263 = ~n28261 & n28262 ;
  assign n28264 = ( n20937 & n22994 ) | ( n20937 & ~n24873 ) | ( n22994 & ~n24873 ) ;
  assign n28265 = ( n4197 & ~n14379 ) | ( n4197 & n28264 ) | ( ~n14379 & n28264 ) ;
  assign n28266 = n28265 ^ n21470 ^ 1'b0 ;
  assign n28267 = n1723 | n28266 ;
  assign n28268 = n20648 ^ n13971 ^ 1'b0 ;
  assign n28269 = n25715 ^ n21623 ^ 1'b0 ;
  assign n28270 = n24254 & ~n28269 ;
  assign n28271 = n1212 & ~n4259 ;
  assign n28272 = ( n4972 & ~n17401 ) | ( n4972 & n28271 ) | ( ~n17401 & n28271 ) ;
  assign n28273 = ( ~n7373 & n13118 ) | ( ~n7373 & n24952 ) | ( n13118 & n24952 ) ;
  assign n28274 = n23256 ^ n8879 ^ 1'b0 ;
  assign n28275 = ( n4933 & ~n5543 ) | ( n4933 & n28274 ) | ( ~n5543 & n28274 ) ;
  assign n28276 = n9183 ^ n7520 ^ 1'b0 ;
  assign n28277 = ~n15754 & n28276 ;
  assign n28278 = ( n2638 & n20094 ) | ( n2638 & n28277 ) | ( n20094 & n28277 ) ;
  assign n28279 = ( n2272 & n26837 ) | ( n2272 & n28278 ) | ( n26837 & n28278 ) ;
  assign n28280 = n9374 & ~n17112 ;
  assign n28281 = ~n11763 & n28280 ;
  assign n28282 = ~n9462 & n13052 ;
  assign n28283 = ~n7397 & n28282 ;
  assign n28284 = n19862 ^ n9032 ^ 1'b0 ;
  assign n28285 = n28283 | n28284 ;
  assign n28286 = n22216 ^ n16265 ^ 1'b0 ;
  assign n28287 = n28286 ^ n25439 ^ 1'b0 ;
  assign n28288 = ~n21552 & n28287 ;
  assign n28289 = ~n6176 & n19510 ;
  assign n28290 = n28289 ^ n2647 ^ 1'b0 ;
  assign n28291 = n5071 | n28290 ;
  assign n28292 = n18756 ^ n4739 ^ 1'b0 ;
  assign n28293 = n15114 & ~n28292 ;
  assign n28294 = n9518 & n11430 ;
  assign n28295 = n21893 & n28294 ;
  assign n28296 = n1129 & n7712 ;
  assign n28297 = ~n1077 & n28296 ;
  assign n28298 = n28297 ^ n14279 ^ n9411 ;
  assign n28299 = ( n1761 & n28295 ) | ( n1761 & ~n28298 ) | ( n28295 & ~n28298 ) ;
  assign n28301 = n13453 ^ n10258 ^ 1'b0 ;
  assign n28300 = n7165 & ~n10233 ;
  assign n28302 = n28301 ^ n28300 ^ n11958 ;
  assign n28303 = ( n10688 & n10698 ) | ( n10688 & ~n24914 ) | ( n10698 & ~n24914 ) ;
  assign n28304 = ( n1053 & n8649 ) | ( n1053 & ~n23977 ) | ( n8649 & ~n23977 ) ;
  assign n28305 = n19313 ^ n8549 ^ n2056 ;
  assign n28306 = ~n139 & n25241 ;
  assign n28307 = n28096 ^ n24253 ^ 1'b0 ;
  assign n28308 = n2728 & ~n28307 ;
  assign n28309 = n16481 ^ n2723 ^ 1'b0 ;
  assign n28310 = n22269 & ~n28309 ;
  assign n28311 = n13802 ^ n833 ^ 1'b0 ;
  assign n28312 = n10364 ^ n10317 ^ n3338 ;
  assign n28313 = ( ~n2187 & n22386 ) | ( ~n2187 & n28312 ) | ( n22386 & n28312 ) ;
  assign n28314 = ( ~n9324 & n9846 ) | ( ~n9324 & n28313 ) | ( n9846 & n28313 ) ;
  assign n28315 = n26628 ^ n1048 ^ 1'b0 ;
  assign n28316 = ~n13472 & n28315 ;
  assign n28317 = n28316 ^ n8368 ^ n6180 ;
  assign n28318 = n7635 ^ n7604 ^ 1'b0 ;
  assign n28319 = n2199 & ~n28318 ;
  assign n28320 = n28319 ^ n14121 ^ n8281 ;
  assign n28321 = ( n9445 & n15138 ) | ( n9445 & n28320 ) | ( n15138 & n28320 ) ;
  assign n28322 = ~n827 & n9598 ;
  assign n28323 = n28322 ^ n11387 ^ n6963 ;
  assign n28324 = n24253 ^ n19956 ^ n6336 ;
  assign n28326 = ( ~n257 & n3521 ) | ( ~n257 & n5949 ) | ( n3521 & n5949 ) ;
  assign n28325 = ~n9719 & n13282 ;
  assign n28327 = n28326 ^ n28325 ^ 1'b0 ;
  assign n28328 = ~n4989 & n21085 ;
  assign n28329 = n19120 & n28328 ;
  assign n28330 = n8163 & n12972 ;
  assign n28331 = n11601 ^ n9145 ^ 1'b0 ;
  assign n28332 = ( n3870 & n5714 ) | ( n3870 & ~n28331 ) | ( n5714 & ~n28331 ) ;
  assign n28333 = n28332 ^ n23869 ^ n14301 ;
  assign n28334 = n17982 ^ n17270 ^ n9814 ;
  assign n28335 = n24061 ^ n4816 ^ n3897 ;
  assign n28336 = n24720 & n28335 ;
  assign n28337 = n13661 ^ n6797 ^ n4882 ;
  assign n28338 = n28337 ^ n20813 ^ 1'b0 ;
  assign n28339 = n11234 & ~n28338 ;
  assign n28340 = ~n5823 & n28339 ;
  assign n28341 = n19841 ^ n13752 ^ 1'b0 ;
  assign n28342 = ~n28340 & n28341 ;
  assign n28343 = x48 & ~n15735 ;
  assign n28344 = ( ~n2271 & n8276 ) | ( ~n2271 & n28343 ) | ( n8276 & n28343 ) ;
  assign n28345 = n28344 ^ n19498 ^ n2911 ;
  assign n28346 = n18082 ^ n11047 ^ n3596 ;
  assign n28347 = n28346 ^ n18521 ^ n10760 ;
  assign n28348 = n16507 | n20897 ;
  assign n28349 = n28347 & ~n28348 ;
  assign n28350 = n2874 & ~n12839 ;
  assign n28351 = n3297 & n7928 ;
  assign n28352 = n25593 & n28351 ;
  assign n28353 = n15764 ^ n11628 ^ 1'b0 ;
  assign n28354 = n5221 | n8690 ;
  assign n28355 = n1828 & ~n28354 ;
  assign n28356 = ~n21906 & n28355 ;
  assign n28357 = ~n6169 & n6739 ;
  assign n28358 = n28357 ^ n6641 ^ 1'b0 ;
  assign n28359 = ( n9906 & ~n28356 ) | ( n9906 & n28358 ) | ( ~n28356 & n28358 ) ;
  assign n28360 = n19156 ^ n7104 ^ n2365 ;
  assign n28361 = ~n680 & n1188 ;
  assign n28362 = ~n12865 & n28361 ;
  assign n28363 = n28362 ^ n9621 ^ 1'b0 ;
  assign n28364 = ( ~n17719 & n28360 ) | ( ~n17719 & n28363 ) | ( n28360 & n28363 ) ;
  assign n28365 = ( ~n15242 & n26584 ) | ( ~n15242 & n28364 ) | ( n26584 & n28364 ) ;
  assign n28366 = ( n6082 & n21359 ) | ( n6082 & ~n26782 ) | ( n21359 & ~n26782 ) ;
  assign n28367 = ( n2050 & n6067 ) | ( n2050 & ~n28366 ) | ( n6067 & ~n28366 ) ;
  assign n28368 = n6133 | n10057 ;
  assign n28369 = ( ~n1726 & n6635 ) | ( ~n1726 & n28368 ) | ( n6635 & n28368 ) ;
  assign n28370 = n5313 & n13485 ;
  assign n28371 = n28370 ^ n17217 ^ 1'b0 ;
  assign n28372 = n3257 | n4294 ;
  assign n28373 = n520 | n28372 ;
  assign n28374 = ~n3986 & n28373 ;
  assign n28375 = n28374 ^ n24999 ^ 1'b0 ;
  assign n28376 = n11441 | n26313 ;
  assign n28377 = n5415 & ~n12950 ;
  assign n28387 = n5262 ^ n4578 ^ 1'b0 ;
  assign n28382 = n13315 ^ n3443 ^ 1'b0 ;
  assign n28383 = ~n4029 & n28382 ;
  assign n28381 = ~n3640 & n11623 ;
  assign n28384 = n28383 ^ n28381 ^ 1'b0 ;
  assign n28378 = n8174 ^ n6390 ^ 1'b0 ;
  assign n28379 = ~n2712 & n28378 ;
  assign n28380 = ~n14554 & n28379 ;
  assign n28385 = n28384 ^ n28380 ^ 1'b0 ;
  assign n28386 = ~n22540 & n28385 ;
  assign n28388 = n28387 ^ n28386 ^ 1'b0 ;
  assign n28389 = n14705 & n28388 ;
  assign n28390 = ( n3642 & ~n6851 ) | ( n3642 & n23482 ) | ( ~n6851 & n23482 ) ;
  assign n28391 = ( n16327 & ~n20217 ) | ( n16327 & n28390 ) | ( ~n20217 & n28390 ) ;
  assign n28392 = n3225 & n3985 ;
  assign n28393 = n28392 ^ n3303 ^ 1'b0 ;
  assign n28394 = ( ~n14651 & n22019 ) | ( ~n14651 & n28393 ) | ( n22019 & n28393 ) ;
  assign n28395 = n13003 & ~n23081 ;
  assign n28396 = n1038 & ~n4741 ;
  assign n28397 = n28396 ^ n5403 ^ 1'b0 ;
  assign n28398 = n20653 ^ n14359 ^ 1'b0 ;
  assign n28399 = n28397 & ~n28398 ;
  assign n28400 = n5025 ^ n455 ^ 1'b0 ;
  assign n28401 = ~n11544 & n28400 ;
  assign n28402 = n2962 & n23757 ;
  assign n28403 = ~n2962 & n28402 ;
  assign n28404 = n14170 & n23415 ;
  assign n28405 = n28404 ^ n6451 ^ 1'b0 ;
  assign n28406 = n28405 ^ n22506 ^ 1'b0 ;
  assign n28407 = ~n28403 & n28406 ;
  assign n28408 = n14912 | n18143 ;
  assign n28409 = n2407 | n28408 ;
  assign n28410 = n19729 ^ n14381 ^ n4283 ;
  assign n28411 = n12005 | n14410 ;
  assign n28412 = n10099 ^ n7042 ^ n570 ;
  assign n28413 = n6085 & n28412 ;
  assign n28414 = n28413 ^ n25483 ^ n15647 ;
  assign n28415 = n23008 ^ n11151 ^ n10019 ;
  assign n28416 = n6797 | n28415 ;
  assign n28417 = n4377 & ~n7840 ;
  assign n28419 = n7969 ^ n3923 ^ 1'b0 ;
  assign n28418 = n4266 | n27011 ;
  assign n28420 = n28419 ^ n28418 ^ 1'b0 ;
  assign n28421 = n15520 ^ n7644 ^ 1'b0 ;
  assign n28422 = n13644 | n28421 ;
  assign n28423 = n26527 ^ n4274 ^ 1'b0 ;
  assign n28424 = ~n6284 & n8049 ;
  assign n28425 = n28423 & n28424 ;
  assign n28426 = n23122 ^ n6941 ^ 1'b0 ;
  assign n28427 = ~n28425 & n28426 ;
  assign n28428 = n28427 ^ n24982 ^ 1'b0 ;
  assign n28429 = n28422 | n28428 ;
  assign n28431 = n10703 | n11331 ;
  assign n28432 = n576 & ~n28431 ;
  assign n28430 = n1020 & ~n10737 ;
  assign n28433 = n28432 ^ n28430 ^ 1'b0 ;
  assign n28434 = n13202 | n20233 ;
  assign n28435 = n25022 ^ n13802 ^ n4049 ;
  assign n28436 = ~n5142 & n5779 ;
  assign n28437 = ( n9365 & n15565 ) | ( n9365 & ~n28436 ) | ( n15565 & ~n28436 ) ;
  assign n28438 = n10304 ^ x33 ^ 1'b0 ;
  assign n28439 = n28438 ^ n5497 ^ n5437 ;
  assign n28442 = n1399 | n26386 ;
  assign n28443 = n10361 & ~n28442 ;
  assign n28444 = n28443 ^ n23352 ^ n4830 ;
  assign n28440 = n13816 ^ n13618 ^ 1'b0 ;
  assign n28441 = ~n7768 & n28440 ;
  assign n28445 = n28444 ^ n28441 ^ n28286 ;
  assign n28446 = ~n5308 & n21170 ;
  assign n28447 = ( n1205 & n8406 ) | ( n1205 & ~n28446 ) | ( n8406 & ~n28446 ) ;
  assign n28448 = n6627 & ~n28447 ;
  assign n28449 = n11201 | n27981 ;
  assign n28450 = n5336 | n28449 ;
  assign n28451 = ~n277 & n2648 ;
  assign n28452 = n10971 & ~n23474 ;
  assign n28453 = n28452 ^ n12663 ^ 1'b0 ;
  assign n28454 = n24512 ^ n19086 ^ n11573 ;
  assign n28455 = n18860 ^ n18676 ^ n2303 ;
  assign n28456 = ( ~n14346 & n28454 ) | ( ~n14346 & n28455 ) | ( n28454 & n28455 ) ;
  assign n28459 = n24853 ^ n1484 ^ 1'b0 ;
  assign n28457 = n17934 ^ n12341 ^ 1'b0 ;
  assign n28458 = ~n13658 & n28457 ;
  assign n28460 = n28459 ^ n28458 ^ n6376 ;
  assign n28461 = ( n6353 & n19393 ) | ( n6353 & ~n23895 ) | ( n19393 & ~n23895 ) ;
  assign n28462 = ( n6835 & ~n17339 ) | ( n6835 & n22037 ) | ( ~n17339 & n22037 ) ;
  assign n28463 = n19743 ^ n5297 ^ n164 ;
  assign n28464 = ( ~n8280 & n19282 ) | ( ~n8280 & n28463 ) | ( n19282 & n28463 ) ;
  assign n28465 = ( n7462 & n10913 ) | ( n7462 & ~n28464 ) | ( n10913 & ~n28464 ) ;
  assign n28466 = n243 | n5030 ;
  assign n28467 = n894 & ~n3131 ;
  assign n28468 = n28467 ^ n5537 ^ 1'b0 ;
  assign n28469 = n4046 & n10381 ;
  assign n28470 = ~n5370 & n28469 ;
  assign n28471 = n4758 | n19648 ;
  assign n28473 = n9717 & ~n14702 ;
  assign n28474 = n28473 ^ n13759 ^ 1'b0 ;
  assign n28475 = n6676 & n28474 ;
  assign n28472 = n3903 ^ n2831 ^ 1'b0 ;
  assign n28476 = n28475 ^ n28472 ^ n6311 ;
  assign n28477 = n5699 & ~n18117 ;
  assign n28478 = n28477 ^ n8672 ^ n1279 ;
  assign n28479 = n5886 | n10677 ;
  assign n28480 = n16701 & n28479 ;
  assign n28481 = n10263 | n28480 ;
  assign n28482 = n10681 | n28481 ;
  assign n28483 = n28482 ^ n17348 ^ n14592 ;
  assign n28484 = n15532 ^ n11981 ^ 1'b0 ;
  assign n28486 = n1976 | n8888 ;
  assign n28487 = n28486 ^ n8249 ^ 1'b0 ;
  assign n28485 = n27793 ^ n16847 ^ 1'b0 ;
  assign n28488 = n28487 ^ n28485 ^ n24808 ;
  assign n28489 = n17879 ^ n16509 ^ 1'b0 ;
  assign n28490 = n2744 ^ n2301 ^ 1'b0 ;
  assign n28491 = ~n8174 & n28490 ;
  assign n28492 = n23126 ^ n5113 ^ 1'b0 ;
  assign n28493 = ~n7241 & n22848 ;
  assign n28494 = n14771 ^ n10787 ^ 1'b0 ;
  assign n28495 = n4778 & n28494 ;
  assign n28496 = n28495 ^ n15704 ^ 1'b0 ;
  assign n28497 = n28496 ^ n17019 ^ n6746 ;
  assign n28498 = n7410 ^ n6376 ^ n2331 ;
  assign n28499 = n17542 ^ n9553 ^ n8839 ;
  assign n28500 = n13702 & ~n14090 ;
  assign n28501 = n25855 ^ n23461 ^ n14644 ;
  assign n28502 = n1482 & n23044 ;
  assign n28503 = n3265 ^ n1244 ^ 1'b0 ;
  assign n28504 = n28502 & n28503 ;
  assign n28505 = n3422 & n16509 ;
  assign n28506 = n28505 ^ n5827 ^ 1'b0 ;
  assign n28507 = n12457 ^ n2808 ^ 1'b0 ;
  assign n28508 = n13727 | n28507 ;
  assign n28509 = n28508 ^ n16047 ^ 1'b0 ;
  assign n28510 = ~n23810 & n24090 ;
  assign n28511 = ( n10763 & n12147 ) | ( n10763 & n28510 ) | ( n12147 & n28510 ) ;
  assign n28512 = n935 & ~n17661 ;
  assign n28513 = ~n28511 & n28512 ;
  assign n28514 = ( n7410 & n12567 ) | ( n7410 & ~n19352 ) | ( n12567 & ~n19352 ) ;
  assign n28515 = ( n447 & n1156 ) | ( n447 & ~n4727 ) | ( n1156 & ~n4727 ) ;
  assign n28516 = n28515 ^ n15756 ^ n14609 ;
  assign n28517 = n21963 ^ n10252 ^ 1'b0 ;
  assign n28518 = n3896 & n28517 ;
  assign n28519 = ( n314 & ~n2325 ) | ( n314 & n25795 ) | ( ~n2325 & n25795 ) ;
  assign n28520 = n11727 ^ n558 ^ 1'b0 ;
  assign n28521 = n6480 | n28520 ;
  assign n28522 = n28521 ^ n9040 ^ n5414 ;
  assign n28523 = n8647 | n28522 ;
  assign n28524 = ~n2336 & n15408 ;
  assign n28525 = ~n1526 & n28524 ;
  assign n28526 = n19581 | n26689 ;
  assign n28527 = n28526 ^ n12089 ^ 1'b0 ;
  assign n28528 = n23871 ^ n18009 ^ 1'b0 ;
  assign n28529 = n18829 & ~n28528 ;
  assign n28530 = ~n16036 & n28529 ;
  assign n28531 = n3022 & n24124 ;
  assign n28532 = ~n17102 & n28531 ;
  assign n28536 = ~n12971 & n14715 ;
  assign n28537 = n17456 & n28536 ;
  assign n28533 = ~n6759 & n15523 ;
  assign n28534 = n7025 | n28533 ;
  assign n28535 = ~n8342 & n28534 ;
  assign n28538 = n28537 ^ n28535 ^ 1'b0 ;
  assign n28539 = n1107 | n2070 ;
  assign n28540 = n13713 ^ n13703 ^ 1'b0 ;
  assign n28541 = ( ~n7263 & n21392 ) | ( ~n7263 & n28540 ) | ( n21392 & n28540 ) ;
  assign n28542 = ( ~n7597 & n22084 ) | ( ~n7597 & n28541 ) | ( n22084 & n28541 ) ;
  assign n28543 = ( n8464 & n10030 ) | ( n8464 & n16661 ) | ( n10030 & n16661 ) ;
  assign n28544 = n28543 ^ n21644 ^ 1'b0 ;
  assign n28545 = n21233 ^ n20894 ^ n10450 ;
  assign n28546 = ( n13857 & ~n22054 ) | ( n13857 & n28545 ) | ( ~n22054 & n28545 ) ;
  assign n28547 = n1781 & ~n6317 ;
  assign n28548 = n28547 ^ n16921 ^ n13214 ;
  assign n28549 = n19317 & n22806 ;
  assign n28550 = n28549 ^ n12954 ^ 1'b0 ;
  assign n28551 = n18670 & ~n28550 ;
  assign n28552 = n12176 & n28551 ;
  assign n28553 = n27432 ^ n16153 ^ 1'b0 ;
  assign n28554 = n8532 ^ n5807 ^ 1'b0 ;
  assign n28555 = ~n5566 & n28554 ;
  assign n28556 = n14427 ^ n10782 ^ n4331 ;
  assign n28557 = ( n255 & ~n15414 ) | ( n255 & n28556 ) | ( ~n15414 & n28556 ) ;
  assign n28558 = n28557 ^ n9581 ^ n1476 ;
  assign n28559 = n327 & n3629 ;
  assign n28560 = n28559 ^ n3527 ^ 1'b0 ;
  assign n28561 = n28558 | n28560 ;
  assign n28562 = n12311 & ~n22174 ;
  assign n28563 = n28562 ^ n20150 ^ n16676 ;
  assign n28564 = n23694 ^ n15443 ^ 1'b0 ;
  assign n28565 = n1295 & ~n28564 ;
  assign n28566 = ( ~n8915 & n11458 ) | ( ~n8915 & n28565 ) | ( n11458 & n28565 ) ;
  assign n28567 = n11770 ^ n1942 ^ 1'b0 ;
  assign n28568 = n19821 ^ n12159 ^ n204 ;
  assign n28569 = n26978 ^ n19740 ^ n18953 ;
  assign n28570 = n3265 & n20228 ;
  assign n28571 = n9245 & n28570 ;
  assign n28572 = n16581 ^ n2749 ^ 1'b0 ;
  assign n28573 = ~n10144 & n28572 ;
  assign n28574 = ~n17846 & n28573 ;
  assign n28576 = n543 & ~n8516 ;
  assign n28575 = n8641 & ~n11848 ;
  assign n28577 = n28576 ^ n28575 ^ 1'b0 ;
  assign n28578 = n15832 ^ n14605 ^ 1'b0 ;
  assign n28579 = ~n21303 & n28578 ;
  assign n28580 = n3209 & ~n15177 ;
  assign n28581 = n20401 & n28580 ;
  assign n28582 = ( n8643 & n16292 ) | ( n8643 & ~n18102 ) | ( n16292 & ~n18102 ) ;
  assign n28583 = n25917 | n28582 ;
  assign n28584 = n28583 ^ n8749 ^ 1'b0 ;
  assign n28585 = ~n28581 & n28584 ;
  assign n28586 = n10568 | n28585 ;
  assign n28587 = n13255 | n24412 ;
  assign n28588 = n28587 ^ n10585 ^ 1'b0 ;
  assign n28589 = n28588 ^ n26482 ^ 1'b0 ;
  assign n28590 = ( n472 & n5662 ) | ( n472 & ~n28589 ) | ( n5662 & ~n28589 ) ;
  assign n28591 = ( n3979 & n20954 ) | ( n3979 & ~n24937 ) | ( n20954 & ~n24937 ) ;
  assign n28592 = n7418 & n16445 ;
  assign n28593 = n5538 & n28592 ;
  assign n28594 = n9805 ^ n7788 ^ n431 ;
  assign n28595 = n28593 & n28594 ;
  assign n28596 = ( n13124 & ~n22733 ) | ( n13124 & n28595 ) | ( ~n22733 & n28595 ) ;
  assign n28599 = n2334 & ~n7289 ;
  assign n28600 = n5751 & n28599 ;
  assign n28601 = n28600 ^ n14758 ^ 1'b0 ;
  assign n28597 = n9045 ^ n7600 ^ 1'b0 ;
  assign n28598 = ~n15747 & n28597 ;
  assign n28602 = n28601 ^ n28598 ^ n16576 ;
  assign n28603 = n6906 | n14908 ;
  assign n28604 = n4049 ^ n3709 ^ 1'b0 ;
  assign n28605 = n10127 & n22148 ;
  assign n28606 = n28604 & n28605 ;
  assign n28607 = n4671 | n18821 ;
  assign n28608 = n14359 | n18195 ;
  assign n28609 = n2713 | n8601 ;
  assign n28610 = n2353 & ~n28609 ;
  assign n28611 = ( n6491 & ~n21579 ) | ( n6491 & n28610 ) | ( ~n21579 & n28610 ) ;
  assign n28612 = n28611 ^ n6926 ^ n5123 ;
  assign n28613 = ~n1586 & n28612 ;
  assign n28614 = ( n154 & ~n4069 ) | ( n154 & n10391 ) | ( ~n4069 & n10391 ) ;
  assign n28615 = ( ~n19901 & n26618 ) | ( ~n19901 & n28614 ) | ( n26618 & n28614 ) ;
  assign n28616 = n25552 ^ n5502 ^ 1'b0 ;
  assign n28617 = n23777 ^ n12715 ^ n4038 ;
  assign n28618 = n23426 ^ n5151 ^ n1851 ;
  assign n28619 = n19476 ^ n7797 ^ n2296 ;
  assign n28620 = n28619 ^ n15788 ^ 1'b0 ;
  assign n28621 = ( n243 & ~n3035 ) | ( n243 & n6845 ) | ( ~n3035 & n6845 ) ;
  assign n28622 = n22820 ^ n8584 ^ n7589 ;
  assign n28623 = n28622 ^ n6345 ^ 1'b0 ;
  assign n28624 = n28621 & ~n28623 ;
  assign n28625 = n7229 & n8706 ;
  assign n28626 = n4671 ^ n2830 ^ 1'b0 ;
  assign n28627 = n28625 & n28626 ;
  assign n28628 = n1761 & n19372 ;
  assign n28629 = n28628 ^ n6786 ^ 1'b0 ;
  assign n28630 = n20519 ^ n8549 ^ 1'b0 ;
  assign n28631 = n17787 & n23463 ;
  assign n28632 = ~n17601 & n23827 ;
  assign n28633 = ~n23188 & n27244 ;
  assign n28634 = ( n11578 & ~n26365 ) | ( n11578 & n28633 ) | ( ~n26365 & n28633 ) ;
  assign n28635 = n4691 ^ x125 ^ 1'b0 ;
  assign n28636 = ~n16818 & n20733 ;
  assign n28637 = n22210 ^ n8582 ^ 1'b0 ;
  assign n28638 = n13212 ^ n162 ^ 1'b0 ;
  assign n28639 = n28637 & ~n28638 ;
  assign n28640 = ~n17022 & n28639 ;
  assign n28641 = n28640 ^ n12167 ^ 1'b0 ;
  assign n28642 = ~n11235 & n21667 ;
  assign n28643 = ~n26856 & n28642 ;
  assign n28644 = ( ~n773 & n4110 ) | ( ~n773 & n4837 ) | ( n4110 & n4837 ) ;
  assign n28645 = n28644 ^ n12270 ^ 1'b0 ;
  assign n28646 = ~n3028 & n6048 ;
  assign n28647 = n7039 & n28646 ;
  assign n28648 = n5891 & ~n28647 ;
  assign n28649 = ( n2808 & n6250 ) | ( n2808 & ~n25940 ) | ( n6250 & ~n25940 ) ;
  assign n28650 = n28648 | n28649 ;
  assign n28651 = n25027 ^ n22386 ^ n9855 ;
  assign n28652 = n13473 & ~n16840 ;
  assign n28653 = ( ~n9922 & n22823 ) | ( ~n9922 & n28652 ) | ( n22823 & n28652 ) ;
  assign n28654 = n27453 ^ n22285 ^ n4836 ;
  assign n28656 = n3149 ^ n673 ^ 1'b0 ;
  assign n28655 = ~n4629 & n6161 ;
  assign n28657 = n28656 ^ n28655 ^ 1'b0 ;
  assign n28658 = ( n1602 & n2106 ) | ( n1602 & n12908 ) | ( n2106 & n12908 ) ;
  assign n28659 = ( n19066 & n24955 ) | ( n19066 & ~n25398 ) | ( n24955 & ~n25398 ) ;
  assign n28660 = ( x49 & x113 ) | ( x49 & ~n9644 ) | ( x113 & ~n9644 ) ;
  assign n28661 = n889 & ~n28660 ;
  assign n28662 = ( n8413 & n10252 ) | ( n8413 & n27332 ) | ( n10252 & n27332 ) ;
  assign n28663 = ( ~n8630 & n28661 ) | ( ~n8630 & n28662 ) | ( n28661 & n28662 ) ;
  assign n28664 = n9040 & n28663 ;
  assign n28665 = ~n28659 & n28664 ;
  assign n28666 = n24288 ^ n19365 ^ 1'b0 ;
  assign n28667 = n27281 ^ n3044 ^ 1'b0 ;
  assign n28668 = n8280 ^ n6434 ^ n2029 ;
  assign n28672 = n4142 ^ n984 ^ n491 ;
  assign n28670 = n7988 & n14760 ;
  assign n28671 = ~n13425 & n28670 ;
  assign n28669 = n15667 ^ n8114 ^ 1'b0 ;
  assign n28673 = n28672 ^ n28671 ^ n28669 ;
  assign n28674 = n755 & ~n851 ;
  assign n28675 = n28674 ^ n26149 ^ n12603 ;
  assign n28676 = n4727 ^ n739 ^ 1'b0 ;
  assign n28677 = n12871 & n24978 ;
  assign n28678 = n14149 & ~n28677 ;
  assign n28679 = ~n1326 & n19204 ;
  assign n28680 = n14654 ^ n2368 ^ 1'b0 ;
  assign n28681 = ( n1580 & n6135 ) | ( n1580 & ~n18589 ) | ( n6135 & ~n18589 ) ;
  assign n28682 = n265 | n11179 ;
  assign n28683 = n28681 & ~n28682 ;
  assign n28684 = n11749 ^ n5302 ^ 1'b0 ;
  assign n28685 = n2707 & ~n3861 ;
  assign n28686 = n28685 ^ n22422 ^ n11339 ;
  assign n28687 = ( n5382 & n6841 ) | ( n5382 & n16993 ) | ( n6841 & n16993 ) ;
  assign n28688 = n13363 ^ n9180 ^ 1'b0 ;
  assign n28689 = n7152 ^ n1463 ^ 1'b0 ;
  assign n28690 = ~n13607 & n28689 ;
  assign n28691 = n28690 ^ n25330 ^ 1'b0 ;
  assign n28692 = n1870 | n28691 ;
  assign n28693 = n18349 ^ n8770 ^ 1'b0 ;
  assign n28694 = n15785 | n28693 ;
  assign n28695 = n19111 ^ n820 ^ 1'b0 ;
  assign n28696 = n22267 & n28695 ;
  assign n28697 = n3806 | n7724 ;
  assign n28698 = n28697 ^ n15462 ^ n4215 ;
  assign n28699 = n28696 & n28698 ;
  assign n28700 = ( n9145 & n11661 ) | ( n9145 & n18857 ) | ( n11661 & n18857 ) ;
  assign n28701 = ( n2136 & n9928 ) | ( n2136 & ~n13499 ) | ( n9928 & ~n13499 ) ;
  assign n28704 = ~n4787 & n13393 ;
  assign n28705 = n28704 ^ n10472 ^ 1'b0 ;
  assign n28706 = ( n10496 & n23749 ) | ( n10496 & ~n28705 ) | ( n23749 & ~n28705 ) ;
  assign n28702 = n8704 & ~n18063 ;
  assign n28703 = n28702 ^ n2776 ^ 1'b0 ;
  assign n28707 = n28706 ^ n28703 ^ n17845 ;
  assign n28708 = n13334 ^ n3229 ^ 1'b0 ;
  assign n28709 = n24468 ^ n2453 ^ 1'b0 ;
  assign n28710 = n16321 ^ n6388 ^ 1'b0 ;
  assign n28711 = n17490 ^ n7771 ^ 1'b0 ;
  assign n28712 = n28711 ^ n15154 ^ 1'b0 ;
  assign n28713 = ~n315 & n28712 ;
  assign n28714 = n21137 ^ n16871 ^ 1'b0 ;
  assign n28715 = n858 & ~n28714 ;
  assign n28716 = ( n17762 & n20444 ) | ( n17762 & ~n21121 ) | ( n20444 & ~n21121 ) ;
  assign n28717 = n11746 ^ n9466 ^ 1'b0 ;
  assign n28718 = n4993 & n28717 ;
  assign n28719 = ( ~n12297 & n27517 ) | ( ~n12297 & n28718 ) | ( n27517 & n28718 ) ;
  assign n28720 = n25783 ^ n22552 ^ n5824 ;
  assign n28721 = n25908 ^ n11881 ^ 1'b0 ;
  assign n28722 = ( n4097 & n5827 ) | ( n4097 & ~n12472 ) | ( n5827 & ~n12472 ) ;
  assign n28724 = n8565 | n21956 ;
  assign n28723 = n14219 & n15165 ;
  assign n28725 = n28724 ^ n28723 ^ 1'b0 ;
  assign n28726 = ( ~n914 & n28722 ) | ( ~n914 & n28725 ) | ( n28722 & n28725 ) ;
  assign n28727 = n6067 & ~n22294 ;
  assign n28728 = n5097 ^ n3224 ^ 1'b0 ;
  assign n28729 = n28727 & n28728 ;
  assign n28730 = n8577 ^ n1968 ^ 1'b0 ;
  assign n28731 = ( ~n1198 & n3641 ) | ( ~n1198 & n15929 ) | ( n3641 & n15929 ) ;
  assign n28732 = ( n5867 & ~n8078 ) | ( n5867 & n28731 ) | ( ~n8078 & n28731 ) ;
  assign n28733 = n5255 & n28732 ;
  assign n28734 = n28733 ^ n14662 ^ 1'b0 ;
  assign n28735 = n7801 | n15563 ;
  assign n28736 = n28735 ^ n13748 ^ 1'b0 ;
  assign n28737 = n12425 & ~n18692 ;
  assign n28738 = n28737 ^ n1277 ^ 1'b0 ;
  assign n28739 = n1060 & ~n21299 ;
  assign n28740 = n18741 & n28739 ;
  assign n28741 = ( n5198 & n28738 ) | ( n5198 & ~n28740 ) | ( n28738 & ~n28740 ) ;
  assign n28742 = n18176 | n20231 ;
  assign n28743 = n18397 & ~n28742 ;
  assign n28744 = n3962 & n14526 ;
  assign n28745 = n13574 & n28744 ;
  assign n28746 = n28745 ^ n5670 ^ n824 ;
  assign n28747 = ~n21449 & n28746 ;
  assign n28748 = n28747 ^ n19264 ^ 1'b0 ;
  assign n28749 = n9186 & n10079 ;
  assign n28750 = ~n21560 & n28749 ;
  assign n28751 = n28750 ^ n5349 ^ 1'b0 ;
  assign n28752 = n23676 & n28751 ;
  assign n28753 = n28752 ^ n23777 ^ 1'b0 ;
  assign n28754 = ~n2779 & n17351 ;
  assign n28755 = n7692 ^ n4426 ^ 1'b0 ;
  assign n28756 = n16038 & ~n28755 ;
  assign n28757 = n3604 & ~n6986 ;
  assign n28758 = ~n18235 & n28757 ;
  assign n28759 = n13406 ^ n9850 ^ 1'b0 ;
  assign n28760 = n23528 ^ n17284 ^ n13353 ;
  assign n28761 = ( n8740 & ~n28759 ) | ( n8740 & n28760 ) | ( ~n28759 & n28760 ) ;
  assign n28762 = n8803 ^ n2417 ^ x69 ;
  assign n28763 = n28762 ^ n23527 ^ n6355 ;
  assign n28764 = n10689 ^ n2701 ^ 1'b0 ;
  assign n28765 = n8026 & ~n25300 ;
  assign n28766 = n28765 ^ n6452 ^ 1'b0 ;
  assign n28767 = n28766 ^ n16277 ^ 1'b0 ;
  assign n28768 = ( n7721 & n26699 ) | ( n7721 & n28767 ) | ( n26699 & n28767 ) ;
  assign n28769 = ( n13961 & ~n14466 ) | ( n13961 & n22722 ) | ( ~n14466 & n22722 ) ;
  assign n28770 = n1333 & ~n5798 ;
  assign n28771 = n10613 & n28770 ;
  assign n28772 = n10230 & ~n13656 ;
  assign n28773 = ~x59 & n28772 ;
  assign n28774 = n12616 ^ n556 ^ 1'b0 ;
  assign n28775 = ~n28773 & n28774 ;
  assign n28776 = n5247 | n12309 ;
  assign n28777 = n28776 ^ x94 ^ 1'b0 ;
  assign n28778 = n171 & n28777 ;
  assign n28779 = n28778 ^ n10381 ^ 1'b0 ;
  assign n28780 = n10504 ^ n2468 ^ 1'b0 ;
  assign n28781 = n25387 ^ n2033 ^ 1'b0 ;
  assign n28782 = ~n13223 & n28781 ;
  assign n28783 = n9411 & n28782 ;
  assign n28784 = n861 & n28783 ;
  assign n28785 = ( ~n12892 & n20598 ) | ( ~n12892 & n20612 ) | ( n20598 & n20612 ) ;
  assign n28786 = n28289 ^ n8735 ^ n154 ;
  assign n28787 = n15014 ^ n14023 ^ 1'b0 ;
  assign n28788 = n1620 & ~n16570 ;
  assign n28789 = n15916 ^ n15547 ^ n6274 ;
  assign n28790 = n24533 ^ n15467 ^ 1'b0 ;
  assign n28791 = n17014 | n28790 ;
  assign n28792 = n2905 | n14691 ;
  assign n28793 = n3264 & ~n8084 ;
  assign n28794 = ~n28792 & n28793 ;
  assign n28795 = n21415 & ~n26447 ;
  assign n28796 = n28795 ^ n1475 ^ 1'b0 ;
  assign n28797 = n8349 & ~n28796 ;
  assign n28798 = n28797 ^ n6841 ^ 1'b0 ;
  assign n28799 = ( n9347 & n15875 ) | ( n9347 & n22919 ) | ( n15875 & n22919 ) ;
  assign n28800 = ( ~n16109 & n25908 ) | ( ~n16109 & n28799 ) | ( n25908 & n28799 ) ;
  assign n28801 = ~n18470 & n23793 ;
  assign n28802 = ( n687 & ~n8058 ) | ( n687 & n24922 ) | ( ~n8058 & n24922 ) ;
  assign n28803 = n6662 & ~n28802 ;
  assign n28804 = n2724 ^ n1732 ^ n1254 ;
  assign n28805 = n28804 ^ n6419 ^ 1'b0 ;
  assign n28806 = n4378 | n7705 ;
  assign n28807 = n5249 & ~n28806 ;
  assign n28808 = n24869 ^ n12045 ^ 1'b0 ;
  assign n28809 = n6886 & ~n24170 ;
  assign n28810 = n28809 ^ n15600 ^ 1'b0 ;
  assign n28811 = n16924 ^ n6196 ^ 1'b0 ;
  assign n28812 = ( n777 & n14023 ) | ( n777 & ~n16268 ) | ( n14023 & ~n16268 ) ;
  assign n28813 = n28812 ^ n2122 ^ 1'b0 ;
  assign n28814 = ~n3214 & n6308 ;
  assign n28815 = n28814 ^ n16647 ^ n1538 ;
  assign n28816 = ( ~n6128 & n7494 ) | ( ~n6128 & n25119 ) | ( n7494 & n25119 ) ;
  assign n28817 = n12497 | n28816 ;
  assign n28818 = n1547 & n4261 ;
  assign n28819 = ( n275 & ~n738 ) | ( n275 & n7335 ) | ( ~n738 & n7335 ) ;
  assign n28820 = n4723 ^ n3437 ^ 1'b0 ;
  assign n28821 = ( n28818 & n28819 ) | ( n28818 & ~n28820 ) | ( n28819 & ~n28820 ) ;
  assign n28822 = n10836 | n22589 ;
  assign n28823 = n28822 ^ n23721 ^ 1'b0 ;
  assign n28824 = n16091 | n28823 ;
  assign n28825 = n28824 ^ n3151 ^ 1'b0 ;
  assign n28826 = n4712 ^ n3511 ^ 1'b0 ;
  assign n28827 = n19189 & n28826 ;
  assign n28829 = n10263 & ~n13595 ;
  assign n28828 = ~n502 & n11198 ;
  assign n28830 = n28829 ^ n28828 ^ 1'b0 ;
  assign n28832 = ( ~n659 & n2774 ) | ( ~n659 & n6730 ) | ( n2774 & n6730 ) ;
  assign n28831 = n5863 | n24866 ;
  assign n28833 = n28832 ^ n28831 ^ 1'b0 ;
  assign n28834 = n28833 ^ n27099 ^ 1'b0 ;
  assign n28835 = n14301 ^ n5450 ^ n1205 ;
  assign n28836 = n20429 ^ n20192 ^ 1'b0 ;
  assign n28837 = n188 & n13295 ;
  assign n28838 = n17839 & ~n21229 ;
  assign n28839 = ( ~n619 & n9092 ) | ( ~n619 & n16167 ) | ( n9092 & n16167 ) ;
  assign n28840 = ( n28837 & n28838 ) | ( n28837 & ~n28839 ) | ( n28838 & ~n28839 ) ;
  assign n28841 = ( ~n3447 & n4148 ) | ( ~n3447 & n10585 ) | ( n4148 & n10585 ) ;
  assign n28842 = ( ~n2718 & n15354 ) | ( ~n2718 & n28841 ) | ( n15354 & n28841 ) ;
  assign n28843 = n12936 ^ n9754 ^ 1'b0 ;
  assign n28844 = n17752 & n28843 ;
  assign n28845 = ~n3273 & n4115 ;
  assign n28846 = n2972 ^ n158 ^ 1'b0 ;
  assign n28847 = n15675 | n25930 ;
  assign n28848 = n28847 ^ n8062 ^ 1'b0 ;
  assign n28849 = n11784 | n28848 ;
  assign n28850 = n24321 ^ n6120 ^ 1'b0 ;
  assign n28851 = n9678 & ~n23339 ;
  assign n28852 = n12779 & n28851 ;
  assign n28853 = n28852 ^ n11423 ^ 1'b0 ;
  assign n28854 = ( n15168 & n25743 ) | ( n15168 & ~n28853 ) | ( n25743 & ~n28853 ) ;
  assign n28855 = n482 & n17602 ;
  assign n28856 = n28855 ^ n1571 ^ 1'b0 ;
  assign n28857 = n26829 ^ n15191 ^ n7913 ;
  assign n28858 = ( n9068 & n14815 ) | ( n9068 & n15026 ) | ( n14815 & n15026 ) ;
  assign n28859 = n6483 & n14420 ;
  assign n28860 = n28859 ^ n18935 ^ 1'b0 ;
  assign n28861 = ( n1723 & n7296 ) | ( n1723 & ~n17228 ) | ( n7296 & ~n17228 ) ;
  assign n28862 = ( n26384 & n28860 ) | ( n26384 & n28861 ) | ( n28860 & n28861 ) ;
  assign n28863 = ( n5323 & ~n15253 ) | ( n5323 & n16233 ) | ( ~n15253 & n16233 ) ;
  assign n28864 = n2217 & n10160 ;
  assign n28865 = n1196 & n25535 ;
  assign n28866 = ( n6426 & ~n8752 ) | ( n6426 & n24227 ) | ( ~n8752 & n24227 ) ;
  assign n28867 = n11992 | n28866 ;
  assign n28868 = n11199 & ~n19425 ;
  assign n28869 = n28679 & n28868 ;
  assign n28870 = n28867 & n28869 ;
  assign n28871 = n2963 & ~n12603 ;
  assign n28872 = n26039 | n28871 ;
  assign n28873 = n20188 ^ n4576 ^ 1'b0 ;
  assign n28874 = n11521 ^ n7249 ^ 1'b0 ;
  assign n28875 = n22654 ^ n13222 ^ n8607 ;
  assign n28877 = n10553 & n28644 ;
  assign n28878 = n15442 & n28877 ;
  assign n28876 = n2929 & ~n17171 ;
  assign n28879 = n28878 ^ n28876 ^ 1'b0 ;
  assign n28880 = n28879 ^ n28475 ^ 1'b0 ;
  assign n28881 = n3167 & ~n16959 ;
  assign n28882 = n13363 & n28881 ;
  assign n28883 = n26542 ^ n10838 ^ 1'b0 ;
  assign n28884 = n1531 & ~n28883 ;
  assign n28885 = n4462 ^ n3004 ^ 1'b0 ;
  assign n28888 = ( n994 & n5071 ) | ( n994 & ~n8957 ) | ( n5071 & ~n8957 ) ;
  assign n28889 = ( n149 & ~n6754 ) | ( n149 & n28888 ) | ( ~n6754 & n28888 ) ;
  assign n28886 = n403 | n27772 ;
  assign n28887 = n28886 ^ n4972 ^ 1'b0 ;
  assign n28890 = n28889 ^ n28887 ^ n17989 ;
  assign n28891 = n28890 ^ n12723 ^ 1'b0 ;
  assign n28892 = n28885 & n28891 ;
  assign n28893 = ( ~n5900 & n9056 ) | ( ~n5900 & n10033 ) | ( n9056 & n10033 ) ;
  assign n28894 = n2239 ^ n1283 ^ n859 ;
  assign n28895 = ~n8746 & n11273 ;
  assign n28896 = n28895 ^ n6710 ^ 1'b0 ;
  assign n28897 = n10678 | n28896 ;
  assign n28898 = n19008 ^ n6317 ^ n4192 ;
  assign n28899 = n28898 ^ n17102 ^ 1'b0 ;
  assign n28900 = n16875 | n20991 ;
  assign n28901 = n28900 ^ n6586 ^ 1'b0 ;
  assign n28902 = n11883 ^ n346 ^ 1'b0 ;
  assign n28904 = n8460 & ~n13933 ;
  assign n28903 = ( n3371 & n5498 ) | ( n3371 & ~n17943 ) | ( n5498 & ~n17943 ) ;
  assign n28905 = n28904 ^ n28903 ^ 1'b0 ;
  assign n28906 = n28902 & n28905 ;
  assign n28907 = n22590 & ~n28906 ;
  assign n28908 = ~n17952 & n25661 ;
  assign n28909 = n21283 ^ n3442 ^ 1'b0 ;
  assign n28910 = n2316 | n28909 ;
  assign n28911 = n18506 ^ n13296 ^ n10306 ;
  assign n28912 = ( n6737 & n22638 ) | ( n6737 & n24661 ) | ( n22638 & n24661 ) ;
  assign n28913 = ~n7449 & n28853 ;
  assign n28914 = n16288 ^ n5488 ^ 1'b0 ;
  assign n28915 = n11234 ^ n4619 ^ 1'b0 ;
  assign n28916 = ~n6918 & n19119 ;
  assign n28917 = n12853 & n28916 ;
  assign n28919 = n14726 ^ n12526 ^ n1082 ;
  assign n28918 = n380 & ~n4064 ;
  assign n28920 = n28919 ^ n28918 ^ 1'b0 ;
  assign n28921 = n16067 | n28920 ;
  assign n28922 = n4771 | n28656 ;
  assign n28923 = n10872 | n28922 ;
  assign n28924 = n18355 & ~n28923 ;
  assign n28925 = n22293 ^ n17536 ^ 1'b0 ;
  assign n28926 = n28924 | n28925 ;
  assign n28927 = n13567 | n15675 ;
  assign n28928 = n28927 ^ n20222 ^ 1'b0 ;
  assign n28929 = n27024 ^ n15231 ^ 1'b0 ;
  assign n28930 = n13525 ^ n7285 ^ 1'b0 ;
  assign n28931 = n17983 ^ n15795 ^ 1'b0 ;
  assign n28932 = ~n8727 & n11339 ;
  assign n28933 = n28932 ^ n8196 ^ 1'b0 ;
  assign n28934 = n28933 ^ n784 ^ n374 ;
  assign n28935 = n12583 ^ n12522 ^ n8830 ;
  assign n28936 = n27198 ^ n7002 ^ n6903 ;
  assign n28937 = n15976 ^ n5932 ^ 1'b0 ;
  assign n28938 = n21397 ^ n20886 ^ 1'b0 ;
  assign n28939 = n4397 | n28938 ;
  assign n28940 = n341 | n28939 ;
  assign n28941 = ~n6227 & n28940 ;
  assign n28942 = n28941 ^ n4677 ^ 1'b0 ;
  assign n28943 = n8495 | n28942 ;
  assign n28944 = ~n6187 & n6981 ;
  assign n28945 = ~n12383 & n15465 ;
  assign n28946 = n8593 | n24887 ;
  assign n28947 = n28946 ^ n5156 ^ 1'b0 ;
  assign n28949 = ( n6624 & n8302 ) | ( n6624 & n25286 ) | ( n8302 & n25286 ) ;
  assign n28948 = n25427 ^ n12747 ^ 1'b0 ;
  assign n28950 = n28949 ^ n28948 ^ n27654 ;
  assign n28951 = ( n3819 & n5728 ) | ( n3819 & n28950 ) | ( n5728 & n28950 ) ;
  assign n28952 = ( n14901 & ~n15462 ) | ( n14901 & n16172 ) | ( ~n15462 & n16172 ) ;
  assign n28953 = n7317 | n7795 ;
  assign n28954 = ( n6532 & n9506 ) | ( n6532 & ~n9875 ) | ( n9506 & ~n9875 ) ;
  assign n28955 = n4628 & ~n28954 ;
  assign n28956 = n28955 ^ n15275 ^ 1'b0 ;
  assign n28957 = n28956 ^ n10242 ^ 1'b0 ;
  assign n28964 = n5633 ^ n783 ^ 1'b0 ;
  assign n28961 = n8162 & n13903 ;
  assign n28962 = n6908 & n28961 ;
  assign n28963 = n28962 ^ n4501 ^ 1'b0 ;
  assign n28965 = n28964 ^ n28963 ^ 1'b0 ;
  assign n28958 = n880 | n23253 ;
  assign n28959 = n4388 & ~n28958 ;
  assign n28960 = n28959 ^ n936 ^ 1'b0 ;
  assign n28966 = n28965 ^ n28960 ^ x35 ;
  assign n28967 = n23734 ^ n17481 ^ n14887 ;
  assign n28968 = n22779 | n28967 ;
  assign n28969 = n16953 | n19986 ;
  assign n28970 = n28968 & ~n28969 ;
  assign n28971 = n17776 | n28970 ;
  assign n28972 = n1702 | n28660 ;
  assign n28973 = n28972 ^ n3858 ^ 1'b0 ;
  assign n28975 = ( n831 & n4094 ) | ( n831 & ~n14469 ) | ( n4094 & ~n14469 ) ;
  assign n28974 = n3027 & ~n14806 ;
  assign n28976 = n28975 ^ n28974 ^ n15493 ;
  assign n28977 = n2561 | n28976 ;
  assign n28978 = n752 & ~n28977 ;
  assign n28979 = n28978 ^ n27158 ^ n4867 ;
  assign n28980 = n14144 ^ n3791 ^ 1'b0 ;
  assign n28981 = n28979 & n28980 ;
  assign n28982 = n23736 ^ n4367 ^ 1'b0 ;
  assign n28983 = ( n3648 & ~n6239 ) | ( n3648 & n11286 ) | ( ~n6239 & n11286 ) ;
  assign n28984 = n28983 ^ n12147 ^ 1'b0 ;
  assign n28987 = n7563 | n9224 ;
  assign n28985 = n1561 ^ n1213 ^ 1'b0 ;
  assign n28986 = n10181 & n28985 ;
  assign n28988 = n28987 ^ n28986 ^ 1'b0 ;
  assign n28989 = n22775 ^ n18827 ^ n16816 ;
  assign n28990 = n1866 & n4733 ;
  assign n28991 = ( n1907 & ~n8560 ) | ( n1907 & n28990 ) | ( ~n8560 & n28990 ) ;
  assign n28992 = ~n5049 & n18366 ;
  assign n28993 = ( n1754 & ~n9319 ) | ( n1754 & n28992 ) | ( ~n9319 & n28992 ) ;
  assign n28994 = n28993 ^ n209 ^ 1'b0 ;
  assign n28995 = n11361 ^ n9651 ^ 1'b0 ;
  assign n28996 = ~n2796 & n28995 ;
  assign n28997 = ~n25670 & n28996 ;
  assign n28998 = n26945 ^ n8574 ^ n367 ;
  assign n28999 = ~n1355 & n28998 ;
  assign n29000 = n28999 ^ n3872 ^ 1'b0 ;
  assign n29001 = n4055 & ~n6030 ;
  assign n29002 = n14233 | n17988 ;
  assign n29003 = n29001 | n29002 ;
  assign n29004 = ~n3720 & n8517 ;
  assign n29005 = n29004 ^ n16418 ^ 1'b0 ;
  assign n29006 = n5598 & ~n29005 ;
  assign n29007 = n516 & ~n28383 ;
  assign n29008 = n1310 & n29007 ;
  assign n29009 = n29008 ^ n11544 ^ 1'b0 ;
  assign n29010 = n29009 ^ n3169 ^ n2421 ;
  assign n29011 = n29010 ^ n26005 ^ 1'b0 ;
  assign n29012 = ( n3533 & n14041 ) | ( n3533 & n18881 ) | ( n14041 & n18881 ) ;
  assign n29013 = ( x120 & ~n11481 ) | ( x120 & n29012 ) | ( ~n11481 & n29012 ) ;
  assign n29014 = n20492 ^ n11871 ^ n8368 ;
  assign n29015 = n11250 ^ n10018 ^ 1'b0 ;
  assign n29016 = n17228 | n22577 ;
  assign n29017 = n29016 ^ n8493 ^ 1'b0 ;
  assign n29018 = ( n1934 & n6668 ) | ( n1934 & n29017 ) | ( n6668 & n29017 ) ;
  assign n29020 = ( n3971 & n17089 ) | ( n3971 & n28661 ) | ( n17089 & n28661 ) ;
  assign n29019 = n8109 ^ n6344 ^ n2715 ;
  assign n29021 = n29020 ^ n29019 ^ 1'b0 ;
  assign n29022 = n3736 | n12772 ;
  assign n29023 = ~n835 & n3631 ;
  assign n29024 = n29023 ^ n363 ^ 1'b0 ;
  assign n29025 = n13337 ^ n7624 ^ n5133 ;
  assign n29026 = n7943 & ~n29025 ;
  assign n29027 = n10067 & ~n29026 ;
  assign n29028 = n29027 ^ n807 ^ 1'b0 ;
  assign n29029 = n11531 | n25772 ;
  assign n29030 = n29028 & ~n29029 ;
  assign n29031 = n7190 & n7774 ;
  assign n29032 = n4766 & ~n18798 ;
  assign n29033 = n29032 ^ n5969 ^ 1'b0 ;
  assign n29034 = n29033 ^ n10539 ^ n2648 ;
  assign n29035 = n8650 & n29034 ;
  assign n29036 = n29035 ^ n12306 ^ 1'b0 ;
  assign n29037 = ~n18550 & n21334 ;
  assign n29038 = n29037 ^ n538 ^ 1'b0 ;
  assign n29039 = ( n1292 & ~n17553 ) | ( n1292 & n28972 ) | ( ~n17553 & n28972 ) ;
  assign n29040 = ~n3206 & n11118 ;
  assign n29041 = ( n4280 & n23149 ) | ( n4280 & ~n29040 ) | ( n23149 & ~n29040 ) ;
  assign n29042 = n17419 ^ n15023 ^ 1'b0 ;
  assign n29043 = ~n27514 & n29042 ;
  assign n29044 = ( n238 & n13560 ) | ( n238 & n29043 ) | ( n13560 & n29043 ) ;
  assign n29045 = n11812 ^ n2449 ^ 1'b0 ;
  assign n29046 = ~n1329 & n29045 ;
  assign n29047 = n19120 ^ n1634 ^ 1'b0 ;
  assign n29048 = n22488 & n29047 ;
  assign n29049 = n2699 & n29048 ;
  assign n29050 = n23748 & n29049 ;
  assign n29051 = n15700 ^ n1674 ^ 1'b0 ;
  assign n29052 = n5213 & n6525 ;
  assign n29053 = n29052 ^ n2462 ^ 1'b0 ;
  assign n29054 = n6455 ^ n6048 ^ 1'b0 ;
  assign n29055 = n27380 ^ n11542 ^ 1'b0 ;
  assign n29056 = n29054 & n29055 ;
  assign n29059 = n8735 & n26323 ;
  assign n29057 = ( ~n1217 & n16944 ) | ( ~n1217 & n17998 ) | ( n16944 & n17998 ) ;
  assign n29058 = n4528 & ~n29057 ;
  assign n29060 = n29059 ^ n29058 ^ 1'b0 ;
  assign n29064 = n3087 & ~n5535 ;
  assign n29062 = n11292 ^ n8757 ^ n6572 ;
  assign n29061 = n2322 | n3132 ;
  assign n29063 = n29062 ^ n29061 ^ n9103 ;
  assign n29065 = n29064 ^ n29063 ^ n12346 ;
  assign n29066 = ( n415 & n4616 ) | ( n415 & ~n21277 ) | ( n4616 & ~n21277 ) ;
  assign n29067 = n2289 & ~n13695 ;
  assign n29068 = ~n8596 & n29067 ;
  assign n29069 = n22590 | n29068 ;
  assign n29070 = n29069 ^ n27946 ^ n18782 ;
  assign n29071 = n12573 | n29070 ;
  assign n29072 = n14213 | n29071 ;
  assign n29073 = ( n29065 & ~n29066 ) | ( n29065 & n29072 ) | ( ~n29066 & n29072 ) ;
  assign n29074 = n12137 ^ n633 ^ 1'b0 ;
  assign n29075 = n13856 | n29074 ;
  assign n29076 = ~n3481 & n6672 ;
  assign n29077 = n29076 ^ n20365 ^ n1447 ;
  assign n29078 = ( n6927 & n29075 ) | ( n6927 & ~n29077 ) | ( n29075 & ~n29077 ) ;
  assign n29079 = n16091 ^ n15527 ^ 1'b0 ;
  assign n29080 = n29079 ^ n21278 ^ n4897 ;
  assign n29081 = n9859 ^ n2738 ^ 1'b0 ;
  assign n29082 = n3152 & n15995 ;
  assign n29083 = ~n11837 & n29082 ;
  assign n29084 = ( n2003 & n29081 ) | ( n2003 & ~n29083 ) | ( n29081 & ~n29083 ) ;
  assign n29085 = n3525 ^ n3198 ^ 1'b0 ;
  assign n29086 = n2428 & n29085 ;
  assign n29087 = n15910 & n29086 ;
  assign n29088 = n7145 & ~n26988 ;
  assign n29089 = n21627 ^ n19310 ^ 1'b0 ;
  assign n29090 = ~n18294 & n29089 ;
  assign n29091 = n7798 ^ n2142 ^ 1'b0 ;
  assign n29092 = n15319 | n29091 ;
  assign n29094 = n16620 ^ n10708 ^ n789 ;
  assign n29093 = n12927 & n13915 ;
  assign n29095 = n29094 ^ n29093 ^ 1'b0 ;
  assign n29096 = ( n4933 & n6065 ) | ( n4933 & ~n10104 ) | ( n6065 & ~n10104 ) ;
  assign n29097 = n3524 & n16378 ;
  assign n29098 = n29096 & n29097 ;
  assign n29099 = ( ~n2867 & n7885 ) | ( ~n2867 & n29098 ) | ( n7885 & n29098 ) ;
  assign n29100 = n18152 & ~n29099 ;
  assign n29102 = n10539 ^ n1534 ^ 1'b0 ;
  assign n29103 = n1040 & n29102 ;
  assign n29101 = ~n11206 & n24843 ;
  assign n29104 = n29103 ^ n29101 ^ 1'b0 ;
  assign n29105 = n29104 ^ n15258 ^ n7838 ;
  assign n29106 = ( n4931 & n7003 ) | ( n4931 & n18688 ) | ( n7003 & n18688 ) ;
  assign n29107 = ~n623 & n9178 ;
  assign n29108 = n29107 ^ n6884 ^ 1'b0 ;
  assign n29109 = n29108 ^ n21227 ^ n18063 ;
  assign n29110 = ( n451 & n5432 ) | ( n451 & ~n15998 ) | ( n5432 & ~n15998 ) ;
  assign n29111 = n29110 ^ n24240 ^ 1'b0 ;
  assign n29112 = n5381 ^ n1003 ^ 1'b0 ;
  assign n29113 = ~n13937 & n25330 ;
  assign n29114 = ~n2191 & n9277 ;
  assign n29115 = n29114 ^ n20845 ^ 1'b0 ;
  assign n29116 = n22141 ^ n9220 ^ 1'b0 ;
  assign n29117 = n21540 ^ n6216 ^ 1'b0 ;
  assign n29118 = n8616 ^ n7882 ^ n4464 ;
  assign n29119 = n29118 ^ n13555 ^ 1'b0 ;
  assign n29120 = n29119 ^ n14560 ^ n6972 ;
  assign n29121 = ( n428 & ~n2434 ) | ( n428 & n10508 ) | ( ~n2434 & n10508 ) ;
  assign n29122 = n16071 ^ n15958 ^ 1'b0 ;
  assign n29124 = n728 & n1542 ;
  assign n29125 = ~n2868 & n29124 ;
  assign n29123 = ~x112 & n9574 ;
  assign n29126 = n29125 ^ n29123 ^ 1'b0 ;
  assign n29127 = n17875 | n29126 ;
  assign n29128 = n1772 ^ n1319 ^ 1'b0 ;
  assign n29129 = n7790 | n29128 ;
  assign n29130 = n23571 & ~n29129 ;
  assign n29131 = n14096 | n21951 ;
  assign n29132 = n29131 ^ n1076 ^ 1'b0 ;
  assign n29133 = ( x21 & n6692 ) | ( x21 & ~n20524 ) | ( n6692 & ~n20524 ) ;
  assign n29134 = n5702 & ~n29133 ;
  assign n29135 = n17894 ^ n598 ^ 1'b0 ;
  assign n29136 = ( x11 & n5941 ) | ( x11 & n19866 ) | ( n5941 & n19866 ) ;
  assign n29137 = ( ~n13433 & n29135 ) | ( ~n13433 & n29136 ) | ( n29135 & n29136 ) ;
  assign n29138 = n17703 ^ n6208 ^ 1'b0 ;
  assign n29139 = ~n19648 & n29138 ;
  assign n29140 = n29139 ^ n5576 ^ n3990 ;
  assign n29141 = n24671 ^ n21434 ^ 1'b0 ;
  assign n29142 = n10300 & ~n25745 ;
  assign n29143 = n3503 | n16879 ;
  assign n29144 = n20867 & ~n29143 ;
  assign n29145 = n9505 ^ n2498 ^ 1'b0 ;
  assign n29146 = n29144 | n29145 ;
  assign n29147 = n16642 ^ n11546 ^ 1'b0 ;
  assign n29148 = n5261 | n29147 ;
  assign n29149 = n3935 ^ n3162 ^ 1'b0 ;
  assign n29150 = n12497 | n29149 ;
  assign n29151 = ( n1693 & n8352 ) | ( n1693 & ~n15466 ) | ( n8352 & ~n15466 ) ;
  assign n29152 = n9108 & n21415 ;
  assign n29153 = ~n6789 & n19495 ;
  assign n29154 = ( n18161 & n25685 ) | ( n18161 & ~n29153 ) | ( n25685 & ~n29153 ) ;
  assign n29155 = ( n29151 & n29152 ) | ( n29151 & ~n29154 ) | ( n29152 & ~n29154 ) ;
  assign n29156 = n11392 & ~n12549 ;
  assign n29157 = n14785 ^ n1779 ^ 1'b0 ;
  assign n29158 = n29157 ^ n13140 ^ n5601 ;
  assign n29159 = n16609 ^ n11100 ^ n468 ;
  assign n29160 = n29159 ^ n10510 ^ n8078 ;
  assign n29161 = n13566 ^ n13413 ^ 1'b0 ;
  assign n29162 = n3314 & n17945 ;
  assign n29163 = n29162 ^ n16706 ^ 1'b0 ;
  assign n29166 = n26149 ^ n13647 ^ 1'b0 ;
  assign n29167 = ~n26430 & n29166 ;
  assign n29168 = ~n26897 & n29167 ;
  assign n29164 = n9149 ^ n4396 ^ n2415 ;
  assign n29165 = n20950 & n29164 ;
  assign n29169 = n29168 ^ n29165 ^ 1'b0 ;
  assign n29170 = n23750 ^ n11526 ^ 1'b0 ;
  assign n29171 = n13201 | n29170 ;
  assign n29172 = n3052 & ~n11267 ;
  assign n29173 = ~n10282 & n29172 ;
  assign n29174 = n29173 ^ n6740 ^ n1090 ;
  assign n29175 = n28264 ^ n18096 ^ 1'b0 ;
  assign n29176 = n10108 ^ n8718 ^ n7943 ;
  assign n29177 = n24059 ^ n10538 ^ n9526 ;
  assign n29178 = n13927 ^ n7002 ^ n6057 ;
  assign n29179 = ( ~n8516 & n16658 ) | ( ~n8516 & n29178 ) | ( n16658 & n29178 ) ;
  assign n29180 = n29179 ^ n13886 ^ 1'b0 ;
  assign n29181 = n23853 ^ n3439 ^ n2017 ;
  assign n29182 = n29180 & n29181 ;
  assign n29183 = ( ~n12223 & n29177 ) | ( ~n12223 & n29182 ) | ( n29177 & n29182 ) ;
  assign n29184 = ( n10219 & n14399 ) | ( n10219 & n29183 ) | ( n14399 & n29183 ) ;
  assign n29185 = n5116 & ~n14868 ;
  assign n29186 = n143 & ~n17124 ;
  assign n29187 = n29186 ^ n5312 ^ n1700 ;
  assign n29188 = ( n5360 & n9098 ) | ( n5360 & ~n21913 ) | ( n9098 & ~n21913 ) ;
  assign n29189 = n9448 | n27498 ;
  assign n29190 = n28528 & ~n29189 ;
  assign n29191 = n29190 ^ n4810 ^ 1'b0 ;
  assign n29192 = n29188 & n29191 ;
  assign n29193 = n12001 | n23024 ;
  assign n29194 = n22151 ^ n18056 ^ n2776 ;
  assign n29195 = n25729 ^ n14842 ^ n2257 ;
  assign n29196 = n11253 & n16987 ;
  assign n29197 = n5857 | n29196 ;
  assign n29198 = ~n12730 & n18447 ;
  assign n29199 = ~n5897 & n29198 ;
  assign n29200 = n8286 & ~n29199 ;
  assign n29201 = ~n24299 & n29200 ;
  assign n29202 = n29201 ^ n8921 ^ 1'b0 ;
  assign n29203 = n26911 ^ n26540 ^ 1'b0 ;
  assign n29204 = ~n264 & n29203 ;
  assign n29205 = n7349 ^ n533 ^ 1'b0 ;
  assign n29206 = ~n12647 & n29205 ;
  assign n29207 = n21583 ^ n20894 ^ 1'b0 ;
  assign n29208 = n29206 & ~n29207 ;
  assign n29209 = n28138 ^ n16153 ^ 1'b0 ;
  assign n29210 = n16378 & n29209 ;
  assign n29211 = n194 & n14346 ;
  assign n29212 = ~n18589 & n29211 ;
  assign n29213 = n17034 ^ n2000 ^ 1'b0 ;
  assign n29214 = ~n5471 & n29213 ;
  assign n29215 = n28792 ^ n4401 ^ 1'b0 ;
  assign n29216 = n308 | n6594 ;
  assign n29217 = n29216 ^ n9862 ^ n7367 ;
  assign n29218 = ~n8029 & n29217 ;
  assign n29219 = ( n8724 & n10440 ) | ( n8724 & ~n29218 ) | ( n10440 & ~n29218 ) ;
  assign n29220 = n19901 ^ n158 ^ 1'b0 ;
  assign n29221 = ~n743 & n9346 ;
  assign n29222 = ( n26165 & ~n27358 ) | ( n26165 & n29221 ) | ( ~n27358 & n29221 ) ;
  assign n29223 = n26745 ^ n291 ^ 1'b0 ;
  assign n29224 = ~n3633 & n29223 ;
  assign n29225 = n10568 ^ n2309 ^ 1'b0 ;
  assign n29226 = n4856 | n29225 ;
  assign n29227 = n15894 ^ n6974 ^ 1'b0 ;
  assign n29228 = n874 | n29227 ;
  assign n29229 = n767 | n29228 ;
  assign n29230 = n16966 ^ n9427 ^ n2423 ;
  assign n29233 = ( ~n13110 & n14758 ) | ( ~n13110 & n27661 ) | ( n14758 & n27661 ) ;
  assign n29231 = n188 ^ n154 ^ 1'b0 ;
  assign n29232 = ~n9268 & n29231 ;
  assign n29234 = n29233 ^ n29232 ^ n1905 ;
  assign n29237 = n20841 ^ n6418 ^ 1'b0 ;
  assign n29235 = n11091 & ~n13797 ;
  assign n29236 = n29235 ^ n27160 ^ 1'b0 ;
  assign n29238 = n29237 ^ n29236 ^ n15995 ;
  assign n29242 = ( n6331 & ~n9914 ) | ( n6331 & n20261 ) | ( ~n9914 & n20261 ) ;
  assign n29241 = ( n7465 & n7744 ) | ( n7465 & n21385 ) | ( n7744 & n21385 ) ;
  assign n29239 = n3943 & n16563 ;
  assign n29240 = n29239 ^ n10954 ^ 1'b0 ;
  assign n29243 = n29242 ^ n29241 ^ n29240 ;
  assign n29244 = n11696 | n29243 ;
  assign n29245 = n8843 ^ n1150 ^ 1'b0 ;
  assign n29246 = ( n6386 & n24931 ) | ( n6386 & n29245 ) | ( n24931 & n29245 ) ;
  assign n29248 = n5251 & n6655 ;
  assign n29249 = n29248 ^ n1617 ^ 1'b0 ;
  assign n29250 = ~x11 & n29249 ;
  assign n29247 = n9149 & ~n9773 ;
  assign n29251 = n29250 ^ n29247 ^ 1'b0 ;
  assign n29252 = n10404 & n29251 ;
  assign n29253 = ~n8748 & n29252 ;
  assign n29254 = n11738 & n19287 ;
  assign n29255 = ~n6625 & n29254 ;
  assign n29256 = n29255 ^ n17000 ^ 1'b0 ;
  assign n29257 = n20270 ^ n4211 ^ 1'b0 ;
  assign n29258 = ~n8318 & n11537 ;
  assign n29259 = ~n13222 & n29258 ;
  assign n29260 = n4048 & ~n28277 ;
  assign n29261 = n29260 ^ n26323 ^ 1'b0 ;
  assign n29262 = n16753 & ~n29261 ;
  assign n29263 = n3491 & n7853 ;
  assign n29264 = n12456 | n19645 ;
  assign n29265 = n18070 & ~n29264 ;
  assign n29266 = ( ~n9036 & n9384 ) | ( ~n9036 & n29265 ) | ( n9384 & n29265 ) ;
  assign n29267 = ( ~n4185 & n29263 ) | ( ~n4185 & n29266 ) | ( n29263 & n29266 ) ;
  assign n29269 = n7180 ^ n2782 ^ 1'b0 ;
  assign n29268 = ( n5832 & ~n26056 ) | ( n5832 & n29260 ) | ( ~n26056 & n29260 ) ;
  assign n29270 = n29269 ^ n29268 ^ n19847 ;
  assign n29271 = n5364 & n14444 ;
  assign n29272 = ~n5116 & n9165 ;
  assign n29273 = ~n7616 & n19510 ;
  assign n29274 = n29273 ^ n23366 ^ 1'b0 ;
  assign n29275 = n1320 | n3888 ;
  assign n29276 = n12183 & ~n29275 ;
  assign n29277 = n13060 & ~n24048 ;
  assign n29278 = n23721 ^ n8501 ^ x100 ;
  assign n29279 = n29278 ^ n20417 ^ n6730 ;
  assign n29280 = n350 & ~n862 ;
  assign n29281 = ( n16746 & ~n19698 ) | ( n16746 & n29280 ) | ( ~n19698 & n29280 ) ;
  assign n29282 = ( n2093 & n3556 ) | ( n2093 & n5641 ) | ( n3556 & n5641 ) ;
  assign n29283 = ~n4561 & n6486 ;
  assign n29284 = n29283 ^ x69 ^ 1'b0 ;
  assign n29285 = ( n1785 & n2639 ) | ( n1785 & ~n29284 ) | ( n2639 & ~n29284 ) ;
  assign n29286 = ( n8805 & n29282 ) | ( n8805 & ~n29285 ) | ( n29282 & ~n29285 ) ;
  assign n29287 = n25551 ^ n23089 ^ n6959 ;
  assign n29288 = ( ~n20988 & n24281 ) | ( ~n20988 & n29287 ) | ( n24281 & n29287 ) ;
  assign n29289 = n3838 | n16323 ;
  assign n29290 = n8049 | n29289 ;
  assign n29291 = n10815 ^ n3761 ^ 1'b0 ;
  assign n29292 = ~n570 & n9902 ;
  assign n29293 = n570 & n29292 ;
  assign n29294 = n2982 & ~n29293 ;
  assign n29295 = ~n2982 & n29294 ;
  assign n29296 = n8265 & ~n29295 ;
  assign n29297 = ( n8061 & n20888 ) | ( n8061 & ~n29296 ) | ( n20888 & ~n29296 ) ;
  assign n29298 = n22593 | n29297 ;
  assign n29300 = ( x40 & ~n10349 ) | ( x40 & n16043 ) | ( ~n10349 & n16043 ) ;
  assign n29299 = n11270 & ~n14207 ;
  assign n29301 = n29300 ^ n29299 ^ 1'b0 ;
  assign n29302 = n9217 ^ n5889 ^ 1'b0 ;
  assign n29303 = ( n2571 & n18354 ) | ( n2571 & ~n27135 ) | ( n18354 & ~n27135 ) ;
  assign n29304 = ~n742 & n6583 ;
  assign n29305 = n1946 & n29304 ;
  assign n29306 = x74 & n29305 ;
  assign n29307 = n29306 ^ n23534 ^ n19986 ;
  assign n29308 = n25027 ^ n9266 ^ n5924 ;
  assign n29312 = n12711 & n12883 ;
  assign n29313 = n20875 & n29312 ;
  assign n29309 = n1507 & n23722 ;
  assign n29310 = n4419 & n29309 ;
  assign n29311 = n29310 ^ n10949 ^ n2296 ;
  assign n29314 = n29313 ^ n29311 ^ n2846 ;
  assign n29315 = n21403 & n25638 ;
  assign n29316 = ( ~n1886 & n4766 ) | ( ~n1886 & n13528 ) | ( n4766 & n13528 ) ;
  assign n29317 = x29 & ~n22206 ;
  assign n29318 = ~n29316 & n29317 ;
  assign n29319 = n5182 | n29318 ;
  assign n29320 = n29319 ^ n19387 ^ 1'b0 ;
  assign n29321 = n10701 | n24104 ;
  assign n29322 = n28565 ^ n23647 ^ n10787 ;
  assign n29323 = n29322 ^ n28930 ^ 1'b0 ;
  assign n29324 = n7390 & ~n29323 ;
  assign n29325 = ( n2277 & n3271 ) | ( n2277 & n5036 ) | ( n3271 & n5036 ) ;
  assign n29326 = n29325 ^ n19918 ^ 1'b0 ;
  assign n29328 = n8821 & n25664 ;
  assign n29327 = n4474 | n14151 ;
  assign n29329 = n29328 ^ n29327 ^ 1'b0 ;
  assign n29330 = ~n24910 & n27841 ;
  assign n29331 = ~n27649 & n29330 ;
  assign n29332 = n23330 ^ n14652 ^ 1'b0 ;
  assign n29333 = ( n3065 & ~n3555 ) | ( n3065 & n29332 ) | ( ~n3555 & n29332 ) ;
  assign n29334 = n22300 & n28767 ;
  assign n29335 = n26588 ^ n5461 ^ 1'b0 ;
  assign n29336 = n18205 ^ n2670 ^ 1'b0 ;
  assign n29337 = n29336 ^ n7686 ^ n432 ;
  assign n29338 = n16307 ^ n15078 ^ n3710 ;
  assign n29339 = n28975 ^ n6290 ^ 1'b0 ;
  assign n29340 = n9508 | n29339 ;
  assign n29341 = n24037 ^ n2404 ^ 1'b0 ;
  assign n29342 = ~n4338 & n13738 ;
  assign n29343 = ~n1437 & n29342 ;
  assign n29344 = n10871 ^ n5863 ^ n2421 ;
  assign n29345 = n25841 | n29344 ;
  assign n29346 = n29345 ^ n12503 ^ 1'b0 ;
  assign n29347 = ~n13600 & n24858 ;
  assign n29348 = ~n3073 & n5635 ;
  assign n29349 = n29348 ^ n6594 ^ 1'b0 ;
  assign n29350 = n20174 & n29349 ;
  assign n29351 = n15351 & n29350 ;
  assign n29352 = n7600 | n7826 ;
  assign n29353 = n29352 ^ n13472 ^ 1'b0 ;
  assign n29354 = ( n16035 & ~n23966 ) | ( n16035 & n29353 ) | ( ~n23966 & n29353 ) ;
  assign n29355 = n5174 & ~n21881 ;
  assign n29356 = n29355 ^ n27929 ^ n23209 ;
  assign n29357 = ( ~n6189 & n29354 ) | ( ~n6189 & n29356 ) | ( n29354 & n29356 ) ;
  assign n29358 = n7138 & n9174 ;
  assign n29359 = n29358 ^ n28550 ^ n16330 ;
  assign n29363 = n28495 ^ n3373 ^ n2215 ;
  assign n29360 = ( n1514 & ~n3293 ) | ( n1514 & n7248 ) | ( ~n3293 & n7248 ) ;
  assign n29361 = n18281 ^ n2956 ^ 1'b0 ;
  assign n29362 = ~n29360 & n29361 ;
  assign n29364 = n29363 ^ n29362 ^ n1056 ;
  assign n29365 = n15910 | n24680 ;
  assign n29366 = n304 & ~n6249 ;
  assign n29367 = n29366 ^ n5776 ^ 1'b0 ;
  assign n29368 = n29367 ^ n28647 ^ n2200 ;
  assign n29369 = n18498 & ~n29368 ;
  assign n29370 = ~n13873 & n29369 ;
  assign n29371 = n20962 ^ n9324 ^ 1'b0 ;
  assign n29372 = ~n27578 & n29371 ;
  assign n29373 = n942 | n14261 ;
  assign n29374 = n3010 & ~n21853 ;
  assign n29375 = n9967 ^ n921 ^ 1'b0 ;
  assign n29376 = ~n29374 & n29375 ;
  assign n29377 = n16045 ^ n11208 ^ 1'b0 ;
  assign n29378 = ~n1863 & n29377 ;
  assign n29379 = ( n1611 & n1699 ) | ( n1611 & ~n14019 ) | ( n1699 & ~n14019 ) ;
  assign n29380 = n29379 ^ n23840 ^ n9233 ;
  assign n29381 = n5924 & ~n9265 ;
  assign n29382 = n28176 ^ n27834 ^ 1'b0 ;
  assign n29383 = n2805 | n27427 ;
  assign n29384 = n28659 | n29383 ;
  assign n29385 = ( n12484 & n14868 ) | ( n12484 & ~n16133 ) | ( n14868 & ~n16133 ) ;
  assign n29386 = n29385 ^ n14659 ^ 1'b0 ;
  assign n29387 = ~n664 & n21424 ;
  assign n29388 = ~n29386 & n29387 ;
  assign n29389 = n29388 ^ n25260 ^ 1'b0 ;
  assign n29390 = n22009 | n29389 ;
  assign n29391 = n6920 & ~n19720 ;
  assign n29392 = n29391 ^ n13945 ^ 1'b0 ;
  assign n29393 = n3587 & ~n10456 ;
  assign n29394 = ( n15258 & n20613 ) | ( n15258 & n29393 ) | ( n20613 & n29393 ) ;
  assign n29395 = n20575 ^ n3439 ^ 1'b0 ;
  assign n29396 = ( n4823 & n15209 ) | ( n4823 & ~n21595 ) | ( n15209 & ~n21595 ) ;
  assign n29397 = n19598 & ~n22679 ;
  assign n29398 = n29397 ^ n6361 ^ 1'b0 ;
  assign n29399 = n3677 ^ n366 ^ 1'b0 ;
  assign n29400 = n1580 | n2114 ;
  assign n29401 = n29400 ^ n17421 ^ n6730 ;
  assign n29402 = n29399 | n29401 ;
  assign n29403 = n26543 ^ n2426 ^ 1'b0 ;
  assign n29404 = n12269 ^ n4175 ^ 1'b0 ;
  assign n29405 = ~n13590 & n29404 ;
  assign n29406 = n20317 & n21640 ;
  assign n29407 = ~n19743 & n29406 ;
  assign n29408 = n5610 ^ n3358 ^ 1'b0 ;
  assign n29409 = ( n4510 & ~n10551 ) | ( n4510 & n12869 ) | ( ~n10551 & n12869 ) ;
  assign n29410 = n14144 ^ n10092 ^ n8039 ;
  assign n29411 = n4595 ^ n3424 ^ 1'b0 ;
  assign n29412 = n24789 ^ n23157 ^ n16737 ;
  assign n29413 = n29411 & n29412 ;
  assign n29414 = n13884 & n15685 ;
  assign n29415 = n11653 & n29414 ;
  assign n29416 = n19016 ^ n6418 ^ 1'b0 ;
  assign n29417 = ~n4593 & n17073 ;
  assign n29418 = ~n754 & n29417 ;
  assign n29419 = n4943 & ~n17912 ;
  assign n29426 = n4704 & n15047 ;
  assign n29420 = n10508 ^ n1145 ^ 1'b0 ;
  assign n29421 = n11258 & n29420 ;
  assign n29422 = n2853 | n22009 ;
  assign n29423 = n2006 ^ n1504 ^ 1'b0 ;
  assign n29424 = n29423 ^ n17446 ^ n4521 ;
  assign n29425 = ( n29421 & ~n29422 ) | ( n29421 & n29424 ) | ( ~n29422 & n29424 ) ;
  assign n29427 = n29426 ^ n29425 ^ 1'b0 ;
  assign n29428 = ( n2442 & ~n18738 ) | ( n2442 & n19744 ) | ( ~n18738 & n19744 ) ;
  assign n29429 = ( n3753 & n12260 ) | ( n3753 & n15209 ) | ( n12260 & n15209 ) ;
  assign n29430 = n9913 | n12479 ;
  assign n29431 = ~n2119 & n29430 ;
  assign n29432 = n9678 & n17447 ;
  assign n29433 = n29432 ^ n8393 ^ 1'b0 ;
  assign n29434 = ~n1976 & n10735 ;
  assign n29435 = n29434 ^ n5010 ^ 1'b0 ;
  assign n29436 = n25194 | n29435 ;
  assign n29437 = n5609 & ~n8390 ;
  assign n29438 = n29437 ^ n17480 ^ 1'b0 ;
  assign n29439 = n29438 ^ n6991 ^ 1'b0 ;
  assign n29440 = n333 & ~n29439 ;
  assign n29441 = n21893 & n29440 ;
  assign n29442 = n29441 ^ n25804 ^ n12330 ;
  assign n29445 = n390 & ~n4157 ;
  assign n29443 = n16842 ^ n3337 ^ n2735 ;
  assign n29444 = n14023 | n29443 ;
  assign n29446 = n29445 ^ n29444 ^ n26473 ;
  assign n29447 = n14657 ^ n9657 ^ n7636 ;
  assign n29448 = n12752 & n23417 ;
  assign n29449 = ~n465 & n21844 ;
  assign n29450 = n19764 & n29449 ;
  assign n29451 = n29450 ^ n10392 ^ 1'b0 ;
  assign n29452 = n19835 ^ n4341 ^ 1'b0 ;
  assign n29453 = n213 | n14586 ;
  assign n29455 = n10042 ^ n3055 ^ n956 ;
  assign n29454 = n11600 | n18758 ;
  assign n29456 = n29455 ^ n29454 ^ 1'b0 ;
  assign n29457 = n28443 ^ n2509 ^ 1'b0 ;
  assign n29458 = n241 | n29457 ;
  assign n29461 = ( n3607 & n3796 ) | ( n3607 & ~n10803 ) | ( n3796 & ~n10803 ) ;
  assign n29459 = n8859 & n13651 ;
  assign n29460 = n29459 ^ n14831 ^ 1'b0 ;
  assign n29462 = n29461 ^ n29460 ^ 1'b0 ;
  assign n29463 = n6583 | n29462 ;
  assign n29464 = n22163 ^ n19779 ^ n5225 ;
  assign n29465 = ( n5894 & ~n24154 ) | ( n5894 & n27287 ) | ( ~n24154 & n27287 ) ;
  assign n29466 = ( ~n304 & n15873 ) | ( ~n304 & n16251 ) | ( n15873 & n16251 ) ;
  assign n29467 = n2340 & ~n25225 ;
  assign n29468 = n8957 & n13461 ;
  assign n29469 = n29468 ^ n10214 ^ 1'b0 ;
  assign n29470 = n5410 & n15376 ;
  assign n29471 = ~n13893 & n29470 ;
  assign n29472 = n29471 ^ n17042 ^ 1'b0 ;
  assign n29473 = n5221 ^ n2822 ^ 1'b0 ;
  assign n29474 = ~n23144 & n29473 ;
  assign n29475 = ~n8310 & n14284 ;
  assign n29476 = n1880 & ~n22414 ;
  assign n29477 = n29476 ^ n10040 ^ 1'b0 ;
  assign n29478 = n2014 | n21249 ;
  assign n29479 = ~n21896 & n29478 ;
  assign n29480 = n29479 ^ n17831 ^ 1'b0 ;
  assign n29486 = n4964 | n5826 ;
  assign n29481 = n18631 ^ n1340 ^ 1'b0 ;
  assign n29482 = n8468 | n29481 ;
  assign n29483 = n29482 ^ n5661 ^ n390 ;
  assign n29484 = n28718 ^ n8562 ^ 1'b0 ;
  assign n29485 = n29483 | n29484 ;
  assign n29487 = n29486 ^ n29485 ^ n1090 ;
  assign n29488 = n29487 ^ n24507 ^ n7251 ;
  assign n29489 = n14629 ^ n10884 ^ 1'b0 ;
  assign n29491 = n2180 ^ n1253 ^ 1'b0 ;
  assign n29492 = n29491 ^ n16091 ^ 1'b0 ;
  assign n29493 = ~n17249 & n29492 ;
  assign n29490 = ~n1717 & n19430 ;
  assign n29494 = n29493 ^ n29490 ^ 1'b0 ;
  assign n29495 = n8471 | n8854 ;
  assign n29496 = n29495 ^ n27812 ^ 1'b0 ;
  assign n29497 = n23783 ^ n9152 ^ 1'b0 ;
  assign n29498 = n29496 & ~n29497 ;
  assign n29500 = ~n933 & n5542 ;
  assign n29501 = n458 & n29500 ;
  assign n29502 = ( ~n4413 & n14083 ) | ( ~n4413 & n29501 ) | ( n14083 & n29501 ) ;
  assign n29499 = n1501 & n15112 ;
  assign n29503 = n29502 ^ n29499 ^ 1'b0 ;
  assign n29504 = n13013 ^ n8218 ^ 1'b0 ;
  assign n29505 = ~n8643 & n29504 ;
  assign n29506 = n29505 ^ n27161 ^ n20470 ;
  assign n29507 = n24498 & ~n29506 ;
  assign n29508 = n29507 ^ n3441 ^ 1'b0 ;
  assign n29509 = ( ~n272 & n2929 ) | ( ~n272 & n3887 ) | ( n2929 & n3887 ) ;
  assign n29510 = n483 & n29509 ;
  assign n29511 = n4827 | n9513 ;
  assign n29512 = n29511 ^ n8307 ^ 1'b0 ;
  assign n29513 = n7563 | n19489 ;
  assign n29514 = n29512 | n29513 ;
  assign n29515 = n1896 & n29514 ;
  assign n29516 = ( n22330 & n22552 ) | ( n22330 & ~n28878 ) | ( n22552 & ~n28878 ) ;
  assign n29517 = ( n9108 & n17389 ) | ( n9108 & n29516 ) | ( n17389 & n29516 ) ;
  assign n29518 = ( n2187 & ~n11533 ) | ( n2187 & n19016 ) | ( ~n11533 & n19016 ) ;
  assign n29519 = n29518 ^ n17604 ^ 1'b0 ;
  assign n29520 = ( n3448 & n9368 ) | ( n3448 & n29519 ) | ( n9368 & n29519 ) ;
  assign n29522 = ( n2160 & ~n3557 ) | ( n2160 & n15294 ) | ( ~n3557 & n15294 ) ;
  assign n29523 = n29522 ^ n27853 ^ n13026 ;
  assign n29521 = n2498 | n26023 ;
  assign n29524 = n29523 ^ n29521 ^ n970 ;
  assign n29525 = n15673 ^ n10076 ^ 1'b0 ;
  assign n29526 = n6675 & n29525 ;
  assign n29527 = n20130 ^ n4944 ^ 1'b0 ;
  assign n29528 = n16662 & n29527 ;
  assign n29529 = n18359 & n19685 ;
  assign n29530 = n4078 & n14084 ;
  assign n29531 = n29530 ^ n28132 ^ 1'b0 ;
  assign n29532 = n10242 & n20641 ;
  assign n29533 = n29532 ^ n15729 ^ n8365 ;
  assign n29534 = n29533 ^ n17808 ^ 1'b0 ;
  assign n29535 = n7211 | n29534 ;
  assign n29536 = ( n9034 & n14879 ) | ( n9034 & ~n29358 ) | ( n14879 & ~n29358 ) ;
  assign n29537 = n28777 | n29536 ;
  assign n29538 = n21170 & ~n28656 ;
  assign n29539 = n29538 ^ n23157 ^ 1'b0 ;
  assign n29540 = ~n26169 & n29539 ;
  assign n29541 = n25128 ^ n15627 ^ 1'b0 ;
  assign n29542 = n22374 ^ n1059 ^ 1'b0 ;
  assign n29543 = n2638 & n29542 ;
  assign n29544 = n6050 | n10903 ;
  assign n29545 = n29544 ^ n28124 ^ 1'b0 ;
  assign n29546 = n4741 | n12152 ;
  assign n29547 = n3625 & ~n29546 ;
  assign n29548 = n6297 & ~n18829 ;
  assign n29549 = n29548 ^ n3181 ^ 1'b0 ;
  assign n29550 = ( n13492 & ~n25702 ) | ( n13492 & n29549 ) | ( ~n25702 & n29549 ) ;
  assign n29551 = ( n208 & n5431 ) | ( n208 & ~n14012 ) | ( n5431 & ~n14012 ) ;
  assign n29552 = n12658 & n29551 ;
  assign n29553 = n10276 & ~n14509 ;
  assign n29554 = n7098 & n29553 ;
  assign n29555 = ( n2071 & n20441 ) | ( n2071 & n29554 ) | ( n20441 & n29554 ) ;
  assign n29556 = n8243 | n13021 ;
  assign n29557 = n29556 ^ n11189 ^ n776 ;
  assign n29558 = n17707 & ~n29557 ;
  assign n29559 = n17182 ^ n12109 ^ n7197 ;
  assign n29560 = ( ~n19585 & n29558 ) | ( ~n19585 & n29559 ) | ( n29558 & n29559 ) ;
  assign n29561 = n14170 & n19507 ;
  assign n29562 = n26930 ^ n16136 ^ 1'b0 ;
  assign n29563 = ~n6122 & n29562 ;
  assign n29564 = n7628 & ~n29563 ;
  assign n29565 = n29564 ^ n25301 ^ 1'b0 ;
  assign n29566 = ~n19488 & n29565 ;
  assign n29567 = ~n8916 & n9979 ;
  assign n29568 = n7622 & n11708 ;
  assign n29569 = n29568 ^ n17387 ^ 1'b0 ;
  assign n29570 = n19821 ^ n11038 ^ n3411 ;
  assign n29571 = n15342 ^ n3110 ^ 1'b0 ;
  assign n29572 = n269 | n12950 ;
  assign n29573 = ( ~n22217 & n29571 ) | ( ~n22217 & n29572 ) | ( n29571 & n29572 ) ;
  assign n29574 = n7832 | n24863 ;
  assign n29575 = n29574 ^ n6057 ^ 1'b0 ;
  assign n29576 = n29575 ^ n18392 ^ n13594 ;
  assign n29577 = ( n174 & n2684 ) | ( n174 & n2984 ) | ( n2684 & n2984 ) ;
  assign n29578 = n29577 ^ n15494 ^ n8984 ;
  assign n29579 = n12035 & n16303 ;
  assign n29580 = n9442 ^ n6911 ^ 1'b0 ;
  assign n29581 = ( n586 & n2965 ) | ( n586 & ~n14353 ) | ( n2965 & ~n14353 ) ;
  assign n29582 = n29581 ^ n27171 ^ 1'b0 ;
  assign n29583 = n23997 | n26440 ;
  assign n29584 = n17287 & ~n29583 ;
  assign n29585 = n4692 & n29426 ;
  assign n29586 = n29585 ^ n28685 ^ 1'b0 ;
  assign n29587 = ( n2706 & n3658 ) | ( n2706 & n15219 ) | ( n3658 & n15219 ) ;
  assign n29588 = n15526 & ~n29587 ;
  assign n29589 = ( n6424 & ~n8225 ) | ( n6424 & n25385 ) | ( ~n8225 & n25385 ) ;
  assign n29590 = n5915 | n8828 ;
  assign n29591 = ( n872 & ~n6609 ) | ( n872 & n7349 ) | ( ~n6609 & n7349 ) ;
  assign n29592 = n29591 ^ n24524 ^ n22187 ;
  assign n29593 = ~n8245 & n29592 ;
  assign n29594 = n29593 ^ n18282 ^ 1'b0 ;
  assign n29595 = n7682 ^ n7572 ^ 1'b0 ;
  assign n29596 = n7874 & ~n29595 ;
  assign n29597 = n1679 & n29596 ;
  assign n29598 = n29597 ^ n2960 ^ 1'b0 ;
  assign n29599 = n4059 ^ x89 ^ 1'b0 ;
  assign n29600 = ~n9217 & n29599 ;
  assign n29601 = n29600 ^ n4367 ^ 1'b0 ;
  assign n29602 = n28422 ^ n12465 ^ n7030 ;
  assign n29603 = ( n5307 & n8600 ) | ( n5307 & n21611 ) | ( n8600 & n21611 ) ;
  assign n29604 = ( ~n1319 & n12938 ) | ( ~n1319 & n25146 ) | ( n12938 & n25146 ) ;
  assign n29605 = ( n5713 & n12889 ) | ( n5713 & ~n19777 ) | ( n12889 & ~n19777 ) ;
  assign n29606 = n16168 ^ n13560 ^ n3328 ;
  assign n29607 = ( n4132 & n12525 ) | ( n4132 & ~n29606 ) | ( n12525 & ~n29606 ) ;
  assign n29608 = n12974 ^ n7643 ^ 1'b0 ;
  assign n29609 = n26441 | n28340 ;
  assign n29610 = n29608 & ~n29609 ;
  assign n29611 = n15151 ^ n11993 ^ 1'b0 ;
  assign n29612 = n8629 | n29611 ;
  assign n29613 = n5267 | n6145 ;
  assign n29614 = n29612 & ~n29613 ;
  assign n29615 = n11636 ^ n7897 ^ 1'b0 ;
  assign n29616 = n7528 ^ n2356 ^ 1'b0 ;
  assign n29617 = n29615 & n29616 ;
  assign n29618 = n8999 ^ n8108 ^ n3086 ;
  assign n29621 = ( ~n826 & n14886 ) | ( ~n826 & n17324 ) | ( n14886 & n17324 ) ;
  assign n29619 = n8557 ^ n6919 ^ 1'b0 ;
  assign n29620 = n18929 | n29619 ;
  assign n29622 = n29621 ^ n29620 ^ n22380 ;
  assign n29624 = n15799 ^ n7733 ^ 1'b0 ;
  assign n29625 = n10670 | n29624 ;
  assign n29623 = n16838 ^ n727 ^ 1'b0 ;
  assign n29626 = n29625 ^ n29623 ^ n19993 ;
  assign n29627 = n1592 | n12327 ;
  assign n29628 = n29627 ^ n16377 ^ n12143 ;
  assign n29629 = ~n18616 & n28178 ;
  assign n29630 = ~n19682 & n29629 ;
  assign n29631 = n3204 ^ n1611 ^ 1'b0 ;
  assign n29632 = n28719 & n29631 ;
  assign n29633 = ~n12667 & n29632 ;
  assign n29634 = n6769 | n12812 ;
  assign n29635 = n5362 & ~n29634 ;
  assign n29636 = n18789 | n29635 ;
  assign n29637 = x77 & n11834 ;
  assign n29638 = ~n9195 & n29637 ;
  assign n29639 = ~n565 & n4346 ;
  assign n29640 = n29639 ^ n27853 ^ 1'b0 ;
  assign n29641 = n29640 ^ n6334 ^ 1'b0 ;
  assign n29642 = ~n23786 & n29641 ;
  assign n29643 = n26895 ^ n10806 ^ 1'b0 ;
  assign n29644 = n16811 & n17100 ;
  assign n29645 = ( n10518 & n21445 ) | ( n10518 & ~n27576 ) | ( n21445 & ~n27576 ) ;
  assign n29646 = n885 | n29645 ;
  assign n29647 = n19531 ^ n13190 ^ n8105 ;
  assign n29648 = n4718 & n19322 ;
  assign n29649 = ( n8450 & ~n29647 ) | ( n8450 & n29648 ) | ( ~n29647 & n29648 ) ;
  assign n29650 = ( n1699 & ~n4194 ) | ( n1699 & n4745 ) | ( ~n4194 & n4745 ) ;
  assign n29651 = n8408 ^ n8398 ^ 1'b0 ;
  assign n29652 = ~n29650 & n29651 ;
  assign n29653 = n29652 ^ n18829 ^ 1'b0 ;
  assign n29654 = n13175 ^ n3698 ^ 1'b0 ;
  assign n29655 = n17046 & n29654 ;
  assign n29656 = ( n12716 & n20275 ) | ( n12716 & ~n23905 ) | ( n20275 & ~n23905 ) ;
  assign n29657 = n29656 ^ n7168 ^ 1'b0 ;
  assign n29658 = ~n4429 & n29657 ;
  assign n29659 = n17989 ^ n11928 ^ 1'b0 ;
  assign n29660 = ~n2317 & n29659 ;
  assign n29661 = n24037 ^ n1234 ^ 1'b0 ;
  assign n29662 = n16463 ^ n8699 ^ 1'b0 ;
  assign n29663 = n10657 | n29662 ;
  assign n29664 = n24194 ^ n2671 ^ 1'b0 ;
  assign n29665 = ( n5184 & n29663 ) | ( n5184 & n29664 ) | ( n29663 & n29664 ) ;
  assign n29667 = n12483 ^ n7422 ^ 1'b0 ;
  assign n29668 = n13219 | n29667 ;
  assign n29666 = n7574 ^ n809 ^ 1'b0 ;
  assign n29669 = n29668 ^ n29666 ^ n27360 ;
  assign n29670 = ( n5759 & ~n8916 ) | ( n5759 & n15482 ) | ( ~n8916 & n15482 ) ;
  assign n29671 = ( n4830 & n21858 ) | ( n4830 & n29670 ) | ( n21858 & n29670 ) ;
  assign n29672 = ~n7280 & n16343 ;
  assign n29673 = n29672 ^ n767 ^ 1'b0 ;
  assign n29674 = n4121 & n13999 ;
  assign n29675 = n29674 ^ n4660 ^ 1'b0 ;
  assign n29676 = ~n1428 & n16188 ;
  assign n29677 = n29676 ^ n1146 ^ 1'b0 ;
  assign n29678 = n29675 | n29677 ;
  assign n29679 = n22647 & ~n25762 ;
  assign n29680 = ( n14057 & n14949 ) | ( n14057 & ~n16757 ) | ( n14949 & ~n16757 ) ;
  assign n29681 = n29680 ^ n9993 ^ 1'b0 ;
  assign n29682 = ( n5086 & ~n21062 ) | ( n5086 & n29681 ) | ( ~n21062 & n29681 ) ;
  assign n29683 = ~n10790 & n20238 ;
  assign n29684 = n24887 | n28234 ;
  assign n29685 = n4786 & n23882 ;
  assign n29686 = ~n7737 & n29685 ;
  assign n29687 = n29686 ^ n7650 ^ 1'b0 ;
  assign n29689 = n5655 & ~n10570 ;
  assign n29688 = n6201 & ~n24391 ;
  assign n29690 = n29689 ^ n29688 ^ 1'b0 ;
  assign n29691 = ~n19524 & n29690 ;
  assign n29692 = n20406 ^ n15518 ^ 1'b0 ;
  assign n29693 = ( n5272 & n5859 ) | ( n5272 & ~n13942 ) | ( n5859 & ~n13942 ) ;
  assign n29694 = ~n4033 & n29693 ;
  assign n29695 = n15526 & n29694 ;
  assign n29696 = n28795 & n29695 ;
  assign n29697 = n18902 ^ n11885 ^ n10419 ;
  assign n29698 = n26464 & ~n29697 ;
  assign n29699 = n29698 ^ n2401 ^ 1'b0 ;
  assign n29700 = n1909 & n29699 ;
  assign n29701 = n16482 ^ n7232 ^ n1018 ;
  assign n29702 = n21794 ^ n11485 ^ 1'b0 ;
  assign n29703 = n12112 ^ n6999 ^ n5178 ;
  assign n29704 = n7112 & n18729 ;
  assign n29705 = n29704 ^ n26380 ^ n7160 ;
  assign n29706 = n205 & ~n5543 ;
  assign n29707 = n29706 ^ n28601 ^ 1'b0 ;
  assign n29708 = ( ~n6324 & n15632 ) | ( ~n6324 & n29707 ) | ( n15632 & n29707 ) ;
  assign n29709 = n22638 ^ n12432 ^ 1'b0 ;
  assign n29710 = n188 & n26653 ;
  assign n29711 = n25676 & n29344 ;
  assign n29712 = n17510 ^ n10716 ^ n8512 ;
  assign n29713 = n14304 ^ n11027 ^ 1'b0 ;
  assign n29714 = n10272 | n29713 ;
  assign n29715 = n5470 | n7087 ;
  assign n29716 = ( n7152 & n7716 ) | ( n7152 & ~n27646 ) | ( n7716 & ~n27646 ) ;
  assign n29717 = ( n8043 & n15962 ) | ( n8043 & n21532 ) | ( n15962 & n21532 ) ;
  assign n29718 = n29717 ^ n16597 ^ 1'b0 ;
  assign n29719 = ~n24776 & n29718 ;
  assign n29720 = ~n12425 & n29719 ;
  assign n29721 = n10213 | n29720 ;
  assign n29722 = n29721 ^ x18 ^ 1'b0 ;
  assign n29723 = n3707 ^ n2934 ^ 1'b0 ;
  assign n29724 = n11189 & ~n29723 ;
  assign n29725 = n29724 ^ n14966 ^ n5510 ;
  assign n29726 = n1990 | n29725 ;
  assign n29727 = n29726 ^ n3883 ^ 1'b0 ;
  assign n29728 = n15097 & n20792 ;
  assign n29729 = n29728 ^ n27783 ^ 1'b0 ;
  assign n29730 = n20078 | n22939 ;
  assign n29731 = ~n7095 & n15376 ;
  assign n29732 = n29731 ^ n6358 ^ 1'b0 ;
  assign n29733 = ~n12323 & n29732 ;
  assign n29734 = ( n3166 & n22825 ) | ( n3166 & n29733 ) | ( n22825 & n29733 ) ;
  assign n29736 = ( n4701 & n15502 ) | ( n4701 & n23119 ) | ( n15502 & n23119 ) ;
  assign n29735 = n12346 & ~n12866 ;
  assign n29737 = n29736 ^ n29735 ^ 1'b0 ;
  assign n29738 = n29737 ^ n25480 ^ n12605 ;
  assign n29739 = n9701 | n21173 ;
  assign n29740 = n17205 ^ n3018 ^ 1'b0 ;
  assign n29741 = n3030 | n29740 ;
  assign n29742 = n29741 ^ n16061 ^ n2360 ;
  assign n29743 = n17430 & ~n26611 ;
  assign n29744 = n4185 & ~n13202 ;
  assign n29745 = n29744 ^ n9193 ^ 1'b0 ;
  assign n29746 = n2937 & n7002 ;
  assign n29747 = ~n14285 & n29746 ;
  assign n29748 = n13886 & ~n21913 ;
  assign n29749 = n29747 & n29748 ;
  assign n29750 = ~n7913 & n11257 ;
  assign n29751 = n1738 | n10456 ;
  assign n29752 = n4705 & ~n29751 ;
  assign n29753 = ( ~n938 & n18950 ) | ( ~n938 & n29612 ) | ( n18950 & n29612 ) ;
  assign n29755 = n13673 ^ n5990 ^ n3441 ;
  assign n29754 = n6393 & n11319 ;
  assign n29756 = n29755 ^ n29754 ^ n18718 ;
  assign n29757 = n15331 & n23238 ;
  assign n29758 = n9699 & ~n25261 ;
  assign n29759 = ( n6319 & n7743 ) | ( n6319 & n9442 ) | ( n7743 & n9442 ) ;
  assign n29760 = ( n8836 & n29758 ) | ( n8836 & n29759 ) | ( n29758 & n29759 ) ;
  assign n29761 = n11312 | n27244 ;
  assign n29762 = ( n7404 & n16208 ) | ( n7404 & ~n22542 ) | ( n16208 & ~n22542 ) ;
  assign n29763 = n29762 ^ n20051 ^ 1'b0 ;
  assign n29764 = n10977 ^ n7499 ^ n6847 ;
  assign n29765 = n29764 ^ n29461 ^ n874 ;
  assign n29766 = ( n29761 & n29763 ) | ( n29761 & n29765 ) | ( n29763 & n29765 ) ;
  assign n29767 = n20186 ^ n3670 ^ 1'b0 ;
  assign n29768 = n19524 ^ n6226 ^ n887 ;
  assign n29769 = n29768 ^ n19547 ^ 1'b0 ;
  assign n29770 = ~n29767 & n29769 ;
  assign n29771 = n10569 & n15110 ;
  assign n29772 = n29771 ^ n7262 ^ n5603 ;
  assign n29773 = n9567 ^ n5355 ^ 1'b0 ;
  assign n29774 = n29772 | n29773 ;
  assign n29775 = ( ~n3440 & n7094 ) | ( ~n3440 & n10770 ) | ( n7094 & n10770 ) ;
  assign n29776 = n19281 ^ n6142 ^ 1'b0 ;
  assign n29777 = ~n29775 & n29776 ;
  assign n29778 = ~n8574 & n29623 ;
  assign n29779 = ~n29777 & n29778 ;
  assign n29780 = ( n2929 & n18296 ) | ( n2929 & n21893 ) | ( n18296 & n21893 ) ;
  assign n29781 = n29780 ^ n3573 ^ 1'b0 ;
  assign y0 = x1 ;
  assign y1 = x3 ;
  assign y2 = x20 ;
  assign y3 = x29 ;
  assign y4 = x34 ;
  assign y5 = x40 ;
  assign y6 = x44 ;
  assign y7 = x45 ;
  assign y8 = x68 ;
  assign y9 = x75 ;
  assign y10 = x78 ;
  assign y11 = x86 ;
  assign y12 = x96 ;
  assign y13 = x97 ;
  assign y14 = x107 ;
  assign y15 = x120 ;
  assign y16 = n129 ;
  assign y17 = n131 ;
  assign y18 = ~n134 ;
  assign y19 = n136 ;
  assign y20 = n137 ;
  assign y21 = ~1'b0 ;
  assign y22 = ~n141 ;
  assign y23 = n143 ;
  assign y24 = n146 ;
  assign y25 = ~n156 ;
  assign y26 = ~n160 ;
  assign y27 = ~n162 ;
  assign y28 = ~n164 ;
  assign y29 = n167 ;
  assign y30 = n168 ;
  assign y31 = n170 ;
  assign y32 = ~1'b0 ;
  assign y33 = ~n171 ;
  assign y34 = n173 ;
  assign y35 = n174 ;
  assign y36 = n178 ;
  assign y37 = ~1'b0 ;
  assign y38 = ~1'b0 ;
  assign y39 = n180 ;
  assign y40 = ~n184 ;
  assign y41 = n187 ;
  assign y42 = ~n192 ;
  assign y43 = ~n194 ;
  assign y44 = ~n196 ;
  assign y45 = ~1'b0 ;
  assign y46 = n199 ;
  assign y47 = n202 ;
  assign y48 = n205 ;
  assign y49 = n221 ;
  assign y50 = n227 ;
  assign y51 = ~n228 ;
  assign y52 = ~1'b0 ;
  assign y53 = ~n234 ;
  assign y54 = n242 ;
  assign y55 = n246 ;
  assign y56 = ~n247 ;
  assign y57 = ~1'b0 ;
  assign y58 = ~n250 ;
  assign y59 = ~n253 ;
  assign y60 = ~n259 ;
  assign y61 = ~n260 ;
  assign y62 = n266 ;
  assign y63 = n267 ;
  assign y64 = ~1'b0 ;
  assign y65 = n270 ;
  assign y66 = ~1'b0 ;
  assign y67 = ~n272 ;
  assign y68 = ~1'b0 ;
  assign y69 = n149 ;
  assign y70 = ~1'b0 ;
  assign y71 = ~n277 ;
  assign y72 = n281 ;
  assign y73 = ~1'b0 ;
  assign y74 = ~1'b0 ;
  assign y75 = n285 ;
  assign y76 = ~n293 ;
  assign y77 = ~1'b0 ;
  assign y78 = ~1'b0 ;
  assign y79 = ~n295 ;
  assign y80 = n305 ;
  assign y81 = ~n308 ;
  assign y82 = n310 ;
  assign y83 = ~n322 ;
  assign y84 = ~1'b0 ;
  assign y85 = ~1'b0 ;
  assign y86 = ~1'b0 ;
  assign y87 = ~n328 ;
  assign y88 = ~n338 ;
  assign y89 = ~n344 ;
  assign y90 = n348 ;
  assign y91 = ~n349 ;
  assign y92 = ~n352 ;
  assign y93 = n366 ;
  assign y94 = n368 ;
  assign y95 = n370 ;
  assign y96 = ~n379 ;
  assign y97 = ~n381 ;
  assign y98 = n171 ;
  assign y99 = ~1'b0 ;
  assign y100 = ~n383 ;
  assign y101 = n386 ;
  assign y102 = n394 ;
  assign y103 = n399 ;
  assign y104 = ~n403 ;
  assign y105 = n406 ;
  assign y106 = n420 ;
  assign y107 = n421 ;
  assign y108 = n445 ;
  assign y109 = n448 ;
  assign y110 = n449 ;
  assign y111 = n455 ;
  assign y112 = ~n456 ;
  assign y113 = ~n458 ;
  assign y114 = ~n462 ;
  assign y115 = x93 ;
  assign y116 = n464 ;
  assign y117 = n470 ;
  assign y118 = ~1'b0 ;
  assign y119 = ~n476 ;
  assign y120 = ~n478 ;
  assign y121 = ~n479 ;
  assign y122 = n482 ;
  assign y123 = ~1'b0 ;
  assign y124 = n492 ;
  assign y125 = n500 ;
  assign y126 = ~n502 ;
  assign y127 = n505 ;
  assign y128 = ~n506 ;
  assign y129 = ~1'b0 ;
  assign y130 = n509 ;
  assign y131 = n512 ;
  assign y132 = n520 ;
  assign y133 = ~n526 ;
  assign y134 = ~n528 ;
  assign y135 = ~1'b0 ;
  assign y136 = ~n182 ;
  assign y137 = ~1'b0 ;
  assign y138 = n537 ;
  assign y139 = ~n539 ;
  assign y140 = 1'b0 ;
  assign y141 = ~n543 ;
  assign y142 = n545 ;
  assign y143 = n549 ;
  assign y144 = n551 ;
  assign y145 = ~n556 ;
  assign y146 = ~n559 ;
  assign y147 = ~n566 ;
  assign y148 = ~n569 ;
  assign y149 = ~n570 ;
  assign y150 = ~n584 ;
  assign y151 = n588 ;
  assign y152 = n594 ;
  assign y153 = ~n599 ;
  assign y154 = ~n604 ;
  assign y155 = ~n610 ;
  assign y156 = n617 ;
  assign y157 = n626 ;
  assign y158 = ~n631 ;
  assign y159 = ~1'b0 ;
  assign y160 = n637 ;
  assign y161 = ~n639 ;
  assign y162 = ~n644 ;
  assign y163 = n650 ;
  assign y164 = ~1'b0 ;
  assign y165 = n656 ;
  assign y166 = ~n664 ;
  assign y167 = ~1'b0 ;
  assign y168 = n666 ;
  assign y169 = ~n667 ;
  assign y170 = ~n676 ;
  assign y171 = ~n680 ;
  assign y172 = ~n685 ;
  assign y173 = n691 ;
  assign y174 = n695 ;
  assign y175 = n699 ;
  assign y176 = n701 ;
  assign y177 = n704 ;
  assign y178 = ~n708 ;
  assign y179 = ~1'b0 ;
  assign y180 = ~1'b0 ;
  assign y181 = n713 ;
  assign y182 = ~1'b0 ;
  assign y183 = ~n715 ;
  assign y184 = ~n721 ;
  assign y185 = n722 ;
  assign y186 = 1'b0 ;
  assign y187 = n728 ;
  assign y188 = ~n736 ;
  assign y189 = n737 ;
  assign y190 = n751 ;
  assign y191 = ~1'b0 ;
  assign y192 = n755 ;
  assign y193 = ~n759 ;
  assign y194 = ~n760 ;
  assign y195 = n761 ;
  assign y196 = n771 ;
  assign y197 = ~1'b0 ;
  assign y198 = n773 ;
  assign y199 = n775 ;
  assign y200 = n779 ;
  assign y201 = ~n803 ;
  assign y202 = ~n804 ;
  assign y203 = n807 ;
  assign y204 = ~1'b0 ;
  assign y205 = ~n808 ;
  assign y206 = n809 ;
  assign y207 = ~n812 ;
  assign y208 = ~n401 ;
  assign y209 = n821 ;
  assign y210 = ~1'b0 ;
  assign y211 = ~n826 ;
  assign y212 = n833 ;
  assign y213 = ~n847 ;
  assign y214 = ~n850 ;
  assign y215 = ~1'b0 ;
  assign y216 = ~1'b0 ;
  assign y217 = n856 ;
  assign y218 = ~1'b0 ;
  assign y219 = n872 ;
  assign y220 = ~1'b0 ;
  assign y221 = ~n873 ;
  assign y222 = n875 ;
  assign y223 = n877 ;
  assign y224 = n878 ;
  assign y225 = ~n889 ;
  assign y226 = ~1'b0 ;
  assign y227 = n891 ;
  assign y228 = n894 ;
  assign y229 = ~n895 ;
  assign y230 = n898 ;
  assign y231 = ~n903 ;
  assign y232 = n905 ;
  assign y233 = ~n906 ;
  assign y234 = n912 ;
  assign y235 = ~1'b0 ;
  assign y236 = n915 ;
  assign y237 = ~1'b0 ;
  assign y238 = ~n916 ;
  assign y239 = n917 ;
  assign y240 = n926 ;
  assign y241 = ~n927 ;
  assign y242 = n932 ;
  assign y243 = ~1'b0 ;
  assign y244 = n935 ;
  assign y245 = n937 ;
  assign y246 = ~n940 ;
  assign y247 = ~n942 ;
  assign y248 = ~1'b0 ;
  assign y249 = ~1'b0 ;
  assign y250 = n943 ;
  assign y251 = n947 ;
  assign y252 = n948 ;
  assign y253 = n955 ;
  assign y254 = ~1'b0 ;
  assign y255 = ~n958 ;
  assign y256 = n965 ;
  assign y257 = ~n967 ;
  assign y258 = n973 ;
  assign y259 = n974 ;
  assign y260 = ~1'b0 ;
  assign y261 = ~n977 ;
  assign y262 = n981 ;
  assign y263 = n983 ;
  assign y264 = ~1'b0 ;
  assign y265 = n986 ;
  assign y266 = n987 ;
  assign y267 = n990 ;
  assign y268 = n991 ;
  assign y269 = ~1'b0 ;
  assign y270 = n992 ;
  assign y271 = ~n993 ;
  assign y272 = ~1'b0 ;
  assign y273 = n998 ;
  assign y274 = n999 ;
  assign y275 = ~n1000 ;
  assign y276 = ~1'b0 ;
  assign y277 = ~1'b0 ;
  assign y278 = ~1'b0 ;
  assign y279 = n1002 ;
  assign y280 = ~n1013 ;
  assign y281 = ~n1016 ;
  assign y282 = ~n1018 ;
  assign y283 = x108 ;
  assign y284 = ~n1030 ;
  assign y285 = n1033 ;
  assign y286 = n1035 ;
  assign y287 = n1038 ;
  assign y288 = n1043 ;
  assign y289 = ~n1046 ;
  assign y290 = n1052 ;
  assign y291 = ~n1055 ;
  assign y292 = n1058 ;
  assign y293 = ~n1059 ;
  assign y294 = ~n1063 ;
  assign y295 = n1065 ;
  assign y296 = n1069 ;
  assign y297 = n1072 ;
  assign y298 = ~n1075 ;
  assign y299 = ~1'b0 ;
  assign y300 = ~n1076 ;
  assign y301 = ~n1080 ;
  assign y302 = n1083 ;
  assign y303 = n1084 ;
  assign y304 = ~1'b0 ;
  assign y305 = n1087 ;
  assign y306 = ~n915 ;
  assign y307 = n1094 ;
  assign y308 = n1095 ;
  assign y309 = n1097 ;
  assign y310 = ~n1098 ;
  assign y311 = ~n1113 ;
  assign y312 = ~1'b0 ;
  assign y313 = ~n1114 ;
  assign y314 = n1116 ;
  assign y315 = n1126 ;
  assign y316 = ~1'b0 ;
  assign y317 = ~1'b0 ;
  assign y318 = ~n1128 ;
  assign y319 = ~n1138 ;
  assign y320 = 1'b0 ;
  assign y321 = ~n1145 ;
  assign y322 = ~1'b0 ;
  assign y323 = ~n1146 ;
  assign y324 = ~n1152 ;
  assign y325 = ~1'b0 ;
  assign y326 = ~1'b0 ;
  assign y327 = n1153 ;
  assign y328 = ~n1170 ;
  assign y329 = n1172 ;
  assign y330 = ~1'b0 ;
  assign y331 = ~n1180 ;
  assign y332 = n1189 ;
  assign y333 = n141 ;
  assign y334 = ~1'b0 ;
  assign y335 = ~n1190 ;
  assign y336 = ~n1201 ;
  assign y337 = ~1'b0 ;
  assign y338 = ~n1202 ;
  assign y339 = ~n1204 ;
  assign y340 = ~n1205 ;
  assign y341 = ~1'b0 ;
  assign y342 = ~n1207 ;
  assign y343 = ~n1215 ;
  assign y344 = n1218 ;
  assign y345 = n1221 ;
  assign y346 = ~n1225 ;
  assign y347 = ~n1227 ;
  assign y348 = n1236 ;
  assign y349 = n1244 ;
  assign y350 = ~n1256 ;
  assign y351 = n1261 ;
  assign y352 = ~1'b0 ;
  assign y353 = ~n1262 ;
  assign y354 = n1264 ;
  assign y355 = ~n1267 ;
  assign y356 = n1271 ;
  assign y357 = ~n1272 ;
  assign y358 = ~n1274 ;
  assign y359 = n1285 ;
  assign y360 = ~n1286 ;
  assign y361 = ~n1288 ;
  assign y362 = ~n1290 ;
  assign y363 = ~n1291 ;
  assign y364 = n1299 ;
  assign y365 = n1310 ;
  assign y366 = ~n1320 ;
  assign y367 = ~n1321 ;
  assign y368 = ~n1323 ;
  assign y369 = n1328 ;
  assign y370 = n1334 ;
  assign y371 = ~1'b0 ;
  assign y372 = ~n1340 ;
  assign y373 = 1'b0 ;
  assign y374 = ~1'b0 ;
  assign y375 = ~n1342 ;
  assign y376 = n1343 ;
  assign y377 = n1350 ;
  assign y378 = ~n1355 ;
  assign y379 = n1357 ;
  assign y380 = n1364 ;
  assign y381 = ~n1369 ;
  assign y382 = n1377 ;
  assign y383 = n1378 ;
  assign y384 = n1388 ;
  assign y385 = n1389 ;
  assign y386 = ~n1390 ;
  assign y387 = ~n1396 ;
  assign y388 = ~n1399 ;
  assign y389 = ~1'b0 ;
  assign y390 = n1404 ;
  assign y391 = n1407 ;
  assign y392 = ~n1417 ;
  assign y393 = ~n1419 ;
  assign y394 = n1432 ;
  assign y395 = n1434 ;
  assign y396 = ~n1439 ;
  assign y397 = ~n1444 ;
  assign y398 = ~n1199 ;
  assign y399 = n1447 ;
  assign y400 = n1449 ;
  assign y401 = ~n1453 ;
  assign y402 = ~n1458 ;
  assign y403 = ~n1460 ;
  assign y404 = ~n1463 ;
  assign y405 = ~n1464 ;
  assign y406 = n1475 ;
  assign y407 = ~n1484 ;
  assign y408 = n1488 ;
  assign y409 = ~n1493 ;
  assign y410 = ~n1498 ;
  assign y411 = n1501 ;
  assign y412 = ~n1504 ;
  assign y413 = n1507 ;
  assign y414 = ~n1509 ;
  assign y415 = ~n1513 ;
  assign y416 = ~n1516 ;
  assign y417 = ~n1519 ;
  assign y418 = ~1'b0 ;
  assign y419 = ~n1520 ;
  assign y420 = n1525 ;
  assign y421 = ~n1537 ;
  assign y422 = n1541 ;
  assign y423 = n1555 ;
  assign y424 = ~n1558 ;
  assign y425 = n1569 ;
  assign y426 = ~n1570 ;
  assign y427 = n1574 ;
  assign y428 = ~1'b0 ;
  assign y429 = n1576 ;
  assign y430 = ~n1580 ;
  assign y431 = ~1'b0 ;
  assign y432 = 1'b0 ;
  assign y433 = ~n1588 ;
  assign y434 = n1591 ;
  assign y435 = ~n1594 ;
  assign y436 = n1598 ;
  assign y437 = ~n1601 ;
  assign y438 = ~1'b0 ;
  assign y439 = ~n1603 ;
  assign y440 = ~n1607 ;
  assign y441 = n1609 ;
  assign y442 = n1612 ;
  assign y443 = ~n1616 ;
  assign y444 = ~n1619 ;
  assign y445 = n1622 ;
  assign y446 = ~1'b0 ;
  assign y447 = n1629 ;
  assign y448 = ~n1639 ;
  assign y449 = n1640 ;
  assign y450 = n1642 ;
  assign y451 = n1643 ;
  assign y452 = n1646 ;
  assign y453 = n1653 ;
  assign y454 = ~n1654 ;
  assign y455 = n1656 ;
  assign y456 = n1660 ;
  assign y457 = ~n1661 ;
  assign y458 = n1664 ;
  assign y459 = ~n1676 ;
  assign y460 = n1679 ;
  assign y461 = ~n1682 ;
  assign y462 = ~1'b0 ;
  assign y463 = n1685 ;
  assign y464 = n1691 ;
  assign y465 = ~n1692 ;
  assign y466 = ~n1698 ;
  assign y467 = n1700 ;
  assign y468 = ~n1701 ;
  assign y469 = ~n1705 ;
  assign y470 = n1711 ;
  assign y471 = ~n1713 ;
  assign y472 = ~n1714 ;
  assign y473 = ~n1717 ;
  assign y474 = ~n1718 ;
  assign y475 = ~n1728 ;
  assign y476 = n1731 ;
  assign y477 = ~n1732 ;
  assign y478 = ~n1735 ;
  assign y479 = 1'b0 ;
  assign y480 = ~n1738 ;
  assign y481 = n1741 ;
  assign y482 = n1744 ;
  assign y483 = ~1'b0 ;
  assign y484 = ~n1749 ;
  assign y485 = n1757 ;
  assign y486 = ~n1760 ;
  assign y487 = n1761 ;
  assign y488 = ~1'b0 ;
  assign y489 = n1765 ;
  assign y490 = n1767 ;
  assign y491 = ~1'b0 ;
  assign y492 = n1771 ;
  assign y493 = n1772 ;
  assign y494 = ~n1773 ;
  assign y495 = n1781 ;
  assign y496 = ~n1794 ;
  assign y497 = ~1'b0 ;
  assign y498 = n1798 ;
  assign y499 = n1800 ;
  assign y500 = ~1'b0 ;
  assign y501 = ~n1803 ;
  assign y502 = ~n1806 ;
  assign y503 = ~n1807 ;
  assign y504 = n1666 ;
  assign y505 = n1808 ;
  assign y506 = ~n1813 ;
  assign y507 = n1816 ;
  assign y508 = n1822 ;
  assign y509 = ~n1824 ;
  assign y510 = n1828 ;
  assign y511 = ~n1830 ;
  assign y512 = n1832 ;
  assign y513 = n1835 ;
  assign y514 = n1840 ;
  assign y515 = ~1'b0 ;
  assign y516 = ~n1845 ;
  assign y517 = ~n1848 ;
  assign y518 = n1850 ;
  assign y519 = ~1'b0 ;
  assign y520 = ~1'b0 ;
  assign y521 = n1852 ;
  assign y522 = ~n1855 ;
  assign y523 = ~n1866 ;
  assign y524 = n1874 ;
  assign y525 = ~n1876 ;
  assign y526 = n1882 ;
  assign y527 = ~n1889 ;
  assign y528 = n1893 ;
  assign y529 = ~1'b0 ;
  assign y530 = ~1'b0 ;
  assign y531 = ~n580 ;
  assign y532 = n1898 ;
  assign y533 = ~n1903 ;
  assign y534 = ~n1911 ;
  assign y535 = ~n1913 ;
  assign y536 = ~n1916 ;
  assign y537 = n1699 ;
  assign y538 = ~1'b0 ;
  assign y539 = ~n1921 ;
  assign y540 = n1922 ;
  assign y541 = ~1'b0 ;
  assign y542 = ~n1924 ;
  assign y543 = n457 ;
  assign y544 = n1925 ;
  assign y545 = ~n1928 ;
  assign y546 = ~n1932 ;
  assign y547 = ~1'b0 ;
  assign y548 = ~n1938 ;
  assign y549 = ~n1940 ;
  assign y550 = ~n1951 ;
  assign y551 = ~n1955 ;
  assign y552 = ~n390 ;
  assign y553 = n1961 ;
  assign y554 = n1968 ;
  assign y555 = ~n1969 ;
  assign y556 = ~n1974 ;
  assign y557 = ~1'b0 ;
  assign y558 = ~1'b0 ;
  assign y559 = n1978 ;
  assign y560 = ~n1979 ;
  assign y561 = ~n1990 ;
  assign y562 = ~n1992 ;
  assign y563 = ~n2000 ;
  assign y564 = ~n2004 ;
  assign y565 = ~n2007 ;
  assign y566 = ~1'b0 ;
  assign y567 = ~n1057 ;
  assign y568 = ~n307 ;
  assign y569 = ~n2013 ;
  assign y570 = n2018 ;
  assign y571 = ~n2020 ;
  assign y572 = n2022 ;
  assign y573 = n2023 ;
  assign y574 = ~n2025 ;
  assign y575 = n2031 ;
  assign y576 = ~1'b0 ;
  assign y577 = ~n2035 ;
  assign y578 = ~1'b0 ;
  assign y579 = n2036 ;
  assign y580 = ~1'b0 ;
  assign y581 = ~n2042 ;
  assign y582 = n2044 ;
  assign y583 = n2038 ;
  assign y584 = ~n2046 ;
  assign y585 = ~n2048 ;
  assign y586 = ~n2051 ;
  assign y587 = ~1'b0 ;
  assign y588 = ~n2053 ;
  assign y589 = ~1'b0 ;
  assign y590 = ~n2059 ;
  assign y591 = n2069 ;
  assign y592 = ~1'b0 ;
  assign y593 = ~n2071 ;
  assign y594 = n2074 ;
  assign y595 = n2076 ;
  assign y596 = n2088 ;
  assign y597 = ~1'b0 ;
  assign y598 = ~n2107 ;
  assign y599 = ~n2108 ;
  assign y600 = ~n2113 ;
  assign y601 = ~1'b0 ;
  assign y602 = ~1'b0 ;
  assign y603 = ~n2115 ;
  assign y604 = n2118 ;
  assign y605 = ~n2127 ;
  assign y606 = ~n2132 ;
  assign y607 = ~1'b0 ;
  assign y608 = n2138 ;
  assign y609 = n2140 ;
  assign y610 = n2141 ;
  assign y611 = n2142 ;
  assign y612 = ~1'b0 ;
  assign y613 = n2146 ;
  assign y614 = ~n2147 ;
  assign y615 = ~n2153 ;
  assign y616 = ~n2167 ;
  assign y617 = ~1'b0 ;
  assign y618 = ~1'b0 ;
  assign y619 = ~n2174 ;
  assign y620 = ~1'b0 ;
  assign y621 = n2177 ;
  assign y622 = ~n2180 ;
  assign y623 = ~1'b0 ;
  assign y624 = n2181 ;
  assign y625 = n2182 ;
  assign y626 = ~1'b0 ;
  assign y627 = n2184 ;
  assign y628 = n2186 ;
  assign y629 = ~n2188 ;
  assign y630 = ~n2191 ;
  assign y631 = n2192 ;
  assign y632 = ~1'b0 ;
  assign y633 = ~n2195 ;
  assign y634 = n2200 ;
  assign y635 = n2205 ;
  assign y636 = ~n2211 ;
  assign y637 = ~n2213 ;
  assign y638 = ~n2220 ;
  assign y639 = ~1'b0 ;
  assign y640 = ~1'b0 ;
  assign y641 = n2222 ;
  assign y642 = n2223 ;
  assign y643 = n2225 ;
  assign y644 = ~n2229 ;
  assign y645 = ~n2231 ;
  assign y646 = ~n2233 ;
  assign y647 = n2235 ;
  assign y648 = ~1'b0 ;
  assign y649 = n2243 ;
  assign y650 = ~n2244 ;
  assign y651 = n2247 ;
  assign y652 = n2254 ;
  assign y653 = ~n2272 ;
  assign y654 = n194 ;
  assign y655 = ~1'b0 ;
  assign y656 = ~1'b0 ;
  assign y657 = n2279 ;
  assign y658 = n2282 ;
  assign y659 = n2286 ;
  assign y660 = n2289 ;
  assign y661 = ~n2299 ;
  assign y662 = ~n2300 ;
  assign y663 = n2301 ;
  assign y664 = n2311 ;
  assign y665 = ~n2316 ;
  assign y666 = ~n2329 ;
  assign y667 = ~n2335 ;
  assign y668 = ~n2337 ;
  assign y669 = ~n2339 ;
  assign y670 = n2344 ;
  assign y671 = n2348 ;
  assign y672 = ~n2352 ;
  assign y673 = ~n2353 ;
  assign y674 = ~1'b0 ;
  assign y675 = ~n2356 ;
  assign y676 = n2361 ;
  assign y677 = ~n2364 ;
  assign y678 = ~1'b0 ;
  assign y679 = ~n2368 ;
  assign y680 = n2369 ;
  assign y681 = ~1'b0 ;
  assign y682 = ~n2370 ;
  assign y683 = ~n2373 ;
  assign y684 = ~n2375 ;
  assign y685 = ~n2380 ;
  assign y686 = n2391 ;
  assign y687 = n2400 ;
  assign y688 = ~n2401 ;
  assign y689 = n2406 ;
  assign y690 = n2408 ;
  assign y691 = ~n2409 ;
  assign y692 = ~1'b0 ;
  assign y693 = ~1'b0 ;
  assign y694 = n2415 ;
  assign y695 = ~n2422 ;
  assign y696 = ~n2426 ;
  assign y697 = n2430 ;
  assign y698 = ~n2433 ;
  assign y699 = ~n2438 ;
  assign y700 = ~1'b0 ;
  assign y701 = n2441 ;
  assign y702 = n2444 ;
  assign y703 = ~n2445 ;
  assign y704 = n2449 ;
  assign y705 = ~1'b0 ;
  assign y706 = n2451 ;
  assign y707 = ~n2454 ;
  assign y708 = n2457 ;
  assign y709 = ~1'b0 ;
  assign y710 = n2458 ;
  assign y711 = n2463 ;
  assign y712 = ~1'b0 ;
  assign y713 = ~1'b0 ;
  assign y714 = n2467 ;
  assign y715 = ~n2470 ;
  assign y716 = n2475 ;
  assign y717 = n2476 ;
  assign y718 = n2486 ;
  assign y719 = n2487 ;
  assign y720 = ~n2490 ;
  assign y721 = ~n2496 ;
  assign y722 = n2498 ;
  assign y723 = n2509 ;
  assign y724 = ~n2520 ;
  assign y725 = n2523 ;
  assign y726 = ~n2527 ;
  assign y727 = ~n2545 ;
  assign y728 = n2550 ;
  assign y729 = ~n1235 ;
  assign y730 = n2552 ;
  assign y731 = ~1'b0 ;
  assign y732 = ~n2553 ;
  assign y733 = ~n2561 ;
  assign y734 = ~n2565 ;
  assign y735 = n2568 ;
  assign y736 = ~1'b0 ;
  assign y737 = ~n2573 ;
  assign y738 = ~1'b0 ;
  assign y739 = ~1'b0 ;
  assign y740 = ~n2579 ;
  assign y741 = ~n2586 ;
  assign y742 = n2589 ;
  assign y743 = n2590 ;
  assign y744 = ~n2598 ;
  assign y745 = n2602 ;
  assign y746 = ~n2612 ;
  assign y747 = ~n2613 ;
  assign y748 = ~n2615 ;
  assign y749 = n2616 ;
  assign y750 = ~1'b0 ;
  assign y751 = ~1'b0 ;
  assign y752 = ~1'b0 ;
  assign y753 = n2624 ;
  assign y754 = ~n2625 ;
  assign y755 = n2629 ;
  assign y756 = ~n2632 ;
  assign y757 = n2638 ;
  assign y758 = ~1'b0 ;
  assign y759 = ~1'b0 ;
  assign y760 = n2639 ;
  assign y761 = n2641 ;
  assign y762 = n2647 ;
  assign y763 = ~1'b0 ;
  assign y764 = n2653 ;
  assign y765 = n2654 ;
  assign y766 = ~1'b0 ;
  assign y767 = n2655 ;
  assign y768 = ~n2657 ;
  assign y769 = n2658 ;
  assign y770 = ~1'b0 ;
  assign y771 = n2665 ;
  assign y772 = n2666 ;
  assign y773 = n2667 ;
  assign y774 = ~n2670 ;
  assign y775 = n2671 ;
  assign y776 = n2676 ;
  assign y777 = n2681 ;
  assign y778 = n2686 ;
  assign y779 = x74 ;
  assign y780 = ~n2688 ;
  assign y781 = n2689 ;
  assign y782 = n2699 ;
  assign y783 = n2703 ;
  assign y784 = ~n2709 ;
  assign y785 = ~n2713 ;
  assign y786 = n2723 ;
  assign y787 = n2729 ;
  assign y788 = n2733 ;
  assign y789 = ~n2738 ;
  assign y790 = n2740 ;
  assign y791 = ~1'b0 ;
  assign y792 = ~n2742 ;
  assign y793 = ~n2743 ;
  assign y794 = ~n2745 ;
  assign y795 = ~1'b0 ;
  assign y796 = n2752 ;
  assign y797 = ~n154 ;
  assign y798 = n2754 ;
  assign y799 = ~n2757 ;
  assign y800 = ~1'b0 ;
  assign y801 = ~n2761 ;
  assign y802 = n2762 ;
  assign y803 = n2764 ;
  assign y804 = ~n2769 ;
  assign y805 = n2783 ;
  assign y806 = ~n2784 ;
  assign y807 = ~1'b0 ;
  assign y808 = ~n2785 ;
  assign y809 = n2788 ;
  assign y810 = ~n2790 ;
  assign y811 = n2802 ;
  assign y812 = n2816 ;
  assign y813 = n2817 ;
  assign y814 = n2821 ;
  assign y815 = n2823 ;
  assign y816 = n2827 ;
  assign y817 = ~1'b0 ;
  assign y818 = n2831 ;
  assign y819 = n2833 ;
  assign y820 = n2842 ;
  assign y821 = n2843 ;
  assign y822 = ~n2844 ;
  assign y823 = ~n2849 ;
  assign y824 = ~n2851 ;
  assign y825 = n2853 ;
  assign y826 = ~n2858 ;
  assign y827 = ~n2863 ;
  assign y828 = ~1'b0 ;
  assign y829 = n2871 ;
  assign y830 = ~n2875 ;
  assign y831 = n2878 ;
  assign y832 = ~n2881 ;
  assign y833 = n2886 ;
  assign y834 = n2887 ;
  assign y835 = ~n2891 ;
  assign y836 = ~n2894 ;
  assign y837 = ~n2896 ;
  assign y838 = n2897 ;
  assign y839 = ~n2899 ;
  assign y840 = n2903 ;
  assign y841 = ~n2908 ;
  assign y842 = ~1'b0 ;
  assign y843 = ~n2910 ;
  assign y844 = n2912 ;
  assign y845 = n2919 ;
  assign y846 = 1'b0 ;
  assign y847 = ~n2925 ;
  assign y848 = ~1'b0 ;
  assign y849 = n2926 ;
  assign y850 = n2929 ;
  assign y851 = ~1'b0 ;
  assign y852 = n306 ;
  assign y853 = ~n2931 ;
  assign y854 = ~1'b0 ;
  assign y855 = n2932 ;
  assign y856 = ~n2941 ;
  assign y857 = n2949 ;
  assign y858 = n2950 ;
  assign y859 = ~n2955 ;
  assign y860 = n1235 ;
  assign y861 = n2964 ;
  assign y862 = n2968 ;
  assign y863 = ~n2975 ;
  assign y864 = n2977 ;
  assign y865 = ~1'b0 ;
  assign y866 = n2980 ;
  assign y867 = n2982 ;
  assign y868 = n2985 ;
  assign y869 = n2989 ;
  assign y870 = n2990 ;
  assign y871 = ~1'b0 ;
  assign y872 = n2993 ;
  assign y873 = ~n2996 ;
  assign y874 = ~1'b0 ;
  assign y875 = n3001 ;
  assign y876 = ~n3004 ;
  assign y877 = ~n3010 ;
  assign y878 = ~n3026 ;
  assign y879 = ~n3028 ;
  assign y880 = ~n3036 ;
  assign y881 = ~n3037 ;
  assign y882 = n3045 ;
  assign y883 = 1'b0 ;
  assign y884 = ~n3047 ;
  assign y885 = n3054 ;
  assign y886 = ~n3056 ;
  assign y887 = ~n3063 ;
  assign y888 = ~1'b0 ;
  assign y889 = ~n3068 ;
  assign y890 = ~n3070 ;
  assign y891 = ~n3071 ;
  assign y892 = ~n3074 ;
  assign y893 = n3076 ;
  assign y894 = ~n3077 ;
  assign y895 = n3081 ;
  assign y896 = n3086 ;
  assign y897 = n3095 ;
  assign y898 = ~1'b0 ;
  assign y899 = ~n3099 ;
  assign y900 = ~1'b0 ;
  assign y901 = n3101 ;
  assign y902 = ~n1762 ;
  assign y903 = ~n3103 ;
  assign y904 = n3105 ;
  assign y905 = ~1'b0 ;
  assign y906 = ~n3110 ;
  assign y907 = n3111 ;
  assign y908 = n3116 ;
  assign y909 = n3118 ;
  assign y910 = ~n3120 ;
  assign y911 = ~n3121 ;
  assign y912 = ~n3123 ;
  assign y913 = ~n3128 ;
  assign y914 = n3133 ;
  assign y915 = n3135 ;
  assign y916 = n1484 ;
  assign y917 = n3142 ;
  assign y918 = n3145 ;
  assign y919 = n3151 ;
  assign y920 = n3152 ;
  assign y921 = ~1'b0 ;
  assign y922 = n3153 ;
  assign y923 = ~n3154 ;
  assign y924 = n3164 ;
  assign y925 = n3167 ;
  assign y926 = n3177 ;
  assign y927 = n3183 ;
  assign y928 = ~1'b0 ;
  assign y929 = n3190 ;
  assign y930 = ~1'b0 ;
  assign y931 = ~n3195 ;
  assign y932 = ~n3207 ;
  assign y933 = n3209 ;
  assign y934 = n3210 ;
  assign y935 = ~n3213 ;
  assign y936 = ~n3222 ;
  assign y937 = ~n3224 ;
  assign y938 = n3225 ;
  assign y939 = n3230 ;
  assign y940 = ~1'b0 ;
  assign y941 = ~n3234 ;
  assign y942 = n3238 ;
  assign y943 = n3242 ;
  assign y944 = n3251 ;
  assign y945 = n3252 ;
  assign y946 = n3262 ;
  assign y947 = n3264 ;
  assign y948 = n3265 ;
  assign y949 = ~n3270 ;
  assign y950 = ~n3276 ;
  assign y951 = n466 ;
  assign y952 = ~n3279 ;
  assign y953 = ~n3282 ;
  assign y954 = n3290 ;
  assign y955 = n3293 ;
  assign y956 = n3297 ;
  assign y957 = n3299 ;
  assign y958 = n3306 ;
  assign y959 = n1333 ;
  assign y960 = n3310 ;
  assign y961 = ~n3311 ;
  assign y962 = n3314 ;
  assign y963 = n3315 ;
  assign y964 = n3318 ;
  assign y965 = ~1'b0 ;
  assign y966 = ~1'b0 ;
  assign y967 = ~n3322 ;
  assign y968 = ~n3330 ;
  assign y969 = ~1'b0 ;
  assign y970 = ~n3334 ;
  assign y971 = ~n3335 ;
  assign y972 = ~n3340 ;
  assign y973 = ~1'b0 ;
  assign y974 = n3346 ;
  assign y975 = n3347 ;
  assign y976 = ~n3355 ;
  assign y977 = ~1'b0 ;
  assign y978 = ~n3360 ;
  assign y979 = n3363 ;
  assign y980 = ~n3364 ;
  assign y981 = ~1'b0 ;
  assign y982 = n3366 ;
  assign y983 = ~n3380 ;
  assign y984 = n3385 ;
  assign y985 = n3388 ;
  assign y986 = ~n3389 ;
  assign y987 = n3391 ;
  assign y988 = n3398 ;
  assign y989 = n3403 ;
  assign y990 = n3407 ;
  assign y991 = n3415 ;
  assign y992 = ~1'b0 ;
  assign y993 = ~1'b0 ;
  assign y994 = ~n3416 ;
  assign y995 = n3417 ;
  assign y996 = n3426 ;
  assign y997 = n3429 ;
  assign y998 = ~n3440 ;
  assign y999 = ~1'b0 ;
  assign y1000 = n3442 ;
  assign y1001 = n3443 ;
  assign y1002 = ~n3446 ;
  assign y1003 = ~n3447 ;
  assign y1004 = n3450 ;
  assign y1005 = n3454 ;
  assign y1006 = n3465 ;
  assign y1007 = ~n3467 ;
  assign y1008 = n3475 ;
  assign y1009 = ~n3476 ;
  assign y1010 = n3480 ;
  assign y1011 = n3486 ;
  assign y1012 = ~n3492 ;
  assign y1013 = ~n3493 ;
  assign y1014 = ~n3499 ;
  assign y1015 = ~n3503 ;
  assign y1016 = n3505 ;
  assign y1017 = n3510 ;
  assign y1018 = ~n3511 ;
  assign y1019 = ~1'b0 ;
  assign y1020 = n3524 ;
  assign y1021 = n3525 ;
  assign y1022 = ~n3527 ;
  assign y1023 = ~1'b0 ;
  assign y1024 = n3529 ;
  assign y1025 = n3530 ;
  assign y1026 = ~n3536 ;
  assign y1027 = n3542 ;
  assign y1028 = n3544 ;
  assign y1029 = ~n3546 ;
  assign y1030 = ~n3548 ;
  assign y1031 = 1'b0 ;
  assign y1032 = ~n3550 ;
  assign y1033 = ~n3559 ;
  assign y1034 = ~n3560 ;
  assign y1035 = n3573 ;
  assign y1036 = n3575 ;
  assign y1037 = n3576 ;
  assign y1038 = ~1'b0 ;
  assign y1039 = ~1'b0 ;
  assign y1040 = ~n3585 ;
  assign y1041 = ~n3587 ;
  assign y1042 = ~n3592 ;
  assign y1043 = n3596 ;
  assign y1044 = n3605 ;
  assign y1045 = ~n3608 ;
  assign y1046 = ~n3610 ;
  assign y1047 = ~n3611 ;
  assign y1048 = ~n3612 ;
  assign y1049 = ~n3620 ;
  assign y1050 = n3622 ;
  assign y1051 = n3629 ;
  assign y1052 = n3630 ;
  assign y1053 = n3631 ;
  assign y1054 = n3644 ;
  assign y1055 = n3646 ;
  assign y1056 = ~n3654 ;
  assign y1057 = n3655 ;
  assign y1058 = n3658 ;
  assign y1059 = ~n3670 ;
  assign y1060 = ~n3672 ;
  assign y1061 = ~n3680 ;
  assign y1062 = ~1'b0 ;
  assign y1063 = ~n3682 ;
  assign y1064 = ~n3687 ;
  assign y1065 = ~n3697 ;
  assign y1066 = ~1'b0 ;
  assign y1067 = n3698 ;
  assign y1068 = n3701 ;
  assign y1069 = ~n3706 ;
  assign y1070 = n3713 ;
  assign y1071 = ~n3719 ;
  assign y1072 = ~n3722 ;
  assign y1073 = ~n3724 ;
  assign y1074 = ~n3734 ;
  assign y1075 = n3737 ;
  assign y1076 = ~n3744 ;
  assign y1077 = ~n3748 ;
  assign y1078 = ~n3752 ;
  assign y1079 = n3754 ;
  assign y1080 = ~n3757 ;
  assign y1081 = ~n3764 ;
  assign y1082 = ~n3769 ;
  assign y1083 = n3775 ;
  assign y1084 = n2732 ;
  assign y1085 = n3777 ;
  assign y1086 = ~n3780 ;
  assign y1087 = ~1'b0 ;
  assign y1088 = ~1'b0 ;
  assign y1089 = ~n3781 ;
  assign y1090 = n3784 ;
  assign y1091 = ~1'b0 ;
  assign y1092 = ~n3637 ;
  assign y1093 = ~1'b0 ;
  assign y1094 = n3786 ;
  assign y1095 = ~n3788 ;
  assign y1096 = 1'b0 ;
  assign y1097 = ~1'b0 ;
  assign y1098 = ~n3790 ;
  assign y1099 = ~1'b0 ;
  assign y1100 = n3791 ;
  assign y1101 = ~n3793 ;
  assign y1102 = n3796 ;
  assign y1103 = n3797 ;
  assign y1104 = n3798 ;
  assign y1105 = ~1'b0 ;
  assign y1106 = ~n3801 ;
  assign y1107 = ~n3806 ;
  assign y1108 = ~n3809 ;
  assign y1109 = ~n3816 ;
  assign y1110 = n3822 ;
  assign y1111 = ~1'b0 ;
  assign y1112 = ~n3823 ;
  assign y1113 = ~n3829 ;
  assign y1114 = n3830 ;
  assign y1115 = ~n3836 ;
  assign y1116 = ~n3838 ;
  assign y1117 = ~n3851 ;
  assign y1118 = ~n3854 ;
  assign y1119 = ~n3856 ;
  assign y1120 = n3865 ;
  assign y1121 = ~n3867 ;
  assign y1122 = n3881 ;
  assign y1123 = ~1'b0 ;
  assign y1124 = ~n3887 ;
  assign y1125 = n3890 ;
  assign y1126 = ~n3893 ;
  assign y1127 = ~n3894 ;
  assign y1128 = ~n3897 ;
  assign y1129 = ~n3907 ;
  assign y1130 = ~n3915 ;
  assign y1131 = n3921 ;
  assign y1132 = n3925 ;
  assign y1133 = n3926 ;
  assign y1134 = n3927 ;
  assign y1135 = n3935 ;
  assign y1136 = n3940 ;
  assign y1137 = n3942 ;
  assign y1138 = n3944 ;
  assign y1139 = ~n3947 ;
  assign y1140 = ~n3949 ;
  assign y1141 = ~n3952 ;
  assign y1142 = ~n3955 ;
  assign y1143 = ~n3961 ;
  assign y1144 = n3962 ;
  assign y1145 = ~n3966 ;
  assign y1146 = ~1'b0 ;
  assign y1147 = n3972 ;
  assign y1148 = n3973 ;
  assign y1149 = n3976 ;
  assign y1150 = ~n3986 ;
  assign y1151 = n3991 ;
  assign y1152 = ~n3992 ;
  assign y1153 = ~1'b0 ;
  assign y1154 = n4000 ;
  assign y1155 = ~n4002 ;
  assign y1156 = ~n4006 ;
  assign y1157 = ~n4008 ;
  assign y1158 = ~1'b0 ;
  assign y1159 = ~1'b0 ;
  assign y1160 = ~n4017 ;
  assign y1161 = ~1'b0 ;
  assign y1162 = ~n4023 ;
  assign y1163 = ~1'b0 ;
  assign y1164 = n4026 ;
  assign y1165 = ~1'b0 ;
  assign y1166 = 1'b0 ;
  assign y1167 = ~n4032 ;
  assign y1168 = ~1'b0 ;
  assign y1169 = n4034 ;
  assign y1170 = ~1'b0 ;
  assign y1171 = n4039 ;
  assign y1172 = ~n4044 ;
  assign y1173 = ~1'b0 ;
  assign y1174 = ~n4050 ;
  assign y1175 = ~n4051 ;
  assign y1176 = ~n4058 ;
  assign y1177 = n4060 ;
  assign y1178 = ~1'b0 ;
  assign y1179 = ~1'b0 ;
  assign y1180 = ~1'b0 ;
  assign y1181 = n4061 ;
  assign y1182 = n4064 ;
  assign y1183 = ~n4071 ;
  assign y1184 = ~1'b0 ;
  assign y1185 = n4072 ;
  assign y1186 = n4075 ;
  assign y1187 = ~n4081 ;
  assign y1188 = ~n4084 ;
  assign y1189 = ~n4087 ;
  assign y1190 = n4092 ;
  assign y1191 = ~n4093 ;
  assign y1192 = n4107 ;
  assign y1193 = ~1'b0 ;
  assign y1194 = ~1'b0 ;
  assign y1195 = n4108 ;
  assign y1196 = n4109 ;
  assign y1197 = n4110 ;
  assign y1198 = ~n4114 ;
  assign y1199 = n4115 ;
  assign y1200 = ~n4116 ;
  assign y1201 = n4125 ;
  assign y1202 = n4129 ;
  assign y1203 = ~n4134 ;
  assign y1204 = n4141 ;
  assign y1205 = ~n4142 ;
  assign y1206 = ~1'b0 ;
  assign y1207 = n4144 ;
  assign y1208 = ~n4145 ;
  assign y1209 = ~n4148 ;
  assign y1210 = n4152 ;
  assign y1211 = ~1'b0 ;
  assign y1212 = n4155 ;
  assign y1213 = ~n4171 ;
  assign y1214 = ~n4175 ;
  assign y1215 = n4193 ;
  assign y1216 = n4198 ;
  assign y1217 = ~n4202 ;
  assign y1218 = ~n4206 ;
  assign y1219 = n4207 ;
  assign y1220 = ~n4210 ;
  assign y1221 = ~n4215 ;
  assign y1222 = n4219 ;
  assign y1223 = ~n4220 ;
  assign y1224 = n4224 ;
  assign y1225 = n4227 ;
  assign y1226 = n4232 ;
  assign y1227 = n4240 ;
  assign y1228 = n4242 ;
  assign y1229 = ~n4245 ;
  assign y1230 = ~n4250 ;
  assign y1231 = n4255 ;
  assign y1232 = n4261 ;
  assign y1233 = ~n4266 ;
  assign y1234 = n4271 ;
  assign y1235 = ~n1695 ;
  assign y1236 = ~n4272 ;
  assign y1237 = n4275 ;
  assign y1238 = n4277 ;
  assign y1239 = ~1'b0 ;
  assign y1240 = n4278 ;
  assign y1241 = ~n4279 ;
  assign y1242 = ~n4281 ;
  assign y1243 = ~1'b0 ;
  assign y1244 = n4282 ;
  assign y1245 = n4297 ;
  assign y1246 = n4305 ;
  assign y1247 = n4306 ;
  assign y1248 = ~n4311 ;
  assign y1249 = ~n4315 ;
  assign y1250 = n4323 ;
  assign y1251 = ~1'b0 ;
  assign y1252 = ~n4325 ;
  assign y1253 = n4334 ;
  assign y1254 = ~1'b0 ;
  assign y1255 = n4335 ;
  assign y1256 = ~n4336 ;
  assign y1257 = n4341 ;
  assign y1258 = ~n4343 ;
  assign y1259 = ~1'b0 ;
  assign y1260 = n4346 ;
  assign y1261 = ~n4347 ;
  assign y1262 = ~1'b0 ;
  assign y1263 = n4361 ;
  assign y1264 = ~1'b0 ;
  assign y1265 = ~n4363 ;
  assign y1266 = n4365 ;
  assign y1267 = n4367 ;
  assign y1268 = ~n4376 ;
  assign y1269 = ~n4378 ;
  assign y1270 = n4379 ;
  assign y1271 = ~n4382 ;
  assign y1272 = ~n4399 ;
  assign y1273 = ~n4403 ;
  assign y1274 = n4406 ;
  assign y1275 = ~n4408 ;
  assign y1276 = n4409 ;
  assign y1277 = ~n4412 ;
  assign y1278 = n4417 ;
  assign y1279 = n4422 ;
  assign y1280 = n4426 ;
  assign y1281 = ~n4427 ;
  assign y1282 = ~n4432 ;
  assign y1283 = ~n4434 ;
  assign y1284 = n4441 ;
  assign y1285 = n4443 ;
  assign y1286 = n4445 ;
  assign y1287 = n4448 ;
  assign y1288 = n4450 ;
  assign y1289 = n4455 ;
  assign y1290 = ~n4456 ;
  assign y1291 = ~n4459 ;
  assign y1292 = ~n4462 ;
  assign y1293 = n4465 ;
  assign y1294 = ~n4472 ;
  assign y1295 = ~n4474 ;
  assign y1296 = n4475 ;
  assign y1297 = n4483 ;
  assign y1298 = n4487 ;
  assign y1299 = n4489 ;
  assign y1300 = n4500 ;
  assign y1301 = ~n270 ;
  assign y1302 = ~n4503 ;
  assign y1303 = n2199 ;
  assign y1304 = ~n4505 ;
  assign y1305 = ~n4511 ;
  assign y1306 = n4513 ;
  assign y1307 = ~n4517 ;
  assign y1308 = n4525 ;
  assign y1309 = ~1'b0 ;
  assign y1310 = ~n620 ;
  assign y1311 = n4526 ;
  assign y1312 = ~n4527 ;
  assign y1313 = n4528 ;
  assign y1314 = ~n4529 ;
  assign y1315 = ~n4532 ;
  assign y1316 = ~1'b0 ;
  assign y1317 = n4543 ;
  assign y1318 = ~n689 ;
  assign y1319 = n4544 ;
  assign y1320 = ~1'b0 ;
  assign y1321 = ~1'b0 ;
  assign y1322 = ~n4545 ;
  assign y1323 = ~n4548 ;
  assign y1324 = ~n4567 ;
  assign y1325 = n4569 ;
  assign y1326 = ~n4572 ;
  assign y1327 = ~n4573 ;
  assign y1328 = ~n4574 ;
  assign y1329 = ~n4578 ;
  assign y1330 = n4585 ;
  assign y1331 = ~1'b0 ;
  assign y1332 = ~1'b0 ;
  assign y1333 = ~1'b0 ;
  assign y1334 = n401 ;
  assign y1335 = n4587 ;
  assign y1336 = n4589 ;
  assign y1337 = ~1'b0 ;
  assign y1338 = n4597 ;
  assign y1339 = ~n4600 ;
  assign y1340 = ~n4605 ;
  assign y1341 = ~n4614 ;
  assign y1342 = n4615 ;
  assign y1343 = n4621 ;
  assign y1344 = n4622 ;
  assign y1345 = ~1'b0 ;
  assign y1346 = n4624 ;
  assign y1347 = ~n4629 ;
  assign y1348 = n4636 ;
  assign y1349 = ~1'b0 ;
  assign y1350 = n4637 ;
  assign y1351 = n1692 ;
  assign y1352 = n4639 ;
  assign y1353 = n4640 ;
  assign y1354 = n4648 ;
  assign y1355 = ~n4656 ;
  assign y1356 = ~1'b0 ;
  assign y1357 = ~n4657 ;
  assign y1358 = ~n4671 ;
  assign y1359 = ~n4678 ;
  assign y1360 = n4679 ;
  assign y1361 = ~n4683 ;
  assign y1362 = n4690 ;
  assign y1363 = ~1'b0 ;
  assign y1364 = ~1'b0 ;
  assign y1365 = n4691 ;
  assign y1366 = n2639 ;
  assign y1367 = ~n4693 ;
  assign y1368 = n4694 ;
  assign y1369 = n4697 ;
  assign y1370 = ~n4700 ;
  assign y1371 = ~1'b0 ;
  assign y1372 = ~n4702 ;
  assign y1373 = ~1'b0 ;
  assign y1374 = ~1'b0 ;
  assign y1375 = n4706 ;
  assign y1376 = n4713 ;
  assign y1377 = ~n4716 ;
  assign y1378 = ~n4718 ;
  assign y1379 = n4719 ;
  assign y1380 = ~1'b0 ;
  assign y1381 = ~n4726 ;
  assign y1382 = ~n4727 ;
  assign y1383 = ~1'b0 ;
  assign y1384 = n4732 ;
  assign y1385 = n4736 ;
  assign y1386 = n4739 ;
  assign y1387 = n4740 ;
  assign y1388 = ~1'b0 ;
  assign y1389 = ~n2934 ;
  assign y1390 = ~n4741 ;
  assign y1391 = n4744 ;
  assign y1392 = n4750 ;
  assign y1393 = ~n4751 ;
  assign y1394 = n4752 ;
  assign y1395 = ~1'b0 ;
  assign y1396 = n4765 ;
  assign y1397 = n4766 ;
  assign y1398 = ~n4771 ;
  assign y1399 = ~n4777 ;
  assign y1400 = n4779 ;
  assign y1401 = ~1'b0 ;
  assign y1402 = ~n4783 ;
  assign y1403 = n4786 ;
  assign y1404 = n4793 ;
  assign y1405 = n4802 ;
  assign y1406 = n4804 ;
  assign y1407 = n4805 ;
  assign y1408 = ~n4810 ;
  assign y1409 = ~n4814 ;
  assign y1410 = ~n4819 ;
  assign y1411 = ~n4831 ;
  assign y1412 = ~n4838 ;
  assign y1413 = ~n4839 ;
  assign y1414 = ~n4842 ;
  assign y1415 = n4848 ;
  assign y1416 = ~n4851 ;
  assign y1417 = ~n4862 ;
  assign y1418 = n4864 ;
  assign y1419 = ~n4870 ;
  assign y1420 = ~1'b0 ;
  assign y1421 = ~n4872 ;
  assign y1422 = ~n4873 ;
  assign y1423 = n4874 ;
  assign y1424 = ~1'b0 ;
  assign y1425 = ~n4876 ;
  assign y1426 = ~n4880 ;
  assign y1427 = ~1'b0 ;
  assign y1428 = ~n4881 ;
  assign y1429 = ~n4882 ;
  assign y1430 = ~n4883 ;
  assign y1431 = n4890 ;
  assign y1432 = n4892 ;
  assign y1433 = n4895 ;
  assign y1434 = ~1'b0 ;
  assign y1435 = ~n4896 ;
  assign y1436 = ~n4900 ;
  assign y1437 = n4902 ;
  assign y1438 = ~n4905 ;
  assign y1439 = ~n2532 ;
  assign y1440 = ~n4907 ;
  assign y1441 = ~n4908 ;
  assign y1442 = n4918 ;
  assign y1443 = ~n4920 ;
  assign y1444 = ~n4927 ;
  assign y1445 = ~1'b0 ;
  assign y1446 = ~n4930 ;
  assign y1447 = ~1'b0 ;
  assign y1448 = ~n4944 ;
  assign y1449 = ~n4946 ;
  assign y1450 = ~1'b0 ;
  assign y1451 = ~n4948 ;
  assign y1452 = n4950 ;
  assign y1453 = n4952 ;
  assign y1454 = ~1'b0 ;
  assign y1455 = n4960 ;
  assign y1456 = ~n4964 ;
  assign y1457 = ~n4970 ;
  assign y1458 = ~n4973 ;
  assign y1459 = ~n4987 ;
  assign y1460 = n4992 ;
  assign y1461 = n4995 ;
  assign y1462 = ~n4996 ;
  assign y1463 = n4999 ;
  assign y1464 = ~n5004 ;
  assign y1465 = ~1'b0 ;
  assign y1466 = ~1'b0 ;
  assign y1467 = ~n5005 ;
  assign y1468 = ~n5006 ;
  assign y1469 = ~n5010 ;
  assign y1470 = n5011 ;
  assign y1471 = n5020 ;
  assign y1472 = n5022 ;
  assign y1473 = n5024 ;
  assign y1474 = ~1'b0 ;
  assign y1475 = ~n5025 ;
  assign y1476 = ~n5035 ;
  assign y1477 = ~1'b0 ;
  assign y1478 = n5042 ;
  assign y1479 = n5051 ;
  assign y1480 = ~n5057 ;
  assign y1481 = n5058 ;
  assign y1482 = ~1'b0 ;
  assign y1483 = n5063 ;
  assign y1484 = ~1'b0 ;
  assign y1485 = n5069 ;
  assign y1486 = ~1'b0 ;
  assign y1487 = n5075 ;
  assign y1488 = ~1'b0 ;
  assign y1489 = ~n5077 ;
  assign y1490 = ~n5081 ;
  assign y1491 = ~n5088 ;
  assign y1492 = n5089 ;
  assign y1493 = n5091 ;
  assign y1494 = n5096 ;
  assign y1495 = ~n5099 ;
  assign y1496 = n5103 ;
  assign y1497 = n5112 ;
  assign y1498 = ~n5115 ;
  assign y1499 = ~1'b0 ;
  assign y1500 = ~n5117 ;
  assign y1501 = ~n5123 ;
  assign y1502 = n5124 ;
  assign y1503 = ~n5128 ;
  assign y1504 = ~1'b0 ;
  assign y1505 = ~n5129 ;
  assign y1506 = ~n5133 ;
  assign y1507 = ~n5142 ;
  assign y1508 = ~n5143 ;
  assign y1509 = n5144 ;
  assign y1510 = ~1'b0 ;
  assign y1511 = ~n5148 ;
  assign y1512 = ~n5152 ;
  assign y1513 = ~n5154 ;
  assign y1514 = ~1'b0 ;
  assign y1515 = ~n5163 ;
  assign y1516 = n5165 ;
  assign y1517 = n5166 ;
  assign y1518 = n5172 ;
  assign y1519 = n5174 ;
  assign y1520 = ~n5176 ;
  assign y1521 = ~n5182 ;
  assign y1522 = n5196 ;
  assign y1523 = ~1'b0 ;
  assign y1524 = ~n5200 ;
  assign y1525 = ~n5201 ;
  assign y1526 = ~1'b0 ;
  assign y1527 = n5202 ;
  assign y1528 = ~n5203 ;
  assign y1529 = n5210 ;
  assign y1530 = n5212 ;
  assign y1531 = n5213 ;
  assign y1532 = ~n5215 ;
  assign y1533 = n5216 ;
  assign y1534 = ~n5221 ;
  assign y1535 = ~n5227 ;
  assign y1536 = ~n5233 ;
  assign y1537 = ~n5237 ;
  assign y1538 = ~n5240 ;
  assign y1539 = n5245 ;
  assign y1540 = n5251 ;
  assign y1541 = ~1'b0 ;
  assign y1542 = n5255 ;
  assign y1543 = n5256 ;
  assign y1544 = n5263 ;
  assign y1545 = n5268 ;
  assign y1546 = ~n5271 ;
  assign y1547 = n5275 ;
  assign y1548 = ~n5276 ;
  assign y1549 = ~n5280 ;
  assign y1550 = ~1'b0 ;
  assign y1551 = ~n5284 ;
  assign y1552 = n5286 ;
  assign y1553 = ~n5290 ;
  assign y1554 = n5295 ;
  assign y1555 = n5297 ;
  assign y1556 = ~1'b0 ;
  assign y1557 = n5300 ;
  assign y1558 = n5312 ;
  assign y1559 = ~1'b0 ;
  assign y1560 = n5313 ;
  assign y1561 = ~n5320 ;
  assign y1562 = ~n5326 ;
  assign y1563 = ~1'b0 ;
  assign y1564 = n5329 ;
  assign y1565 = n5331 ;
  assign y1566 = ~1'b0 ;
  assign y1567 = ~n5338 ;
  assign y1568 = n5343 ;
  assign y1569 = ~n5345 ;
  assign y1570 = ~n5354 ;
  assign y1571 = n5355 ;
  assign y1572 = ~1'b0 ;
  assign y1573 = n5362 ;
  assign y1574 = n5366 ;
  assign y1575 = ~n5369 ;
  assign y1576 = n2539 ;
  assign y1577 = ~n5376 ;
  assign y1578 = ~n5379 ;
  assign y1579 = ~1'b0 ;
  assign y1580 = ~n5381 ;
  assign y1581 = n5384 ;
  assign y1582 = ~1'b0 ;
  assign y1583 = n5388 ;
  assign y1584 = n291 ;
  assign y1585 = ~n5394 ;
  assign y1586 = n5405 ;
  assign y1587 = n5410 ;
  assign y1588 = ~1'b0 ;
  assign y1589 = n5412 ;
  assign y1590 = n5416 ;
  assign y1591 = ~n5417 ;
  assign y1592 = ~1'b0 ;
  assign y1593 = ~n5427 ;
  assign y1594 = ~n5429 ;
  assign y1595 = ~n5446 ;
  assign y1596 = ~n5447 ;
  assign y1597 = ~n5451 ;
  assign y1598 = n5461 ;
  assign y1599 = ~n5466 ;
  assign y1600 = n5472 ;
  assign y1601 = n5475 ;
  assign y1602 = ~n5479 ;
  assign y1603 = ~n5486 ;
  assign y1604 = n5490 ;
  assign y1605 = ~1'b0 ;
  assign y1606 = ~1'b0 ;
  assign y1607 = ~n5492 ;
  assign y1608 = ~1'b0 ;
  assign y1609 = n5498 ;
  assign y1610 = ~1'b0 ;
  assign y1611 = n5503 ;
  assign y1612 = n5506 ;
  assign y1613 = ~1'b0 ;
  assign y1614 = n5508 ;
  assign y1615 = n5509 ;
  assign y1616 = ~n5510 ;
  assign y1617 = ~n5511 ;
  assign y1618 = ~n5513 ;
  assign y1619 = ~n5516 ;
  assign y1620 = ~n5526 ;
  assign y1621 = ~n5538 ;
  assign y1622 = 1'b0 ;
  assign y1623 = n5541 ;
  assign y1624 = n5545 ;
  assign y1625 = n5546 ;
  assign y1626 = n5554 ;
  assign y1627 = n5559 ;
  assign y1628 = ~n5560 ;
  assign y1629 = ~n5561 ;
  assign y1630 = ~n5562 ;
  assign y1631 = ~n5579 ;
  assign y1632 = ~n5580 ;
  assign y1633 = ~1'b0 ;
  assign y1634 = ~n5585 ;
  assign y1635 = n5586 ;
  assign y1636 = ~n5587 ;
  assign y1637 = ~1'b0 ;
  assign y1638 = ~n5600 ;
  assign y1639 = ~n5604 ;
  assign y1640 = n5605 ;
  assign y1641 = n5608 ;
  assign y1642 = n5612 ;
  assign y1643 = ~1'b0 ;
  assign y1644 = ~1'b0 ;
  assign y1645 = ~n5623 ;
  assign y1646 = ~n5625 ;
  assign y1647 = n5626 ;
  assign y1648 = ~n5633 ;
  assign y1649 = n5635 ;
  assign y1650 = ~1'b0 ;
  assign y1651 = n5640 ;
  assign y1652 = n5645 ;
  assign y1653 = n5654 ;
  assign y1654 = n5657 ;
  assign y1655 = ~n5660 ;
  assign y1656 = ~n5663 ;
  assign y1657 = ~n5675 ;
  assign y1658 = ~1'b0 ;
  assign y1659 = n5676 ;
  assign y1660 = ~n5683 ;
  assign y1661 = n5685 ;
  assign y1662 = n5687 ;
  assign y1663 = ~n5691 ;
  assign y1664 = ~n5692 ;
  assign y1665 = n5694 ;
  assign y1666 = ~n5701 ;
  assign y1667 = n5705 ;
  assign y1668 = n4285 ;
  assign y1669 = n5706 ;
  assign y1670 = ~n5708 ;
  assign y1671 = ~1'b0 ;
  assign y1672 = ~1'b0 ;
  assign y1673 = n5709 ;
  assign y1674 = ~n5711 ;
  assign y1675 = ~n5715 ;
  assign y1676 = ~n5716 ;
  assign y1677 = ~n4022 ;
  assign y1678 = n5720 ;
  assign y1679 = ~n5724 ;
  assign y1680 = n5730 ;
  assign y1681 = n5732 ;
  assign y1682 = n5734 ;
  assign y1683 = n5735 ;
  assign y1684 = ~n5738 ;
  assign y1685 = n5743 ;
  assign y1686 = ~1'b0 ;
  assign y1687 = ~n5746 ;
  assign y1688 = n5751 ;
  assign y1689 = ~n5769 ;
  assign y1690 = ~1'b0 ;
  assign y1691 = ~1'b0 ;
  assign y1692 = n5772 ;
  assign y1693 = ~n5778 ;
  assign y1694 = ~n5780 ;
  assign y1695 = ~n3734 ;
  assign y1696 = n5784 ;
  assign y1697 = ~n5789 ;
  assign y1698 = ~1'b0 ;
  assign y1699 = ~n5793 ;
  assign y1700 = ~n5802 ;
  assign y1701 = n5803 ;
  assign y1702 = n5804 ;
  assign y1703 = ~1'b0 ;
  assign y1704 = ~n5807 ;
  assign y1705 = ~n5808 ;
  assign y1706 = ~n5812 ;
  assign y1707 = ~n5814 ;
  assign y1708 = n5817 ;
  assign y1709 = ~n5818 ;
  assign y1710 = n2413 ;
  assign y1711 = ~n5821 ;
  assign y1712 = ~n5823 ;
  assign y1713 = n5826 ;
  assign y1714 = n5827 ;
  assign y1715 = ~n5829 ;
  assign y1716 = ~1'b0 ;
  assign y1717 = ~n5833 ;
  assign y1718 = n4185 ;
  assign y1719 = ~n5837 ;
  assign y1720 = n5846 ;
  assign y1721 = ~n5851 ;
  assign y1722 = ~n5855 ;
  assign y1723 = ~n5863 ;
  assign y1724 = n5864 ;
  assign y1725 = n5867 ;
  assign y1726 = n5868 ;
  assign y1727 = ~n5872 ;
  assign y1728 = ~1'b0 ;
  assign y1729 = n5875 ;
  assign y1730 = n5881 ;
  assign y1731 = ~n5883 ;
  assign y1732 = ~n5887 ;
  assign y1733 = ~1'b0 ;
  assign y1734 = n5896 ;
  assign y1735 = ~1'b0 ;
  assign y1736 = ~n5900 ;
  assign y1737 = ~n5911 ;
  assign y1738 = ~n5913 ;
  assign y1739 = n5917 ;
  assign y1740 = n5925 ;
  assign y1741 = ~1'b0 ;
  assign y1742 = n5933 ;
  assign y1743 = ~1'b0 ;
  assign y1744 = n5936 ;
  assign y1745 = n5937 ;
  assign y1746 = n5938 ;
  assign y1747 = ~1'b0 ;
  assign y1748 = n752 ;
  assign y1749 = n5939 ;
  assign y1750 = n5949 ;
  assign y1751 = ~n5951 ;
  assign y1752 = n5953 ;
  assign y1753 = ~n5954 ;
  assign y1754 = ~1'b0 ;
  assign y1755 = n5955 ;
  assign y1756 = n5956 ;
  assign y1757 = n5958 ;
  assign y1758 = ~1'b0 ;
  assign y1759 = n5960 ;
  assign y1760 = n5963 ;
  assign y1761 = n5970 ;
  assign y1762 = n5971 ;
  assign y1763 = n5973 ;
  assign y1764 = n5976 ;
  assign y1765 = n5977 ;
  assign y1766 = n5988 ;
  assign y1767 = ~n5990 ;
  assign y1768 = ~1'b0 ;
  assign y1769 = n5992 ;
  assign y1770 = n5999 ;
  assign y1771 = n6003 ;
  assign y1772 = n6004 ;
  assign y1773 = n6005 ;
  assign y1774 = ~n6014 ;
  assign y1775 = ~n6022 ;
  assign y1776 = ~n6023 ;
  assign y1777 = ~1'b0 ;
  assign y1778 = ~n6026 ;
  assign y1779 = ~1'b0 ;
  assign y1780 = ~n6029 ;
  assign y1781 = n6035 ;
  assign y1782 = ~n6036 ;
  assign y1783 = ~1'b0 ;
  assign y1784 = n6040 ;
  assign y1785 = ~n6043 ;
  assign y1786 = ~n6062 ;
  assign y1787 = ~1'b0 ;
  assign y1788 = n6078 ;
  assign y1789 = n6080 ;
  assign y1790 = 1'b0 ;
  assign y1791 = ~n6088 ;
  assign y1792 = ~1'b0 ;
  assign y1793 = ~n6091 ;
  assign y1794 = ~n6102 ;
  assign y1795 = ~n6112 ;
  assign y1796 = ~n6116 ;
  assign y1797 = ~n6121 ;
  assign y1798 = n6126 ;
  assign y1799 = ~n696 ;
  assign y1800 = n6127 ;
  assign y1801 = ~n6128 ;
  assign y1802 = ~n6134 ;
  assign y1803 = n6135 ;
  assign y1804 = ~n6142 ;
  assign y1805 = n6143 ;
  assign y1806 = ~n6145 ;
  assign y1807 = ~n6148 ;
  assign y1808 = ~n6153 ;
  assign y1809 = ~1'b0 ;
  assign y1810 = n6154 ;
  assign y1811 = n6158 ;
  assign y1812 = ~1'b0 ;
  assign y1813 = n6161 ;
  assign y1814 = n6167 ;
  assign y1815 = ~n6175 ;
  assign y1816 = ~n6182 ;
  assign y1817 = ~n6183 ;
  assign y1818 = ~n6187 ;
  assign y1819 = n6194 ;
  assign y1820 = ~n6199 ;
  assign y1821 = n6201 ;
  assign y1822 = n6202 ;
  assign y1823 = n6203 ;
  assign y1824 = ~1'b0 ;
  assign y1825 = ~1'b0 ;
  assign y1826 = ~1'b0 ;
  assign y1827 = ~n6204 ;
  assign y1828 = ~n6207 ;
  assign y1829 = ~1'b0 ;
  assign y1830 = n6208 ;
  assign y1831 = n6209 ;
  assign y1832 = ~1'b0 ;
  assign y1833 = n6212 ;
  assign y1834 = n6215 ;
  assign y1835 = ~n6217 ;
  assign y1836 = ~n6223 ;
  assign y1837 = ~1'b0 ;
  assign y1838 = ~1'b0 ;
  assign y1839 = ~n6227 ;
  assign y1840 = ~1'b0 ;
  assign y1841 = ~n6229 ;
  assign y1842 = n6230 ;
  assign y1843 = n6231 ;
  assign y1844 = ~n6232 ;
  assign y1845 = ~n6235 ;
  assign y1846 = n6240 ;
  assign y1847 = ~n6244 ;
  assign y1848 = ~1'b0 ;
  assign y1849 = n6245 ;
  assign y1850 = ~n6252 ;
  assign y1851 = n6260 ;
  assign y1852 = ~n6267 ;
  assign y1853 = ~n4133 ;
  assign y1854 = n6268 ;
  assign y1855 = 1'b0 ;
  assign y1856 = n6275 ;
  assign y1857 = n6277 ;
  assign y1858 = ~1'b0 ;
  assign y1859 = ~n6280 ;
  assign y1860 = ~n6284 ;
  assign y1861 = ~n6286 ;
  assign y1862 = ~n6289 ;
  assign y1863 = n6290 ;
  assign y1864 = ~n6303 ;
  assign y1865 = ~n6315 ;
  assign y1866 = ~n6320 ;
  assign y1867 = n6321 ;
  assign y1868 = n6326 ;
  assign y1869 = n6334 ;
  assign y1870 = n6337 ;
  assign y1871 = ~1'b0 ;
  assign y1872 = ~n6341 ;
  assign y1873 = n6342 ;
  assign y1874 = ~n6345 ;
  assign y1875 = n6350 ;
  assign y1876 = ~1'b0 ;
  assign y1877 = n6354 ;
  assign y1878 = ~1'b0 ;
  assign y1879 = ~n6357 ;
  assign y1880 = n6359 ;
  assign y1881 = ~n6360 ;
  assign y1882 = ~n6362 ;
  assign y1883 = ~n6373 ;
  assign y1884 = ~n6380 ;
  assign y1885 = ~1'b0 ;
  assign y1886 = ~n6396 ;
  assign y1887 = ~n6399 ;
  assign y1888 = ~n6401 ;
  assign y1889 = n6408 ;
  assign y1890 = n6412 ;
  assign y1891 = ~n6415 ;
  assign y1892 = ~n6417 ;
  assign y1893 = ~1'b0 ;
  assign y1894 = ~1'b0 ;
  assign y1895 = ~n6418 ;
  assign y1896 = ~n6419 ;
  assign y1897 = ~1'b0 ;
  assign y1898 = n6420 ;
  assign y1899 = ~1'b0 ;
  assign y1900 = n6422 ;
  assign y1901 = ~n4320 ;
  assign y1902 = ~1'b0 ;
  assign y1903 = ~1'b0 ;
  assign y1904 = n6425 ;
  assign y1905 = ~n6428 ;
  assign y1906 = ~n6433 ;
  assign y1907 = ~n6437 ;
  assign y1908 = ~n6438 ;
  assign y1909 = n6439 ;
  assign y1910 = n6442 ;
  assign y1911 = ~n6445 ;
  assign y1912 = n6447 ;
  assign y1913 = ~n6451 ;
  assign y1914 = ~n6453 ;
  assign y1915 = ~n6459 ;
  assign y1916 = ~n6462 ;
  assign y1917 = ~n6463 ;
  assign y1918 = n6472 ;
  assign y1919 = n6483 ;
  assign y1920 = n6488 ;
  assign y1921 = ~n6496 ;
  assign y1922 = ~n6501 ;
  assign y1923 = n6508 ;
  assign y1924 = ~n6510 ;
  assign y1925 = ~n6518 ;
  assign y1926 = ~n6519 ;
  assign y1927 = ~n6520 ;
  assign y1928 = n6523 ;
  assign y1929 = n6525 ;
  assign y1930 = n6533 ;
  assign y1931 = ~1'b0 ;
  assign y1932 = n6535 ;
  assign y1933 = ~1'b0 ;
  assign y1934 = ~1'b0 ;
  assign y1935 = n6542 ;
  assign y1936 = n6549 ;
  assign y1937 = ~n6564 ;
  assign y1938 = n6568 ;
  assign y1939 = ~1'b0 ;
  assign y1940 = ~1'b0 ;
  assign y1941 = n6569 ;
  assign y1942 = n6571 ;
  assign y1943 = ~n6578 ;
  assign y1944 = ~n6580 ;
  assign y1945 = ~n6582 ;
  assign y1946 = ~n6587 ;
  assign y1947 = ~n6593 ;
  assign y1948 = ~n3575 ;
  assign y1949 = ~n6613 ;
  assign y1950 = n6614 ;
  assign y1951 = n6624 ;
  assign y1952 = n6625 ;
  assign y1953 = ~1'b0 ;
  assign y1954 = 1'b0 ;
  assign y1955 = n2897 ;
  assign y1956 = n6627 ;
  assign y1957 = n6629 ;
  assign y1958 = n6630 ;
  assign y1959 = n6632 ;
  assign y1960 = ~n6633 ;
  assign y1961 = n1934 ;
  assign y1962 = n6641 ;
  assign y1963 = ~n6647 ;
  assign y1964 = n6651 ;
  assign y1965 = n6653 ;
  assign y1966 = n6655 ;
  assign y1967 = ~n6657 ;
  assign y1968 = ~1'b0 ;
  assign y1969 = ~n6663 ;
  assign y1970 = ~n6666 ;
  assign y1971 = ~n6673 ;
  assign y1972 = ~1'b0 ;
  assign y1973 = n6674 ;
  assign y1974 = n6677 ;
  assign y1975 = ~1'b0 ;
  assign y1976 = ~1'b0 ;
  assign y1977 = ~n6679 ;
  assign y1978 = ~1'b0 ;
  assign y1979 = n6681 ;
  assign y1980 = ~n6685 ;
  assign y1981 = ~1'b0 ;
  assign y1982 = ~n6687 ;
  assign y1983 = n6689 ;
  assign y1984 = n6695 ;
  assign y1985 = ~n6702 ;
  assign y1986 = ~n6705 ;
  assign y1987 = n6706 ;
  assign y1988 = n6709 ;
  assign y1989 = ~n6717 ;
  assign y1990 = ~n6719 ;
  assign y1991 = ~1'b0 ;
  assign y1992 = ~n6721 ;
  assign y1993 = ~1'b0 ;
  assign y1994 = ~n6722 ;
  assign y1995 = ~1'b0 ;
  assign y1996 = ~n6723 ;
  assign y1997 = ~n6732 ;
  assign y1998 = ~n6733 ;
  assign y1999 = n6739 ;
  assign y2000 = ~1'b0 ;
  assign y2001 = n6742 ;
  assign y2002 = ~n6743 ;
  assign y2003 = n6744 ;
  assign y2004 = ~1'b0 ;
  assign y2005 = ~n6748 ;
  assign y2006 = ~n6749 ;
  assign y2007 = ~n6752 ;
  assign y2008 = n6758 ;
  assign y2009 = ~n6767 ;
  assign y2010 = ~n6769 ;
  assign y2011 = ~1'b0 ;
  assign y2012 = n6774 ;
  assign y2013 = ~n6784 ;
  assign y2014 = 1'b0 ;
  assign y2015 = ~n6789 ;
  assign y2016 = ~1'b0 ;
  assign y2017 = n6791 ;
  assign y2018 = ~n6802 ;
  assign y2019 = n6804 ;
  assign y2020 = n6808 ;
  assign y2021 = n6813 ;
  assign y2022 = n6815 ;
  assign y2023 = n6817 ;
  assign y2024 = ~n6825 ;
  assign y2025 = n6831 ;
  assign y2026 = ~n6834 ;
  assign y2027 = n6837 ;
  assign y2028 = n2730 ;
  assign y2029 = ~1'b0 ;
  assign y2030 = n6839 ;
  assign y2031 = ~n6842 ;
  assign y2032 = n6843 ;
  assign y2033 = ~n6849 ;
  assign y2034 = ~n6851 ;
  assign y2035 = ~n6861 ;
  assign y2036 = n6869 ;
  assign y2037 = n6870 ;
  assign y2038 = ~n6875 ;
  assign y2039 = n6882 ;
  assign y2040 = ~n6883 ;
  assign y2041 = ~n6888 ;
  assign y2042 = n6894 ;
  assign y2043 = n2242 ;
  assign y2044 = ~1'b0 ;
  assign y2045 = ~n6899 ;
  assign y2046 = ~n6902 ;
  assign y2047 = n6905 ;
  assign y2048 = n6906 ;
  assign y2049 = n6907 ;
  assign y2050 = n6908 ;
  assign y2051 = ~n6911 ;
  assign y2052 = n6912 ;
  assign y2053 = ~1'b0 ;
  assign y2054 = ~n6916 ;
  assign y2055 = ~n6919 ;
  assign y2056 = n6921 ;
  assign y2057 = ~n6922 ;
  assign y2058 = n6923 ;
  assign y2059 = n6924 ;
  assign y2060 = ~n6929 ;
  assign y2061 = n6930 ;
  assign y2062 = n6932 ;
  assign y2063 = n6937 ;
  assign y2064 = ~1'b0 ;
  assign y2065 = n6940 ;
  assign y2066 = n6943 ;
  assign y2067 = ~1'b0 ;
  assign y2068 = ~1'b0 ;
  assign y2069 = ~n6946 ;
  assign y2070 = ~n6947 ;
  assign y2071 = ~n6950 ;
  assign y2072 = n6952 ;
  assign y2073 = ~n6954 ;
  assign y2074 = ~n6955 ;
  assign y2075 = ~n6957 ;
  assign y2076 = ~n6962 ;
  assign y2077 = n6964 ;
  assign y2078 = ~n6966 ;
  assign y2079 = ~n6970 ;
  assign y2080 = ~1'b0 ;
  assign y2081 = ~n6971 ;
  assign y2082 = ~n6976 ;
  assign y2083 = n6977 ;
  assign y2084 = ~1'b0 ;
  assign y2085 = ~1'b0 ;
  assign y2086 = ~n6985 ;
  assign y2087 = ~n6986 ;
  assign y2088 = ~1'b0 ;
  assign y2089 = n6987 ;
  assign y2090 = ~1'b0 ;
  assign y2091 = n6991 ;
  assign y2092 = ~1'b0 ;
  assign y2093 = n6997 ;
  assign y2094 = n7008 ;
  assign y2095 = n7009 ;
  assign y2096 = n7011 ;
  assign y2097 = ~1'b0 ;
  assign y2098 = ~n7021 ;
  assign y2099 = ~n7031 ;
  assign y2100 = ~n7035 ;
  assign y2101 = ~n7036 ;
  assign y2102 = n7038 ;
  assign y2103 = ~n7041 ;
  assign y2104 = ~n1138 ;
  assign y2105 = n7044 ;
  assign y2106 = ~n7045 ;
  assign y2107 = n7051 ;
  assign y2108 = ~1'b0 ;
  assign y2109 = n7056 ;
  assign y2110 = ~n7057 ;
  assign y2111 = n7061 ;
  assign y2112 = n7066 ;
  assign y2113 = n7072 ;
  assign y2114 = ~n7075 ;
  assign y2115 = n7079 ;
  assign y2116 = ~n7083 ;
  assign y2117 = ~n7086 ;
  assign y2118 = n7088 ;
  assign y2119 = ~n7090 ;
  assign y2120 = ~n7091 ;
  assign y2121 = ~n7093 ;
  assign y2122 = ~n7095 ;
  assign y2123 = ~n7096 ;
  assign y2124 = ~1'b0 ;
  assign y2125 = ~n7099 ;
  assign y2126 = ~1'b0 ;
  assign y2127 = ~n7104 ;
  assign y2128 = ~1'b0 ;
  assign y2129 = ~n7109 ;
  assign y2130 = ~1'b0 ;
  assign y2131 = ~n7117 ;
  assign y2132 = n7118 ;
  assign y2133 = ~n7123 ;
  assign y2134 = ~n7124 ;
  assign y2135 = ~1'b0 ;
  assign y2136 = n7125 ;
  assign y2137 = ~n7128 ;
  assign y2138 = ~1'b0 ;
  assign y2139 = n7130 ;
  assign y2140 = ~n7135 ;
  assign y2141 = n7140 ;
  assign y2142 = ~n7150 ;
  assign y2143 = ~n7154 ;
  assign y2144 = ~1'b0 ;
  assign y2145 = n7158 ;
  assign y2146 = n7163 ;
  assign y2147 = ~n7165 ;
  assign y2148 = n7167 ;
  assign y2149 = ~n7168 ;
  assign y2150 = n7169 ;
  assign y2151 = ~n7177 ;
  assign y2152 = ~n7178 ;
  assign y2153 = ~n7182 ;
  assign y2154 = ~1'b0 ;
  assign y2155 = ~n7185 ;
  assign y2156 = n7191 ;
  assign y2157 = ~n7197 ;
  assign y2158 = ~1'b0 ;
  assign y2159 = ~n7201 ;
  assign y2160 = n7206 ;
  assign y2161 = ~n7211 ;
  assign y2162 = n7214 ;
  assign y2163 = n7215 ;
  assign y2164 = n7216 ;
  assign y2165 = 1'b0 ;
  assign y2166 = ~n7221 ;
  assign y2167 = n7223 ;
  assign y2168 = ~n7226 ;
  assign y2169 = ~1'b0 ;
  assign y2170 = n7229 ;
  assign y2171 = ~1'b0 ;
  assign y2172 = ~1'b0 ;
  assign y2173 = ~n7233 ;
  assign y2174 = n7238 ;
  assign y2175 = ~n7240 ;
  assign y2176 = n7246 ;
  assign y2177 = n7247 ;
  assign y2178 = ~n7249 ;
  assign y2179 = ~n7254 ;
  assign y2180 = n7257 ;
  assign y2181 = n7263 ;
  assign y2182 = ~n7265 ;
  assign y2183 = ~1'b0 ;
  assign y2184 = n7266 ;
  assign y2185 = ~n7268 ;
  assign y2186 = ~n7269 ;
  assign y2187 = ~1'b0 ;
  assign y2188 = ~n7273 ;
  assign y2189 = ~n7277 ;
  assign y2190 = ~n7279 ;
  assign y2191 = ~n7280 ;
  assign y2192 = ~1'b0 ;
  assign y2193 = n7282 ;
  assign y2194 = ~n7286 ;
  assign y2195 = ~n7287 ;
  assign y2196 = n7289 ;
  assign y2197 = ~n7291 ;
  assign y2198 = ~1'b0 ;
  assign y2199 = n7294 ;
  assign y2200 = ~n7301 ;
  assign y2201 = ~n7307 ;
  assign y2202 = n7309 ;
  assign y2203 = n7315 ;
  assign y2204 = n7320 ;
  assign y2205 = x113 ;
  assign y2206 = n7327 ;
  assign y2207 = ~1'b0 ;
  assign y2208 = n7328 ;
  assign y2209 = n7331 ;
  assign y2210 = ~n7333 ;
  assign y2211 = n7338 ;
  assign y2212 = ~n7343 ;
  assign y2213 = ~n7348 ;
  assign y2214 = n7351 ;
  assign y2215 = ~1'b0 ;
  assign y2216 = ~n7354 ;
  assign y2217 = n7361 ;
  assign y2218 = n7362 ;
  assign y2219 = n428 ;
  assign y2220 = ~1'b0 ;
  assign y2221 = ~n7364 ;
  assign y2222 = n7367 ;
  assign y2223 = n7372 ;
  assign y2224 = ~n7377 ;
  assign y2225 = n7382 ;
  assign y2226 = n7383 ;
  assign y2227 = ~n5154 ;
  assign y2228 = ~n7384 ;
  assign y2229 = ~1'b0 ;
  assign y2230 = ~n7387 ;
  assign y2231 = ~1'b0 ;
  assign y2232 = ~n7394 ;
  assign y2233 = n7396 ;
  assign y2234 = n7399 ;
  assign y2235 = n7403 ;
  assign y2236 = n7424 ;
  assign y2237 = ~n7429 ;
  assign y2238 = ~n7436 ;
  assign y2239 = n7437 ;
  assign y2240 = n7453 ;
  assign y2241 = ~n7458 ;
  assign y2242 = n7461 ;
  assign y2243 = ~1'b0 ;
  assign y2244 = ~1'b0 ;
  assign y2245 = n7464 ;
  assign y2246 = n7467 ;
  assign y2247 = n7468 ;
  assign y2248 = ~n7470 ;
  assign y2249 = n7471 ;
  assign y2250 = n7475 ;
  assign y2251 = ~1'b0 ;
  assign y2252 = ~n7476 ;
  assign y2253 = n7478 ;
  assign y2254 = ~n1080 ;
  assign y2255 = ~n7490 ;
  assign y2256 = n7497 ;
  assign y2257 = ~1'b0 ;
  assign y2258 = ~n7498 ;
  assign y2259 = n7506 ;
  assign y2260 = n7515 ;
  assign y2261 = ~n7516 ;
  assign y2262 = ~1'b0 ;
  assign y2263 = n7519 ;
  assign y2264 = ~n7521 ;
  assign y2265 = n7534 ;
  assign y2266 = n7543 ;
  assign y2267 = n7545 ;
  assign y2268 = ~n7561 ;
  assign y2269 = n7562 ;
  assign y2270 = ~1'b0 ;
  assign y2271 = ~n7563 ;
  assign y2272 = ~n7569 ;
  assign y2273 = ~n7576 ;
  assign y2274 = ~n7582 ;
  assign y2275 = n7585 ;
  assign y2276 = n7589 ;
  assign y2277 = ~n7591 ;
  assign y2278 = ~n7593 ;
  assign y2279 = n7595 ;
  assign y2280 = ~n7596 ;
  assign y2281 = ~1'b0 ;
  assign y2282 = n7599 ;
  assign y2283 = n7604 ;
  assign y2284 = n7605 ;
  assign y2285 = ~1'b0 ;
  assign y2286 = n7608 ;
  assign y2287 = n7612 ;
  assign y2288 = ~n7617 ;
  assign y2289 = n7619 ;
  assign y2290 = n7622 ;
  assign y2291 = ~1'b0 ;
  assign y2292 = n7628 ;
  assign y2293 = n7630 ;
  assign y2294 = ~n7633 ;
  assign y2295 = ~n7634 ;
  assign y2296 = n7644 ;
  assign y2297 = n7652 ;
  assign y2298 = ~n7659 ;
  assign y2299 = n7664 ;
  assign y2300 = ~n7665 ;
  assign y2301 = n7671 ;
  assign y2302 = ~1'b0 ;
  assign y2303 = ~1'b0 ;
  assign y2304 = n7676 ;
  assign y2305 = ~n7679 ;
  assign y2306 = ~n7680 ;
  assign y2307 = ~n7683 ;
  assign y2308 = ~n7685 ;
  assign y2309 = ~n7689 ;
  assign y2310 = ~n7692 ;
  assign y2311 = ~n7693 ;
  assign y2312 = ~1'b0 ;
  assign y2313 = ~n7708 ;
  assign y2314 = ~n7711 ;
  assign y2315 = n7714 ;
  assign y2316 = n7722 ;
  assign y2317 = n7724 ;
  assign y2318 = ~n7725 ;
  assign y2319 = ~1'b0 ;
  assign y2320 = ~1'b0 ;
  assign y2321 = ~n7727 ;
  assign y2322 = n7734 ;
  assign y2323 = ~1'b0 ;
  assign y2324 = ~n7741 ;
  assign y2325 = ~1'b0 ;
  assign y2326 = ~n7744 ;
  assign y2327 = ~n7747 ;
  assign y2328 = ~n7751 ;
  assign y2329 = n7753 ;
  assign y2330 = n7760 ;
  assign y2331 = ~n7762 ;
  assign y2332 = ~n7765 ;
  assign y2333 = ~1'b0 ;
  assign y2334 = n7766 ;
  assign y2335 = n7769 ;
  assign y2336 = ~1'b0 ;
  assign y2337 = ~1'b0 ;
  assign y2338 = ~n7773 ;
  assign y2339 = ~n7784 ;
  assign y2340 = ~1'b0 ;
  assign y2341 = ~n7790 ;
  assign y2342 = ~n7801 ;
  assign y2343 = ~n7804 ;
  assign y2344 = n7805 ;
  assign y2345 = n7807 ;
  assign y2346 = n7815 ;
  assign y2347 = ~1'b0 ;
  assign y2348 = ~n7817 ;
  assign y2349 = n7819 ;
  assign y2350 = n7820 ;
  assign y2351 = ~n7826 ;
  assign y2352 = n7836 ;
  assign y2353 = n7845 ;
  assign y2354 = n7846 ;
  assign y2355 = n7861 ;
  assign y2356 = ~n7864 ;
  assign y2357 = n7868 ;
  assign y2358 = n7871 ;
  assign y2359 = ~n7873 ;
  assign y2360 = n7879 ;
  assign y2361 = ~n7881 ;
  assign y2362 = n7886 ;
  assign y2363 = n7890 ;
  assign y2364 = n7898 ;
  assign y2365 = n7899 ;
  assign y2366 = n7900 ;
  assign y2367 = ~1'b0 ;
  assign y2368 = ~1'b0 ;
  assign y2369 = n7903 ;
  assign y2370 = ~1'b0 ;
  assign y2371 = ~n7908 ;
  assign y2372 = ~n7916 ;
  assign y2373 = ~n7919 ;
  assign y2374 = n7920 ;
  assign y2375 = n7924 ;
  assign y2376 = ~n7930 ;
  assign y2377 = ~n7933 ;
  assign y2378 = ~n7935 ;
  assign y2379 = n7938 ;
  assign y2380 = n7939 ;
  assign y2381 = ~n7946 ;
  assign y2382 = n7947 ;
  assign y2383 = ~n7957 ;
  assign y2384 = ~n7961 ;
  assign y2385 = n7963 ;
  assign y2386 = n7971 ;
  assign y2387 = ~n7976 ;
  assign y2388 = n7983 ;
  assign y2389 = ~n7984 ;
  assign y2390 = n7987 ;
  assign y2391 = ~n7997 ;
  assign y2392 = ~n7999 ;
  assign y2393 = n8000 ;
  assign y2394 = ~1'b0 ;
  assign y2395 = ~1'b0 ;
  assign y2396 = n8003 ;
  assign y2397 = ~1'b0 ;
  assign y2398 = ~n8004 ;
  assign y2399 = ~1'b0 ;
  assign y2400 = ~1'b0 ;
  assign y2401 = n8005 ;
  assign y2402 = n8009 ;
  assign y2403 = ~n7853 ;
  assign y2404 = n8011 ;
  assign y2405 = ~n8012 ;
  assign y2406 = n8014 ;
  assign y2407 = ~1'b0 ;
  assign y2408 = ~n7338 ;
  assign y2409 = ~n8015 ;
  assign y2410 = ~n8019 ;
  assign y2411 = ~1'b0 ;
  assign y2412 = ~n8022 ;
  assign y2413 = ~n8024 ;
  assign y2414 = ~n8025 ;
  assign y2415 = n8026 ;
  assign y2416 = n8040 ;
  assign y2417 = ~n8045 ;
  assign y2418 = ~n8046 ;
  assign y2419 = ~n8048 ;
  assign y2420 = ~n8052 ;
  assign y2421 = ~n8055 ;
  assign y2422 = ~1'b0 ;
  assign y2423 = ~1'b0 ;
  assign y2424 = ~n8056 ;
  assign y2425 = n8062 ;
  assign y2426 = ~n8064 ;
  assign y2427 = ~n8068 ;
  assign y2428 = ~n8083 ;
  assign y2429 = ~n8086 ;
  assign y2430 = n8088 ;
  assign y2431 = n8092 ;
  assign y2432 = ~n8095 ;
  assign y2433 = ~n8105 ;
  assign y2434 = ~n8110 ;
  assign y2435 = n8115 ;
  assign y2436 = ~1'b0 ;
  assign y2437 = ~n8123 ;
  assign y2438 = ~1'b0 ;
  assign y2439 = ~n8124 ;
  assign y2440 = ~n8128 ;
  assign y2441 = ~n8129 ;
  assign y2442 = ~n8132 ;
  assign y2443 = ~n8137 ;
  assign y2444 = ~1'b0 ;
  assign y2445 = ~1'b0 ;
  assign y2446 = ~n8140 ;
  assign y2447 = 1'b0 ;
  assign y2448 = n8145 ;
  assign y2449 = ~1'b0 ;
  assign y2450 = ~n8146 ;
  assign y2451 = n8149 ;
  assign y2452 = ~1'b0 ;
  assign y2453 = ~1'b0 ;
  assign y2454 = n8156 ;
  assign y2455 = ~1'b0 ;
  assign y2456 = n8157 ;
  assign y2457 = ~n8159 ;
  assign y2458 = ~1'b0 ;
  assign y2459 = ~n8160 ;
  assign y2460 = n8161 ;
  assign y2461 = ~n8168 ;
  assign y2462 = ~1'b0 ;
  assign y2463 = ~n8175 ;
  assign y2464 = n8177 ;
  assign y2465 = ~n8180 ;
  assign y2466 = ~n8181 ;
  assign y2467 = ~n8182 ;
  assign y2468 = ~n8183 ;
  assign y2469 = ~1'b0 ;
  assign y2470 = ~n8187 ;
  assign y2471 = ~n8191 ;
  assign y2472 = n8193 ;
  assign y2473 = ~n8201 ;
  assign y2474 = ~n8203 ;
  assign y2475 = n8207 ;
  assign y2476 = n8208 ;
  assign y2477 = n8210 ;
  assign y2478 = ~n8211 ;
  assign y2479 = n8216 ;
  assign y2480 = ~n8217 ;
  assign y2481 = n8219 ;
  assign y2482 = ~1'b0 ;
  assign y2483 = ~1'b0 ;
  assign y2484 = n8231 ;
  assign y2485 = n6275 ;
  assign y2486 = n8232 ;
  assign y2487 = ~1'b0 ;
  assign y2488 = ~n8233 ;
  assign y2489 = n8235 ;
  assign y2490 = ~1'b0 ;
  assign y2491 = ~n8237 ;
  assign y2492 = ~n8239 ;
  assign y2493 = n8242 ;
  assign y2494 = ~n8245 ;
  assign y2495 = ~n8247 ;
  assign y2496 = ~n8254 ;
  assign y2497 = ~n8261 ;
  assign y2498 = ~n8267 ;
  assign y2499 = n8269 ;
  assign y2500 = ~n8270 ;
  assign y2501 = ~n8271 ;
  assign y2502 = ~n8277 ;
  assign y2503 = n8284 ;
  assign y2504 = n8286 ;
  assign y2505 = ~1'b0 ;
  assign y2506 = ~1'b0 ;
  assign y2507 = ~n8291 ;
  assign y2508 = ~n8295 ;
  assign y2509 = ~n8302 ;
  assign y2510 = n8303 ;
  assign y2511 = ~n8306 ;
  assign y2512 = n8309 ;
  assign y2513 = ~1'b0 ;
  assign y2514 = ~n8312 ;
  assign y2515 = n8317 ;
  assign y2516 = ~1'b0 ;
  assign y2517 = 1'b0 ;
  assign y2518 = ~n8322 ;
  assign y2519 = ~n8327 ;
  assign y2520 = n8328 ;
  assign y2521 = n8330 ;
  assign y2522 = ~n8333 ;
  assign y2523 = ~1'b0 ;
  assign y2524 = n8337 ;
  assign y2525 = n8338 ;
  assign y2526 = n8339 ;
  assign y2527 = n8341 ;
  assign y2528 = n658 ;
  assign y2529 = ~n8342 ;
  assign y2530 = ~n8343 ;
  assign y2531 = ~n8344 ;
  assign y2532 = ~n8348 ;
  assign y2533 = n8349 ;
  assign y2534 = ~n8355 ;
  assign y2535 = ~1'b0 ;
  assign y2536 = ~n8357 ;
  assign y2537 = n8360 ;
  assign y2538 = n8362 ;
  assign y2539 = ~n8364 ;
  assign y2540 = ~n5890 ;
  assign y2541 = ~n8365 ;
  assign y2542 = ~n8369 ;
  assign y2543 = n8372 ;
  assign y2544 = ~n8377 ;
  assign y2545 = ~n8380 ;
  assign y2546 = ~n8383 ;
  assign y2547 = ~n8385 ;
  assign y2548 = ~n8388 ;
  assign y2549 = n8404 ;
  assign y2550 = ~n8405 ;
  assign y2551 = ~1'b0 ;
  assign y2552 = ~1'b0 ;
  assign y2553 = n8408 ;
  assign y2554 = ~n8412 ;
  assign y2555 = n8419 ;
  assign y2556 = ~n8421 ;
  assign y2557 = ~n8430 ;
  assign y2558 = ~n8431 ;
  assign y2559 = ~n8433 ;
  assign y2560 = n8434 ;
  assign y2561 = ~1'b0 ;
  assign y2562 = ~n8437 ;
  assign y2563 = n8438 ;
  assign y2564 = ~n8445 ;
  assign y2565 = n8453 ;
  assign y2566 = n8456 ;
  assign y2567 = n8458 ;
  assign y2568 = ~1'b0 ;
  assign y2569 = n8461 ;
  assign y2570 = ~1'b0 ;
  assign y2571 = n8462 ;
  assign y2572 = n8466 ;
  assign y2573 = ~1'b0 ;
  assign y2574 = ~n8472 ;
  assign y2575 = ~n8480 ;
  assign y2576 = ~1'b0 ;
  assign y2577 = n8483 ;
  assign y2578 = ~n8485 ;
  assign y2579 = ~1'b0 ;
  assign y2580 = ~n8489 ;
  assign y2581 = ~n8494 ;
  assign y2582 = ~n8495 ;
  assign y2583 = ~1'b0 ;
  assign y2584 = n8500 ;
  assign y2585 = n8501 ;
  assign y2586 = ~n8503 ;
  assign y2587 = n8507 ;
  assign y2588 = ~1'b0 ;
  assign y2589 = ~n8520 ;
  assign y2590 = ~n8521 ;
  assign y2591 = ~1'b0 ;
  assign y2592 = ~1'b0 ;
  assign y2593 = ~n8523 ;
  assign y2594 = ~n8527 ;
  assign y2595 = ~n8530 ;
  assign y2596 = ~1'b0 ;
  assign y2597 = n8532 ;
  assign y2598 = ~n8539 ;
  assign y2599 = ~n8543 ;
  assign y2600 = ~1'b0 ;
  assign y2601 = ~n8544 ;
  assign y2602 = ~n8550 ;
  assign y2603 = ~n8558 ;
  assign y2604 = n8565 ;
  assign y2605 = ~n8568 ;
  assign y2606 = ~n8570 ;
  assign y2607 = ~n8574 ;
  assign y2608 = n8575 ;
  assign y2609 = ~1'b0 ;
  assign y2610 = n8578 ;
  assign y2611 = ~n8581 ;
  assign y2612 = n8583 ;
  assign y2613 = ~n8587 ;
  assign y2614 = n8591 ;
  assign y2615 = ~n8593 ;
  assign y2616 = ~n8595 ;
  assign y2617 = ~1'b0 ;
  assign y2618 = ~n8598 ;
  assign y2619 = ~n8605 ;
  assign y2620 = n8608 ;
  assign y2621 = n8609 ;
  assign y2622 = ~n8610 ;
  assign y2623 = ~n8613 ;
  assign y2624 = ~n8618 ;
  assign y2625 = n8619 ;
  assign y2626 = 1'b0 ;
  assign y2627 = ~n8624 ;
  assign y2628 = ~n8644 ;
  assign y2629 = ~n8647 ;
  assign y2630 = n8648 ;
  assign y2631 = n8650 ;
  assign y2632 = ~1'b0 ;
  assign y2633 = ~n8654 ;
  assign y2634 = ~n8656 ;
  assign y2635 = ~n8657 ;
  assign y2636 = ~1'b0 ;
  assign y2637 = ~n8658 ;
  assign y2638 = ~1'b0 ;
  assign y2639 = n8665 ;
  assign y2640 = n8666 ;
  assign y2641 = n8667 ;
  assign y2642 = n8670 ;
  assign y2643 = ~n8673 ;
  assign y2644 = n8674 ;
  assign y2645 = n8680 ;
  assign y2646 = n8681 ;
  assign y2647 = ~1'b0 ;
  assign y2648 = ~1'b0 ;
  assign y2649 = n8682 ;
  assign y2650 = n7947 ;
  assign y2651 = ~1'b0 ;
  assign y2652 = ~1'b0 ;
  assign y2653 = ~1'b0 ;
  assign y2654 = ~1'b0 ;
  assign y2655 = n8688 ;
  assign y2656 = ~n8693 ;
  assign y2657 = ~1'b0 ;
  assign y2658 = n8704 ;
  assign y2659 = ~1'b0 ;
  assign y2660 = ~n8710 ;
  assign y2661 = n8716 ;
  assign y2662 = ~n8719 ;
  assign y2663 = n8720 ;
  assign y2664 = ~1'b0 ;
  assign y2665 = n8723 ;
  assign y2666 = n8726 ;
  assign y2667 = ~n8727 ;
  assign y2668 = n8734 ;
  assign y2669 = n8736 ;
  assign y2670 = n8750 ;
  assign y2671 = ~1'b0 ;
  assign y2672 = n8756 ;
  assign y2673 = ~n8758 ;
  assign y2674 = ~1'b0 ;
  assign y2675 = ~n8766 ;
  assign y2676 = ~n8767 ;
  assign y2677 = ~n8768 ;
  assign y2678 = ~n8770 ;
  assign y2679 = ~n8774 ;
  assign y2680 = ~n8776 ;
  assign y2681 = ~1'b0 ;
  assign y2682 = n8784 ;
  assign y2683 = ~n8786 ;
  assign y2684 = 1'b0 ;
  assign y2685 = ~n8789 ;
  assign y2686 = n8796 ;
  assign y2687 = ~n8798 ;
  assign y2688 = ~n8807 ;
  assign y2689 = n8808 ;
  assign y2690 = ~n8809 ;
  assign y2691 = n8810 ;
  assign y2692 = n8811 ;
  assign y2693 = ~n8814 ;
  assign y2694 = ~1'b0 ;
  assign y2695 = ~n8816 ;
  assign y2696 = n8818 ;
  assign y2697 = n8821 ;
  assign y2698 = n8826 ;
  assign y2699 = n8833 ;
  assign y2700 = n8837 ;
  assign y2701 = ~n8841 ;
  assign y2702 = ~1'b0 ;
  assign y2703 = ~1'b0 ;
  assign y2704 = ~n8843 ;
  assign y2705 = ~1'b0 ;
  assign y2706 = ~n8845 ;
  assign y2707 = ~n8846 ;
  assign y2708 = n8847 ;
  assign y2709 = ~n8849 ;
  assign y2710 = ~n8854 ;
  assign y2711 = ~1'b0 ;
  assign y2712 = ~n8855 ;
  assign y2713 = ~1'b0 ;
  assign y2714 = n8858 ;
  assign y2715 = ~n8861 ;
  assign y2716 = n8862 ;
  assign y2717 = ~n8863 ;
  assign y2718 = n8864 ;
  assign y2719 = ~1'b0 ;
  assign y2720 = ~1'b0 ;
  assign y2721 = n8868 ;
  assign y2722 = n8871 ;
  assign y2723 = ~n8873 ;
  assign y2724 = ~n8876 ;
  assign y2725 = ~n8879 ;
  assign y2726 = n8884 ;
  assign y2727 = ~1'b0 ;
  assign y2728 = ~n8890 ;
  assign y2729 = ~n8893 ;
  assign y2730 = ~n8894 ;
  assign y2731 = n8896 ;
  assign y2732 = ~1'b0 ;
  assign y2733 = ~n8898 ;
  assign y2734 = ~n8901 ;
  assign y2735 = n8903 ;
  assign y2736 = n8904 ;
  assign y2737 = ~n8905 ;
  assign y2738 = ~1'b0 ;
  assign y2739 = ~n8907 ;
  assign y2740 = n8909 ;
  assign y2741 = ~n8916 ;
  assign y2742 = ~n8919 ;
  assign y2743 = n8922 ;
  assign y2744 = ~n8925 ;
  assign y2745 = n8926 ;
  assign y2746 = ~n8929 ;
  assign y2747 = n8930 ;
  assign y2748 = n8932 ;
  assign y2749 = ~n8936 ;
  assign y2750 = n8938 ;
  assign y2751 = n8939 ;
  assign y2752 = n8941 ;
  assign y2753 = ~1'b0 ;
  assign y2754 = ~n8944 ;
  assign y2755 = ~n8948 ;
  assign y2756 = n8951 ;
  assign y2757 = n8955 ;
  assign y2758 = n8957 ;
  assign y2759 = ~1'b0 ;
  assign y2760 = ~1'b0 ;
  assign y2761 = ~n8959 ;
  assign y2762 = ~n3131 ;
  assign y2763 = ~1'b0 ;
  assign y2764 = ~1'b0 ;
  assign y2765 = ~n8961 ;
  assign y2766 = n8963 ;
  assign y2767 = ~n8964 ;
  assign y2768 = ~1'b0 ;
  assign y2769 = n8965 ;
  assign y2770 = n8966 ;
  assign y2771 = n8973 ;
  assign y2772 = n8979 ;
  assign y2773 = ~n8985 ;
  assign y2774 = n8999 ;
  assign y2775 = ~1'b0 ;
  assign y2776 = ~n9012 ;
  assign y2777 = ~n9017 ;
  assign y2778 = ~n9021 ;
  assign y2779 = ~n9025 ;
  assign y2780 = n7398 ;
  assign y2781 = ~1'b0 ;
  assign y2782 = ~n9030 ;
  assign y2783 = ~n9032 ;
  assign y2784 = ~n9033 ;
  assign y2785 = ~n9034 ;
  assign y2786 = ~1'b0 ;
  assign y2787 = n9040 ;
  assign y2788 = ~n9041 ;
  assign y2789 = ~n3602 ;
  assign y2790 = ~n9044 ;
  assign y2791 = ~n9049 ;
  assign y2792 = ~1'b0 ;
  assign y2793 = n9050 ;
  assign y2794 = n9052 ;
  assign y2795 = ~n9061 ;
  assign y2796 = n9062 ;
  assign y2797 = n9067 ;
  assign y2798 = ~n9069 ;
  assign y2799 = ~n9071 ;
  assign y2800 = ~n9074 ;
  assign y2801 = n9075 ;
  assign y2802 = ~n9077 ;
  assign y2803 = ~n9079 ;
  assign y2804 = 1'b0 ;
  assign y2805 = ~n9086 ;
  assign y2806 = ~n3272 ;
  assign y2807 = n9088 ;
  assign y2808 = ~n9093 ;
  assign y2809 = ~1'b0 ;
  assign y2810 = n9095 ;
  assign y2811 = n9097 ;
  assign y2812 = ~n9104 ;
  assign y2813 = n9105 ;
  assign y2814 = ~n9106 ;
  assign y2815 = ~n9107 ;
  assign y2816 = n9109 ;
  assign y2817 = n9110 ;
  assign y2818 = n9115 ;
  assign y2819 = n9117 ;
  assign y2820 = ~1'b0 ;
  assign y2821 = ~n9119 ;
  assign y2822 = 1'b0 ;
  assign y2823 = n9126 ;
  assign y2824 = n9135 ;
  assign y2825 = ~1'b0 ;
  assign y2826 = n9138 ;
  assign y2827 = n9141 ;
  assign y2828 = n9143 ;
  assign y2829 = ~n9144 ;
  assign y2830 = n9149 ;
  assign y2831 = n9154 ;
  assign y2832 = ~n9157 ;
  assign y2833 = n9159 ;
  assign y2834 = ~n9166 ;
  assign y2835 = ~1'b0 ;
  assign y2836 = n9168 ;
  assign y2837 = ~n9173 ;
  assign y2838 = ~n9176 ;
  assign y2839 = ~n9177 ;
  assign y2840 = n9178 ;
  assign y2841 = n9181 ;
  assign y2842 = ~n383 ;
  assign y2843 = n9189 ;
  assign y2844 = ~n9199 ;
  assign y2845 = n9200 ;
  assign y2846 = n9201 ;
  assign y2847 = ~n9203 ;
  assign y2848 = n9204 ;
  assign y2849 = ~1'b0 ;
  assign y2850 = n9205 ;
  assign y2851 = n9206 ;
  assign y2852 = n9207 ;
  assign y2853 = ~1'b0 ;
  assign y2854 = ~n9210 ;
  assign y2855 = n9211 ;
  assign y2856 = ~n9213 ;
  assign y2857 = ~n9215 ;
  assign y2858 = ~n9217 ;
  assign y2859 = ~n9224 ;
  assign y2860 = n9229 ;
  assign y2861 = ~1'b0 ;
  assign y2862 = n9230 ;
  assign y2863 = ~n9235 ;
  assign y2864 = ~n9237 ;
  assign y2865 = n9240 ;
  assign y2866 = n9241 ;
  assign y2867 = ~n9247 ;
  assign y2868 = n9250 ;
  assign y2869 = n9251 ;
  assign y2870 = ~n2227 ;
  assign y2871 = ~n9252 ;
  assign y2872 = n9257 ;
  assign y2873 = ~n9259 ;
  assign y2874 = ~n9260 ;
  assign y2875 = n9261 ;
  assign y2876 = ~n9267 ;
  assign y2877 = ~n9268 ;
  assign y2878 = ~n9271 ;
  assign y2879 = ~n9273 ;
  assign y2880 = n9275 ;
  assign y2881 = ~n9280 ;
  assign y2882 = ~n3858 ;
  assign y2883 = n9282 ;
  assign y2884 = ~1'b0 ;
  assign y2885 = ~n9283 ;
  assign y2886 = ~n9286 ;
  assign y2887 = n9287 ;
  assign y2888 = ~n9292 ;
  assign y2889 = n9294 ;
  assign y2890 = ~1'b0 ;
  assign y2891 = n9299 ;
  assign y2892 = ~n9300 ;
  assign y2893 = ~n9301 ;
  assign y2894 = ~n9302 ;
  assign y2895 = ~n9304 ;
  assign y2896 = ~n9305 ;
  assign y2897 = n9306 ;
  assign y2898 = ~n9309 ;
  assign y2899 = ~n9310 ;
  assign y2900 = n8340 ;
  assign y2901 = ~n9317 ;
  assign y2902 = ~n9321 ;
  assign y2903 = n3338 ;
  assign y2904 = n9323 ;
  assign y2905 = ~n9339 ;
  assign y2906 = ~n9344 ;
  assign y2907 = ~n9349 ;
  assign y2908 = ~n9355 ;
  assign y2909 = ~n9359 ;
  assign y2910 = ~1'b0 ;
  assign y2911 = ~n9360 ;
  assign y2912 = n9361 ;
  assign y2913 = ~1'b0 ;
  assign y2914 = ~n9362 ;
  assign y2915 = n9366 ;
  assign y2916 = ~n9377 ;
  assign y2917 = ~1'b0 ;
  assign y2918 = n9379 ;
  assign y2919 = ~n9381 ;
  assign y2920 = n9383 ;
  assign y2921 = n9385 ;
  assign y2922 = ~n9389 ;
  assign y2923 = ~1'b0 ;
  assign y2924 = n9397 ;
  assign y2925 = n7903 ;
  assign y2926 = n9400 ;
  assign y2927 = ~n9408 ;
  assign y2928 = ~1'b0 ;
  assign y2929 = n9411 ;
  assign y2930 = ~1'b0 ;
  assign y2931 = n9413 ;
  assign y2932 = ~n9414 ;
  assign y2933 = ~n9420 ;
  assign y2934 = ~n9421 ;
  assign y2935 = ~n9430 ;
  assign y2936 = n9431 ;
  assign y2937 = ~1'b0 ;
  assign y2938 = ~n9433 ;
  assign y2939 = ~n9436 ;
  assign y2940 = ~n9437 ;
  assign y2941 = n9441 ;
  assign y2942 = ~n9448 ;
  assign y2943 = 1'b0 ;
  assign y2944 = ~n9449 ;
  assign y2945 = ~n9450 ;
  assign y2946 = ~n9454 ;
  assign y2947 = ~n9455 ;
  assign y2948 = ~n9458 ;
  assign y2949 = ~1'b0 ;
  assign y2950 = n9460 ;
  assign y2951 = n9466 ;
  assign y2952 = ~1'b0 ;
  assign y2953 = n9469 ;
  assign y2954 = n9470 ;
  assign y2955 = ~n9479 ;
  assign y2956 = n9480 ;
  assign y2957 = ~n9484 ;
  assign y2958 = n9491 ;
  assign y2959 = ~1'b0 ;
  assign y2960 = n9493 ;
  assign y2961 = n9494 ;
  assign y2962 = n9500 ;
  assign y2963 = ~n9504 ;
  assign y2964 = ~n9513 ;
  assign y2965 = ~1'b0 ;
  assign y2966 = n9518 ;
  assign y2967 = n9520 ;
  assign y2968 = ~1'b0 ;
  assign y2969 = ~1'b0 ;
  assign y2970 = ~1'b0 ;
  assign y2971 = ~n9521 ;
  assign y2972 = ~1'b0 ;
  assign y2973 = ~n9524 ;
  assign y2974 = ~1'b0 ;
  assign y2975 = ~n9526 ;
  assign y2976 = ~n9544 ;
  assign y2977 = ~1'b0 ;
  assign y2978 = ~1'b0 ;
  assign y2979 = ~n9548 ;
  assign y2980 = ~n9550 ;
  assign y2981 = ~n9554 ;
  assign y2982 = n9559 ;
  assign y2983 = n9561 ;
  assign y2984 = n1922 ;
  assign y2985 = n9565 ;
  assign y2986 = n9566 ;
  assign y2987 = ~n9571 ;
  assign y2988 = ~n9577 ;
  assign y2989 = n9578 ;
  assign y2990 = n9582 ;
  assign y2991 = n9588 ;
  assign y2992 = ~1'b0 ;
  assign y2993 = ~n9589 ;
  assign y2994 = n9593 ;
  assign y2995 = n9603 ;
  assign y2996 = n9612 ;
  assign y2997 = ~1'b0 ;
  assign y2998 = n9614 ;
  assign y2999 = ~n9618 ;
  assign y3000 = ~n9624 ;
  assign y3001 = ~n9632 ;
  assign y3002 = ~n9634 ;
  assign y3003 = n9637 ;
  assign y3004 = ~n9638 ;
  assign y3005 = n9645 ;
  assign y3006 = ~n9648 ;
  assign y3007 = ~n9653 ;
  assign y3008 = ~n9666 ;
  assign y3009 = ~1'b0 ;
  assign y3010 = n9678 ;
  assign y3011 = n9681 ;
  assign y3012 = ~n9689 ;
  assign y3013 = ~n9696 ;
  assign y3014 = ~n9700 ;
  assign y3015 = n9705 ;
  assign y3016 = ~1'b0 ;
  assign y3017 = n9710 ;
  assign y3018 = ~1'b0 ;
  assign y3019 = ~n9711 ;
  assign y3020 = n9714 ;
  assign y3021 = ~n9723 ;
  assign y3022 = ~1'b0 ;
  assign y3023 = ~1'b0 ;
  assign y3024 = ~n9725 ;
  assign y3025 = ~n9734 ;
  assign y3026 = ~n9737 ;
  assign y3027 = n9739 ;
  assign y3028 = ~1'b0 ;
  assign y3029 = ~1'b0 ;
  assign y3030 = n9745 ;
  assign y3031 = ~n9754 ;
  assign y3032 = n9758 ;
  assign y3033 = ~1'b0 ;
  assign y3034 = n9764 ;
  assign y3035 = ~n9765 ;
  assign y3036 = ~n9768 ;
  assign y3037 = n9770 ;
  assign y3038 = ~1'b0 ;
  assign y3039 = n9771 ;
  assign y3040 = n9780 ;
  assign y3041 = n9781 ;
  assign y3042 = ~1'b0 ;
  assign y3043 = ~n9787 ;
  assign y3044 = n9790 ;
  assign y3045 = n9792 ;
  assign y3046 = ~1'b0 ;
  assign y3047 = ~n9793 ;
  assign y3048 = ~n9795 ;
  assign y3049 = n9797 ;
  assign y3050 = ~n9809 ;
  assign y3051 = ~n9810 ;
  assign y3052 = n9816 ;
  assign y3053 = n9822 ;
  assign y3054 = ~1'b0 ;
  assign y3055 = ~n9823 ;
  assign y3056 = ~n9826 ;
  assign y3057 = n9830 ;
  assign y3058 = ~1'b0 ;
  assign y3059 = ~1'b0 ;
  assign y3060 = ~n9834 ;
  assign y3061 = ~n9839 ;
  assign y3062 = ~n9843 ;
  assign y3063 = n9853 ;
  assign y3064 = 1'b0 ;
  assign y3065 = n9863 ;
  assign y3066 = ~n9865 ;
  assign y3067 = n9871 ;
  assign y3068 = n9875 ;
  assign y3069 = n209 ;
  assign y3070 = n9883 ;
  assign y3071 = ~n9884 ;
  assign y3072 = ~1'b0 ;
  assign y3073 = n9885 ;
  assign y3074 = ~n911 ;
  assign y3075 = ~1'b0 ;
  assign y3076 = n9888 ;
  assign y3077 = ~n9890 ;
  assign y3078 = n9892 ;
  assign y3079 = n9907 ;
  assign y3080 = ~n9912 ;
  assign y3081 = n9917 ;
  assign y3082 = n9923 ;
  assign y3083 = ~1'b0 ;
  assign y3084 = n9924 ;
  assign y3085 = ~n9929 ;
  assign y3086 = n9932 ;
  assign y3087 = n9940 ;
  assign y3088 = ~1'b0 ;
  assign y3089 = ~n9942 ;
  assign y3090 = ~n9943 ;
  assign y3091 = ~n9948 ;
  assign y3092 = ~1'b0 ;
  assign y3093 = ~n9956 ;
  assign y3094 = n9959 ;
  assign y3095 = n9964 ;
  assign y3096 = ~n9966 ;
  assign y3097 = ~n9968 ;
  assign y3098 = ~n9969 ;
  assign y3099 = n9970 ;
  assign y3100 = n9979 ;
  assign y3101 = n9982 ;
  assign y3102 = n9985 ;
  assign y3103 = ~n9987 ;
  assign y3104 = n9989 ;
  assign y3105 = ~n9994 ;
  assign y3106 = n9995 ;
  assign y3107 = ~1'b0 ;
  assign y3108 = ~n9996 ;
  assign y3109 = n9998 ;
  assign y3110 = ~n10002 ;
  assign y3111 = ~n10005 ;
  assign y3112 = ~n10013 ;
  assign y3113 = ~n10014 ;
  assign y3114 = ~n10031 ;
  assign y3115 = ~n10032 ;
  assign y3116 = ~n10044 ;
  assign y3117 = 1'b0 ;
  assign y3118 = ~n10045 ;
  assign y3119 = n10050 ;
  assign y3120 = n10052 ;
  assign y3121 = ~n10064 ;
  assign y3122 = n10067 ;
  assign y3123 = ~n10071 ;
  assign y3124 = n10073 ;
  assign y3125 = 1'b0 ;
  assign y3126 = ~n7100 ;
  assign y3127 = ~n10075 ;
  assign y3128 = ~1'b0 ;
  assign y3129 = n10076 ;
  assign y3130 = ~n10077 ;
  assign y3131 = ~n10082 ;
  assign y3132 = ~n10090 ;
  assign y3133 = ~n10096 ;
  assign y3134 = n10100 ;
  assign y3135 = ~1'b0 ;
  assign y3136 = ~n10106 ;
  assign y3137 = n10112 ;
  assign y3138 = n10114 ;
  assign y3139 = ~n10117 ;
  assign y3140 = ~n10120 ;
  assign y3141 = n10124 ;
  assign y3142 = ~n10129 ;
  assign y3143 = n10130 ;
  assign y3144 = ~n10131 ;
  assign y3145 = n10132 ;
  assign y3146 = n10135 ;
  assign y3147 = n10136 ;
  assign y3148 = n10138 ;
  assign y3149 = ~n10139 ;
  assign y3150 = ~n10144 ;
  assign y3151 = n10145 ;
  assign y3152 = ~1'b0 ;
  assign y3153 = ~n10147 ;
  assign y3154 = ~1'b0 ;
  assign y3155 = ~1'b0 ;
  assign y3156 = ~n10150 ;
  assign y3157 = ~n10158 ;
  assign y3158 = ~n10164 ;
  assign y3159 = ~n10169 ;
  assign y3160 = n1289 ;
  assign y3161 = ~n10177 ;
  assign y3162 = ~n10178 ;
  assign y3163 = ~n10184 ;
  assign y3164 = ~n10185 ;
  assign y3165 = n10186 ;
  assign y3166 = ~n10189 ;
  assign y3167 = ~n10191 ;
  assign y3168 = ~1'b0 ;
  assign y3169 = ~1'b0 ;
  assign y3170 = n10197 ;
  assign y3171 = ~1'b0 ;
  assign y3172 = n10199 ;
  assign y3173 = ~n10203 ;
  assign y3174 = n10205 ;
  assign y3175 = n10207 ;
  assign y3176 = ~n10209 ;
  assign y3177 = ~1'b0 ;
  assign y3178 = ~n10213 ;
  assign y3179 = ~n10222 ;
  assign y3180 = n10227 ;
  assign y3181 = n10229 ;
  assign y3182 = n10230 ;
  assign y3183 = ~n10232 ;
  assign y3184 = n10236 ;
  assign y3185 = ~n2433 ;
  assign y3186 = ~1'b0 ;
  assign y3187 = ~n10237 ;
  assign y3188 = ~n10238 ;
  assign y3189 = n5284 ;
  assign y3190 = n10244 ;
  assign y3191 = ~n10251 ;
  assign y3192 = n10257 ;
  assign y3193 = ~1'b0 ;
  assign y3194 = n10265 ;
  assign y3195 = ~1'b0 ;
  assign y3196 = ~1'b0 ;
  assign y3197 = n10267 ;
  assign y3198 = ~1'b0 ;
  assign y3199 = ~n10269 ;
  assign y3200 = ~1'b0 ;
  assign y3201 = n10277 ;
  assign y3202 = n10278 ;
  assign y3203 = n10279 ;
  assign y3204 = ~n10280 ;
  assign y3205 = ~1'b0 ;
  assign y3206 = n10281 ;
  assign y3207 = n10282 ;
  assign y3208 = n10283 ;
  assign y3209 = ~n10284 ;
  assign y3210 = n10293 ;
  assign y3211 = n10300 ;
  assign y3212 = n10301 ;
  assign y3213 = ~n10302 ;
  assign y3214 = n10304 ;
  assign y3215 = n10313 ;
  assign y3216 = ~n10315 ;
  assign y3217 = n10316 ;
  assign y3218 = ~n10324 ;
  assign y3219 = ~n10326 ;
  assign y3220 = ~n10332 ;
  assign y3221 = n10333 ;
  assign y3222 = n10337 ;
  assign y3223 = ~n10339 ;
  assign y3224 = n10345 ;
  assign y3225 = ~n10352 ;
  assign y3226 = ~n10361 ;
  assign y3227 = ~n10362 ;
  assign y3228 = ~n10366 ;
  assign y3229 = ~n10378 ;
  assign y3230 = n10379 ;
  assign y3231 = ~n796 ;
  assign y3232 = ~1'b0 ;
  assign y3233 = n10390 ;
  assign y3234 = n10393 ;
  assign y3235 = ~n10396 ;
  assign y3236 = ~n10401 ;
  assign y3237 = ~1'b0 ;
  assign y3238 = ~n10402 ;
  assign y3239 = n10404 ;
  assign y3240 = n10405 ;
  assign y3241 = n10410 ;
  assign y3242 = n10413 ;
  assign y3243 = n10049 ;
  assign y3244 = ~n10416 ;
  assign y3245 = ~1'b0 ;
  assign y3246 = ~n10417 ;
  assign y3247 = n10424 ;
  assign y3248 = ~1'b0 ;
  assign y3249 = ~n10435 ;
  assign y3250 = n10436 ;
  assign y3251 = n10437 ;
  assign y3252 = ~n10442 ;
  assign y3253 = ~1'b0 ;
  assign y3254 = n10454 ;
  assign y3255 = n10457 ;
  assign y3256 = ~n10466 ;
  assign y3257 = n10471 ;
  assign y3258 = n10472 ;
  assign y3259 = ~1'b0 ;
  assign y3260 = n10476 ;
  assign y3261 = ~n10478 ;
  assign y3262 = ~n10483 ;
  assign y3263 = n10486 ;
  assign y3264 = ~1'b0 ;
  assign y3265 = ~n10495 ;
  assign y3266 = ~n10501 ;
  assign y3267 = 1'b0 ;
  assign y3268 = n10504 ;
  assign y3269 = n10512 ;
  assign y3270 = n10515 ;
  assign y3271 = ~n10521 ;
  assign y3272 = n10522 ;
  assign y3273 = n10523 ;
  assign y3274 = ~n10524 ;
  assign y3275 = ~1'b0 ;
  assign y3276 = n10525 ;
  assign y3277 = ~n10532 ;
  assign y3278 = n10542 ;
  assign y3279 = n10544 ;
  assign y3280 = n10548 ;
  assign y3281 = n10552 ;
  assign y3282 = n10553 ;
  assign y3283 = n10556 ;
  assign y3284 = ~n10560 ;
  assign y3285 = ~1'b0 ;
  assign y3286 = n10566 ;
  assign y3287 = n10567 ;
  assign y3288 = ~1'b0 ;
  assign y3289 = ~n10568 ;
  assign y3290 = ~n10569 ;
  assign y3291 = n10570 ;
  assign y3292 = ~1'b0 ;
  assign y3293 = ~n10572 ;
  assign y3294 = n10573 ;
  assign y3295 = n10577 ;
  assign y3296 = n10578 ;
  assign y3297 = ~n10582 ;
  assign y3298 = ~1'b0 ;
  assign y3299 = n10591 ;
  assign y3300 = ~n10594 ;
  assign y3301 = n10598 ;
  assign y3302 = n10604 ;
  assign y3303 = ~1'b0 ;
  assign y3304 = n10615 ;
  assign y3305 = ~n10617 ;
  assign y3306 = ~1'b0 ;
  assign y3307 = ~n10621 ;
  assign y3308 = n10631 ;
  assign y3309 = n10632 ;
  assign y3310 = n10635 ;
  assign y3311 = ~n10638 ;
  assign y3312 = ~n10641 ;
  assign y3313 = n10648 ;
  assign y3314 = ~n10651 ;
  assign y3315 = n10652 ;
  assign y3316 = ~n10655 ;
  assign y3317 = ~n10656 ;
  assign y3318 = ~n10501 ;
  assign y3319 = ~1'b0 ;
  assign y3320 = ~n10657 ;
  assign y3321 = n9827 ;
  assign y3322 = ~n10659 ;
  assign y3323 = ~n10660 ;
  assign y3324 = n10662 ;
  assign y3325 = n10664 ;
  assign y3326 = ~n10676 ;
  assign y3327 = ~n10679 ;
  assign y3328 = n10684 ;
  assign y3329 = n10685 ;
  assign y3330 = n10686 ;
  assign y3331 = ~1'b0 ;
  assign y3332 = ~n10690 ;
  assign y3333 = ~1'b0 ;
  assign y3334 = ~n10692 ;
  assign y3335 = n10695 ;
  assign y3336 = ~n5793 ;
  assign y3337 = ~n10696 ;
  assign y3338 = ~n10703 ;
  assign y3339 = n10709 ;
  assign y3340 = n2762 ;
  assign y3341 = ~n10710 ;
  assign y3342 = ~n10717 ;
  assign y3343 = n10718 ;
  assign y3344 = n10726 ;
  assign y3345 = ~n10727 ;
  assign y3346 = ~n10729 ;
  assign y3347 = ~n10733 ;
  assign y3348 = ~n10734 ;
  assign y3349 = ~1'b0 ;
  assign y3350 = n10736 ;
  assign y3351 = n10738 ;
  assign y3352 = n10740 ;
  assign y3353 = ~1'b0 ;
  assign y3354 = n10745 ;
  assign y3355 = n10746 ;
  assign y3356 = ~n10748 ;
  assign y3357 = ~n10750 ;
  assign y3358 = ~n10752 ;
  assign y3359 = n10753 ;
  assign y3360 = n10754 ;
  assign y3361 = n10757 ;
  assign y3362 = ~n10759 ;
  assign y3363 = ~1'b0 ;
  assign y3364 = ~1'b0 ;
  assign y3365 = ~n10774 ;
  assign y3366 = ~n10782 ;
  assign y3367 = ~1'b0 ;
  assign y3368 = n10784 ;
  assign y3369 = ~1'b0 ;
  assign y3370 = ~n7691 ;
  assign y3371 = n10791 ;
  assign y3372 = n10797 ;
  assign y3373 = ~n10798 ;
  assign y3374 = ~1'b0 ;
  assign y3375 = 1'b0 ;
  assign y3376 = ~n3377 ;
  assign y3377 = ~1'b0 ;
  assign y3378 = n10804 ;
  assign y3379 = n10809 ;
  assign y3380 = n10814 ;
  assign y3381 = ~1'b0 ;
  assign y3382 = n10816 ;
  assign y3383 = n10819 ;
  assign y3384 = n10820 ;
  assign y3385 = n10821 ;
  assign y3386 = n10828 ;
  assign y3387 = ~n10829 ;
  assign y3388 = n5450 ;
  assign y3389 = n10833 ;
  assign y3390 = ~n10835 ;
  assign y3391 = n10845 ;
  assign y3392 = ~n10847 ;
  assign y3393 = ~n10854 ;
  assign y3394 = ~n10855 ;
  assign y3395 = n10858 ;
  assign y3396 = n10864 ;
  assign y3397 = ~n10878 ;
  assign y3398 = ~n10882 ;
  assign y3399 = ~n10886 ;
  assign y3400 = ~n10888 ;
  assign y3401 = ~n10890 ;
  assign y3402 = n10891 ;
  assign y3403 = ~n10892 ;
  assign y3404 = n10893 ;
  assign y3405 = ~n9111 ;
  assign y3406 = ~n10894 ;
  assign y3407 = ~1'b0 ;
  assign y3408 = ~1'b0 ;
  assign y3409 = n10896 ;
  assign y3410 = ~n10903 ;
  assign y3411 = ~1'b0 ;
  assign y3412 = n10906 ;
  assign y3413 = ~n10909 ;
  assign y3414 = n10920 ;
  assign y3415 = ~n10921 ;
  assign y3416 = ~n10922 ;
  assign y3417 = n10924 ;
  assign y3418 = n10925 ;
  assign y3419 = ~n10930 ;
  assign y3420 = n10931 ;
  assign y3421 = n10936 ;
  assign y3422 = ~n10947 ;
  assign y3423 = ~n10948 ;
  assign y3424 = ~n10953 ;
  assign y3425 = ~n10960 ;
  assign y3426 = ~n10963 ;
  assign y3427 = ~n10965 ;
  assign y3428 = ~1'b0 ;
  assign y3429 = ~1'b0 ;
  assign y3430 = ~n10967 ;
  assign y3431 = n10968 ;
  assign y3432 = n10971 ;
  assign y3433 = n10973 ;
  assign y3434 = n10975 ;
  assign y3435 = ~n10978 ;
  assign y3436 = n10986 ;
  assign y3437 = ~1'b0 ;
  assign y3438 = ~1'b0 ;
  assign y3439 = ~n10987 ;
  assign y3440 = ~n10992 ;
  assign y3441 = n10999 ;
  assign y3442 = ~n11000 ;
  assign y3443 = n11002 ;
  assign y3444 = ~n11005 ;
  assign y3445 = ~n11006 ;
  assign y3446 = ~n11014 ;
  assign y3447 = ~1'b0 ;
  assign y3448 = ~n11016 ;
  assign y3449 = ~n11018 ;
  assign y3450 = ~n11019 ;
  assign y3451 = n11022 ;
  assign y3452 = n11036 ;
  assign y3453 = n11037 ;
  assign y3454 = n11042 ;
  assign y3455 = ~1'b0 ;
  assign y3456 = ~n11043 ;
  assign y3457 = ~n11044 ;
  assign y3458 = n11045 ;
  assign y3459 = ~n11046 ;
  assign y3460 = n11057 ;
  assign y3461 = ~1'b0 ;
  assign y3462 = ~n11060 ;
  assign y3463 = ~n11061 ;
  assign y3464 = ~1'b0 ;
  assign y3465 = ~n11064 ;
  assign y3466 = ~n11065 ;
  assign y3467 = n11073 ;
  assign y3468 = ~n11075 ;
  assign y3469 = ~1'b0 ;
  assign y3470 = ~n11077 ;
  assign y3471 = ~n11078 ;
  assign y3472 = n11079 ;
  assign y3473 = ~n11080 ;
  assign y3474 = n479 ;
  assign y3475 = n11088 ;
  assign y3476 = ~1'b0 ;
  assign y3477 = n11090 ;
  assign y3478 = n11096 ;
  assign y3479 = ~n11099 ;
  assign y3480 = ~n11102 ;
  assign y3481 = ~n11107 ;
  assign y3482 = ~1'b0 ;
  assign y3483 = ~n11110 ;
  assign y3484 = n3631 ;
  assign y3485 = n11118 ;
  assign y3486 = ~1'b0 ;
  assign y3487 = n11119 ;
  assign y3488 = ~n11122 ;
  assign y3489 = n11124 ;
  assign y3490 = ~n11125 ;
  assign y3491 = ~1'b0 ;
  assign y3492 = ~n1615 ;
  assign y3493 = ~n11126 ;
  assign y3494 = ~1'b0 ;
  assign y3495 = n11129 ;
  assign y3496 = ~n11130 ;
  assign y3497 = n3077 ;
  assign y3498 = n11133 ;
  assign y3499 = ~n9517 ;
  assign y3500 = 1'b0 ;
  assign y3501 = ~n11136 ;
  assign y3502 = n11142 ;
  assign y3503 = n11148 ;
  assign y3504 = n11153 ;
  assign y3505 = ~n11157 ;
  assign y3506 = ~n11162 ;
  assign y3507 = ~1'b0 ;
  assign y3508 = n4493 ;
  assign y3509 = ~n11170 ;
  assign y3510 = n11171 ;
  assign y3511 = ~n10000 ;
  assign y3512 = n11173 ;
  assign y3513 = ~n11179 ;
  assign y3514 = n11180 ;
  assign y3515 = n11182 ;
  assign y3516 = ~n11186 ;
  assign y3517 = n11189 ;
  assign y3518 = ~n11197 ;
  assign y3519 = ~n11201 ;
  assign y3520 = n11205 ;
  assign y3521 = ~n11207 ;
  assign y3522 = ~n11214 ;
  assign y3523 = n11216 ;
  assign y3524 = ~1'b0 ;
  assign y3525 = n11217 ;
  assign y3526 = ~n11221 ;
  assign y3527 = ~1'b0 ;
  assign y3528 = ~1'b0 ;
  assign y3529 = n11225 ;
  assign y3530 = ~n11227 ;
  assign y3531 = n11231 ;
  assign y3532 = ~n11232 ;
  assign y3533 = ~n11235 ;
  assign y3534 = ~n11237 ;
  assign y3535 = ~1'b0 ;
  assign y3536 = ~1'b0 ;
  assign y3537 = ~n11247 ;
  assign y3538 = n11251 ;
  assign y3539 = ~n11255 ;
  assign y3540 = ~n11260 ;
  assign y3541 = ~1'b0 ;
  assign y3542 = ~n11261 ;
  assign y3543 = 1'b0 ;
  assign y3544 = n11264 ;
  assign y3545 = ~n11265 ;
  assign y3546 = ~n11267 ;
  assign y3547 = n11268 ;
  assign y3548 = n11277 ;
  assign y3549 = ~n11278 ;
  assign y3550 = n11283 ;
  assign y3551 = ~1'b0 ;
  assign y3552 = ~n11284 ;
  assign y3553 = ~n11291 ;
  assign y3554 = ~n11295 ;
  assign y3555 = n11298 ;
  assign y3556 = ~n11301 ;
  assign y3557 = ~1'b0 ;
  assign y3558 = n11305 ;
  assign y3559 = ~1'b0 ;
  assign y3560 = ~n10700 ;
  assign y3561 = ~n11311 ;
  assign y3562 = n11316 ;
  assign y3563 = ~1'b0 ;
  assign y3564 = n11318 ;
  assign y3565 = n11322 ;
  assign y3566 = ~1'b0 ;
  assign y3567 = ~n11323 ;
  assign y3568 = n11327 ;
  assign y3569 = ~n11329 ;
  assign y3570 = ~n11330 ;
  assign y3571 = ~n11337 ;
  assign y3572 = ~1'b0 ;
  assign y3573 = n11344 ;
  assign y3574 = n11347 ;
  assign y3575 = ~n11350 ;
  assign y3576 = n11352 ;
  assign y3577 = ~1'b0 ;
  assign y3578 = ~n11358 ;
  assign y3579 = n11366 ;
  assign y3580 = n11375 ;
  assign y3581 = ~n11379 ;
  assign y3582 = ~1'b0 ;
  assign y3583 = ~1'b0 ;
  assign y3584 = ~n11389 ;
  assign y3585 = n11395 ;
  assign y3586 = ~n11402 ;
  assign y3587 = ~n11412 ;
  assign y3588 = n11413 ;
  assign y3589 = ~n11423 ;
  assign y3590 = ~1'b0 ;
  assign y3591 = n11425 ;
  assign y3592 = n11427 ;
  assign y3593 = n11435 ;
  assign y3594 = n11438 ;
  assign y3595 = ~1'b0 ;
  assign y3596 = ~1'b0 ;
  assign y3597 = n11445 ;
  assign y3598 = n11448 ;
  assign y3599 = n11450 ;
  assign y3600 = n11457 ;
  assign y3601 = ~n11460 ;
  assign y3602 = ~n11463 ;
  assign y3603 = n11465 ;
  assign y3604 = ~1'b0 ;
  assign y3605 = ~n11471 ;
  assign y3606 = ~1'b0 ;
  assign y3607 = ~n11475 ;
  assign y3608 = ~1'b0 ;
  assign y3609 = n11486 ;
  assign y3610 = ~n11497 ;
  assign y3611 = n11502 ;
  assign y3612 = ~n11504 ;
  assign y3613 = n11505 ;
  assign y3614 = ~1'b0 ;
  assign y3615 = ~n11506 ;
  assign y3616 = n11507 ;
  assign y3617 = n11509 ;
  assign y3618 = n11513 ;
  assign y3619 = ~n11514 ;
  assign y3620 = n11516 ;
  assign y3621 = ~1'b0 ;
  assign y3622 = n11523 ;
  assign y3623 = ~n11527 ;
  assign y3624 = ~n11531 ;
  assign y3625 = ~n11537 ;
  assign y3626 = ~n11542 ;
  assign y3627 = n11545 ;
  assign y3628 = n11549 ;
  assign y3629 = ~1'b0 ;
  assign y3630 = n8051 ;
  assign y3631 = ~n4115 ;
  assign y3632 = n11558 ;
  assign y3633 = ~1'b0 ;
  assign y3634 = n11560 ;
  assign y3635 = ~1'b0 ;
  assign y3636 = n11564 ;
  assign y3637 = n11565 ;
  assign y3638 = ~n11566 ;
  assign y3639 = ~n11568 ;
  assign y3640 = n11571 ;
  assign y3641 = n11573 ;
  assign y3642 = ~1'b0 ;
  assign y3643 = n11574 ;
  assign y3644 = ~1'b0 ;
  assign y3645 = ~1'b0 ;
  assign y3646 = n11575 ;
  assign y3647 = n11576 ;
  assign y3648 = n11579 ;
  assign y3649 = ~1'b0 ;
  assign y3650 = 1'b0 ;
  assign y3651 = ~1'b0 ;
  assign y3652 = ~1'b0 ;
  assign y3653 = n11580 ;
  assign y3654 = ~1'b0 ;
  assign y3655 = n11583 ;
  assign y3656 = ~n11593 ;
  assign y3657 = ~n2114 ;
  assign y3658 = ~n11598 ;
  assign y3659 = n11602 ;
  assign y3660 = ~1'b0 ;
  assign y3661 = ~n11603 ;
  assign y3662 = n6261 ;
  assign y3663 = ~1'b0 ;
  assign y3664 = ~n11609 ;
  assign y3665 = ~n11614 ;
  assign y3666 = n11617 ;
  assign y3667 = n11620 ;
  assign y3668 = n11623 ;
  assign y3669 = ~1'b0 ;
  assign y3670 = n11627 ;
  assign y3671 = n11629 ;
  assign y3672 = ~n11631 ;
  assign y3673 = n11634 ;
  assign y3674 = ~1'b0 ;
  assign y3675 = n11635 ;
  assign y3676 = ~n11636 ;
  assign y3677 = ~n11640 ;
  assign y3678 = ~n11642 ;
  assign y3679 = ~n11652 ;
  assign y3680 = ~n11655 ;
  assign y3681 = ~n11662 ;
  assign y3682 = ~1'b0 ;
  assign y3683 = n11663 ;
  assign y3684 = n11666 ;
  assign y3685 = ~n11667 ;
  assign y3686 = ~1'b0 ;
  assign y3687 = ~n11668 ;
  assign y3688 = n11669 ;
  assign y3689 = ~n11670 ;
  assign y3690 = n11673 ;
  assign y3691 = n11675 ;
  assign y3692 = ~n11676 ;
  assign y3693 = n11682 ;
  assign y3694 = ~1'b0 ;
  assign y3695 = ~n11684 ;
  assign y3696 = n11688 ;
  assign y3697 = n11697 ;
  assign y3698 = ~1'b0 ;
  assign y3699 = ~n11699 ;
  assign y3700 = ~n11702 ;
  assign y3701 = n11703 ;
  assign y3702 = n11707 ;
  assign y3703 = ~1'b0 ;
  assign y3704 = n11710 ;
  assign y3705 = ~n11711 ;
  assign y3706 = ~n11715 ;
  assign y3707 = n11716 ;
  assign y3708 = ~n11719 ;
  assign y3709 = ~n11724 ;
  assign y3710 = ~1'b0 ;
  assign y3711 = n11729 ;
  assign y3712 = ~n11732 ;
  assign y3713 = ~n11735 ;
  assign y3714 = ~n11743 ;
  assign y3715 = n11744 ;
  assign y3716 = n11746 ;
  assign y3717 = n11753 ;
  assign y3718 = ~n11764 ;
  assign y3719 = n11772 ;
  assign y3720 = n11773 ;
  assign y3721 = ~1'b0 ;
  assign y3722 = n11775 ;
  assign y3723 = ~n11778 ;
  assign y3724 = ~n11785 ;
  assign y3725 = n11788 ;
  assign y3726 = n11792 ;
  assign y3727 = n11796 ;
  assign y3728 = ~n11798 ;
  assign y3729 = ~n11803 ;
  assign y3730 = ~n11805 ;
  assign y3731 = n11806 ;
  assign y3732 = ~n11811 ;
  assign y3733 = ~n11813 ;
  assign y3734 = ~n5714 ;
  assign y3735 = ~n7279 ;
  assign y3736 = ~n11817 ;
  assign y3737 = n11821 ;
  assign y3738 = ~1'b0 ;
  assign y3739 = ~1'b0 ;
  assign y3740 = n11824 ;
  assign y3741 = n11825 ;
  assign y3742 = ~n11828 ;
  assign y3743 = ~1'b0 ;
  assign y3744 = n11832 ;
  assign y3745 = n11834 ;
  assign y3746 = ~n11839 ;
  assign y3747 = n11840 ;
  assign y3748 = ~n11848 ;
  assign y3749 = n11851 ;
  assign y3750 = ~1'b0 ;
  assign y3751 = n11856 ;
  assign y3752 = ~n11857 ;
  assign y3753 = ~1'b0 ;
  assign y3754 = n11862 ;
  assign y3755 = n11864 ;
  assign y3756 = n11865 ;
  assign y3757 = ~n11872 ;
  assign y3758 = n11873 ;
  assign y3759 = n11875 ;
  assign y3760 = n11883 ;
  assign y3761 = ~n11896 ;
  assign y3762 = ~1'b0 ;
  assign y3763 = n11897 ;
  assign y3764 = ~n11899 ;
  assign y3765 = n11901 ;
  assign y3766 = n11903 ;
  assign y3767 = ~n11904 ;
  assign y3768 = ~n11907 ;
  assign y3769 = n11910 ;
  assign y3770 = ~n11912 ;
  assign y3771 = ~1'b0 ;
  assign y3772 = ~1'b0 ;
  assign y3773 = ~n11916 ;
  assign y3774 = ~n11920 ;
  assign y3775 = ~n11923 ;
  assign y3776 = ~n11928 ;
  assign y3777 = n11930 ;
  assign y3778 = n11932 ;
  assign y3779 = ~n11940 ;
  assign y3780 = ~1'b0 ;
  assign y3781 = ~1'b0 ;
  assign y3782 = ~n11944 ;
  assign y3783 = n11945 ;
  assign y3784 = n11946 ;
  assign y3785 = ~n11948 ;
  assign y3786 = n11951 ;
  assign y3787 = n11952 ;
  assign y3788 = ~n11970 ;
  assign y3789 = n11976 ;
  assign y3790 = ~n11979 ;
  assign y3791 = n11987 ;
  assign y3792 = n11992 ;
  assign y3793 = n11994 ;
  assign y3794 = ~n11995 ;
  assign y3795 = ~n11999 ;
  assign y3796 = ~n12000 ;
  assign y3797 = n12003 ;
  assign y3798 = n12007 ;
  assign y3799 = ~n12011 ;
  assign y3800 = n11053 ;
  assign y3801 = ~n12014 ;
  assign y3802 = n12016 ;
  assign y3803 = ~n12020 ;
  assign y3804 = n11844 ;
  assign y3805 = n12023 ;
  assign y3806 = ~n12025 ;
  assign y3807 = n12027 ;
  assign y3808 = n12029 ;
  assign y3809 = ~n12031 ;
  assign y3810 = n12049 ;
  assign y3811 = ~1'b0 ;
  assign y3812 = ~1'b0 ;
  assign y3813 = ~1'b0 ;
  assign y3814 = n12051 ;
  assign y3815 = ~1'b0 ;
  assign y3816 = ~n12053 ;
  assign y3817 = n12061 ;
  assign y3818 = n12065 ;
  assign y3819 = ~n12067 ;
  assign y3820 = n12069 ;
  assign y3821 = ~n12072 ;
  assign y3822 = ~1'b0 ;
  assign y3823 = ~n9492 ;
  assign y3824 = n12075 ;
  assign y3825 = ~n12076 ;
  assign y3826 = ~n12078 ;
  assign y3827 = ~n12084 ;
  assign y3828 = n12086 ;
  assign y3829 = ~n12087 ;
  assign y3830 = n12091 ;
  assign y3831 = n12094 ;
  assign y3832 = ~n11115 ;
  assign y3833 = ~1'b0 ;
  assign y3834 = ~n12096 ;
  assign y3835 = n12100 ;
  assign y3836 = ~n12102 ;
  assign y3837 = ~1'b0 ;
  assign y3838 = n12103 ;
  assign y3839 = ~n12106 ;
  assign y3840 = ~n12113 ;
  assign y3841 = ~n12122 ;
  assign y3842 = ~n12127 ;
  assign y3843 = ~1'b0 ;
  assign y3844 = ~1'b0 ;
  assign y3845 = ~n12130 ;
  assign y3846 = n12138 ;
  assign y3847 = ~n12139 ;
  assign y3848 = n12141 ;
  assign y3849 = ~n12150 ;
  assign y3850 = ~n12153 ;
  assign y3851 = n12161 ;
  assign y3852 = ~n12163 ;
  assign y3853 = n12164 ;
  assign y3854 = ~n12165 ;
  assign y3855 = ~n12172 ;
  assign y3856 = ~1'b0 ;
  assign y3857 = n12174 ;
  assign y3858 = n12177 ;
  assign y3859 = n12179 ;
  assign y3860 = ~n12185 ;
  assign y3861 = ~n12186 ;
  assign y3862 = n12188 ;
  assign y3863 = n12190 ;
  assign y3864 = n12192 ;
  assign y3865 = n12196 ;
  assign y3866 = ~n12206 ;
  assign y3867 = n12210 ;
  assign y3868 = ~n12215 ;
  assign y3869 = ~1'b0 ;
  assign y3870 = ~n12220 ;
  assign y3871 = ~1'b0 ;
  assign y3872 = ~n5730 ;
  assign y3873 = ~n12221 ;
  assign y3874 = n12224 ;
  assign y3875 = n12228 ;
  assign y3876 = n12229 ;
  assign y3877 = n12231 ;
  assign y3878 = ~n12238 ;
  assign y3879 = n12241 ;
  assign y3880 = ~n12246 ;
  assign y3881 = n12257 ;
  assign y3882 = ~1'b0 ;
  assign y3883 = ~n12263 ;
  assign y3884 = ~n12265 ;
  assign y3885 = n12267 ;
  assign y3886 = n12279 ;
  assign y3887 = n12280 ;
  assign y3888 = ~n12282 ;
  assign y3889 = ~n12293 ;
  assign y3890 = ~n12294 ;
  assign y3891 = n12299 ;
  assign y3892 = ~n12300 ;
  assign y3893 = ~n12302 ;
  assign y3894 = n12312 ;
  assign y3895 = n12317 ;
  assign y3896 = n10304 ;
  assign y3897 = n12320 ;
  assign y3898 = ~n12322 ;
  assign y3899 = ~n12325 ;
  assign y3900 = ~n9544 ;
  assign y3901 = ~n12327 ;
  assign y3902 = n12338 ;
  assign y3903 = n12341 ;
  assign y3904 = ~1'b0 ;
  assign y3905 = ~n12342 ;
  assign y3906 = n12351 ;
  assign y3907 = n12353 ;
  assign y3908 = ~1'b0 ;
  assign y3909 = n12356 ;
  assign y3910 = ~n12365 ;
  assign y3911 = ~n12369 ;
  assign y3912 = ~n12378 ;
  assign y3913 = ~n12384 ;
  assign y3914 = n12387 ;
  assign y3915 = ~n12390 ;
  assign y3916 = ~n2422 ;
  assign y3917 = ~n12391 ;
  assign y3918 = n12393 ;
  assign y3919 = ~1'b0 ;
  assign y3920 = ~n12399 ;
  assign y3921 = ~n12400 ;
  assign y3922 = n12401 ;
  assign y3923 = ~n12407 ;
  assign y3924 = n12411 ;
  assign y3925 = ~1'b0 ;
  assign y3926 = n12412 ;
  assign y3927 = ~1'b0 ;
  assign y3928 = ~n12417 ;
  assign y3929 = n12421 ;
  assign y3930 = ~n12423 ;
  assign y3931 = ~n12424 ;
  assign y3932 = ~n12430 ;
  assign y3933 = n12435 ;
  assign y3934 = ~n12437 ;
  assign y3935 = n12438 ;
  assign y3936 = ~n12443 ;
  assign y3937 = n12444 ;
  assign y3938 = ~n12458 ;
  assign y3939 = ~n12462 ;
  assign y3940 = ~n12467 ;
  assign y3941 = 1'b0 ;
  assign y3942 = ~n12471 ;
  assign y3943 = n12478 ;
  assign y3944 = ~1'b0 ;
  assign y3945 = ~n12479 ;
  assign y3946 = n12482 ;
  assign y3947 = n12483 ;
  assign y3948 = ~n12485 ;
  assign y3949 = n12488 ;
  assign y3950 = ~n12502 ;
  assign y3951 = ~n12506 ;
  assign y3952 = ~n12507 ;
  assign y3953 = ~n12511 ;
  assign y3954 = ~n12517 ;
  assign y3955 = ~n5736 ;
  assign y3956 = ~1'b0 ;
  assign y3957 = ~1'b0 ;
  assign y3958 = ~1'b0 ;
  assign y3959 = ~n12519 ;
  assign y3960 = n12530 ;
  assign y3961 = n12533 ;
  assign y3962 = n1925 ;
  assign y3963 = n12538 ;
  assign y3964 = ~n12544 ;
  assign y3965 = ~n12546 ;
  assign y3966 = ~1'b0 ;
  assign y3967 = ~n12548 ;
  assign y3968 = n12552 ;
  assign y3969 = ~1'b0 ;
  assign y3970 = ~n12556 ;
  assign y3971 = ~1'b0 ;
  assign y3972 = ~n12557 ;
  assign y3973 = n10917 ;
  assign y3974 = n12561 ;
  assign y3975 = n12562 ;
  assign y3976 = ~n12568 ;
  assign y3977 = n12569 ;
  assign y3978 = ~n12571 ;
  assign y3979 = ~n12573 ;
  assign y3980 = n12574 ;
  assign y3981 = n12575 ;
  assign y3982 = n12580 ;
  assign y3983 = ~1'b0 ;
  assign y3984 = ~n12582 ;
  assign y3985 = ~1'b0 ;
  assign y3986 = ~n12586 ;
  assign y3987 = n12587 ;
  assign y3988 = ~n12592 ;
  assign y3989 = n12594 ;
  assign y3990 = ~n12600 ;
  assign y3991 = ~1'b0 ;
  assign y3992 = n1110 ;
  assign y3993 = n12602 ;
  assign y3994 = ~1'b0 ;
  assign y3995 = ~1'b0 ;
  assign y3996 = ~n12609 ;
  assign y3997 = n12613 ;
  assign y3998 = ~n12620 ;
  assign y3999 = ~n12624 ;
  assign y4000 = n12626 ;
  assign y4001 = ~n12627 ;
  assign y4002 = n12629 ;
  assign y4003 = ~1'b0 ;
  assign y4004 = ~n12634 ;
  assign y4005 = n12636 ;
  assign y4006 = n12640 ;
  assign y4007 = ~n12641 ;
  assign y4008 = ~1'b0 ;
  assign y4009 = ~n5526 ;
  assign y4010 = ~n12643 ;
  assign y4011 = n12644 ;
  assign y4012 = ~n12645 ;
  assign y4013 = ~n12652 ;
  assign y4014 = ~1'b0 ;
  assign y4015 = ~1'b0 ;
  assign y4016 = n12653 ;
  assign y4017 = n12654 ;
  assign y4018 = ~n12655 ;
  assign y4019 = n12660 ;
  assign y4020 = x24 ;
  assign y4021 = ~n12661 ;
  assign y4022 = ~n12668 ;
  assign y4023 = n12672 ;
  assign y4024 = n12673 ;
  assign y4025 = ~1'b0 ;
  assign y4026 = ~n12676 ;
  assign y4027 = ~1'b0 ;
  assign y4028 = ~1'b0 ;
  assign y4029 = ~n12678 ;
  assign y4030 = ~n12681 ;
  assign y4031 = ~1'b0 ;
  assign y4032 = ~n12688 ;
  assign y4033 = ~n12689 ;
  assign y4034 = ~n12694 ;
  assign y4035 = ~n12695 ;
  assign y4036 = n12702 ;
  assign y4037 = n12705 ;
  assign y4038 = ~n12706 ;
  assign y4039 = ~1'b0 ;
  assign y4040 = ~n12709 ;
  assign y4041 = ~1'b0 ;
  assign y4042 = n12711 ;
  assign y4043 = ~1'b0 ;
  assign y4044 = ~n12712 ;
  assign y4045 = n12718 ;
  assign y4046 = ~1'b0 ;
  assign y4047 = ~1'b0 ;
  assign y4048 = ~n12723 ;
  assign y4049 = n12724 ;
  assign y4050 = n12728 ;
  assign y4051 = n12733 ;
  assign y4052 = n12738 ;
  assign y4053 = n12741 ;
  assign y4054 = ~n12742 ;
  assign y4055 = n12744 ;
  assign y4056 = ~1'b0 ;
  assign y4057 = n12748 ;
  assign y4058 = n12750 ;
  assign y4059 = ~n12753 ;
  assign y4060 = n12755 ;
  assign y4061 = n12760 ;
  assign y4062 = ~n12765 ;
  assign y4063 = n12767 ;
  assign y4064 = ~n12770 ;
  assign y4065 = n12772 ;
  assign y4066 = n12776 ;
  assign y4067 = ~n12780 ;
  assign y4068 = n12786 ;
  assign y4069 = ~n12788 ;
  assign y4070 = ~n12796 ;
  assign y4071 = n12799 ;
  assign y4072 = ~n12801 ;
  assign y4073 = n12804 ;
  assign y4074 = ~n12810 ;
  assign y4075 = ~n12813 ;
  assign y4076 = n12815 ;
  assign y4077 = ~n12816 ;
  assign y4078 = ~1'b0 ;
  assign y4079 = n12817 ;
  assign y4080 = n12826 ;
  assign y4081 = ~n12830 ;
  assign y4082 = ~n12834 ;
  assign y4083 = ~n12837 ;
  assign y4084 = ~n12839 ;
  assign y4085 = n12840 ;
  assign y4086 = ~n12845 ;
  assign y4087 = ~n12846 ;
  assign y4088 = ~n12847 ;
  assign y4089 = n12848 ;
  assign y4090 = ~1'b0 ;
  assign y4091 = ~1'b0 ;
  assign y4092 = ~n12852 ;
  assign y4093 = n12854 ;
  assign y4094 = ~n12859 ;
  assign y4095 = n12862 ;
  assign y4096 = ~1'b0 ;
  assign y4097 = ~n12863 ;
  assign y4098 = ~n12865 ;
  assign y4099 = ~n12866 ;
  assign y4100 = n12871 ;
  assign y4101 = ~1'b0 ;
  assign y4102 = n12873 ;
  assign y4103 = n12880 ;
  assign y4104 = ~1'b0 ;
  assign y4105 = ~n12882 ;
  assign y4106 = n12885 ;
  assign y4107 = n12891 ;
  assign y4108 = n12894 ;
  assign y4109 = ~1'b0 ;
  assign y4110 = n12901 ;
  assign y4111 = n12902 ;
  assign y4112 = ~n12908 ;
  assign y4113 = n12915 ;
  assign y4114 = n12918 ;
  assign y4115 = ~n12920 ;
  assign y4116 = ~n12921 ;
  assign y4117 = n12927 ;
  assign y4118 = n1543 ;
  assign y4119 = ~n12930 ;
  assign y4120 = n12937 ;
  assign y4121 = ~1'b0 ;
  assign y4122 = ~n12940 ;
  assign y4123 = ~n12942 ;
  assign y4124 = ~1'b0 ;
  assign y4125 = n12943 ;
  assign y4126 = ~n12950 ;
  assign y4127 = ~1'b0 ;
  assign y4128 = n12951 ;
  assign y4129 = n12956 ;
  assign y4130 = ~1'b0 ;
  assign y4131 = n12957 ;
  assign y4132 = n12959 ;
  assign y4133 = ~1'b0 ;
  assign y4134 = n12962 ;
  assign y4135 = ~1'b0 ;
  assign y4136 = ~x37 ;
  assign y4137 = n12972 ;
  assign y4138 = ~1'b0 ;
  assign y4139 = ~n12977 ;
  assign y4140 = ~n12980 ;
  assign y4141 = ~n12986 ;
  assign y4142 = ~n12988 ;
  assign y4143 = n12989 ;
  assign y4144 = 1'b0 ;
  assign y4145 = n12993 ;
  assign y4146 = n12994 ;
  assign y4147 = n12997 ;
  assign y4148 = n12998 ;
  assign y4149 = ~n12999 ;
  assign y4150 = ~n11340 ;
  assign y4151 = n13007 ;
  assign y4152 = n13008 ;
  assign y4153 = ~n13009 ;
  assign y4154 = n13011 ;
  assign y4155 = ~1'b0 ;
  assign y4156 = n13013 ;
  assign y4157 = ~1'b0 ;
  assign y4158 = ~n13014 ;
  assign y4159 = ~n13015 ;
  assign y4160 = ~1'b0 ;
  assign y4161 = ~1'b0 ;
  assign y4162 = n13016 ;
  assign y4163 = ~n13018 ;
  assign y4164 = ~n13023 ;
  assign y4165 = n13026 ;
  assign y4166 = n13028 ;
  assign y4167 = ~n13030 ;
  assign y4168 = ~n13031 ;
  assign y4169 = ~n13032 ;
  assign y4170 = ~1'b0 ;
  assign y4171 = ~1'b0 ;
  assign y4172 = n13035 ;
  assign y4173 = ~1'b0 ;
  assign y4174 = ~1'b0 ;
  assign y4175 = n13036 ;
  assign y4176 = ~n13040 ;
  assign y4177 = ~n13042 ;
  assign y4178 = n13046 ;
  assign y4179 = n13052 ;
  assign y4180 = ~n13057 ;
  assign y4181 = ~n13066 ;
  assign y4182 = ~n13071 ;
  assign y4183 = ~1'b0 ;
  assign y4184 = n13076 ;
  assign y4185 = n13078 ;
  assign y4186 = n13082 ;
  assign y4187 = ~n13084 ;
  assign y4188 = ~1'b0 ;
  assign y4189 = ~1'b0 ;
  assign y4190 = ~1'b0 ;
  assign y4191 = n13086 ;
  assign y4192 = ~n13097 ;
  assign y4193 = n13102 ;
  assign y4194 = ~1'b0 ;
  assign y4195 = ~1'b0 ;
  assign y4196 = ~n13105 ;
  assign y4197 = n1762 ;
  assign y4198 = ~1'b0 ;
  assign y4199 = n13108 ;
  assign y4200 = ~n13115 ;
  assign y4201 = ~n13121 ;
  assign y4202 = n13122 ;
  assign y4203 = n13129 ;
  assign y4204 = ~n13132 ;
  assign y4205 = ~n13151 ;
  assign y4206 = 1'b0 ;
  assign y4207 = n13156 ;
  assign y4208 = n13157 ;
  assign y4209 = n13164 ;
  assign y4210 = ~1'b0 ;
  assign y4211 = ~n13167 ;
  assign y4212 = ~n13173 ;
  assign y4213 = n13174 ;
  assign y4214 = n13180 ;
  assign y4215 = ~n13185 ;
  assign y4216 = ~n13189 ;
  assign y4217 = ~n13199 ;
  assign y4218 = ~n13207 ;
  assign y4219 = n13213 ;
  assign y4220 = n13218 ;
  assign y4221 = ~n13225 ;
  assign y4222 = ~1'b0 ;
  assign y4223 = n13228 ;
  assign y4224 = ~n13230 ;
  assign y4225 = ~1'b0 ;
  assign y4226 = ~n13236 ;
  assign y4227 = n13238 ;
  assign y4228 = ~1'b0 ;
  assign y4229 = ~n13240 ;
  assign y4230 = ~n13248 ;
  assign y4231 = n13249 ;
  assign y4232 = n13251 ;
  assign y4233 = ~n13253 ;
  assign y4234 = n12832 ;
  assign y4235 = ~n13256 ;
  assign y4236 = ~1'b0 ;
  assign y4237 = ~1'b0 ;
  assign y4238 = ~1'b0 ;
  assign y4239 = ~1'b0 ;
  assign y4240 = ~n13258 ;
  assign y4241 = n13259 ;
  assign y4242 = ~1'b0 ;
  assign y4243 = n13260 ;
  assign y4244 = ~n13268 ;
  assign y4245 = ~n13269 ;
  assign y4246 = n13270 ;
  assign y4247 = ~n13271 ;
  assign y4248 = ~n13274 ;
  assign y4249 = n13275 ;
  assign y4250 = n13276 ;
  assign y4251 = ~n13279 ;
  assign y4252 = n13282 ;
  assign y4253 = ~n13284 ;
  assign y4254 = ~n13287 ;
  assign y4255 = ~1'b0 ;
  assign y4256 = ~1'b0 ;
  assign y4257 = n13291 ;
  assign y4258 = ~1'b0 ;
  assign y4259 = ~n13292 ;
  assign y4260 = ~1'b0 ;
  assign y4261 = ~n13293 ;
  assign y4262 = ~n13294 ;
  assign y4263 = ~n13297 ;
  assign y4264 = ~n1482 ;
  assign y4265 = ~n13301 ;
  assign y4266 = n13302 ;
  assign y4267 = ~n13304 ;
  assign y4268 = ~n13306 ;
  assign y4269 = n13309 ;
  assign y4270 = ~1'b0 ;
  assign y4271 = ~n13311 ;
  assign y4272 = n13313 ;
  assign y4273 = n13316 ;
  assign y4274 = n13317 ;
  assign y4275 = ~n13320 ;
  assign y4276 = ~n13322 ;
  assign y4277 = ~n1612 ;
  assign y4278 = n13326 ;
  assign y4279 = n13327 ;
  assign y4280 = ~n13328 ;
  assign y4281 = ~n13336 ;
  assign y4282 = n13341 ;
  assign y4283 = ~n13346 ;
  assign y4284 = ~n13348 ;
  assign y4285 = n13349 ;
  assign y4286 = ~n13352 ;
  assign y4287 = ~n13356 ;
  assign y4288 = ~n13357 ;
  assign y4289 = ~n13223 ;
  assign y4290 = ~1'b0 ;
  assign y4291 = ~n13358 ;
  assign y4292 = ~n13361 ;
  assign y4293 = ~1'b0 ;
  assign y4294 = ~n13365 ;
  assign y4295 = n13369 ;
  assign y4296 = ~n13373 ;
  assign y4297 = ~n13375 ;
  assign y4298 = ~n13378 ;
  assign y4299 = n13380 ;
  assign y4300 = n13383 ;
  assign y4301 = ~n13385 ;
  assign y4302 = ~n12862 ;
  assign y4303 = n13386 ;
  assign y4304 = ~n13387 ;
  assign y4305 = n13391 ;
  assign y4306 = ~n13395 ;
  assign y4307 = ~n13402 ;
  assign y4308 = n13403 ;
  assign y4309 = n13405 ;
  assign y4310 = n13408 ;
  assign y4311 = ~1'b0 ;
  assign y4312 = ~n13409 ;
  assign y4313 = n13411 ;
  assign y4314 = ~n13420 ;
  assign y4315 = ~1'b0 ;
  assign y4316 = n13429 ;
  assign y4317 = ~n13430 ;
  assign y4318 = ~n13432 ;
  assign y4319 = n13436 ;
  assign y4320 = ~1'b0 ;
  assign y4321 = n13438 ;
  assign y4322 = ~n13439 ;
  assign y4323 = ~n13446 ;
  assign y4324 = ~1'b0 ;
  assign y4325 = ~n13452 ;
  assign y4326 = n13459 ;
  assign y4327 = n13463 ;
  assign y4328 = ~1'b0 ;
  assign y4329 = ~n13464 ;
  assign y4330 = n13465 ;
  assign y4331 = n13467 ;
  assign y4332 = n13471 ;
  assign y4333 = n13473 ;
  assign y4334 = ~n13475 ;
  assign y4335 = n13482 ;
  assign y4336 = ~n8972 ;
  assign y4337 = ~1'b0 ;
  assign y4338 = ~1'b0 ;
  assign y4339 = n13483 ;
  assign y4340 = ~n13484 ;
  assign y4341 = ~n13491 ;
  assign y4342 = ~n13492 ;
  assign y4343 = n13501 ;
  assign y4344 = n13502 ;
  assign y4345 = n13508 ;
  assign y4346 = n13509 ;
  assign y4347 = ~n13513 ;
  assign y4348 = n13517 ;
  assign y4349 = ~1'b0 ;
  assign y4350 = ~n13520 ;
  assign y4351 = n13527 ;
  assign y4352 = 1'b0 ;
  assign y4353 = n13532 ;
  assign y4354 = ~1'b0 ;
  assign y4355 = n13533 ;
  assign y4356 = ~n8754 ;
  assign y4357 = ~n13536 ;
  assign y4358 = ~n13537 ;
  assign y4359 = n13538 ;
  assign y4360 = n13543 ;
  assign y4361 = ~n13546 ;
  assign y4362 = ~n13552 ;
  assign y4363 = n13557 ;
  assign y4364 = n13562 ;
  assign y4365 = ~n13565 ;
  assign y4366 = ~n13567 ;
  assign y4367 = ~n13569 ;
  assign y4368 = ~n13575 ;
  assign y4369 = n13581 ;
  assign y4370 = n13586 ;
  assign y4371 = ~1'b0 ;
  assign y4372 = ~n13589 ;
  assign y4373 = ~1'b0 ;
  assign y4374 = ~1'b0 ;
  assign y4375 = ~n13593 ;
  assign y4376 = n13596 ;
  assign y4377 = n13598 ;
  assign y4378 = ~1'b0 ;
  assign y4379 = ~1'b0 ;
  assign y4380 = ~n13599 ;
  assign y4381 = ~1'b0 ;
  assign y4382 = ~n13602 ;
  assign y4383 = n13605 ;
  assign y4384 = ~n13609 ;
  assign y4385 = ~1'b0 ;
  assign y4386 = n13610 ;
  assign y4387 = ~n13618 ;
  assign y4388 = ~n13622 ;
  assign y4389 = n13623 ;
  assign y4390 = ~n13626 ;
  assign y4391 = ~n13630 ;
  assign y4392 = n13635 ;
  assign y4393 = n13648 ;
  assign y4394 = n13650 ;
  assign y4395 = n13651 ;
  assign y4396 = n13652 ;
  assign y4397 = ~n13659 ;
  assign y4398 = n13662 ;
  assign y4399 = n13665 ;
  assign y4400 = n13666 ;
  assign y4401 = n13669 ;
  assign y4402 = ~1'b0 ;
  assign y4403 = ~n13670 ;
  assign y4404 = ~n13675 ;
  assign y4405 = ~1'b0 ;
  assign y4406 = n13677 ;
  assign y4407 = ~n5821 ;
  assign y4408 = n13679 ;
  assign y4409 = n13682 ;
  assign y4410 = n13683 ;
  assign y4411 = ~n13689 ;
  assign y4412 = ~n13691 ;
  assign y4413 = n13697 ;
  assign y4414 = ~n13698 ;
  assign y4415 = n13708 ;
  assign y4416 = ~n13710 ;
  assign y4417 = ~n13711 ;
  assign y4418 = ~n13715 ;
  assign y4419 = n7542 ;
  assign y4420 = ~n13723 ;
  assign y4421 = ~1'b0 ;
  assign y4422 = ~n13724 ;
  assign y4423 = ~n13727 ;
  assign y4424 = ~n13126 ;
  assign y4425 = ~1'b0 ;
  assign y4426 = n13730 ;
  assign y4427 = ~n13731 ;
  assign y4428 = n13735 ;
  assign y4429 = ~n13736 ;
  assign y4430 = ~1'b0 ;
  assign y4431 = n13738 ;
  assign y4432 = n13745 ;
  assign y4433 = ~n13747 ;
  assign y4434 = ~n13749 ;
  assign y4435 = n13750 ;
  assign y4436 = n13755 ;
  assign y4437 = ~1'b0 ;
  assign y4438 = n13756 ;
  assign y4439 = n13757 ;
  assign y4440 = n13762 ;
  assign y4441 = n13766 ;
  assign y4442 = n13767 ;
  assign y4443 = ~n13771 ;
  assign y4444 = ~n13772 ;
  assign y4445 = ~n13775 ;
  assign y4446 = ~n13776 ;
  assign y4447 = ~n13778 ;
  assign y4448 = n13780 ;
  assign y4449 = ~n13785 ;
  assign y4450 = n13789 ;
  assign y4451 = ~n13791 ;
  assign y4452 = ~n13793 ;
  assign y4453 = n13796 ;
  assign y4454 = ~n13797 ;
  assign y4455 = ~1'b0 ;
  assign y4456 = ~n13801 ;
  assign y4457 = ~1'b0 ;
  assign y4458 = ~n13805 ;
  assign y4459 = ~1'b0 ;
  assign y4460 = ~n13806 ;
  assign y4461 = ~n13808 ;
  assign y4462 = n13809 ;
  assign y4463 = ~1'b0 ;
  assign y4464 = ~1'b0 ;
  assign y4465 = ~1'b0 ;
  assign y4466 = n13811 ;
  assign y4467 = ~n13812 ;
  assign y4468 = ~n1311 ;
  assign y4469 = ~1'b0 ;
  assign y4470 = n13813 ;
  assign y4471 = ~1'b0 ;
  assign y4472 = ~n13818 ;
  assign y4473 = ~n13819 ;
  assign y4474 = ~n13822 ;
  assign y4475 = ~n13825 ;
  assign y4476 = ~1'b0 ;
  assign y4477 = n13826 ;
  assign y4478 = ~n13830 ;
  assign y4479 = n13835 ;
  assign y4480 = ~n13839 ;
  assign y4481 = n13842 ;
  assign y4482 = n13843 ;
  assign y4483 = n13844 ;
  assign y4484 = n13846 ;
  assign y4485 = ~1'b0 ;
  assign y4486 = n13847 ;
  assign y4487 = ~1'b0 ;
  assign y4488 = n13849 ;
  assign y4489 = ~1'b0 ;
  assign y4490 = n13851 ;
  assign y4491 = ~n13854 ;
  assign y4492 = ~n13858 ;
  assign y4493 = ~n13860 ;
  assign y4494 = ~n13863 ;
  assign y4495 = n13866 ;
  assign y4496 = n13867 ;
  assign y4497 = ~n13880 ;
  assign y4498 = ~1'b0 ;
  assign y4499 = n13884 ;
  assign y4500 = ~1'b0 ;
  assign y4501 = n13886 ;
  assign y4502 = ~n13887 ;
  assign y4503 = ~n13890 ;
  assign y4504 = ~1'b0 ;
  assign y4505 = ~n13897 ;
  assign y4506 = ~n13901 ;
  assign y4507 = n13905 ;
  assign y4508 = n13907 ;
  assign y4509 = ~n13913 ;
  assign y4510 = n13918 ;
  assign y4511 = n13919 ;
  assign y4512 = n13920 ;
  assign y4513 = n13923 ;
  assign y4514 = ~n13925 ;
  assign y4515 = ~1'b0 ;
  assign y4516 = ~1'b0 ;
  assign y4517 = ~n13926 ;
  assign y4518 = n13932 ;
  assign y4519 = n13934 ;
  assign y4520 = ~1'b0 ;
  assign y4521 = ~1'b0 ;
  assign y4522 = n13940 ;
  assign y4523 = n13946 ;
  assign y4524 = ~n13947 ;
  assign y4525 = n13948 ;
  assign y4526 = ~n13949 ;
  assign y4527 = n13953 ;
  assign y4528 = ~n13957 ;
  assign y4529 = ~1'b0 ;
  assign y4530 = ~1'b0 ;
  assign y4531 = ~n13959 ;
  assign y4532 = ~n13966 ;
  assign y4533 = n13968 ;
  assign y4534 = ~1'b0 ;
  assign y4535 = ~1'b0 ;
  assign y4536 = n13969 ;
  assign y4537 = n13970 ;
  assign y4538 = n13971 ;
  assign y4539 = ~n13976 ;
  assign y4540 = n13978 ;
  assign y4541 = ~n13982 ;
  assign y4542 = n13990 ;
  assign y4543 = ~n13992 ;
  assign y4544 = ~n13996 ;
  assign y4545 = n14000 ;
  assign y4546 = n14002 ;
  assign y4547 = ~n14004 ;
  assign y4548 = ~n14005 ;
  assign y4549 = ~1'b0 ;
  assign y4550 = ~n14008 ;
  assign y4551 = ~n14012 ;
  assign y4552 = ~n14015 ;
  assign y4553 = ~n14016 ;
  assign y4554 = ~n14017 ;
  assign y4555 = ~n14021 ;
  assign y4556 = ~1'b0 ;
  assign y4557 = ~n14025 ;
  assign y4558 = n14030 ;
  assign y4559 = ~n14031 ;
  assign y4560 = ~n14036 ;
  assign y4561 = n14039 ;
  assign y4562 = n14042 ;
  assign y4563 = ~n14044 ;
  assign y4564 = n14046 ;
  assign y4565 = n14047 ;
  assign y4566 = ~n14050 ;
  assign y4567 = 1'b0 ;
  assign y4568 = ~1'b0 ;
  assign y4569 = n14061 ;
  assign y4570 = n14063 ;
  assign y4571 = ~1'b0 ;
  assign y4572 = ~n10135 ;
  assign y4573 = ~n14070 ;
  assign y4574 = ~n14072 ;
  assign y4575 = ~n14074 ;
  assign y4576 = ~n14080 ;
  assign y4577 = n14086 ;
  assign y4578 = n1802 ;
  assign y4579 = ~n14087 ;
  assign y4580 = ~n14091 ;
  assign y4581 = ~1'b0 ;
  assign y4582 = ~n14096 ;
  assign y4583 = n14099 ;
  assign y4584 = n14103 ;
  assign y4585 = ~1'b0 ;
  assign y4586 = n14104 ;
  assign y4587 = ~n14105 ;
  assign y4588 = ~n14107 ;
  assign y4589 = ~n14111 ;
  assign y4590 = n14114 ;
  assign y4591 = ~1'b0 ;
  assign y4592 = ~1'b0 ;
  assign y4593 = ~n14115 ;
  assign y4594 = n14116 ;
  assign y4595 = n14118 ;
  assign y4596 = n14120 ;
  assign y4597 = ~n14124 ;
  assign y4598 = ~1'b0 ;
  assign y4599 = n14125 ;
  assign y4600 = n14129 ;
  assign y4601 = n14130 ;
  assign y4602 = ~n14134 ;
  assign y4603 = ~n14135 ;
  assign y4604 = n14138 ;
  assign y4605 = ~n14139 ;
  assign y4606 = n14143 ;
  assign y4607 = n14153 ;
  assign y4608 = n14154 ;
  assign y4609 = ~n14156 ;
  assign y4610 = n14160 ;
  assign y4611 = ~n14165 ;
  assign y4612 = n14167 ;
  assign y4613 = n14169 ;
  assign y4614 = n14171 ;
  assign y4615 = n14173 ;
  assign y4616 = n14180 ;
  assign y4617 = n14184 ;
  assign y4618 = n14192 ;
  assign y4619 = ~1'b0 ;
  assign y4620 = ~1'b0 ;
  assign y4621 = ~n14194 ;
  assign y4622 = ~n14195 ;
  assign y4623 = n14196 ;
  assign y4624 = ~n14197 ;
  assign y4625 = ~1'b0 ;
  assign y4626 = ~n14200 ;
  assign y4627 = ~1'b0 ;
  assign y4628 = ~n14201 ;
  assign y4629 = ~n14202 ;
  assign y4630 = n14205 ;
  assign y4631 = ~n14207 ;
  assign y4632 = ~n14208 ;
  assign y4633 = ~1'b0 ;
  assign y4634 = ~n14214 ;
  assign y4635 = n14217 ;
  assign y4636 = n2496 ;
  assign y4637 = n14219 ;
  assign y4638 = ~1'b0 ;
  assign y4639 = ~n14223 ;
  assign y4640 = ~1'b0 ;
  assign y4641 = ~n14228 ;
  assign y4642 = ~n14234 ;
  assign y4643 = ~1'b0 ;
  assign y4644 = n14239 ;
  assign y4645 = n14241 ;
  assign y4646 = n14245 ;
  assign y4647 = ~1'b0 ;
  assign y4648 = ~n14246 ;
  assign y4649 = n14248 ;
  assign y4650 = ~n14250 ;
  assign y4651 = ~1'b0 ;
  assign y4652 = n14258 ;
  assign y4653 = n14263 ;
  assign y4654 = ~1'b0 ;
  assign y4655 = ~n14264 ;
  assign y4656 = ~n14267 ;
  assign y4657 = n14269 ;
  assign y4658 = n14275 ;
  assign y4659 = n14276 ;
  assign y4660 = ~n14277 ;
  assign y4661 = ~n14280 ;
  assign y4662 = n14281 ;
  assign y4663 = n14282 ;
  assign y4664 = ~n14283 ;
  assign y4665 = n14288 ;
  assign y4666 = ~n14291 ;
  assign y4667 = ~n14294 ;
  assign y4668 = n14295 ;
  assign y4669 = n14302 ;
  assign y4670 = ~n14303 ;
  assign y4671 = ~n14304 ;
  assign y4672 = n14306 ;
  assign y4673 = ~n14307 ;
  assign y4674 = ~1'b0 ;
  assign y4675 = n14311 ;
  assign y4676 = ~n14315 ;
  assign y4677 = n14316 ;
  assign y4678 = ~n14317 ;
  assign y4679 = 1'b0 ;
  assign y4680 = ~1'b0 ;
  assign y4681 = ~1'b0 ;
  assign y4682 = ~n14329 ;
  assign y4683 = n14334 ;
  assign y4684 = ~n14336 ;
  assign y4685 = n14340 ;
  assign y4686 = n14349 ;
  assign y4687 = n14351 ;
  assign y4688 = ~n14352 ;
  assign y4689 = ~n14353 ;
  assign y4690 = n14355 ;
  assign y4691 = ~n14358 ;
  assign y4692 = n14364 ;
  assign y4693 = n14366 ;
  assign y4694 = n14370 ;
  assign y4695 = n14380 ;
  assign y4696 = ~n14383 ;
  assign y4697 = n14384 ;
  assign y4698 = n14386 ;
  assign y4699 = n14393 ;
  assign y4700 = ~1'b0 ;
  assign y4701 = n14394 ;
  assign y4702 = ~n14395 ;
  assign y4703 = ~n14397 ;
  assign y4704 = ~n14405 ;
  assign y4705 = ~n14407 ;
  assign y4706 = ~n14411 ;
  assign y4707 = n14417 ;
  assign y4708 = n14421 ;
  assign y4709 = ~n14424 ;
  assign y4710 = ~n14427 ;
  assign y4711 = n14430 ;
  assign y4712 = ~1'b0 ;
  assign y4713 = ~n14434 ;
  assign y4714 = n14436 ;
  assign y4715 = ~n14437 ;
  assign y4716 = n14438 ;
  assign y4717 = n14440 ;
  assign y4718 = ~1'b0 ;
  assign y4719 = n12041 ;
  assign y4720 = ~1'b0 ;
  assign y4721 = n14451 ;
  assign y4722 = n14452 ;
  assign y4723 = ~1'b0 ;
  assign y4724 = ~1'b0 ;
  assign y4725 = n14454 ;
  assign y4726 = n14455 ;
  assign y4727 = ~n14456 ;
  assign y4728 = ~1'b0 ;
  assign y4729 = ~n14458 ;
  assign y4730 = ~n14459 ;
  assign y4731 = n14464 ;
  assign y4732 = ~n14468 ;
  assign y4733 = ~n14471 ;
  assign y4734 = ~n14479 ;
  assign y4735 = ~n14481 ;
  assign y4736 = n14483 ;
  assign y4737 = n14486 ;
  assign y4738 = ~n5774 ;
  assign y4739 = ~1'b0 ;
  assign y4740 = ~n14487 ;
  assign y4741 = n14491 ;
  assign y4742 = ~n10729 ;
  assign y4743 = ~n14495 ;
  assign y4744 = ~n14498 ;
  assign y4745 = ~n14499 ;
  assign y4746 = ~n14505 ;
  assign y4747 = ~1'b0 ;
  assign y4748 = ~n14507 ;
  assign y4749 = n14517 ;
  assign y4750 = n14529 ;
  assign y4751 = ~1'b0 ;
  assign y4752 = ~n14536 ;
  assign y4753 = ~1'b0 ;
  assign y4754 = ~n14538 ;
  assign y4755 = n14539 ;
  assign y4756 = n14546 ;
  assign y4757 = ~n14547 ;
  assign y4758 = ~1'b0 ;
  assign y4759 = ~n14552 ;
  assign y4760 = n14555 ;
  assign y4761 = n14558 ;
  assign y4762 = n14565 ;
  assign y4763 = n7273 ;
  assign y4764 = n14566 ;
  assign y4765 = ~n14570 ;
  assign y4766 = ~n14571 ;
  assign y4767 = n14573 ;
  assign y4768 = n11620 ;
  assign y4769 = n14584 ;
  assign y4770 = ~n14586 ;
  assign y4771 = ~n14587 ;
  assign y4772 = ~n14595 ;
  assign y4773 = n14596 ;
  assign y4774 = n14604 ;
  assign y4775 = ~1'b0 ;
  assign y4776 = n14606 ;
  assign y4777 = n14607 ;
  assign y4778 = ~n14611 ;
  assign y4779 = ~1'b0 ;
  assign y4780 = ~n14613 ;
  assign y4781 = n14614 ;
  assign y4782 = n14616 ;
  assign y4783 = ~1'b0 ;
  assign y4784 = n14621 ;
  assign y4785 = n14622 ;
  assign y4786 = ~n14624 ;
  assign y4787 = n14626 ;
  assign y4788 = ~1'b0 ;
  assign y4789 = ~n14638 ;
  assign y4790 = ~n14642 ;
  assign y4791 = ~n14647 ;
  assign y4792 = n14648 ;
  assign y4793 = ~n14649 ;
  assign y4794 = ~1'b0 ;
  assign y4795 = ~1'b0 ;
  assign y4796 = ~n14652 ;
  assign y4797 = ~n14655 ;
  assign y4798 = n14661 ;
  assign y4799 = ~1'b0 ;
  assign y4800 = n11231 ;
  assign y4801 = ~n14665 ;
  assign y4802 = n14674 ;
  assign y4803 = ~n14676 ;
  assign y4804 = ~n5173 ;
  assign y4805 = ~n3766 ;
  assign y4806 = ~n14680 ;
  assign y4807 = ~n14684 ;
  assign y4808 = n14686 ;
  assign y4809 = n14687 ;
  assign y4810 = ~n14690 ;
  assign y4811 = ~1'b0 ;
  assign y4812 = ~n14693 ;
  assign y4813 = n14694 ;
  assign y4814 = n14695 ;
  assign y4815 = ~n14696 ;
  assign y4816 = ~1'b0 ;
  assign y4817 = ~1'b0 ;
  assign y4818 = n14699 ;
  assign y4819 = n14704 ;
  assign y4820 = ~n14706 ;
  assign y4821 = ~n14707 ;
  assign y4822 = n14711 ;
  assign y4823 = ~n14713 ;
  assign y4824 = n14716 ;
  assign y4825 = ~n14720 ;
  assign y4826 = ~n14725 ;
  assign y4827 = n14730 ;
  assign y4828 = ~n14733 ;
  assign y4829 = ~1'b0 ;
  assign y4830 = ~n14737 ;
  assign y4831 = n14739 ;
  assign y4832 = ~n14742 ;
  assign y4833 = ~n14748 ;
  assign y4834 = n14758 ;
  assign y4835 = n14760 ;
  assign y4836 = 1'b0 ;
  assign y4837 = ~1'b0 ;
  assign y4838 = ~n14761 ;
  assign y4839 = ~n14763 ;
  assign y4840 = n14764 ;
  assign y4841 = n14765 ;
  assign y4842 = ~1'b0 ;
  assign y4843 = n14768 ;
  assign y4844 = ~n14770 ;
  assign y4845 = n14774 ;
  assign y4846 = ~1'b0 ;
  assign y4847 = n14779 ;
  assign y4848 = ~n14781 ;
  assign y4849 = n14783 ;
  assign y4850 = n14789 ;
  assign y4851 = n14791 ;
  assign y4852 = n14797 ;
  assign y4853 = ~1'b0 ;
  assign y4854 = ~1'b0 ;
  assign y4855 = ~1'b0 ;
  assign y4856 = ~1'b0 ;
  assign y4857 = n14800 ;
  assign y4858 = ~1'b0 ;
  assign y4859 = ~1'b0 ;
  assign y4860 = ~n14801 ;
  assign y4861 = ~n14802 ;
  assign y4862 = ~n14804 ;
  assign y4863 = ~n14809 ;
  assign y4864 = n14811 ;
  assign y4865 = n14816 ;
  assign y4866 = n14820 ;
  assign y4867 = ~n14824 ;
  assign y4868 = ~1'b0 ;
  assign y4869 = n14826 ;
  assign y4870 = ~n14828 ;
  assign y4871 = ~n14830 ;
  assign y4872 = ~1'b0 ;
  assign y4873 = ~n14836 ;
  assign y4874 = n14838 ;
  assign y4875 = ~n14840 ;
  assign y4876 = n14843 ;
  assign y4877 = n14845 ;
  assign y4878 = ~1'b0 ;
  assign y4879 = ~n14848 ;
  assign y4880 = ~n14853 ;
  assign y4881 = n14854 ;
  assign y4882 = n14857 ;
  assign y4883 = ~n14859 ;
  assign y4884 = ~n14860 ;
  assign y4885 = ~n14864 ;
  assign y4886 = ~n14869 ;
  assign y4887 = n14870 ;
  assign y4888 = n14873 ;
  assign y4889 = ~1'b0 ;
  assign y4890 = ~n14874 ;
  assign y4891 = n14876 ;
  assign y4892 = n14877 ;
  assign y4893 = ~n14881 ;
  assign y4894 = ~n14884 ;
  assign y4895 = ~n14889 ;
  assign y4896 = n14892 ;
  assign y4897 = ~1'b0 ;
  assign y4898 = ~n14896 ;
  assign y4899 = ~n14903 ;
  assign y4900 = ~n14906 ;
  assign y4901 = n14910 ;
  assign y4902 = ~n14912 ;
  assign y4903 = n14917 ;
  assign y4904 = ~1'b0 ;
  assign y4905 = ~n14920 ;
  assign y4906 = ~n14922 ;
  assign y4907 = ~n14924 ;
  assign y4908 = ~1'b0 ;
  assign y4909 = n14926 ;
  assign y4910 = ~n14929 ;
  assign y4911 = ~n14935 ;
  assign y4912 = n14937 ;
  assign y4913 = ~1'b0 ;
  assign y4914 = n14939 ;
  assign y4915 = n14941 ;
  assign y4916 = ~n14946 ;
  assign y4917 = ~n14957 ;
  assign y4918 = n14959 ;
  assign y4919 = ~1'b0 ;
  assign y4920 = n14963 ;
  assign y4921 = n14964 ;
  assign y4922 = n14969 ;
  assign y4923 = n14973 ;
  assign y4924 = ~n14975 ;
  assign y4925 = ~n14977 ;
  assign y4926 = n14982 ;
  assign y4927 = n14987 ;
  assign y4928 = n14988 ;
  assign y4929 = ~1'b0 ;
  assign y4930 = ~1'b0 ;
  assign y4931 = ~n14989 ;
  assign y4932 = ~n14991 ;
  assign y4933 = ~n14992 ;
  assign y4934 = ~1'b0 ;
  assign y4935 = n14995 ;
  assign y4936 = ~1'b0 ;
  assign y4937 = ~1'b0 ;
  assign y4938 = n15002 ;
  assign y4939 = ~n15005 ;
  assign y4940 = ~n15006 ;
  assign y4941 = ~1'b0 ;
  assign y4942 = n15008 ;
  assign y4943 = ~n15010 ;
  assign y4944 = ~n15011 ;
  assign y4945 = n15012 ;
  assign y4946 = ~n15017 ;
  assign y4947 = ~1'b0 ;
  assign y4948 = ~n15024 ;
  assign y4949 = ~n15033 ;
  assign y4950 = n15034 ;
  assign y4951 = ~n15037 ;
  assign y4952 = ~n15044 ;
  assign y4953 = ~n15046 ;
  assign y4954 = ~n15048 ;
  assign y4955 = ~n15050 ;
  assign y4956 = ~n15055 ;
  assign y4957 = n15057 ;
  assign y4958 = ~n15060 ;
  assign y4959 = ~n15062 ;
  assign y4960 = ~1'b0 ;
  assign y4961 = n15066 ;
  assign y4962 = n15073 ;
  assign y4963 = n15076 ;
  assign y4964 = ~1'b0 ;
  assign y4965 = ~n15077 ;
  assign y4966 = ~n15080 ;
  assign y4967 = n15083 ;
  assign y4968 = n15084 ;
  assign y4969 = ~n15088 ;
  assign y4970 = ~1'b0 ;
  assign y4971 = ~1'b0 ;
  assign y4972 = ~n15090 ;
  assign y4973 = n15092 ;
  assign y4974 = n15094 ;
  assign y4975 = n15101 ;
  assign y4976 = ~n15105 ;
  assign y4977 = ~1'b0 ;
  assign y4978 = ~n15109 ;
  assign y4979 = n15113 ;
  assign y4980 = ~n15117 ;
  assign y4981 = n15121 ;
  assign y4982 = n15125 ;
  assign y4983 = ~n15134 ;
  assign y4984 = ~n15140 ;
  assign y4985 = n15141 ;
  assign y4986 = ~n15142 ;
  assign y4987 = n15146 ;
  assign y4988 = n15147 ;
  assign y4989 = ~1'b0 ;
  assign y4990 = n15149 ;
  assign y4991 = ~n15152 ;
  assign y4992 = n15154 ;
  assign y4993 = n15155 ;
  assign y4994 = ~1'b0 ;
  assign y4995 = ~n15157 ;
  assign y4996 = ~1'b0 ;
  assign y4997 = n15158 ;
  assign y4998 = ~n8586 ;
  assign y4999 = ~n15159 ;
  assign y5000 = n15163 ;
  assign y5001 = ~n15170 ;
  assign y5002 = n15171 ;
  assign y5003 = n15174 ;
  assign y5004 = n15179 ;
  assign y5005 = n15180 ;
  assign y5006 = ~1'b0 ;
  assign y5007 = n15181 ;
  assign y5008 = ~n15185 ;
  assign y5009 = ~n15193 ;
  assign y5010 = n15195 ;
  assign y5011 = ~1'b0 ;
  assign y5012 = n15198 ;
  assign y5013 = ~n15204 ;
  assign y5014 = ~n15208 ;
  assign y5015 = n15214 ;
  assign y5016 = n15215 ;
  assign y5017 = n15216 ;
  assign y5018 = ~n15223 ;
  assign y5019 = ~n15225 ;
  assign y5020 = n15230 ;
  assign y5021 = ~1'b0 ;
  assign y5022 = n15234 ;
  assign y5023 = ~n15235 ;
  assign y5024 = ~1'b0 ;
  assign y5025 = ~1'b0 ;
  assign y5026 = ~n15241 ;
  assign y5027 = n15243 ;
  assign y5028 = ~1'b0 ;
  assign y5029 = ~1'b0 ;
  assign y5030 = ~1'b0 ;
  assign y5031 = ~n15244 ;
  assign y5032 = ~1'b0 ;
  assign y5033 = n15247 ;
  assign y5034 = n15252 ;
  assign y5035 = n15255 ;
  assign y5036 = ~n15259 ;
  assign y5037 = ~n15262 ;
  assign y5038 = ~n15263 ;
  assign y5039 = n15267 ;
  assign y5040 = ~1'b0 ;
  assign y5041 = ~1'b0 ;
  assign y5042 = n15269 ;
  assign y5043 = ~n15270 ;
  assign y5044 = n15276 ;
  assign y5045 = ~n15277 ;
  assign y5046 = n15278 ;
  assign y5047 = ~n15279 ;
  assign y5048 = ~1'b0 ;
  assign y5049 = ~n15281 ;
  assign y5050 = ~1'b0 ;
  assign y5051 = ~1'b0 ;
  assign y5052 = n15282 ;
  assign y5053 = ~1'b0 ;
  assign y5054 = ~n15283 ;
  assign y5055 = n15286 ;
  assign y5056 = n15287 ;
  assign y5057 = ~n15289 ;
  assign y5058 = n15292 ;
  assign y5059 = n15296 ;
  assign y5060 = ~n15298 ;
  assign y5061 = ~1'b0 ;
  assign y5062 = ~n15302 ;
  assign y5063 = n15303 ;
  assign y5064 = ~n15304 ;
  assign y5065 = n15308 ;
  assign y5066 = ~n15310 ;
  assign y5067 = ~1'b0 ;
  assign y5068 = n15311 ;
  assign y5069 = n11022 ;
  assign y5070 = ~n15312 ;
  assign y5071 = n15314 ;
  assign y5072 = n15316 ;
  assign y5073 = n15320 ;
  assign y5074 = n15321 ;
  assign y5075 = n15322 ;
  assign y5076 = ~n15323 ;
  assign y5077 = ~1'b0 ;
  assign y5078 = ~1'b0 ;
  assign y5079 = ~n15327 ;
  assign y5080 = n15329 ;
  assign y5081 = ~n15334 ;
  assign y5082 = ~n15338 ;
  assign y5083 = n15339 ;
  assign y5084 = n15343 ;
  assign y5085 = ~1'b0 ;
  assign y5086 = ~n15349 ;
  assign y5087 = ~n15352 ;
  assign y5088 = n15355 ;
  assign y5089 = ~1'b0 ;
  assign y5090 = ~1'b0 ;
  assign y5091 = n15357 ;
  assign y5092 = ~n15359 ;
  assign y5093 = n15360 ;
  assign y5094 = n13330 ;
  assign y5095 = n15364 ;
  assign y5096 = ~1'b0 ;
  assign y5097 = n15367 ;
  assign y5098 = n15372 ;
  assign y5099 = ~1'b0 ;
  assign y5100 = n15379 ;
  assign y5101 = ~n15382 ;
  assign y5102 = ~n15388 ;
  assign y5103 = n15389 ;
  assign y5104 = n15394 ;
  assign y5105 = n15396 ;
  assign y5106 = ~n15401 ;
  assign y5107 = n15403 ;
  assign y5108 = n15407 ;
  assign y5109 = n15408 ;
  assign y5110 = ~n15409 ;
  assign y5111 = n15411 ;
  assign y5112 = ~1'b0 ;
  assign y5113 = ~n15419 ;
  assign y5114 = n15424 ;
  assign y5115 = n15426 ;
  assign y5116 = n15429 ;
  assign y5117 = ~n15432 ;
  assign y5118 = ~n15435 ;
  assign y5119 = ~1'b0 ;
  assign y5120 = ~n15439 ;
  assign y5121 = ~n15441 ;
  assign y5122 = n15444 ;
  assign y5123 = ~n15445 ;
  assign y5124 = ~1'b0 ;
  assign y5125 = n15446 ;
  assign y5126 = ~n15448 ;
  assign y5127 = ~1'b0 ;
  assign y5128 = ~n15450 ;
  assign y5129 = ~n13784 ;
  assign y5130 = ~n15451 ;
  assign y5131 = n15452 ;
  assign y5132 = n15455 ;
  assign y5133 = ~1'b0 ;
  assign y5134 = ~n15457 ;
  assign y5135 = ~n15467 ;
  assign y5136 = ~n15469 ;
  assign y5137 = n15470 ;
  assign y5138 = ~1'b0 ;
  assign y5139 = n15471 ;
  assign y5140 = ~1'b0 ;
  assign y5141 = ~n15472 ;
  assign y5142 = n15473 ;
  assign y5143 = n15484 ;
  assign y5144 = ~1'b0 ;
  assign y5145 = ~n15488 ;
  assign y5146 = ~n15498 ;
  assign y5147 = n15500 ;
  assign y5148 = ~1'b0 ;
  assign y5149 = n15504 ;
  assign y5150 = ~n15506 ;
  assign y5151 = ~n15510 ;
  assign y5152 = ~n15511 ;
  assign y5153 = n15513 ;
  assign y5154 = ~1'b0 ;
  assign y5155 = ~n15514 ;
  assign y5156 = ~n15515 ;
  assign y5157 = ~n15520 ;
  assign y5158 = n15522 ;
  assign y5159 = ~n15523 ;
  assign y5160 = n15524 ;
  assign y5161 = ~n15525 ;
  assign y5162 = n15526 ;
  assign y5163 = ~n15530 ;
  assign y5164 = ~1'b0 ;
  assign y5165 = ~n15536 ;
  assign y5166 = n15537 ;
  assign y5167 = ~n15540 ;
  assign y5168 = n15542 ;
  assign y5169 = ~n15544 ;
  assign y5170 = ~1'b0 ;
  assign y5171 = n15555 ;
  assign y5172 = n15557 ;
  assign y5173 = n15560 ;
  assign y5174 = ~n15571 ;
  assign y5175 = n15572 ;
  assign y5176 = ~1'b0 ;
  assign y5177 = n15578 ;
  assign y5178 = n15586 ;
  assign y5179 = n15587 ;
  assign y5180 = ~n15589 ;
  assign y5181 = ~n15591 ;
  assign y5182 = n15598 ;
  assign y5183 = ~1'b0 ;
  assign y5184 = n15601 ;
  assign y5185 = n15603 ;
  assign y5186 = n15605 ;
  assign y5187 = n15609 ;
  assign y5188 = ~n15616 ;
  assign y5189 = ~n15621 ;
  assign y5190 = ~1'b0 ;
  assign y5191 = n15623 ;
  assign y5192 = ~n15628 ;
  assign y5193 = ~n6482 ;
  assign y5194 = ~n15629 ;
  assign y5195 = n15630 ;
  assign y5196 = n15633 ;
  assign y5197 = n15634 ;
  assign y5198 = n15635 ;
  assign y5199 = n3422 ;
  assign y5200 = n15636 ;
  assign y5201 = ~1'b0 ;
  assign y5202 = ~1'b0 ;
  assign y5203 = ~n15637 ;
  assign y5204 = ~n15638 ;
  assign y5205 = ~n15642 ;
  assign y5206 = n15644 ;
  assign y5207 = n15656 ;
  assign y5208 = ~1'b0 ;
  assign y5209 = n15657 ;
  assign y5210 = n15660 ;
  assign y5211 = n15665 ;
  assign y5212 = n15667 ;
  assign y5213 = 1'b0 ;
  assign y5214 = ~1'b0 ;
  assign y5215 = ~n15668 ;
  assign y5216 = ~1'b0 ;
  assign y5217 = ~1'b0 ;
  assign y5218 = ~n15672 ;
  assign y5219 = ~n15674 ;
  assign y5220 = n15678 ;
  assign y5221 = ~n15683 ;
  assign y5222 = n15686 ;
  assign y5223 = ~1'b0 ;
  assign y5224 = ~n15687 ;
  assign y5225 = ~n15688 ;
  assign y5226 = n15689 ;
  assign y5227 = n15690 ;
  assign y5228 = n15695 ;
  assign y5229 = ~n15697 ;
  assign y5230 = ~1'b0 ;
  assign y5231 = ~n15702 ;
  assign y5232 = n15710 ;
  assign y5233 = ~n15711 ;
  assign y5234 = n15713 ;
  assign y5235 = n15715 ;
  assign y5236 = ~n15720 ;
  assign y5237 = ~n15721 ;
  assign y5238 = ~n15725 ;
  assign y5239 = ~n15730 ;
  assign y5240 = n15738 ;
  assign y5241 = ~n15744 ;
  assign y5242 = n15745 ;
  assign y5243 = ~n15748 ;
  assign y5244 = ~n15750 ;
  assign y5245 = ~n15760 ;
  assign y5246 = ~1'b0 ;
  assign y5247 = ~n15761 ;
  assign y5248 = ~n15762 ;
  assign y5249 = n15767 ;
  assign y5250 = ~n15772 ;
  assign y5251 = ~n15774 ;
  assign y5252 = n15779 ;
  assign y5253 = ~n15784 ;
  assign y5254 = ~n15789 ;
  assign y5255 = n15792 ;
  assign y5256 = n15794 ;
  assign y5257 = ~n15799 ;
  assign y5258 = ~n15800 ;
  assign y5259 = ~n15805 ;
  assign y5260 = ~n15807 ;
  assign y5261 = n15808 ;
  assign y5262 = n15809 ;
  assign y5263 = ~n15811 ;
  assign y5264 = n15814 ;
  assign y5265 = ~1'b0 ;
  assign y5266 = ~1'b0 ;
  assign y5267 = ~1'b0 ;
  assign y5268 = ~n15819 ;
  assign y5269 = ~n15821 ;
  assign y5270 = n15830 ;
  assign y5271 = ~1'b0 ;
  assign y5272 = n15832 ;
  assign y5273 = n15835 ;
  assign y5274 = ~1'b0 ;
  assign y5275 = n15839 ;
  assign y5276 = ~1'b0 ;
  assign y5277 = n15841 ;
  assign y5278 = ~n15844 ;
  assign y5279 = n15845 ;
  assign y5280 = n15849 ;
  assign y5281 = ~1'b0 ;
  assign y5282 = n15852 ;
  assign y5283 = n15856 ;
  assign y5284 = ~n15861 ;
  assign y5285 = n15866 ;
  assign y5286 = n15867 ;
  assign y5287 = ~1'b0 ;
  assign y5288 = ~1'b0 ;
  assign y5289 = ~n15872 ;
  assign y5290 = ~n15874 ;
  assign y5291 = ~n15877 ;
  assign y5292 = n15878 ;
  assign y5293 = ~n15885 ;
  assign y5294 = ~1'b0 ;
  assign y5295 = ~n15889 ;
  assign y5296 = ~n9819 ;
  assign y5297 = n15890 ;
  assign y5298 = n15900 ;
  assign y5299 = n15903 ;
  assign y5300 = n15905 ;
  assign y5301 = ~n15907 ;
  assign y5302 = ~n15908 ;
  assign y5303 = n15911 ;
  assign y5304 = ~n15912 ;
  assign y5305 = ~1'b0 ;
  assign y5306 = ~n15915 ;
  assign y5307 = ~n15917 ;
  assign y5308 = n15922 ;
  assign y5309 = ~1'b0 ;
  assign y5310 = ~1'b0 ;
  assign y5311 = ~n15927 ;
  assign y5312 = ~n15931 ;
  assign y5313 = n15933 ;
  assign y5314 = ~1'b0 ;
  assign y5315 = ~n15935 ;
  assign y5316 = ~1'b0 ;
  assign y5317 = ~n15939 ;
  assign y5318 = ~n15941 ;
  assign y5319 = n15943 ;
  assign y5320 = ~1'b0 ;
  assign y5321 = n15945 ;
  assign y5322 = ~n15953 ;
  assign y5323 = ~1'b0 ;
  assign y5324 = ~n15956 ;
  assign y5325 = ~n15962 ;
  assign y5326 = ~1'b0 ;
  assign y5327 = ~n15964 ;
  assign y5328 = n15965 ;
  assign y5329 = ~n149 ;
  assign y5330 = ~n15969 ;
  assign y5331 = ~n15973 ;
  assign y5332 = n15976 ;
  assign y5333 = ~n15980 ;
  assign y5334 = ~n15988 ;
  assign y5335 = n15997 ;
  assign y5336 = n16003 ;
  assign y5337 = n16004 ;
  assign y5338 = ~1'b0 ;
  assign y5339 = ~1'b0 ;
  assign y5340 = ~n16008 ;
  assign y5341 = ~n16011 ;
  assign y5342 = n16020 ;
  assign y5343 = ~n16028 ;
  assign y5344 = ~n16033 ;
  assign y5345 = n16038 ;
  assign y5346 = ~1'b0 ;
  assign y5347 = ~1'b0 ;
  assign y5348 = ~n16040 ;
  assign y5349 = ~n16046 ;
  assign y5350 = n16047 ;
  assign y5351 = ~n16054 ;
  assign y5352 = n16056 ;
  assign y5353 = n16059 ;
  assign y5354 = n16061 ;
  assign y5355 = n16064 ;
  assign y5356 = ~n16065 ;
  assign y5357 = n16066 ;
  assign y5358 = ~n5387 ;
  assign y5359 = ~n16073 ;
  assign y5360 = ~n16074 ;
  assign y5361 = n16075 ;
  assign y5362 = ~n16079 ;
  assign y5363 = n16080 ;
  assign y5364 = n16081 ;
  assign y5365 = ~n16083 ;
  assign y5366 = n16084 ;
  assign y5367 = ~n16088 ;
  assign y5368 = ~n16091 ;
  assign y5369 = n16092 ;
  assign y5370 = ~1'b0 ;
  assign y5371 = ~1'b0 ;
  assign y5372 = ~1'b0 ;
  assign y5373 = ~n16098 ;
  assign y5374 = ~n16099 ;
  assign y5375 = ~n16100 ;
  assign y5376 = ~n16103 ;
  assign y5377 = ~1'b0 ;
  assign y5378 = ~1'b0 ;
  assign y5379 = ~n16104 ;
  assign y5380 = n16105 ;
  assign y5381 = ~n16107 ;
  assign y5382 = ~n16113 ;
  assign y5383 = ~n16116 ;
  assign y5384 = n16118 ;
  assign y5385 = ~n16124 ;
  assign y5386 = ~1'b0 ;
  assign y5387 = ~1'b0 ;
  assign y5388 = n16129 ;
  assign y5389 = n16130 ;
  assign y5390 = ~n16134 ;
  assign y5391 = ~n16142 ;
  assign y5392 = ~1'b0 ;
  assign y5393 = ~n16144 ;
  assign y5394 = ~n16148 ;
  assign y5395 = ~n16152 ;
  assign y5396 = n16155 ;
  assign y5397 = ~n16160 ;
  assign y5398 = n16164 ;
  assign y5399 = ~n3538 ;
  assign y5400 = ~n16169 ;
  assign y5401 = n11406 ;
  assign y5402 = n16173 ;
  assign y5403 = ~1'b0 ;
  assign y5404 = ~n16176 ;
  assign y5405 = n16184 ;
  assign y5406 = ~n16194 ;
  assign y5407 = ~n16196 ;
  assign y5408 = n16198 ;
  assign y5409 = ~n16202 ;
  assign y5410 = ~n16204 ;
  assign y5411 = n16206 ;
  assign y5412 = n16208 ;
  assign y5413 = ~1'b0 ;
  assign y5414 = ~n16210 ;
  assign y5415 = ~n16213 ;
  assign y5416 = n16215 ;
  assign y5417 = n16216 ;
  assign y5418 = ~n16217 ;
  assign y5419 = ~n16219 ;
  assign y5420 = ~n16220 ;
  assign y5421 = ~n16221 ;
  assign y5422 = ~n16222 ;
  assign y5423 = ~1'b0 ;
  assign y5424 = n16223 ;
  assign y5425 = ~1'b0 ;
  assign y5426 = n16224 ;
  assign y5427 = ~n16226 ;
  assign y5428 = ~n16228 ;
  assign y5429 = ~n16231 ;
  assign y5430 = n16235 ;
  assign y5431 = ~n16237 ;
  assign y5432 = ~1'b0 ;
  assign y5433 = ~n16243 ;
  assign y5434 = n16246 ;
  assign y5435 = n16247 ;
  assign y5436 = ~n16249 ;
  assign y5437 = n16257 ;
  assign y5438 = ~n16260 ;
  assign y5439 = ~1'b0 ;
  assign y5440 = ~n16263 ;
  assign y5441 = ~n16271 ;
  assign y5442 = n16274 ;
  assign y5443 = n16278 ;
  assign y5444 = ~n16284 ;
  assign y5445 = ~1'b0 ;
  assign y5446 = 1'b0 ;
  assign y5447 = n16285 ;
  assign y5448 = ~n16293 ;
  assign y5449 = ~n16296 ;
  assign y5450 = ~1'b0 ;
  assign y5451 = n7912 ;
  assign y5452 = ~n16297 ;
  assign y5453 = ~n16298 ;
  assign y5454 = ~1'b0 ;
  assign y5455 = ~n16300 ;
  assign y5456 = n16309 ;
  assign y5457 = n16321 ;
  assign y5458 = ~n16322 ;
  assign y5459 = n16329 ;
  assign y5460 = ~n16332 ;
  assign y5461 = n16334 ;
  assign y5462 = ~1'b0 ;
  assign y5463 = ~n16347 ;
  assign y5464 = ~n16352 ;
  assign y5465 = n16354 ;
  assign y5466 = 1'b0 ;
  assign y5467 = 1'b0 ;
  assign y5468 = n16357 ;
  assign y5469 = n7104 ;
  assign y5470 = n16358 ;
  assign y5471 = ~n16359 ;
  assign y5472 = ~n16368 ;
  assign y5473 = ~1'b0 ;
  assign y5474 = n16375 ;
  assign y5475 = n16381 ;
  assign y5476 = ~1'b0 ;
  assign y5477 = ~n16382 ;
  assign y5478 = n16383 ;
  assign y5479 = n16389 ;
  assign y5480 = ~n16390 ;
  assign y5481 = n16392 ;
  assign y5482 = n16393 ;
  assign y5483 = n16395 ;
  assign y5484 = ~1'b0 ;
  assign y5485 = ~1'b0 ;
  assign y5486 = ~1'b0 ;
  assign y5487 = n16401 ;
  assign y5488 = n16402 ;
  assign y5489 = ~n16403 ;
  assign y5490 = ~n16405 ;
  assign y5491 = ~n16406 ;
  assign y5492 = n16409 ;
  assign y5493 = ~n16413 ;
  assign y5494 = ~1'b0 ;
  assign y5495 = ~1'b0 ;
  assign y5496 = ~n16417 ;
  assign y5497 = n6575 ;
  assign y5498 = ~n16418 ;
  assign y5499 = ~1'b0 ;
  assign y5500 = n16420 ;
  assign y5501 = n16423 ;
  assign y5502 = ~n16425 ;
  assign y5503 = n16427 ;
  assign y5504 = ~1'b0 ;
  assign y5505 = ~1'b0 ;
  assign y5506 = ~1'b0 ;
  assign y5507 = n16429 ;
  assign y5508 = ~1'b0 ;
  assign y5509 = ~n16437 ;
  assign y5510 = n16439 ;
  assign y5511 = ~1'b0 ;
  assign y5512 = n16441 ;
  assign y5513 = ~n16444 ;
  assign y5514 = ~n16449 ;
  assign y5515 = ~n16451 ;
  assign y5516 = n16453 ;
  assign y5517 = ~1'b0 ;
  assign y5518 = n16454 ;
  assign y5519 = ~n16457 ;
  assign y5520 = ~1'b0 ;
  assign y5521 = n16458 ;
  assign y5522 = ~1'b0 ;
  assign y5523 = ~1'b0 ;
  assign y5524 = ~n16460 ;
  assign y5525 = n16463 ;
  assign y5526 = ~n16471 ;
  assign y5527 = ~n16472 ;
  assign y5528 = n1701 ;
  assign y5529 = ~1'b0 ;
  assign y5530 = n16479 ;
  assign y5531 = ~1'b0 ;
  assign y5532 = n16486 ;
  assign y5533 = ~n16489 ;
  assign y5534 = ~n16491 ;
  assign y5535 = ~n16493 ;
  assign y5536 = ~n16495 ;
  assign y5537 = n16497 ;
  assign y5538 = ~n16503 ;
  assign y5539 = ~n16504 ;
  assign y5540 = ~1'b0 ;
  assign y5541 = ~1'b0 ;
  assign y5542 = ~n16505 ;
  assign y5543 = ~n16506 ;
  assign y5544 = n16510 ;
  assign y5545 = ~n16511 ;
  assign y5546 = n16513 ;
  assign y5547 = ~n16515 ;
  assign y5548 = n16516 ;
  assign y5549 = ~1'b0 ;
  assign y5550 = ~1'b0 ;
  assign y5551 = ~1'b0 ;
  assign y5552 = ~n16518 ;
  assign y5553 = n16524 ;
  assign y5554 = ~n16528 ;
  assign y5555 = n16529 ;
  assign y5556 = ~1'b0 ;
  assign y5557 = ~n16532 ;
  assign y5558 = n16534 ;
  assign y5559 = n16535 ;
  assign y5560 = ~n16536 ;
  assign y5561 = n16539 ;
  assign y5562 = ~n16542 ;
  assign y5563 = 1'b0 ;
  assign y5564 = ~1'b0 ;
  assign y5565 = ~n16545 ;
  assign y5566 = ~n16551 ;
  assign y5567 = ~n16552 ;
  assign y5568 = n16561 ;
  assign y5569 = ~n16566 ;
  assign y5570 = ~n16568 ;
  assign y5571 = ~n16569 ;
  assign y5572 = ~n16571 ;
  assign y5573 = ~n16572 ;
  assign y5574 = n16580 ;
  assign y5575 = ~n16581 ;
  assign y5576 = ~1'b0 ;
  assign y5577 = ~n13460 ;
  assign y5578 = ~n16582 ;
  assign y5579 = n16586 ;
  assign y5580 = n16590 ;
  assign y5581 = ~1'b0 ;
  assign y5582 = ~n16592 ;
  assign y5583 = ~n16599 ;
  assign y5584 = n16600 ;
  assign y5585 = ~1'b0 ;
  assign y5586 = ~n16603 ;
  assign y5587 = n16605 ;
  assign y5588 = n16615 ;
  assign y5589 = ~1'b0 ;
  assign y5590 = ~1'b0 ;
  assign y5591 = n16623 ;
  assign y5592 = n16626 ;
  assign y5593 = n1838 ;
  assign y5594 = ~n16628 ;
  assign y5595 = ~n16632 ;
  assign y5596 = ~n16635 ;
  assign y5597 = n16637 ;
  assign y5598 = ~n16638 ;
  assign y5599 = n16640 ;
  assign y5600 = ~n16642 ;
  assign y5601 = ~n16644 ;
  assign y5602 = ~n16645 ;
  assign y5603 = ~1'b0 ;
  assign y5604 = ~1'b0 ;
  assign y5605 = ~1'b0 ;
  assign y5606 = n16649 ;
  assign y5607 = ~n16650 ;
  assign y5608 = n16655 ;
  assign y5609 = ~n16663 ;
  assign y5610 = ~1'b0 ;
  assign y5611 = ~1'b0 ;
  assign y5612 = ~n16669 ;
  assign y5613 = ~1'b0 ;
  assign y5614 = n16671 ;
  assign y5615 = ~n16674 ;
  assign y5616 = n16678 ;
  assign y5617 = ~n16686 ;
  assign y5618 = ~n16687 ;
  assign y5619 = ~n16688 ;
  assign y5620 = ~n16695 ;
  assign y5621 = ~1'b0 ;
  assign y5622 = ~1'b0 ;
  assign y5623 = n16701 ;
  assign y5624 = n16702 ;
  assign y5625 = ~n16707 ;
  assign y5626 = n16710 ;
  assign y5627 = n16712 ;
  assign y5628 = ~1'b0 ;
  assign y5629 = ~n16713 ;
  assign y5630 = ~n16716 ;
  assign y5631 = n16720 ;
  assign y5632 = ~n16724 ;
  assign y5633 = n16734 ;
  assign y5634 = n16740 ;
  assign y5635 = n16743 ;
  assign y5636 = n16747 ;
  assign y5637 = n16748 ;
  assign y5638 = ~n16752 ;
  assign y5639 = n16761 ;
  assign y5640 = 1'b0 ;
  assign y5641 = ~n16768 ;
  assign y5642 = ~1'b0 ;
  assign y5643 = ~n16770 ;
  assign y5644 = ~n16771 ;
  assign y5645 = n16773 ;
  assign y5646 = ~n16775 ;
  assign y5647 = ~n16776 ;
  assign y5648 = ~1'b0 ;
  assign y5649 = ~n16780 ;
  assign y5650 = n16783 ;
  assign y5651 = n16784 ;
  assign y5652 = ~1'b0 ;
  assign y5653 = ~1'b0 ;
  assign y5654 = ~n16788 ;
  assign y5655 = n16789 ;
  assign y5656 = ~n16790 ;
  assign y5657 = ~n16793 ;
  assign y5658 = n16796 ;
  assign y5659 = n16798 ;
  assign y5660 = n16801 ;
  assign y5661 = n16804 ;
  assign y5662 = ~1'b0 ;
  assign y5663 = ~1'b0 ;
  assign y5664 = n16820 ;
  assign y5665 = n16821 ;
  assign y5666 = ~n16823 ;
  assign y5667 = n16825 ;
  assign y5668 = ~n16829 ;
  assign y5669 = n16835 ;
  assign y5670 = ~n16836 ;
  assign y5671 = ~n16848 ;
  assign y5672 = n16849 ;
  assign y5673 = n16851 ;
  assign y5674 = n16852 ;
  assign y5675 = n16853 ;
  assign y5676 = ~n16855 ;
  assign y5677 = ~n16859 ;
  assign y5678 = ~n16861 ;
  assign y5679 = ~1'b0 ;
  assign y5680 = ~n16868 ;
  assign y5681 = ~n16873 ;
  assign y5682 = ~n16874 ;
  assign y5683 = ~n16875 ;
  assign y5684 = ~1'b0 ;
  assign y5685 = n16876 ;
  assign y5686 = ~1'b0 ;
  assign y5687 = ~n16883 ;
  assign y5688 = ~n16887 ;
  assign y5689 = n16893 ;
  assign y5690 = ~n16897 ;
  assign y5691 = ~n16899 ;
  assign y5692 = ~n16900 ;
  assign y5693 = ~1'b0 ;
  assign y5694 = ~n16905 ;
  assign y5695 = n16906 ;
  assign y5696 = ~n16907 ;
  assign y5697 = ~n16911 ;
  assign y5698 = n16913 ;
  assign y5699 = ~n16917 ;
  assign y5700 = ~n16925 ;
  assign y5701 = n16926 ;
  assign y5702 = ~n16927 ;
  assign y5703 = ~n16936 ;
  assign y5704 = ~n16938 ;
  assign y5705 = ~n16939 ;
  assign y5706 = ~n16942 ;
  assign y5707 = ~n16949 ;
  assign y5708 = ~n16951 ;
  assign y5709 = ~n16953 ;
  assign y5710 = ~n16957 ;
  assign y5711 = ~n1217 ;
  assign y5712 = ~n16958 ;
  assign y5713 = n16964 ;
  assign y5714 = n16969 ;
  assign y5715 = n16971 ;
  assign y5716 = n16974 ;
  assign y5717 = ~n16977 ;
  assign y5718 = n16984 ;
  assign y5719 = ~n16985 ;
  assign y5720 = ~n16988 ;
  assign y5721 = n16997 ;
  assign y5722 = ~1'b0 ;
  assign y5723 = ~n16999 ;
  assign y5724 = ~n17002 ;
  assign y5725 = ~n17004 ;
  assign y5726 = ~n17007 ;
  assign y5727 = ~n7874 ;
  assign y5728 = ~n17009 ;
  assign y5729 = ~1'b0 ;
  assign y5730 = ~n12601 ;
  assign y5731 = ~n17010 ;
  assign y5732 = ~n17021 ;
  assign y5733 = ~n17022 ;
  assign y5734 = n17023 ;
  assign y5735 = n17026 ;
  assign y5736 = ~n17028 ;
  assign y5737 = 1'b0 ;
  assign y5738 = ~n17030 ;
  assign y5739 = n17032 ;
  assign y5740 = ~n17036 ;
  assign y5741 = 1'b0 ;
  assign y5742 = ~n17037 ;
  assign y5743 = n17042 ;
  assign y5744 = ~n17044 ;
  assign y5745 = n17045 ;
  assign y5746 = n17051 ;
  assign y5747 = ~1'b0 ;
  assign y5748 = ~1'b0 ;
  assign y5749 = ~n17052 ;
  assign y5750 = n17053 ;
  assign y5751 = n17055 ;
  assign y5752 = ~n17056 ;
  assign y5753 = ~n17062 ;
  assign y5754 = n17067 ;
  assign y5755 = ~n17072 ;
  assign y5756 = n17073 ;
  assign y5757 = n17077 ;
  assign y5758 = n17080 ;
  assign y5759 = n17084 ;
  assign y5760 = n17085 ;
  assign y5761 = 1'b0 ;
  assign y5762 = ~1'b0 ;
  assign y5763 = ~n17088 ;
  assign y5764 = ~n17090 ;
  assign y5765 = n17092 ;
  assign y5766 = n17094 ;
  assign y5767 = n4515 ;
  assign y5768 = n17096 ;
  assign y5769 = ~n17098 ;
  assign y5770 = n17099 ;
  assign y5771 = n17106 ;
  assign y5772 = ~n17110 ;
  assign y5773 = ~n17111 ;
  assign y5774 = ~n17112 ;
  assign y5775 = ~n17114 ;
  assign y5776 = ~n17115 ;
  assign y5777 = ~n17118 ;
  assign y5778 = ~1'b0 ;
  assign y5779 = n17119 ;
  assign y5780 = n10214 ;
  assign y5781 = ~n17121 ;
  assign y5782 = ~n17122 ;
  assign y5783 = ~n17125 ;
  assign y5784 = ~1'b0 ;
  assign y5785 = ~1'b0 ;
  assign y5786 = ~1'b0 ;
  assign y5787 = n17127 ;
  assign y5788 = n17128 ;
  assign y5789 = n17129 ;
  assign y5790 = n17130 ;
  assign y5791 = ~n17135 ;
  assign y5792 = ~n17137 ;
  assign y5793 = ~n17142 ;
  assign y5794 = n17143 ;
  assign y5795 = n17145 ;
  assign y5796 = ~n17146 ;
  assign y5797 = ~1'b0 ;
  assign y5798 = n17150 ;
  assign y5799 = ~1'b0 ;
  assign y5800 = n17158 ;
  assign y5801 = ~n17163 ;
  assign y5802 = ~1'b0 ;
  assign y5803 = ~1'b0 ;
  assign y5804 = n17166 ;
  assign y5805 = n17168 ;
  assign y5806 = ~n17171 ;
  assign y5807 = ~n17173 ;
  assign y5808 = ~n17178 ;
  assign y5809 = ~n4118 ;
  assign y5810 = ~1'b0 ;
  assign y5811 = n17180 ;
  assign y5812 = n17188 ;
  assign y5813 = ~1'b0 ;
  assign y5814 = ~n17190 ;
  assign y5815 = ~1'b0 ;
  assign y5816 = n17192 ;
  assign y5817 = n17193 ;
  assign y5818 = n17194 ;
  assign y5819 = n17196 ;
  assign y5820 = ~1'b0 ;
  assign y5821 = ~n17199 ;
  assign y5822 = ~n17200 ;
  assign y5823 = n17201 ;
  assign y5824 = n17202 ;
  assign y5825 = ~n17203 ;
  assign y5826 = ~n17208 ;
  assign y5827 = ~n17209 ;
  assign y5828 = ~1'b0 ;
  assign y5829 = ~n17214 ;
  assign y5830 = n6953 ;
  assign y5831 = n17215 ;
  assign y5832 = n17224 ;
  assign y5833 = n17227 ;
  assign y5834 = n17232 ;
  assign y5835 = ~n17236 ;
  assign y5836 = n17240 ;
  assign y5837 = n17243 ;
  assign y5838 = n17253 ;
  assign y5839 = ~1'b0 ;
  assign y5840 = ~1'b0 ;
  assign y5841 = n17254 ;
  assign y5842 = ~n17258 ;
  assign y5843 = ~n17263 ;
  assign y5844 = n17265 ;
  assign y5845 = ~n17268 ;
  assign y5846 = n17269 ;
  assign y5847 = ~n17272 ;
  assign y5848 = ~n17273 ;
  assign y5849 = ~n17279 ;
  assign y5850 = ~n17288 ;
  assign y5851 = ~1'b0 ;
  assign y5852 = ~1'b0 ;
  assign y5853 = ~n17292 ;
  assign y5854 = n17295 ;
  assign y5855 = ~1'b0 ;
  assign y5856 = ~1'b0 ;
  assign y5857 = n17297 ;
  assign y5858 = n17298 ;
  assign y5859 = ~1'b0 ;
  assign y5860 = ~n17300 ;
  assign y5861 = ~n17303 ;
  assign y5862 = n17305 ;
  assign y5863 = n17308 ;
  assign y5864 = n17309 ;
  assign y5865 = n17316 ;
  assign y5866 = ~n17322 ;
  assign y5867 = n17323 ;
  assign y5868 = n17326 ;
  assign y5869 = n17327 ;
  assign y5870 = ~n17329 ;
  assign y5871 = ~n17334 ;
  assign y5872 = n17335 ;
  assign y5873 = ~n17337 ;
  assign y5874 = ~1'b0 ;
  assign y5875 = n17338 ;
  assign y5876 = n17341 ;
  assign y5877 = n17344 ;
  assign y5878 = ~n17347 ;
  assign y5879 = ~n17353 ;
  assign y5880 = ~1'b0 ;
  assign y5881 = n9728 ;
  assign y5882 = n17356 ;
  assign y5883 = n17357 ;
  assign y5884 = ~n17358 ;
  assign y5885 = ~n17360 ;
  assign y5886 = ~n17365 ;
  assign y5887 = ~n17366 ;
  assign y5888 = ~1'b0 ;
  assign y5889 = ~n629 ;
  assign y5890 = ~n17369 ;
  assign y5891 = ~n17373 ;
  assign y5892 = ~n17377 ;
  assign y5893 = n17381 ;
  assign y5894 = ~n17383 ;
  assign y5895 = n17384 ;
  assign y5896 = ~n17386 ;
  assign y5897 = ~1'b0 ;
  assign y5898 = ~1'b0 ;
  assign y5899 = n17388 ;
  assign y5900 = n17391 ;
  assign y5901 = ~n17392 ;
  assign y5902 = ~1'b0 ;
  assign y5903 = ~n17396 ;
  assign y5904 = ~1'b0 ;
  assign y5905 = n17398 ;
  assign y5906 = ~n17399 ;
  assign y5907 = ~n17402 ;
  assign y5908 = ~n17416 ;
  assign y5909 = ~n17419 ;
  assign y5910 = ~n17424 ;
  assign y5911 = ~1'b0 ;
  assign y5912 = n17426 ;
  assign y5913 = n17429 ;
  assign y5914 = n17432 ;
  assign y5915 = ~1'b0 ;
  assign y5916 = n17435 ;
  assign y5917 = ~1'b0 ;
  assign y5918 = n17441 ;
  assign y5919 = ~n17443 ;
  assign y5920 = n17444 ;
  assign y5921 = n17449 ;
  assign y5922 = n17450 ;
  assign y5923 = ~n17452 ;
  assign y5924 = ~1'b0 ;
  assign y5925 = ~n17454 ;
  assign y5926 = n17456 ;
  assign y5927 = n9857 ;
  assign y5928 = n17457 ;
  assign y5929 = ~n17460 ;
  assign y5930 = ~n17461 ;
  assign y5931 = ~1'b0 ;
  assign y5932 = ~n17463 ;
  assign y5933 = ~n17466 ;
  assign y5934 = n17467 ;
  assign y5935 = ~1'b0 ;
  assign y5936 = ~1'b0 ;
  assign y5937 = n17468 ;
  assign y5938 = ~n17469 ;
  assign y5939 = n17471 ;
  assign y5940 = ~1'b0 ;
  assign y5941 = n17474 ;
  assign y5942 = ~n17478 ;
  assign y5943 = n17479 ;
  assign y5944 = ~n17486 ;
  assign y5945 = n17488 ;
  assign y5946 = ~n17491 ;
  assign y5947 = n17495 ;
  assign y5948 = ~n17498 ;
  assign y5949 = n17502 ;
  assign y5950 = ~n17506 ;
  assign y5951 = n17508 ;
  assign y5952 = ~n17512 ;
  assign y5953 = n17514 ;
  assign y5954 = ~1'b0 ;
  assign y5955 = ~n17515 ;
  assign y5956 = ~n17518 ;
  assign y5957 = n17520 ;
  assign y5958 = n17521 ;
  assign y5959 = n17528 ;
  assign y5960 = ~n17530 ;
  assign y5961 = ~n17532 ;
  assign y5962 = n17533 ;
  assign y5963 = ~n17534 ;
  assign y5964 = ~n17538 ;
  assign y5965 = ~n17545 ;
  assign y5966 = n17549 ;
  assign y5967 = n7611 ;
  assign y5968 = n17550 ;
  assign y5969 = n17551 ;
  assign y5970 = ~n17556 ;
  assign y5971 = ~n17558 ;
  assign y5972 = n17560 ;
  assign y5973 = ~n17564 ;
  assign y5974 = n17565 ;
  assign y5975 = ~n17567 ;
  assign y5976 = n17569 ;
  assign y5977 = n17581 ;
  assign y5978 = n17588 ;
  assign y5979 = ~n17589 ;
  assign y5980 = ~1'b0 ;
  assign y5981 = ~n17590 ;
  assign y5982 = ~n17594 ;
  assign y5983 = ~n17600 ;
  assign y5984 = ~n17605 ;
  assign y5985 = n17616 ;
  assign y5986 = n17620 ;
  assign y5987 = ~1'b0 ;
  assign y5988 = ~1'b0 ;
  assign y5989 = ~1'b0 ;
  assign y5990 = n17624 ;
  assign y5991 = n17625 ;
  assign y5992 = n17628 ;
  assign y5993 = n17630 ;
  assign y5994 = ~1'b0 ;
  assign y5995 = ~n17632 ;
  assign y5996 = ~1'b0 ;
  assign y5997 = ~n17634 ;
  assign y5998 = ~n17636 ;
  assign y5999 = n17638 ;
  assign y6000 = ~n17639 ;
  assign y6001 = n17640 ;
  assign y6002 = n17642 ;
  assign y6003 = ~n17643 ;
  assign y6004 = n17644 ;
  assign y6005 = n17645 ;
  assign y6006 = n17648 ;
  assign y6007 = n17651 ;
  assign y6008 = ~n17653 ;
  assign y6009 = ~n17654 ;
  assign y6010 = n17655 ;
  assign y6011 = n17657 ;
  assign y6012 = ~n17658 ;
  assign y6013 = ~n17660 ;
  assign y6014 = n17663 ;
  assign y6015 = ~n17665 ;
  assign y6016 = ~1'b0 ;
  assign y6017 = n17667 ;
  assign y6018 = ~n17668 ;
  assign y6019 = ~n17671 ;
  assign y6020 = ~1'b0 ;
  assign y6021 = ~n17675 ;
  assign y6022 = ~n17676 ;
  assign y6023 = ~1'b0 ;
  assign y6024 = ~n17683 ;
  assign y6025 = ~n17685 ;
  assign y6026 = ~n17691 ;
  assign y6027 = ~n17694 ;
  assign y6028 = ~n17697 ;
  assign y6029 = ~1'b0 ;
  assign y6030 = n17700 ;
  assign y6031 = n17704 ;
  assign y6032 = ~n17706 ;
  assign y6033 = n17710 ;
  assign y6034 = ~n3224 ;
  assign y6035 = ~n17716 ;
  assign y6036 = n17717 ;
  assign y6037 = ~n17722 ;
  assign y6038 = ~n17726 ;
  assign y6039 = ~n17727 ;
  assign y6040 = ~n17733 ;
  assign y6041 = n17735 ;
  assign y6042 = ~n17739 ;
  assign y6043 = n17742 ;
  assign y6044 = n17744 ;
  assign y6045 = ~n17748 ;
  assign y6046 = ~n17754 ;
  assign y6047 = ~n17756 ;
  assign y6048 = ~n17759 ;
  assign y6049 = ~n8872 ;
  assign y6050 = n17760 ;
  assign y6051 = ~n17765 ;
  assign y6052 = ~n17767 ;
  assign y6053 = ~n17769 ;
  assign y6054 = ~n17770 ;
  assign y6055 = ~n17771 ;
  assign y6056 = ~n17772 ;
  assign y6057 = n17774 ;
  assign y6058 = n17775 ;
  assign y6059 = n17780 ;
  assign y6060 = n17782 ;
  assign y6061 = ~n17785 ;
  assign y6062 = n17790 ;
  assign y6063 = ~n17791 ;
  assign y6064 = ~n17796 ;
  assign y6065 = ~n11135 ;
  assign y6066 = n17798 ;
  assign y6067 = ~n17802 ;
  assign y6068 = ~1'b0 ;
  assign y6069 = n17803 ;
  assign y6070 = ~1'b0 ;
  assign y6071 = ~n17806 ;
  assign y6072 = n17807 ;
  assign y6073 = ~n17812 ;
  assign y6074 = ~1'b0 ;
  assign y6075 = ~n17819 ;
  assign y6076 = ~n17824 ;
  assign y6077 = ~n17826 ;
  assign y6078 = n17829 ;
  assign y6079 = ~n17830 ;
  assign y6080 = ~n17833 ;
  assign y6081 = n17838 ;
  assign y6082 = ~n17839 ;
  assign y6083 = n17841 ;
  assign y6084 = n17844 ;
  assign y6085 = ~n17846 ;
  assign y6086 = n17847 ;
  assign y6087 = ~n17854 ;
  assign y6088 = n17856 ;
  assign y6089 = n17857 ;
  assign y6090 = n17858 ;
  assign y6091 = ~n17859 ;
  assign y6092 = ~n17860 ;
  assign y6093 = n17862 ;
  assign y6094 = n17863 ;
  assign y6095 = n17865 ;
  assign y6096 = n17867 ;
  assign y6097 = ~n17871 ;
  assign y6098 = ~n17872 ;
  assign y6099 = ~n17873 ;
  assign y6100 = n17883 ;
  assign y6101 = ~1'b0 ;
  assign y6102 = n17885 ;
  assign y6103 = ~1'b0 ;
  assign y6104 = n17886 ;
  assign y6105 = ~n17887 ;
  assign y6106 = n17888 ;
  assign y6107 = n17892 ;
  assign y6108 = 1'b0 ;
  assign y6109 = n17895 ;
  assign y6110 = n17898 ;
  assign y6111 = n17900 ;
  assign y6112 = ~1'b0 ;
  assign y6113 = ~1'b0 ;
  assign y6114 = ~n17902 ;
  assign y6115 = n17903 ;
  assign y6116 = ~n17904 ;
  assign y6117 = ~n17908 ;
  assign y6118 = ~1'b0 ;
  assign y6119 = ~1'b0 ;
  assign y6120 = ~n17909 ;
  assign y6121 = ~n17910 ;
  assign y6122 = n17913 ;
  assign y6123 = ~n17917 ;
  assign y6124 = ~n17921 ;
  assign y6125 = ~1'b0 ;
  assign y6126 = ~n17923 ;
  assign y6127 = n17924 ;
  assign y6128 = ~n17925 ;
  assign y6129 = ~n17928 ;
  assign y6130 = ~1'b0 ;
  assign y6131 = ~1'b0 ;
  assign y6132 = ~n17933 ;
  assign y6133 = ~1'b0 ;
  assign y6134 = n17934 ;
  assign y6135 = ~n17935 ;
  assign y6136 = ~n17936 ;
  assign y6137 = ~n17938 ;
  assign y6138 = ~n17947 ;
  assign y6139 = ~n17952 ;
  assign y6140 = ~n17954 ;
  assign y6141 = n17955 ;
  assign y6142 = ~n17960 ;
  assign y6143 = ~n17962 ;
  assign y6144 = ~1'b0 ;
  assign y6145 = n17964 ;
  assign y6146 = ~n17971 ;
  assign y6147 = ~1'b0 ;
  assign y6148 = n17973 ;
  assign y6149 = n17978 ;
  assign y6150 = n17985 ;
  assign y6151 = ~n17988 ;
  assign y6152 = ~n17991 ;
  assign y6153 = ~n17993 ;
  assign y6154 = n17994 ;
  assign y6155 = n17995 ;
  assign y6156 = n17996 ;
  assign y6157 = n17997 ;
  assign y6158 = ~n18000 ;
  assign y6159 = ~n18003 ;
  assign y6160 = ~n18007 ;
  assign y6161 = ~n18009 ;
  assign y6162 = n18011 ;
  assign y6163 = 1'b0 ;
  assign y6164 = ~n18012 ;
  assign y6165 = n18013 ;
  assign y6166 = ~n18018 ;
  assign y6167 = ~n18021 ;
  assign y6168 = ~n18025 ;
  assign y6169 = ~n18028 ;
  assign y6170 = n18029 ;
  assign y6171 = n18032 ;
  assign y6172 = ~n18033 ;
  assign y6173 = ~1'b0 ;
  assign y6174 = n18035 ;
  assign y6175 = n18039 ;
  assign y6176 = ~n18046 ;
  assign y6177 = n18050 ;
  assign y6178 = ~n18061 ;
  assign y6179 = n18067 ;
  assign y6180 = ~1'b0 ;
  assign y6181 = n18068 ;
  assign y6182 = n18071 ;
  assign y6183 = ~n18077 ;
  assign y6184 = n18079 ;
  assign y6185 = ~1'b0 ;
  assign y6186 = n18080 ;
  assign y6187 = ~n18086 ;
  assign y6188 = ~1'b0 ;
  assign y6189 = ~n18094 ;
  assign y6190 = ~n3699 ;
  assign y6191 = ~n18101 ;
  assign y6192 = ~1'b0 ;
  assign y6193 = ~n18111 ;
  assign y6194 = ~n18112 ;
  assign y6195 = ~n18115 ;
  assign y6196 = ~n18116 ;
  assign y6197 = n18120 ;
  assign y6198 = n18122 ;
  assign y6199 = n18123 ;
  assign y6200 = ~n18125 ;
  assign y6201 = ~n18126 ;
  assign y6202 = n18127 ;
  assign y6203 = n18128 ;
  assign y6204 = ~n18132 ;
  assign y6205 = ~1'b0 ;
  assign y6206 = n18135 ;
  assign y6207 = n18140 ;
  assign y6208 = n18144 ;
  assign y6209 = n7611 ;
  assign y6210 = ~1'b0 ;
  assign y6211 = ~1'b0 ;
  assign y6212 = n18146 ;
  assign y6213 = ~n18151 ;
  assign y6214 = n18154 ;
  assign y6215 = n18155 ;
  assign y6216 = n18156 ;
  assign y6217 = n18157 ;
  assign y6218 = n18159 ;
  assign y6219 = ~1'b0 ;
  assign y6220 = n18163 ;
  assign y6221 = n18165 ;
  assign y6222 = n18169 ;
  assign y6223 = n18170 ;
  assign y6224 = ~1'b0 ;
  assign y6225 = ~1'b0 ;
  assign y6226 = ~1'b0 ;
  assign y6227 = n17786 ;
  assign y6228 = ~1'b0 ;
  assign y6229 = n18173 ;
  assign y6230 = n18179 ;
  assign y6231 = ~n18185 ;
  assign y6232 = n18191 ;
  assign y6233 = ~n18194 ;
  assign y6234 = ~n18195 ;
  assign y6235 = n18196 ;
  assign y6236 = ~n18199 ;
  assign y6237 = ~n18203 ;
  assign y6238 = ~1'b0 ;
  assign y6239 = ~n18205 ;
  assign y6240 = n18209 ;
  assign y6241 = ~n18210 ;
  assign y6242 = n18211 ;
  assign y6243 = ~1'b0 ;
  assign y6244 = n18217 ;
  assign y6245 = ~1'b0 ;
  assign y6246 = n18218 ;
  assign y6247 = n18223 ;
  assign y6248 = ~n18227 ;
  assign y6249 = ~n18228 ;
  assign y6250 = n18231 ;
  assign y6251 = ~n18233 ;
  assign y6252 = ~n18234 ;
  assign y6253 = ~n18237 ;
  assign y6254 = ~n18241 ;
  assign y6255 = n18242 ;
  assign y6256 = ~n18247 ;
  assign y6257 = ~n18248 ;
  assign y6258 = n18249 ;
  assign y6259 = ~1'b0 ;
  assign y6260 = n18253 ;
  assign y6261 = n18256 ;
  assign y6262 = ~n18258 ;
  assign y6263 = ~1'b0 ;
  assign y6264 = 1'b0 ;
  assign y6265 = n18259 ;
  assign y6266 = n18263 ;
  assign y6267 = ~n18265 ;
  assign y6268 = n18269 ;
  assign y6269 = n18270 ;
  assign y6270 = ~1'b0 ;
  assign y6271 = ~n18271 ;
  assign y6272 = n18272 ;
  assign y6273 = ~n18273 ;
  assign y6274 = ~n18276 ;
  assign y6275 = n18278 ;
  assign y6276 = n18281 ;
  assign y6277 = ~1'b0 ;
  assign y6278 = n18283 ;
  assign y6279 = n18285 ;
  assign y6280 = n18286 ;
  assign y6281 = n18287 ;
  assign y6282 = n18289 ;
  assign y6283 = ~1'b0 ;
  assign y6284 = ~n18292 ;
  assign y6285 = ~n18299 ;
  assign y6286 = n18301 ;
  assign y6287 = n18303 ;
  assign y6288 = ~n18305 ;
  assign y6289 = ~1'b0 ;
  assign y6290 = ~n1799 ;
  assign y6291 = ~n18309 ;
  assign y6292 = n18316 ;
  assign y6293 = ~1'b0 ;
  assign y6294 = n18320 ;
  assign y6295 = ~1'b0 ;
  assign y6296 = n18323 ;
  assign y6297 = n18324 ;
  assign y6298 = n18327 ;
  assign y6299 = ~n18328 ;
  assign y6300 = n18331 ;
  assign y6301 = ~1'b0 ;
  assign y6302 = n18332 ;
  assign y6303 = ~n18335 ;
  assign y6304 = ~n18336 ;
  assign y6305 = ~n18337 ;
  assign y6306 = n18341 ;
  assign y6307 = n18342 ;
  assign y6308 = ~n18345 ;
  assign y6309 = n18348 ;
  assign y6310 = ~1'b0 ;
  assign y6311 = n18353 ;
  assign y6312 = ~n18357 ;
  assign y6313 = ~1'b0 ;
  assign y6314 = ~n18361 ;
  assign y6315 = ~n18365 ;
  assign y6316 = ~n18367 ;
  assign y6317 = n18372 ;
  assign y6318 = n18376 ;
  assign y6319 = ~n18378 ;
  assign y6320 = n18380 ;
  assign y6321 = n18383 ;
  assign y6322 = ~n18384 ;
  assign y6323 = ~n18387 ;
  assign y6324 = ~n18388 ;
  assign y6325 = n18390 ;
  assign y6326 = n18397 ;
  assign y6327 = n18398 ;
  assign y6328 = ~n18402 ;
  assign y6329 = ~n18412 ;
  assign y6330 = ~n18413 ;
  assign y6331 = n18414 ;
  assign y6332 = n18418 ;
  assign y6333 = ~1'b0 ;
  assign y6334 = n18420 ;
  assign y6335 = ~n18422 ;
  assign y6336 = ~n10623 ;
  assign y6337 = n18423 ;
  assign y6338 = ~n18424 ;
  assign y6339 = ~n18426 ;
  assign y6340 = n18428 ;
  assign y6341 = ~n18430 ;
  assign y6342 = ~n18433 ;
  assign y6343 = n18436 ;
  assign y6344 = ~n18439 ;
  assign y6345 = n18440 ;
  assign y6346 = n18442 ;
  assign y6347 = n18444 ;
  assign y6348 = ~1'b0 ;
  assign y6349 = n18447 ;
  assign y6350 = ~n18451 ;
  assign y6351 = ~n18452 ;
  assign y6352 = ~1'b0 ;
  assign y6353 = n18454 ;
  assign y6354 = ~n18458 ;
  assign y6355 = ~n18462 ;
  assign y6356 = ~1'b0 ;
  assign y6357 = ~n18463 ;
  assign y6358 = ~n1426 ;
  assign y6359 = ~n18464 ;
  assign y6360 = ~n18465 ;
  assign y6361 = n18467 ;
  assign y6362 = n18469 ;
  assign y6363 = n18481 ;
  assign y6364 = n18487 ;
  assign y6365 = ~n18491 ;
  assign y6366 = ~n18494 ;
  assign y6367 = ~n18497 ;
  assign y6368 = n18498 ;
  assign y6369 = ~1'b0 ;
  assign y6370 = ~1'b0 ;
  assign y6371 = ~1'b0 ;
  assign y6372 = ~n18502 ;
  assign y6373 = n11560 ;
  assign y6374 = n18504 ;
  assign y6375 = ~n18510 ;
  assign y6376 = n18512 ;
  assign y6377 = n18517 ;
  assign y6378 = n18520 ;
  assign y6379 = ~n18523 ;
  assign y6380 = ~n18526 ;
  assign y6381 = n18527 ;
  assign y6382 = n18528 ;
  assign y6383 = ~n18530 ;
  assign y6384 = ~n18533 ;
  assign y6385 = n18536 ;
  assign y6386 = n18537 ;
  assign y6387 = ~n18539 ;
  assign y6388 = n18540 ;
  assign y6389 = n18541 ;
  assign y6390 = ~1'b0 ;
  assign y6391 = ~n18544 ;
  assign y6392 = ~1'b0 ;
  assign y6393 = ~1'b0 ;
  assign y6394 = ~n18546 ;
  assign y6395 = ~n18548 ;
  assign y6396 = ~n18551 ;
  assign y6397 = n18554 ;
  assign y6398 = ~n18560 ;
  assign y6399 = ~1'b0 ;
  assign y6400 = n18562 ;
  assign y6401 = n18564 ;
  assign y6402 = n18566 ;
  assign y6403 = n18571 ;
  assign y6404 = n18572 ;
  assign y6405 = n18574 ;
  assign y6406 = ~n18576 ;
  assign y6407 = n18577 ;
  assign y6408 = n18578 ;
  assign y6409 = n18579 ;
  assign y6410 = ~n18580 ;
  assign y6411 = ~1'b0 ;
  assign y6412 = ~1'b0 ;
  assign y6413 = n18581 ;
  assign y6414 = n16572 ;
  assign y6415 = n18586 ;
  assign y6416 = n18590 ;
  assign y6417 = ~1'b0 ;
  assign y6418 = n18592 ;
  assign y6419 = ~n18594 ;
  assign y6420 = n18595 ;
  assign y6421 = ~n18598 ;
  assign y6422 = n18602 ;
  assign y6423 = ~n18609 ;
  assign y6424 = n18611 ;
  assign y6425 = ~n18613 ;
  assign y6426 = n18614 ;
  assign y6427 = n18618 ;
  assign y6428 = ~n18620 ;
  assign y6429 = n18622 ;
  assign y6430 = ~n18625 ;
  assign y6431 = ~n18626 ;
  assign y6432 = n18629 ;
  assign y6433 = n18632 ;
  assign y6434 = ~1'b0 ;
  assign y6435 = ~1'b0 ;
  assign y6436 = n18635 ;
  assign y6437 = ~n18641 ;
  assign y6438 = ~n18642 ;
  assign y6439 = n18643 ;
  assign y6440 = n18646 ;
  assign y6441 = n18653 ;
  assign y6442 = ~1'b0 ;
  assign y6443 = ~n18656 ;
  assign y6444 = ~n18657 ;
  assign y6445 = ~n18663 ;
  assign y6446 = n18671 ;
  assign y6447 = ~1'b0 ;
  assign y6448 = ~n18674 ;
  assign y6449 = ~n18675 ;
  assign y6450 = ~n18680 ;
  assign y6451 = ~1'b0 ;
  assign y6452 = ~n18684 ;
  assign y6453 = ~n18690 ;
  assign y6454 = ~n18695 ;
  assign y6455 = n18697 ;
  assign y6456 = ~1'b0 ;
  assign y6457 = ~n18700 ;
  assign y6458 = n18702 ;
  assign y6459 = n18705 ;
  assign y6460 = ~n18707 ;
  assign y6461 = n18715 ;
  assign y6462 = n18721 ;
  assign y6463 = ~1'b0 ;
  assign y6464 = ~n18722 ;
  assign y6465 = ~n18725 ;
  assign y6466 = ~n18726 ;
  assign y6467 = n18731 ;
  assign y6468 = ~n18734 ;
  assign y6469 = ~1'b0 ;
  assign y6470 = ~n18737 ;
  assign y6471 = n18740 ;
  assign y6472 = ~n18750 ;
  assign y6473 = ~n18754 ;
  assign y6474 = ~1'b0 ;
  assign y6475 = 1'b0 ;
  assign y6476 = ~1'b0 ;
  assign y6477 = ~n18758 ;
  assign y6478 = n18759 ;
  assign y6479 = ~n18760 ;
  assign y6480 = ~1'b0 ;
  assign y6481 = n18765 ;
  assign y6482 = ~1'b0 ;
  assign y6483 = ~n18766 ;
  assign y6484 = ~n18767 ;
  assign y6485 = ~n18771 ;
  assign y6486 = n18772 ;
  assign y6487 = ~1'b0 ;
  assign y6488 = n18774 ;
  assign y6489 = ~1'b0 ;
  assign y6490 = n18775 ;
  assign y6491 = n18777 ;
  assign y6492 = n18789 ;
  assign y6493 = n18792 ;
  assign y6494 = n18796 ;
  assign y6495 = ~n18800 ;
  assign y6496 = n18802 ;
  assign y6497 = ~n18803 ;
  assign y6498 = ~1'b0 ;
  assign y6499 = ~n18807 ;
  assign y6500 = ~n18808 ;
  assign y6501 = ~n17707 ;
  assign y6502 = n18813 ;
  assign y6503 = ~1'b0 ;
  assign y6504 = ~n18816 ;
  assign y6505 = ~1'b0 ;
  assign y6506 = n18822 ;
  assign y6507 = ~n18826 ;
  assign y6508 = ~1'b0 ;
  assign y6509 = ~n18830 ;
  assign y6510 = ~n18833 ;
  assign y6511 = ~1'b0 ;
  assign y6512 = n18836 ;
  assign y6513 = ~n18840 ;
  assign y6514 = ~1'b0 ;
  assign y6515 = ~1'b0 ;
  assign y6516 = n18842 ;
  assign y6517 = n18847 ;
  assign y6518 = n18851 ;
  assign y6519 = ~n18853 ;
  assign y6520 = n18858 ;
  assign y6521 = ~n18863 ;
  assign y6522 = ~n13222 ;
  assign y6523 = ~1'b0 ;
  assign y6524 = ~n18865 ;
  assign y6525 = n18867 ;
  assign y6526 = n18869 ;
  assign y6527 = ~n18870 ;
  assign y6528 = ~n18871 ;
  assign y6529 = n18872 ;
  assign y6530 = n18878 ;
  assign y6531 = ~n18880 ;
  assign y6532 = ~1'b0 ;
  assign y6533 = ~1'b0 ;
  assign y6534 = ~n18889 ;
  assign y6535 = n18890 ;
  assign y6536 = n18892 ;
  assign y6537 = n18893 ;
  assign y6538 = n4180 ;
  assign y6539 = n18897 ;
  assign y6540 = ~1'b0 ;
  assign y6541 = ~1'b0 ;
  assign y6542 = n18903 ;
  assign y6543 = ~n17497 ;
  assign y6544 = ~n18908 ;
  assign y6545 = ~1'b0 ;
  assign y6546 = ~n18910 ;
  assign y6547 = ~n18911 ;
  assign y6548 = ~n18918 ;
  assign y6549 = ~1'b0 ;
  assign y6550 = n18921 ;
  assign y6551 = n18924 ;
  assign y6552 = ~n18928 ;
  assign y6553 = ~n18932 ;
  assign y6554 = n18934 ;
  assign y6555 = ~1'b0 ;
  assign y6556 = n18937 ;
  assign y6557 = n18942 ;
  assign y6558 = ~n18943 ;
  assign y6559 = ~n18944 ;
  assign y6560 = ~1'b0 ;
  assign y6561 = n18954 ;
  assign y6562 = n18955 ;
  assign y6563 = ~n14863 ;
  assign y6564 = ~n18958 ;
  assign y6565 = ~1'b0 ;
  assign y6566 = ~n18960 ;
  assign y6567 = ~n18964 ;
  assign y6568 = n18967 ;
  assign y6569 = ~n18970 ;
  assign y6570 = n18973 ;
  assign y6571 = ~n18977 ;
  assign y6572 = ~n18980 ;
  assign y6573 = n18983 ;
  assign y6574 = n18985 ;
  assign y6575 = ~1'b0 ;
  assign y6576 = n18986 ;
  assign y6577 = n18988 ;
  assign y6578 = n18991 ;
  assign y6579 = n18992 ;
  assign y6580 = n18994 ;
  assign y6581 = ~1'b0 ;
  assign y6582 = ~1'b0 ;
  assign y6583 = ~n18995 ;
  assign y6584 = ~n18996 ;
  assign y6585 = ~n19000 ;
  assign y6586 = ~1'b0 ;
  assign y6587 = n19003 ;
  assign y6588 = ~1'b0 ;
  assign y6589 = ~n19006 ;
  assign y6590 = ~n19009 ;
  assign y6591 = ~1'b0 ;
  assign y6592 = n19010 ;
  assign y6593 = ~n19015 ;
  assign y6594 = ~n19025 ;
  assign y6595 = ~n19027 ;
  assign y6596 = n19029 ;
  assign y6597 = n19033 ;
  assign y6598 = n19035 ;
  assign y6599 = n19037 ;
  assign y6600 = ~n19038 ;
  assign y6601 = ~n19040 ;
  assign y6602 = ~1'b0 ;
  assign y6603 = ~n19043 ;
  assign y6604 = n19044 ;
  assign y6605 = ~n19045 ;
  assign y6606 = ~n19050 ;
  assign y6607 = ~1'b0 ;
  assign y6608 = n19053 ;
  assign y6609 = n19055 ;
  assign y6610 = ~n19057 ;
  assign y6611 = ~n19062 ;
  assign y6612 = ~n19067 ;
  assign y6613 = ~n19068 ;
  assign y6614 = ~1'b0 ;
  assign y6615 = ~1'b0 ;
  assign y6616 = n19070 ;
  assign y6617 = ~n19071 ;
  assign y6618 = n19081 ;
  assign y6619 = ~n19083 ;
  assign y6620 = n19085 ;
  assign y6621 = ~n19087 ;
  assign y6622 = n19089 ;
  assign y6623 = n19090 ;
  assign y6624 = ~n19092 ;
  assign y6625 = ~1'b0 ;
  assign y6626 = ~1'b0 ;
  assign y6627 = ~n19098 ;
  assign y6628 = ~n19103 ;
  assign y6629 = n19104 ;
  assign y6630 = ~1'b0 ;
  assign y6631 = ~1'b0 ;
  assign y6632 = ~n19108 ;
  assign y6633 = ~n19109 ;
  assign y6634 = n19114 ;
  assign y6635 = ~1'b0 ;
  assign y6636 = n19119 ;
  assign y6637 = n19121 ;
  assign y6638 = n19124 ;
  assign y6639 = ~1'b0 ;
  assign y6640 = n19125 ;
  assign y6641 = n19127 ;
  assign y6642 = n4578 ;
  assign y6643 = n19133 ;
  assign y6644 = n19134 ;
  assign y6645 = n19143 ;
  assign y6646 = n19149 ;
  assign y6647 = ~1'b0 ;
  assign y6648 = n19150 ;
  assign y6649 = ~n19151 ;
  assign y6650 = ~n19152 ;
  assign y6651 = n19153 ;
  assign y6652 = n19155 ;
  assign y6653 = ~n19158 ;
  assign y6654 = n19160 ;
  assign y6655 = ~n19164 ;
  assign y6656 = n19167 ;
  assign y6657 = ~n19168 ;
  assign y6658 = ~n19170 ;
  assign y6659 = n19171 ;
  assign y6660 = ~n19172 ;
  assign y6661 = ~n19176 ;
  assign y6662 = ~n19182 ;
  assign y6663 = ~1'b0 ;
  assign y6664 = n19183 ;
  assign y6665 = n10451 ;
  assign y6666 = n19185 ;
  assign y6667 = n19186 ;
  assign y6668 = ~n19190 ;
  assign y6669 = ~1'b0 ;
  assign y6670 = 1'b0 ;
  assign y6671 = n19196 ;
  assign y6672 = n19197 ;
  assign y6673 = n19201 ;
  assign y6674 = n19202 ;
  assign y6675 = n19203 ;
  assign y6676 = ~1'b0 ;
  assign y6677 = ~1'b0 ;
  assign y6678 = ~n19204 ;
  assign y6679 = ~n19210 ;
  assign y6680 = ~n19212 ;
  assign y6681 = n19213 ;
  assign y6682 = ~n19215 ;
  assign y6683 = ~1'b0 ;
  assign y6684 = ~1'b0 ;
  assign y6685 = ~1'b0 ;
  assign y6686 = ~n19218 ;
  assign y6687 = n19219 ;
  assign y6688 = ~n14893 ;
  assign y6689 = ~n19221 ;
  assign y6690 = ~1'b0 ;
  assign y6691 = n19223 ;
  assign y6692 = ~1'b0 ;
  assign y6693 = ~1'b0 ;
  assign y6694 = ~n19224 ;
  assign y6695 = n19225 ;
  assign y6696 = n19230 ;
  assign y6697 = ~1'b0 ;
  assign y6698 = ~1'b0 ;
  assign y6699 = ~n19232 ;
  assign y6700 = ~n19233 ;
  assign y6701 = ~n19236 ;
  assign y6702 = ~n19239 ;
  assign y6703 = n19246 ;
  assign y6704 = n19251 ;
  assign y6705 = ~1'b0 ;
  assign y6706 = ~n19252 ;
  assign y6707 = n19254 ;
  assign y6708 = ~n19255 ;
  assign y6709 = n19257 ;
  assign y6710 = ~1'b0 ;
  assign y6711 = ~1'b0 ;
  assign y6712 = ~n19259 ;
  assign y6713 = n19260 ;
  assign y6714 = n19261 ;
  assign y6715 = ~n19268 ;
  assign y6716 = n19270 ;
  assign y6717 = ~n19271 ;
  assign y6718 = ~n19272 ;
  assign y6719 = ~n19275 ;
  assign y6720 = n19280 ;
  assign y6721 = ~1'b0 ;
  assign y6722 = ~n19285 ;
  assign y6723 = n19289 ;
  assign y6724 = n19292 ;
  assign y6725 = n19295 ;
  assign y6726 = ~n19299 ;
  assign y6727 = ~n19302 ;
  assign y6728 = n4073 ;
  assign y6729 = ~n19307 ;
  assign y6730 = ~1'b0 ;
  assign y6731 = n19308 ;
  assign y6732 = ~n19310 ;
  assign y6733 = ~n19312 ;
  assign y6734 = ~n19314 ;
  assign y6735 = ~n19318 ;
  assign y6736 = ~n19320 ;
  assign y6737 = ~n19324 ;
  assign y6738 = n19325 ;
  assign y6739 = n19327 ;
  assign y6740 = ~n19330 ;
  assign y6741 = ~n19333 ;
  assign y6742 = ~1'b0 ;
  assign y6743 = ~1'b0 ;
  assign y6744 = ~1'b0 ;
  assign y6745 = ~n19336 ;
  assign y6746 = ~n19338 ;
  assign y6747 = ~1'b0 ;
  assign y6748 = n19340 ;
  assign y6749 = ~n19345 ;
  assign y6750 = ~n19346 ;
  assign y6751 = n19347 ;
  assign y6752 = ~n19354 ;
  assign y6753 = n19356 ;
  assign y6754 = ~n19360 ;
  assign y6755 = ~n19362 ;
  assign y6756 = ~n19364 ;
  assign y6757 = n19365 ;
  assign y6758 = n19373 ;
  assign y6759 = n19374 ;
  assign y6760 = n19376 ;
  assign y6761 = ~n19377 ;
  assign y6762 = ~n19378 ;
  assign y6763 = n19379 ;
  assign y6764 = ~n19382 ;
  assign y6765 = n19391 ;
  assign y6766 = n19396 ;
  assign y6767 = ~1'b0 ;
  assign y6768 = n19397 ;
  assign y6769 = ~n19399 ;
  assign y6770 = ~1'b0 ;
  assign y6771 = ~n19402 ;
  assign y6772 = ~n19407 ;
  assign y6773 = n19412 ;
  assign y6774 = n19413 ;
  assign y6775 = ~1'b0 ;
  assign y6776 = n19418 ;
  assign y6777 = ~n19421 ;
  assign y6778 = n19422 ;
  assign y6779 = n19424 ;
  assign y6780 = ~n19426 ;
  assign y6781 = n19431 ;
  assign y6782 = n19437 ;
  assign y6783 = ~1'b0 ;
  assign y6784 = n19438 ;
  assign y6785 = ~n19447 ;
  assign y6786 = ~1'b0 ;
  assign y6787 = n19451 ;
  assign y6788 = ~n19453 ;
  assign y6789 = ~n19456 ;
  assign y6790 = ~1'b0 ;
  assign y6791 = ~1'b0 ;
  assign y6792 = ~n19457 ;
  assign y6793 = ~n19465 ;
  assign y6794 = n19466 ;
  assign y6795 = n19467 ;
  assign y6796 = n19470 ;
  assign y6797 = ~n19479 ;
  assign y6798 = ~n19483 ;
  assign y6799 = ~n19484 ;
  assign y6800 = ~n19486 ;
  assign y6801 = ~n19494 ;
  assign y6802 = ~n19497 ;
  assign y6803 = n19500 ;
  assign y6804 = ~n19509 ;
  assign y6805 = n19511 ;
  assign y6806 = ~n19514 ;
  assign y6807 = ~n19519 ;
  assign y6808 = ~1'b0 ;
  assign y6809 = ~1'b0 ;
  assign y6810 = ~1'b0 ;
  assign y6811 = ~n19520 ;
  assign y6812 = ~n19521 ;
  assign y6813 = ~1'b0 ;
  assign y6814 = ~n19523 ;
  assign y6815 = n19526 ;
  assign y6816 = n19528 ;
  assign y6817 = ~n19539 ;
  assign y6818 = ~n19541 ;
  assign y6819 = ~n19547 ;
  assign y6820 = ~n19549 ;
  assign y6821 = n19550 ;
  assign y6822 = ~n19555 ;
  assign y6823 = 1'b0 ;
  assign y6824 = ~n19559 ;
  assign y6825 = ~n19564 ;
  assign y6826 = ~n19565 ;
  assign y6827 = ~1'b0 ;
  assign y6828 = ~1'b0 ;
  assign y6829 = ~1'b0 ;
  assign y6830 = n19573 ;
  assign y6831 = n19576 ;
  assign y6832 = ~n19584 ;
  assign y6833 = ~n19586 ;
  assign y6834 = ~1'b0 ;
  assign y6835 = ~n19587 ;
  assign y6836 = n19591 ;
  assign y6837 = n19595 ;
  assign y6838 = ~n19596 ;
  assign y6839 = n19598 ;
  assign y6840 = n19599 ;
  assign y6841 = ~n19603 ;
  assign y6842 = ~1'b0 ;
  assign y6843 = ~n19606 ;
  assign y6844 = n19607 ;
  assign y6845 = ~n19610 ;
  assign y6846 = ~1'b0 ;
  assign y6847 = ~n14903 ;
  assign y6848 = ~1'b0 ;
  assign y6849 = ~n19612 ;
  assign y6850 = ~n19613 ;
  assign y6851 = ~n19618 ;
  assign y6852 = ~n19619 ;
  assign y6853 = ~n19620 ;
  assign y6854 = n19623 ;
  assign y6855 = ~1'b0 ;
  assign y6856 = ~n19626 ;
  assign y6857 = n19628 ;
  assign y6858 = n19630 ;
  assign y6859 = n19634 ;
  assign y6860 = ~n19637 ;
  assign y6861 = n19640 ;
  assign y6862 = n19641 ;
  assign y6863 = ~1'b0 ;
  assign y6864 = ~n19643 ;
  assign y6865 = ~n19646 ;
  assign y6866 = n19650 ;
  assign y6867 = ~1'b0 ;
  assign y6868 = ~n19654 ;
  assign y6869 = n19658 ;
  assign y6870 = ~1'b0 ;
  assign y6871 = n19660 ;
  assign y6872 = ~n19661 ;
  assign y6873 = ~n19662 ;
  assign y6874 = n19663 ;
  assign y6875 = n19673 ;
  assign y6876 = n19674 ;
  assign y6877 = ~n19676 ;
  assign y6878 = ~n19678 ;
  assign y6879 = ~n19679 ;
  assign y6880 = ~n19680 ;
  assign y6881 = n19681 ;
  assign y6882 = n19683 ;
  assign y6883 = ~1'b0 ;
  assign y6884 = ~n19685 ;
  assign y6885 = ~n19688 ;
  assign y6886 = n19692 ;
  assign y6887 = n19693 ;
  assign y6888 = ~n19694 ;
  assign y6889 = n19696 ;
  assign y6890 = n19701 ;
  assign y6891 = ~1'b0 ;
  assign y6892 = n19706 ;
  assign y6893 = ~n19713 ;
  assign y6894 = n19715 ;
  assign y6895 = n19716 ;
  assign y6896 = ~n19717 ;
  assign y6897 = ~n19720 ;
  assign y6898 = ~n19721 ;
  assign y6899 = n19722 ;
  assign y6900 = n19726 ;
  assign y6901 = ~1'b0 ;
  assign y6902 = n19728 ;
  assign y6903 = n19737 ;
  assign y6904 = ~n19738 ;
  assign y6905 = ~1'b0 ;
  assign y6906 = n19746 ;
  assign y6907 = ~n19748 ;
  assign y6908 = n19749 ;
  assign y6909 = n19752 ;
  assign y6910 = ~n19756 ;
  assign y6911 = ~n19759 ;
  assign y6912 = ~1'b0 ;
  assign y6913 = n19762 ;
  assign y6914 = ~1'b0 ;
  assign y6915 = n19770 ;
  assign y6916 = n19771 ;
  assign y6917 = n19773 ;
  assign y6918 = ~1'b0 ;
  assign y6919 = n19774 ;
  assign y6920 = n19775 ;
  assign y6921 = ~n19778 ;
  assign y6922 = n19781 ;
  assign y6923 = n19782 ;
  assign y6924 = ~n19784 ;
  assign y6925 = ~n19786 ;
  assign y6926 = ~n19789 ;
  assign y6927 = ~n19800 ;
  assign y6928 = n19802 ;
  assign y6929 = n19804 ;
  assign y6930 = n946 ;
  assign y6931 = n19807 ;
  assign y6932 = n19808 ;
  assign y6933 = ~n19810 ;
  assign y6934 = ~n19813 ;
  assign y6935 = ~n19817 ;
  assign y6936 = n19820 ;
  assign y6937 = n19823 ;
  assign y6938 = ~n19826 ;
  assign y6939 = ~n19827 ;
  assign y6940 = n19828 ;
  assign y6941 = n19830 ;
  assign y6942 = ~n19832 ;
  assign y6943 = ~n19839 ;
  assign y6944 = ~n8135 ;
  assign y6945 = n19844 ;
  assign y6946 = n972 ;
  assign y6947 = n19851 ;
  assign y6948 = ~n19853 ;
  assign y6949 = n19856 ;
  assign y6950 = n19859 ;
  assign y6951 = n19861 ;
  assign y6952 = ~n19863 ;
  assign y6953 = ~n19868 ;
  assign y6954 = ~1'b0 ;
  assign y6955 = ~n19869 ;
  assign y6956 = ~n19874 ;
  assign y6957 = ~n19882 ;
  assign y6958 = n19893 ;
  assign y6959 = ~n19896 ;
  assign y6960 = ~n19900 ;
  assign y6961 = n19906 ;
  assign y6962 = ~1'b0 ;
  assign y6963 = n19910 ;
  assign y6964 = n19914 ;
  assign y6965 = ~n1209 ;
  assign y6966 = ~n19916 ;
  assign y6967 = n19918 ;
  assign y6968 = n19921 ;
  assign y6969 = ~n19923 ;
  assign y6970 = ~1'b0 ;
  assign y6971 = n19926 ;
  assign y6972 = ~1'b0 ;
  assign y6973 = ~1'b0 ;
  assign y6974 = ~1'b0 ;
  assign y6975 = ~1'b0 ;
  assign y6976 = ~n19928 ;
  assign y6977 = ~n8822 ;
  assign y6978 = n19930 ;
  assign y6979 = ~n19933 ;
  assign y6980 = ~1'b0 ;
  assign y6981 = ~n19936 ;
  assign y6982 = n19941 ;
  assign y6983 = ~n19942 ;
  assign y6984 = ~n19947 ;
  assign y6985 = ~n19948 ;
  assign y6986 = n19949 ;
  assign y6987 = n19952 ;
  assign y6988 = ~n19958 ;
  assign y6989 = ~n19960 ;
  assign y6990 = ~n19969 ;
  assign y6991 = ~n11245 ;
  assign y6992 = ~n19972 ;
  assign y6993 = n19974 ;
  assign y6994 = ~n19975 ;
  assign y6995 = n19976 ;
  assign y6996 = ~n19977 ;
  assign y6997 = ~1'b0 ;
  assign y6998 = ~n19980 ;
  assign y6999 = n19982 ;
  assign y7000 = ~n19984 ;
  assign y7001 = ~n19987 ;
  assign y7002 = n19994 ;
  assign y7003 = ~n19995 ;
  assign y7004 = n20000 ;
  assign y7005 = ~n20006 ;
  assign y7006 = ~1'b0 ;
  assign y7007 = ~1'b0 ;
  assign y7008 = ~1'b0 ;
  assign y7009 = n20007 ;
  assign y7010 = ~n20010 ;
  assign y7011 = ~n20011 ;
  assign y7012 = ~n20013 ;
  assign y7013 = ~1'b0 ;
  assign y7014 = n17245 ;
  assign y7015 = n20026 ;
  assign y7016 = n20029 ;
  assign y7017 = n20032 ;
  assign y7018 = n20035 ;
  assign y7019 = ~n20036 ;
  assign y7020 = ~n20039 ;
  assign y7021 = n20047 ;
  assign y7022 = ~n20049 ;
  assign y7023 = ~n20062 ;
  assign y7024 = ~n20063 ;
  assign y7025 = ~n20069 ;
  assign y7026 = n20077 ;
  assign y7027 = ~n20082 ;
  assign y7028 = n20084 ;
  assign y7029 = ~n20085 ;
  assign y7030 = 1'b0 ;
  assign y7031 = ~n20089 ;
  assign y7032 = ~n20090 ;
  assign y7033 = n20098 ;
  assign y7034 = n20102 ;
  assign y7035 = ~n20106 ;
  assign y7036 = ~n20107 ;
  assign y7037 = ~1'b0 ;
  assign y7038 = n20110 ;
  assign y7039 = ~n20114 ;
  assign y7040 = ~n20117 ;
  assign y7041 = n20121 ;
  assign y7042 = ~n20123 ;
  assign y7043 = ~1'b0 ;
  assign y7044 = ~n20124 ;
  assign y7045 = n20125 ;
  assign y7046 = n20129 ;
  assign y7047 = ~n20135 ;
  assign y7048 = ~n20138 ;
  assign y7049 = n8582 ;
  assign y7050 = ~1'b0 ;
  assign y7051 = ~n20139 ;
  assign y7052 = ~n20145 ;
  assign y7053 = ~n20147 ;
  assign y7054 = ~n20148 ;
  assign y7055 = ~n20154 ;
  assign y7056 = n20155 ;
  assign y7057 = 1'b0 ;
  assign y7058 = ~1'b0 ;
  assign y7059 = n20156 ;
  assign y7060 = ~n20157 ;
  assign y7061 = n20159 ;
  assign y7062 = ~1'b0 ;
  assign y7063 = ~1'b0 ;
  assign y7064 = ~1'b0 ;
  assign y7065 = ~n20163 ;
  assign y7066 = ~n12039 ;
  assign y7067 = n20164 ;
  assign y7068 = n20174 ;
  assign y7069 = ~n20178 ;
  assign y7070 = ~n20179 ;
  assign y7071 = ~n20183 ;
  assign y7072 = ~n20184 ;
  assign y7073 = ~n20193 ;
  assign y7074 = ~n20196 ;
  assign y7075 = ~1'b0 ;
  assign y7076 = n20199 ;
  assign y7077 = n20202 ;
  assign y7078 = ~1'b0 ;
  assign y7079 = ~1'b0 ;
  assign y7080 = ~n20203 ;
  assign y7081 = ~1'b0 ;
  assign y7082 = n20205 ;
  assign y7083 = ~n20207 ;
  assign y7084 = ~n20209 ;
  assign y7085 = n20210 ;
  assign y7086 = n20211 ;
  assign y7087 = ~n20215 ;
  assign y7088 = n20220 ;
  assign y7089 = ~1'b0 ;
  assign y7090 = ~1'b0 ;
  assign y7091 = n7684 ;
  assign y7092 = n20221 ;
  assign y7093 = ~n20224 ;
  assign y7094 = ~1'b0 ;
  assign y7095 = ~1'b0 ;
  assign y7096 = n20229 ;
  assign y7097 = ~x79 ;
  assign y7098 = ~1'b0 ;
  assign y7099 = ~n20236 ;
  assign y7100 = ~1'b0 ;
  assign y7101 = n20239 ;
  assign y7102 = n20241 ;
  assign y7103 = n20245 ;
  assign y7104 = ~n20249 ;
  assign y7105 = n20255 ;
  assign y7106 = ~n20257 ;
  assign y7107 = n20259 ;
  assign y7108 = n20266 ;
  assign y7109 = ~n20270 ;
  assign y7110 = ~n20273 ;
  assign y7111 = ~n20276 ;
  assign y7112 = n20277 ;
  assign y7113 = ~n20282 ;
  assign y7114 = ~1'b0 ;
  assign y7115 = ~n20283 ;
  assign y7116 = ~n20285 ;
  assign y7117 = n20287 ;
  assign y7118 = ~n14523 ;
  assign y7119 = ~n20288 ;
  assign y7120 = n20289 ;
  assign y7121 = ~n20290 ;
  assign y7122 = n20291 ;
  assign y7123 = ~1'b0 ;
  assign y7124 = ~n20293 ;
  assign y7125 = ~n20295 ;
  assign y7126 = ~n20298 ;
  assign y7127 = ~n20299 ;
  assign y7128 = n20303 ;
  assign y7129 = ~1'b0 ;
  assign y7130 = ~1'b0 ;
  assign y7131 = ~1'b0 ;
  assign y7132 = ~n20304 ;
  assign y7133 = n20306 ;
  assign y7134 = n20310 ;
  assign y7135 = ~n20311 ;
  assign y7136 = n20314 ;
  assign y7137 = n20317 ;
  assign y7138 = n20319 ;
  assign y7139 = n17527 ;
  assign y7140 = ~n20320 ;
  assign y7141 = ~1'b0 ;
  assign y7142 = ~1'b0 ;
  assign y7143 = ~1'b0 ;
  assign y7144 = ~1'b0 ;
  assign y7145 = n20323 ;
  assign y7146 = n20324 ;
  assign y7147 = n7409 ;
  assign y7148 = ~n20326 ;
  assign y7149 = n20328 ;
  assign y7150 = ~n20332 ;
  assign y7151 = ~n20333 ;
  assign y7152 = ~1'b0 ;
  assign y7153 = ~n20334 ;
  assign y7154 = n20342 ;
  assign y7155 = ~1'b0 ;
  assign y7156 = n20348 ;
  assign y7157 = ~n20349 ;
  assign y7158 = n20351 ;
  assign y7159 = ~n20359 ;
  assign y7160 = n20361 ;
  assign y7161 = n20363 ;
  assign y7162 = ~1'b0 ;
  assign y7163 = ~n20365 ;
  assign y7164 = n20370 ;
  assign y7165 = ~1'b0 ;
  assign y7166 = ~n20379 ;
  assign y7167 = ~1'b0 ;
  assign y7168 = ~n20381 ;
  assign y7169 = n20387 ;
  assign y7170 = ~n20389 ;
  assign y7171 = n20390 ;
  assign y7172 = ~n20396 ;
  assign y7173 = n20398 ;
  assign y7174 = ~n20399 ;
  assign y7175 = ~n20400 ;
  assign y7176 = n20403 ;
  assign y7177 = ~n20404 ;
  assign y7178 = n20406 ;
  assign y7179 = ~n20411 ;
  assign y7180 = 1'b0 ;
  assign y7181 = ~1'b0 ;
  assign y7182 = ~n20412 ;
  assign y7183 = ~n20413 ;
  assign y7184 = n20414 ;
  assign y7185 = ~n20419 ;
  assign y7186 = ~1'b0 ;
  assign y7187 = n20421 ;
  assign y7188 = ~1'b0 ;
  assign y7189 = n20423 ;
  assign y7190 = n20424 ;
  assign y7191 = n20426 ;
  assign y7192 = ~n20427 ;
  assign y7193 = ~n20431 ;
  assign y7194 = ~n20439 ;
  assign y7195 = n20443 ;
  assign y7196 = ~n20446 ;
  assign y7197 = ~1'b0 ;
  assign y7198 = ~1'b0 ;
  assign y7199 = n20447 ;
  assign y7200 = n20448 ;
  assign y7201 = n20453 ;
  assign y7202 = ~n20454 ;
  assign y7203 = n20456 ;
  assign y7204 = ~n20459 ;
  assign y7205 = n20466 ;
  assign y7206 = ~1'b0 ;
  assign y7207 = n20469 ;
  assign y7208 = ~n20471 ;
  assign y7209 = n20473 ;
  assign y7210 = ~n20475 ;
  assign y7211 = ~1'b0 ;
  assign y7212 = ~n20478 ;
  assign y7213 = ~n20481 ;
  assign y7214 = ~n20483 ;
  assign y7215 = ~n20487 ;
  assign y7216 = n20489 ;
  assign y7217 = ~n20493 ;
  assign y7218 = n20496 ;
  assign y7219 = ~1'b0 ;
  assign y7220 = n20497 ;
  assign y7221 = ~n20500 ;
  assign y7222 = ~n20502 ;
  assign y7223 = n20509 ;
  assign y7224 = ~1'b0 ;
  assign y7225 = n20513 ;
  assign y7226 = n20515 ;
  assign y7227 = n20518 ;
  assign y7228 = n20522 ;
  assign y7229 = n20529 ;
  assign y7230 = ~n20532 ;
  assign y7231 = ~n20535 ;
  assign y7232 = ~n20540 ;
  assign y7233 = ~1'b0 ;
  assign y7234 = n20542 ;
  assign y7235 = ~n20549 ;
  assign y7236 = ~n20553 ;
  assign y7237 = ~n20555 ;
  assign y7238 = ~n20557 ;
  assign y7239 = ~1'b0 ;
  assign y7240 = n20558 ;
  assign y7241 = ~n20569 ;
  assign y7242 = ~n3259 ;
  assign y7243 = ~n20573 ;
  assign y7244 = ~1'b0 ;
  assign y7245 = n20576 ;
  assign y7246 = ~1'b0 ;
  assign y7247 = ~n20577 ;
  assign y7248 = n20578 ;
  assign y7249 = ~n20579 ;
  assign y7250 = ~n20588 ;
  assign y7251 = n20592 ;
  assign y7252 = ~1'b0 ;
  assign y7253 = ~n20594 ;
  assign y7254 = n20599 ;
  assign y7255 = n20602 ;
  assign y7256 = ~n20617 ;
  assign y7257 = ~n20619 ;
  assign y7258 = n20620 ;
  assign y7259 = n14084 ;
  assign y7260 = ~n20622 ;
  assign y7261 = ~1'b0 ;
  assign y7262 = ~n20624 ;
  assign y7263 = ~n20626 ;
  assign y7264 = n20627 ;
  assign y7265 = n20628 ;
  assign y7266 = ~1'b0 ;
  assign y7267 = n20631 ;
  assign y7268 = n20632 ;
  assign y7269 = ~n20635 ;
  assign y7270 = ~n20638 ;
  assign y7271 = n20640 ;
  assign y7272 = ~n20642 ;
  assign y7273 = n20643 ;
  assign y7274 = ~n10448 ;
  assign y7275 = n20647 ;
  assign y7276 = ~n20649 ;
  assign y7277 = n20650 ;
  assign y7278 = n20653 ;
  assign y7279 = n20654 ;
  assign y7280 = n20655 ;
  assign y7281 = ~1'b0 ;
  assign y7282 = ~n20659 ;
  assign y7283 = n20660 ;
  assign y7284 = ~n20661 ;
  assign y7285 = ~n20662 ;
  assign y7286 = ~n20666 ;
  assign y7287 = ~n20668 ;
  assign y7288 = ~n20671 ;
  assign y7289 = n20673 ;
  assign y7290 = ~n20675 ;
  assign y7291 = n20678 ;
  assign y7292 = ~1'b0 ;
  assign y7293 = ~n20679 ;
  assign y7294 = ~n20680 ;
  assign y7295 = ~n20681 ;
  assign y7296 = n20682 ;
  assign y7297 = n20685 ;
  assign y7298 = n20688 ;
  assign y7299 = ~1'b0 ;
  assign y7300 = ~1'b0 ;
  assign y7301 = n20689 ;
  assign y7302 = n20690 ;
  assign y7303 = ~n20691 ;
  assign y7304 = n20694 ;
  assign y7305 = ~n20696 ;
  assign y7306 = ~1'b0 ;
  assign y7307 = n20699 ;
  assign y7308 = ~n20700 ;
  assign y7309 = n20703 ;
  assign y7310 = ~n20705 ;
  assign y7311 = ~n20706 ;
  assign y7312 = ~1'b0 ;
  assign y7313 = n20708 ;
  assign y7314 = ~1'b0 ;
  assign y7315 = n20715 ;
  assign y7316 = n20722 ;
  assign y7317 = n20726 ;
  assign y7318 = ~1'b0 ;
  assign y7319 = ~1'b0 ;
  assign y7320 = ~1'b0 ;
  assign y7321 = ~1'b0 ;
  assign y7322 = ~1'b0 ;
  assign y7323 = n20730 ;
  assign y7324 = ~n20731 ;
  assign y7325 = ~n20734 ;
  assign y7326 = n20736 ;
  assign y7327 = n20738 ;
  assign y7328 = n20740 ;
  assign y7329 = ~n20741 ;
  assign y7330 = n20743 ;
  assign y7331 = ~n20746 ;
  assign y7332 = ~n20748 ;
  assign y7333 = ~n20750 ;
  assign y7334 = ~1'b0 ;
  assign y7335 = n20751 ;
  assign y7336 = ~n20752 ;
  assign y7337 = n20754 ;
  assign y7338 = n20760 ;
  assign y7339 = ~n20762 ;
  assign y7340 = ~n20769 ;
  assign y7341 = n20770 ;
  assign y7342 = n20771 ;
  assign y7343 = ~1'b0 ;
  assign y7344 = n20773 ;
  assign y7345 = ~1'b0 ;
  assign y7346 = ~1'b0 ;
  assign y7347 = 1'b0 ;
  assign y7348 = ~n20774 ;
  assign y7349 = n17803 ;
  assign y7350 = n20776 ;
  assign y7351 = ~n20779 ;
  assign y7352 = ~n20781 ;
  assign y7353 = n20787 ;
  assign y7354 = ~1'b0 ;
  assign y7355 = ~n20789 ;
  assign y7356 = n20790 ;
  assign y7357 = ~n20791 ;
  assign y7358 = n20792 ;
  assign y7359 = ~1'b0 ;
  assign y7360 = ~n20794 ;
  assign y7361 = n20801 ;
  assign y7362 = ~n3295 ;
  assign y7363 = n20802 ;
  assign y7364 = ~n20803 ;
  assign y7365 = n20808 ;
  assign y7366 = ~n20811 ;
  assign y7367 = n20814 ;
  assign y7368 = ~n20816 ;
  assign y7369 = ~n20818 ;
  assign y7370 = ~n20821 ;
  assign y7371 = ~1'b0 ;
  assign y7372 = n20825 ;
  assign y7373 = ~1'b0 ;
  assign y7374 = ~1'b0 ;
  assign y7375 = n20831 ;
  assign y7376 = ~1'b0 ;
  assign y7377 = ~n20833 ;
  assign y7378 = n20835 ;
  assign y7379 = n20837 ;
  assign y7380 = n20839 ;
  assign y7381 = ~1'b0 ;
  assign y7382 = ~n20843 ;
  assign y7383 = n20848 ;
  assign y7384 = ~n20849 ;
  assign y7385 = ~n20852 ;
  assign y7386 = ~1'b0 ;
  assign y7387 = n20858 ;
  assign y7388 = n20859 ;
  assign y7389 = ~n20862 ;
  assign y7390 = n20864 ;
  assign y7391 = ~n20865 ;
  assign y7392 = ~n20878 ;
  assign y7393 = ~n20880 ;
  assign y7394 = n20882 ;
  assign y7395 = ~n20883 ;
  assign y7396 = n20890 ;
  assign y7397 = n20891 ;
  assign y7398 = ~n20892 ;
  assign y7399 = ~n20896 ;
  assign y7400 = ~n20897 ;
  assign y7401 = ~1'b0 ;
  assign y7402 = ~1'b0 ;
  assign y7403 = n20906 ;
  assign y7404 = ~n20909 ;
  assign y7405 = ~n20910 ;
  assign y7406 = n20911 ;
  assign y7407 = ~n20914 ;
  assign y7408 = ~n20919 ;
  assign y7409 = n20920 ;
  assign y7410 = n20921 ;
  assign y7411 = ~n20922 ;
  assign y7412 = ~n20927 ;
  assign y7413 = ~n20931 ;
  assign y7414 = 1'b0 ;
  assign y7415 = ~n20933 ;
  assign y7416 = n20936 ;
  assign y7417 = ~n20941 ;
  assign y7418 = ~1'b0 ;
  assign y7419 = ~1'b0 ;
  assign y7420 = n20942 ;
  assign y7421 = ~n20944 ;
  assign y7422 = n20945 ;
  assign y7423 = n20946 ;
  assign y7424 = n20950 ;
  assign y7425 = ~n20952 ;
  assign y7426 = ~1'b0 ;
  assign y7427 = n7472 ;
  assign y7428 = ~n20956 ;
  assign y7429 = n20959 ;
  assign y7430 = n20960 ;
  assign y7431 = n14353 ;
  assign y7432 = n20964 ;
  assign y7433 = n20967 ;
  assign y7434 = ~n20968 ;
  assign y7435 = ~n20971 ;
  assign y7436 = ~n20975 ;
  assign y7437 = n20983 ;
  assign y7438 = n20985 ;
  assign y7439 = n20990 ;
  assign y7440 = ~n20992 ;
  assign y7441 = n20993 ;
  assign y7442 = ~1'b0 ;
  assign y7443 = n20995 ;
  assign y7444 = ~1'b0 ;
  assign y7445 = ~n20997 ;
  assign y7446 = n20998 ;
  assign y7447 = ~n21003 ;
  assign y7448 = n21007 ;
  assign y7449 = ~1'b0 ;
  assign y7450 = n21008 ;
  assign y7451 = n21009 ;
  assign y7452 = ~n21011 ;
  assign y7453 = ~n21012 ;
  assign y7454 = ~1'b0 ;
  assign y7455 = ~n21016 ;
  assign y7456 = ~n21027 ;
  assign y7457 = ~n7955 ;
  assign y7458 = n21030 ;
  assign y7459 = n21035 ;
  assign y7460 = n21041 ;
  assign y7461 = n21043 ;
  assign y7462 = ~1'b0 ;
  assign y7463 = ~1'b0 ;
  assign y7464 = n21049 ;
  assign y7465 = ~n21051 ;
  assign y7466 = n21056 ;
  assign y7467 = ~1'b0 ;
  assign y7468 = ~1'b0 ;
  assign y7469 = ~n21057 ;
  assign y7470 = n21059 ;
  assign y7471 = n21061 ;
  assign y7472 = ~n21067 ;
  assign y7473 = n21076 ;
  assign y7474 = ~n21079 ;
  assign y7475 = n21085 ;
  assign y7476 = n21087 ;
  assign y7477 = ~n21088 ;
  assign y7478 = ~1'b0 ;
  assign y7479 = ~n21090 ;
  assign y7480 = ~n21092 ;
  assign y7481 = n21093 ;
  assign y7482 = ~n21096 ;
  assign y7483 = n21098 ;
  assign y7484 = ~n21100 ;
  assign y7485 = ~1'b0 ;
  assign y7486 = n21102 ;
  assign y7487 = n21105 ;
  assign y7488 = ~n21107 ;
  assign y7489 = n21108 ;
  assign y7490 = ~n21109 ;
  assign y7491 = ~n21112 ;
  assign y7492 = ~n21119 ;
  assign y7493 = ~1'b0 ;
  assign y7494 = ~1'b0 ;
  assign y7495 = ~n21123 ;
  assign y7496 = n21124 ;
  assign y7497 = n21126 ;
  assign y7498 = ~n21129 ;
  assign y7499 = ~n21132 ;
  assign y7500 = ~n21134 ;
  assign y7501 = n607 ;
  assign y7502 = ~n21137 ;
  assign y7503 = n21138 ;
  assign y7504 = ~n21139 ;
  assign y7505 = ~n21143 ;
  assign y7506 = ~n21145 ;
  assign y7507 = ~n21147 ;
  assign y7508 = ~1'b0 ;
  assign y7509 = ~n21150 ;
  assign y7510 = n21154 ;
  assign y7511 = n8217 ;
  assign y7512 = ~n21157 ;
  assign y7513 = ~n21160 ;
  assign y7514 = n21161 ;
  assign y7515 = n21162 ;
  assign y7516 = n21165 ;
  assign y7517 = n21166 ;
  assign y7518 = ~n21168 ;
  assign y7519 = ~n21169 ;
  assign y7520 = ~n21174 ;
  assign y7521 = ~n21181 ;
  assign y7522 = n21186 ;
  assign y7523 = ~1'b0 ;
  assign y7524 = ~1'b0 ;
  assign y7525 = n21191 ;
  assign y7526 = ~n19084 ;
  assign y7527 = n21192 ;
  assign y7528 = ~n21193 ;
  assign y7529 = ~n21194 ;
  assign y7530 = ~n21195 ;
  assign y7531 = ~1'b0 ;
  assign y7532 = ~n21197 ;
  assign y7533 = n21199 ;
  assign y7534 = ~1'b0 ;
  assign y7535 = ~n21205 ;
  assign y7536 = ~n21209 ;
  assign y7537 = ~n21211 ;
  assign y7538 = n21212 ;
  assign y7539 = n21215 ;
  assign y7540 = ~1'b0 ;
  assign y7541 = n21220 ;
  assign y7542 = ~n21223 ;
  assign y7543 = ~n21230 ;
  assign y7544 = n21237 ;
  assign y7545 = ~1'b0 ;
  assign y7546 = ~n21243 ;
  assign y7547 = ~n21244 ;
  assign y7548 = ~n21247 ;
  assign y7549 = ~n5800 ;
  assign y7550 = ~n21250 ;
  assign y7551 = n21252 ;
  assign y7552 = n21253 ;
  assign y7553 = n21254 ;
  assign y7554 = n21255 ;
  assign y7555 = n21256 ;
  assign y7556 = n21260 ;
  assign y7557 = ~n21264 ;
  assign y7558 = n21265 ;
  assign y7559 = n21267 ;
  assign y7560 = ~n21269 ;
  assign y7561 = ~n21271 ;
  assign y7562 = ~n21275 ;
  assign y7563 = n21279 ;
  assign y7564 = ~n21280 ;
  assign y7565 = n21285 ;
  assign y7566 = ~1'b0 ;
  assign y7567 = ~1'b0 ;
  assign y7568 = ~n21287 ;
  assign y7569 = ~n21289 ;
  assign y7570 = ~n21291 ;
  assign y7571 = n21292 ;
  assign y7572 = n21295 ;
  assign y7573 = ~1'b0 ;
  assign y7574 = n21297 ;
  assign y7575 = ~n21298 ;
  assign y7576 = ~n21299 ;
  assign y7577 = ~n21301 ;
  assign y7578 = n21302 ;
  assign y7579 = n21304 ;
  assign y7580 = ~n21306 ;
  assign y7581 = ~n21307 ;
  assign y7582 = ~1'b0 ;
  assign y7583 = ~n21311 ;
  assign y7584 = n21312 ;
  assign y7585 = n21313 ;
  assign y7586 = ~1'b0 ;
  assign y7587 = ~1'b0 ;
  assign y7588 = ~n21317 ;
  assign y7589 = n21320 ;
  assign y7590 = ~n21321 ;
  assign y7591 = n21323 ;
  assign y7592 = ~n21325 ;
  assign y7593 = n21327 ;
  assign y7594 = 1'b0 ;
  assign y7595 = n21333 ;
  assign y7596 = ~n4179 ;
  assign y7597 = n21335 ;
  assign y7598 = n21337 ;
  assign y7599 = ~1'b0 ;
  assign y7600 = ~n21338 ;
  assign y7601 = n21342 ;
  assign y7602 = n21347 ;
  assign y7603 = n21350 ;
  assign y7604 = n21351 ;
  assign y7605 = n21352 ;
  assign y7606 = ~1'b0 ;
  assign y7607 = n21354 ;
  assign y7608 = ~1'b0 ;
  assign y7609 = n21357 ;
  assign y7610 = n21361 ;
  assign y7611 = ~n21366 ;
  assign y7612 = n21368 ;
  assign y7613 = ~n21370 ;
  assign y7614 = n21372 ;
  assign y7615 = ~1'b0 ;
  assign y7616 = ~1'b0 ;
  assign y7617 = n21376 ;
  assign y7618 = ~n21377 ;
  assign y7619 = n21383 ;
  assign y7620 = ~n21387 ;
  assign y7621 = n21393 ;
  assign y7622 = n21395 ;
  assign y7623 = ~n21396 ;
  assign y7624 = ~n21401 ;
  assign y7625 = ~1'b0 ;
  assign y7626 = n21404 ;
  assign y7627 = n21405 ;
  assign y7628 = n21406 ;
  assign y7629 = ~1'b0 ;
  assign y7630 = ~1'b0 ;
  assign y7631 = n21407 ;
  assign y7632 = ~1'b0 ;
  assign y7633 = n21410 ;
  assign y7634 = ~n21411 ;
  assign y7635 = n9389 ;
  assign y7636 = n21413 ;
  assign y7637 = ~n21418 ;
  assign y7638 = ~1'b0 ;
  assign y7639 = ~n21419 ;
  assign y7640 = n21420 ;
  assign y7641 = ~n21422 ;
  assign y7642 = n21425 ;
  assign y7643 = ~n21428 ;
  assign y7644 = n21440 ;
  assign y7645 = ~n21443 ;
  assign y7646 = ~n21444 ;
  assign y7647 = n21446 ;
  assign y7648 = ~1'b0 ;
  assign y7649 = 1'b0 ;
  assign y7650 = ~1'b0 ;
  assign y7651 = ~n21449 ;
  assign y7652 = n21450 ;
  assign y7653 = ~n21457 ;
  assign y7654 = ~n21458 ;
  assign y7655 = ~n2401 ;
  assign y7656 = ~n21459 ;
  assign y7657 = n21461 ;
  assign y7658 = ~1'b0 ;
  assign y7659 = ~1'b0 ;
  assign y7660 = ~1'b0 ;
  assign y7661 = ~1'b0 ;
  assign y7662 = ~n21462 ;
  assign y7663 = ~n21465 ;
  assign y7664 = n21470 ;
  assign y7665 = n21472 ;
  assign y7666 = ~1'b0 ;
  assign y7667 = ~1'b0 ;
  assign y7668 = ~n21475 ;
  assign y7669 = ~n21479 ;
  assign y7670 = n21485 ;
  assign y7671 = n21486 ;
  assign y7672 = n21487 ;
  assign y7673 = 1'b0 ;
  assign y7674 = ~1'b0 ;
  assign y7675 = ~1'b0 ;
  assign y7676 = ~n21489 ;
  assign y7677 = n18150 ;
  assign y7678 = n21493 ;
  assign y7679 = ~n21495 ;
  assign y7680 = ~n21496 ;
  assign y7681 = n21497 ;
  assign y7682 = ~1'b0 ;
  assign y7683 = n21502 ;
  assign y7684 = ~1'b0 ;
  assign y7685 = ~n7987 ;
  assign y7686 = ~n21503 ;
  assign y7687 = n21505 ;
  assign y7688 = ~n21506 ;
  assign y7689 = n21510 ;
  assign y7690 = ~n21512 ;
  assign y7691 = ~n21515 ;
  assign y7692 = ~n21516 ;
  assign y7693 = ~1'b0 ;
  assign y7694 = ~1'b0 ;
  assign y7695 = ~n21517 ;
  assign y7696 = ~n21520 ;
  assign y7697 = ~n21521 ;
  assign y7698 = ~n21523 ;
  assign y7699 = n21525 ;
  assign y7700 = n21529 ;
  assign y7701 = ~n21530 ;
  assign y7702 = ~n21534 ;
  assign y7703 = ~n14956 ;
  assign y7704 = n21541 ;
  assign y7705 = ~n21542 ;
  assign y7706 = n21544 ;
  assign y7707 = n21547 ;
  assign y7708 = n21550 ;
  assign y7709 = ~n21555 ;
  assign y7710 = n21558 ;
  assign y7711 = n21562 ;
  assign y7712 = n21563 ;
  assign y7713 = n21567 ;
  assign y7714 = n21568 ;
  assign y7715 = n21569 ;
  assign y7716 = ~n21572 ;
  assign y7717 = ~n21575 ;
  assign y7718 = n21577 ;
  assign y7719 = ~n21582 ;
  assign y7720 = n21585 ;
  assign y7721 = ~n21586 ;
  assign y7722 = ~n21588 ;
  assign y7723 = n21591 ;
  assign y7724 = ~1'b0 ;
  assign y7725 = ~1'b0 ;
  assign y7726 = ~n21597 ;
  assign y7727 = n21600 ;
  assign y7728 = ~n21603 ;
  assign y7729 = n21605 ;
  assign y7730 = ~n21606 ;
  assign y7731 = ~n21607 ;
  assign y7732 = ~n21612 ;
  assign y7733 = n21613 ;
  assign y7734 = ~n21616 ;
  assign y7735 = ~1'b0 ;
  assign y7736 = n21618 ;
  assign y7737 = ~n15333 ;
  assign y7738 = n21623 ;
  assign y7739 = ~n21626 ;
  assign y7740 = n21628 ;
  assign y7741 = n21630 ;
  assign y7742 = n21631 ;
  assign y7743 = n17277 ;
  assign y7744 = ~1'b0 ;
  assign y7745 = ~n21632 ;
  assign y7746 = n21636 ;
  assign y7747 = n21638 ;
  assign y7748 = ~n21642 ;
  assign y7749 = n21645 ;
  assign y7750 = n21646 ;
  assign y7751 = n21648 ;
  assign y7752 = ~n21649 ;
  assign y7753 = ~n21651 ;
  assign y7754 = ~n21653 ;
  assign y7755 = ~1'b0 ;
  assign y7756 = ~n21654 ;
  assign y7757 = ~n21655 ;
  assign y7758 = ~n21658 ;
  assign y7759 = ~n8704 ;
  assign y7760 = n21661 ;
  assign y7761 = ~1'b0 ;
  assign y7762 = ~n21663 ;
  assign y7763 = n9423 ;
  assign y7764 = n21664 ;
  assign y7765 = n21665 ;
  assign y7766 = n21666 ;
  assign y7767 = ~1'b0 ;
  assign y7768 = ~n21670 ;
  assign y7769 = ~n21672 ;
  assign y7770 = n21674 ;
  assign y7771 = ~n21675 ;
  assign y7772 = n17280 ;
  assign y7773 = n21678 ;
  assign y7774 = n21681 ;
  assign y7775 = ~n21682 ;
  assign y7776 = n18233 ;
  assign y7777 = ~n21687 ;
  assign y7778 = ~1'b0 ;
  assign y7779 = ~1'b0 ;
  assign y7780 = ~1'b0 ;
  assign y7781 = n21688 ;
  assign y7782 = ~n2122 ;
  assign y7783 = ~n21689 ;
  assign y7784 = ~n12589 ;
  assign y7785 = n21692 ;
  assign y7786 = n21693 ;
  assign y7787 = n21695 ;
  assign y7788 = n21696 ;
  assign y7789 = ~n21699 ;
  assign y7790 = ~1'b0 ;
  assign y7791 = n21703 ;
  assign y7792 = n21704 ;
  assign y7793 = ~n21705 ;
  assign y7794 = n21707 ;
  assign y7795 = ~n21711 ;
  assign y7796 = ~n21713 ;
  assign y7797 = ~n21716 ;
  assign y7798 = ~n21717 ;
  assign y7799 = n21718 ;
  assign y7800 = ~n4021 ;
  assign y7801 = n21720 ;
  assign y7802 = ~n21727 ;
  assign y7803 = ~n21728 ;
  assign y7804 = n21729 ;
  assign y7805 = n21730 ;
  assign y7806 = n21736 ;
  assign y7807 = ~n21737 ;
  assign y7808 = n21739 ;
  assign y7809 = n21743 ;
  assign y7810 = n21744 ;
  assign y7811 = n21745 ;
  assign y7812 = ~n21746 ;
  assign y7813 = ~1'b0 ;
  assign y7814 = ~1'b0 ;
  assign y7815 = ~1'b0 ;
  assign y7816 = ~1'b0 ;
  assign y7817 = ~n21749 ;
  assign y7818 = n21750 ;
  assign y7819 = ~n21755 ;
  assign y7820 = n21756 ;
  assign y7821 = ~n21760 ;
  assign y7822 = 1'b0 ;
  assign y7823 = n21767 ;
  assign y7824 = n21768 ;
  assign y7825 = ~n21772 ;
  assign y7826 = ~1'b0 ;
  assign y7827 = n21773 ;
  assign y7828 = ~1'b0 ;
  assign y7829 = ~n21776 ;
  assign y7830 = ~n21782 ;
  assign y7831 = ~1'b0 ;
  assign y7832 = ~n21783 ;
  assign y7833 = n21786 ;
  assign y7834 = n21787 ;
  assign y7835 = ~1'b0 ;
  assign y7836 = n21788 ;
  assign y7837 = n21789 ;
  assign y7838 = ~n8746 ;
  assign y7839 = ~1'b0 ;
  assign y7840 = n21790 ;
  assign y7841 = ~1'b0 ;
  assign y7842 = n21791 ;
  assign y7843 = ~n21797 ;
  assign y7844 = n21799 ;
  assign y7845 = n21800 ;
  assign y7846 = ~n21804 ;
  assign y7847 = n21806 ;
  assign y7848 = n21811 ;
  assign y7849 = n21813 ;
  assign y7850 = n21815 ;
  assign y7851 = ~1'b0 ;
  assign y7852 = ~1'b0 ;
  assign y7853 = n21820 ;
  assign y7854 = ~1'b0 ;
  assign y7855 = n21827 ;
  assign y7856 = n21830 ;
  assign y7857 = n21831 ;
  assign y7858 = ~n21832 ;
  assign y7859 = ~n21836 ;
  assign y7860 = ~n21838 ;
  assign y7861 = n21840 ;
  assign y7862 = ~1'b0 ;
  assign y7863 = n21843 ;
  assign y7864 = n21844 ;
  assign y7865 = n21845 ;
  assign y7866 = ~n21849 ;
  assign y7867 = ~1'b0 ;
  assign y7868 = ~n21850 ;
  assign y7869 = ~n21851 ;
  assign y7870 = ~n21855 ;
  assign y7871 = n21859 ;
  assign y7872 = n21863 ;
  assign y7873 = n21866 ;
  assign y7874 = ~1'b0 ;
  assign y7875 = n21867 ;
  assign y7876 = n21868 ;
  assign y7877 = n21869 ;
  assign y7878 = ~1'b0 ;
  assign y7879 = ~n21871 ;
  assign y7880 = ~n21873 ;
  assign y7881 = ~n21877 ;
  assign y7882 = ~n21878 ;
  assign y7883 = ~n21883 ;
  assign y7884 = n4046 ;
  assign y7885 = n21889 ;
  assign y7886 = ~n21891 ;
  assign y7887 = ~n21896 ;
  assign y7888 = n21897 ;
  assign y7889 = n21903 ;
  assign y7890 = ~n21907 ;
  assign y7891 = n21910 ;
  assign y7892 = n21911 ;
  assign y7893 = n21917 ;
  assign y7894 = ~1'b0 ;
  assign y7895 = ~n21921 ;
  assign y7896 = ~n21929 ;
  assign y7897 = ~1'b0 ;
  assign y7898 = n21931 ;
  assign y7899 = ~n21939 ;
  assign y7900 = ~n21941 ;
  assign y7901 = n21943 ;
  assign y7902 = n21944 ;
  assign y7903 = n21946 ;
  assign y7904 = ~n21947 ;
  assign y7905 = ~n21948 ;
  assign y7906 = n21949 ;
  assign y7907 = ~1'b0 ;
  assign y7908 = n21957 ;
  assign y7909 = ~1'b0 ;
  assign y7910 = n21959 ;
  assign y7911 = ~n21960 ;
  assign y7912 = ~n21961 ;
  assign y7913 = ~n21962 ;
  assign y7914 = n8702 ;
  assign y7915 = n21963 ;
  assign y7916 = n21965 ;
  assign y7917 = ~n21968 ;
  assign y7918 = n21969 ;
  assign y7919 = ~n21970 ;
  assign y7920 = n21972 ;
  assign y7921 = ~1'b0 ;
  assign y7922 = n21973 ;
  assign y7923 = ~1'b0 ;
  assign y7924 = n21974 ;
  assign y7925 = n21977 ;
  assign y7926 = ~n21978 ;
  assign y7927 = ~n21980 ;
  assign y7928 = ~1'b0 ;
  assign y7929 = ~1'b0 ;
  assign y7930 = ~1'b0 ;
  assign y7931 = ~n21982 ;
  assign y7932 = n21984 ;
  assign y7933 = n21985 ;
  assign y7934 = ~n21989 ;
  assign y7935 = n21995 ;
  assign y7936 = ~n21999 ;
  assign y7937 = ~n22000 ;
  assign y7938 = ~n22004 ;
  assign y7939 = ~n22008 ;
  assign y7940 = ~n22012 ;
  assign y7941 = ~n22013 ;
  assign y7942 = n22014 ;
  assign y7943 = ~1'b0 ;
  assign y7944 = ~n22017 ;
  assign y7945 = n22018 ;
  assign y7946 = n22021 ;
  assign y7947 = n22022 ;
  assign y7948 = ~n22025 ;
  assign y7949 = ~n22030 ;
  assign y7950 = n22038 ;
  assign y7951 = n22042 ;
  assign y7952 = ~1'b0 ;
  assign y7953 = ~n22044 ;
  assign y7954 = ~n22046 ;
  assign y7955 = ~n22047 ;
  assign y7956 = ~n22049 ;
  assign y7957 = n22051 ;
  assign y7958 = n22053 ;
  assign y7959 = ~n22058 ;
  assign y7960 = n22061 ;
  assign y7961 = ~n22062 ;
  assign y7962 = n22066 ;
  assign y7963 = ~1'b0 ;
  assign y7964 = n22067 ;
  assign y7965 = n22069 ;
  assign y7966 = ~1'b0 ;
  assign y7967 = n22073 ;
  assign y7968 = ~n13738 ;
  assign y7969 = n22076 ;
  assign y7970 = ~n22078 ;
  assign y7971 = n22085 ;
  assign y7972 = ~1'b0 ;
  assign y7973 = ~n22087 ;
  assign y7974 = ~n22090 ;
  assign y7975 = ~1'b0 ;
  assign y7976 = n22094 ;
  assign y7977 = ~n22098 ;
  assign y7978 = ~n22099 ;
  assign y7979 = n22100 ;
  assign y7980 = ~1'b0 ;
  assign y7981 = ~n22102 ;
  assign y7982 = ~n22104 ;
  assign y7983 = ~n22105 ;
  assign y7984 = ~1'b0 ;
  assign y7985 = ~n22106 ;
  assign y7986 = ~n22107 ;
  assign y7987 = n22108 ;
  assign y7988 = n22109 ;
  assign y7989 = n22111 ;
  assign y7990 = n22114 ;
  assign y7991 = n22119 ;
  assign y7992 = ~n22120 ;
  assign y7993 = n22122 ;
  assign y7994 = ~n22125 ;
  assign y7995 = ~1'b0 ;
  assign y7996 = ~n22126 ;
  assign y7997 = ~n22128 ;
  assign y7998 = ~n22131 ;
  assign y7999 = ~n22132 ;
  assign y8000 = ~n22133 ;
  assign y8001 = n22134 ;
  assign y8002 = n22138 ;
  assign y8003 = ~n22139 ;
  assign y8004 = ~1'b0 ;
  assign y8005 = n22141 ;
  assign y8006 = n22143 ;
  assign y8007 = ~n22147 ;
  assign y8008 = ~n11972 ;
  assign y8009 = n22148 ;
  assign y8010 = ~1'b0 ;
  assign y8011 = ~n22150 ;
  assign y8012 = ~n22156 ;
  assign y8013 = n22157 ;
  assign y8014 = n22160 ;
  assign y8015 = ~n22162 ;
  assign y8016 = n22170 ;
  assign y8017 = ~n22181 ;
  assign y8018 = n22182 ;
  assign y8019 = n22185 ;
  assign y8020 = n22186 ;
  assign y8021 = n22190 ;
  assign y8022 = ~n22194 ;
  assign y8023 = ~n22197 ;
  assign y8024 = ~n22201 ;
  assign y8025 = ~n22205 ;
  assign y8026 = ~n22209 ;
  assign y8027 = ~n22210 ;
  assign y8028 = ~n22219 ;
  assign y8029 = ~n18529 ;
  assign y8030 = n22226 ;
  assign y8031 = n22232 ;
  assign y8032 = ~n22236 ;
  assign y8033 = n22243 ;
  assign y8034 = ~n22244 ;
  assign y8035 = ~1'b0 ;
  assign y8036 = ~n22249 ;
  assign y8037 = n540 ;
  assign y8038 = n22251 ;
  assign y8039 = ~1'b0 ;
  assign y8040 = n22255 ;
  assign y8041 = n22257 ;
  assign y8042 = ~n22260 ;
  assign y8043 = ~n22261 ;
  assign y8044 = n22268 ;
  assign y8045 = ~1'b0 ;
  assign y8046 = ~n22276 ;
  assign y8047 = ~n22280 ;
  assign y8048 = n22289 ;
  assign y8049 = ~n22290 ;
  assign y8050 = n22291 ;
  assign y8051 = n22292 ;
  assign y8052 = n22293 ;
  assign y8053 = ~n22296 ;
  assign y8054 = n22297 ;
  assign y8055 = ~1'b0 ;
  assign y8056 = ~1'b0 ;
  assign y8057 = ~n22298 ;
  assign y8058 = n22301 ;
  assign y8059 = n22303 ;
  assign y8060 = ~1'b0 ;
  assign y8061 = n22307 ;
  assign y8062 = ~n22309 ;
  assign y8063 = ~n22311 ;
  assign y8064 = n22312 ;
  assign y8065 = ~n22313 ;
  assign y8066 = ~n22315 ;
  assign y8067 = ~n22323 ;
  assign y8068 = n22336 ;
  assign y8069 = n22340 ;
  assign y8070 = n22343 ;
  assign y8071 = n22344 ;
  assign y8072 = ~n22346 ;
  assign y8073 = n22347 ;
  assign y8074 = n22348 ;
  assign y8075 = ~n22349 ;
  assign y8076 = ~n22351 ;
  assign y8077 = n22352 ;
  assign y8078 = ~n22363 ;
  assign y8079 = ~1'b0 ;
  assign y8080 = ~1'b0 ;
  assign y8081 = ~n22366 ;
  assign y8082 = ~n22369 ;
  assign y8083 = ~n22370 ;
  assign y8084 = ~n22371 ;
  assign y8085 = ~n22376 ;
  assign y8086 = ~n22377 ;
  assign y8087 = ~1'b0 ;
  assign y8088 = ~n22378 ;
  assign y8089 = ~n22381 ;
  assign y8090 = ~n22382 ;
  assign y8091 = n22384 ;
  assign y8092 = ~n22385 ;
  assign y8093 = ~n22390 ;
  assign y8094 = ~1'b0 ;
  assign y8095 = n22393 ;
  assign y8096 = ~n22398 ;
  assign y8097 = ~n22399 ;
  assign y8098 = ~n22400 ;
  assign y8099 = ~n22403 ;
  assign y8100 = n22408 ;
  assign y8101 = ~n22411 ;
  assign y8102 = ~1'b0 ;
  assign y8103 = ~1'b0 ;
  assign y8104 = ~n22413 ;
  assign y8105 = ~n22416 ;
  assign y8106 = ~n22418 ;
  assign y8107 = ~n22425 ;
  assign y8108 = n22430 ;
  assign y8109 = ~n22431 ;
  assign y8110 = ~1'b0 ;
  assign y8111 = ~1'b0 ;
  assign y8112 = ~1'b0 ;
  assign y8113 = n22436 ;
  assign y8114 = ~n22437 ;
  assign y8115 = ~n22440 ;
  assign y8116 = n22441 ;
  assign y8117 = ~n22445 ;
  assign y8118 = ~n22448 ;
  assign y8119 = ~1'b0 ;
  assign y8120 = n22453 ;
  assign y8121 = ~1'b0 ;
  assign y8122 = ~n22454 ;
  assign y8123 = ~n22459 ;
  assign y8124 = ~n22464 ;
  assign y8125 = ~n22467 ;
  assign y8126 = n22473 ;
  assign y8127 = n22475 ;
  assign y8128 = ~1'b0 ;
  assign y8129 = ~1'b0 ;
  assign y8130 = n134 ;
  assign y8131 = n22480 ;
  assign y8132 = ~n3833 ;
  assign y8133 = n22484 ;
  assign y8134 = ~n22486 ;
  assign y8135 = ~n22489 ;
  assign y8136 = n22491 ;
  assign y8137 = ~1'b0 ;
  assign y8138 = ~n22493 ;
  assign y8139 = n22494 ;
  assign y8140 = ~n22496 ;
  assign y8141 = ~n22500 ;
  assign y8142 = ~n22501 ;
  assign y8143 = ~n22503 ;
  assign y8144 = ~1'b0 ;
  assign y8145 = ~n22504 ;
  assign y8146 = n22506 ;
  assign y8147 = n22509 ;
  assign y8148 = n22513 ;
  assign y8149 = ~n22515 ;
  assign y8150 = ~n22520 ;
  assign y8151 = ~1'b0 ;
  assign y8152 = n22521 ;
  assign y8153 = n7324 ;
  assign y8154 = n22525 ;
  assign y8155 = ~n22527 ;
  assign y8156 = ~n22534 ;
  assign y8157 = ~n22535 ;
  assign y8158 = ~n22540 ;
  assign y8159 = n22541 ;
  assign y8160 = ~n22544 ;
  assign y8161 = ~1'b0 ;
  assign y8162 = ~1'b0 ;
  assign y8163 = n22545 ;
  assign y8164 = n22546 ;
  assign y8165 = ~n22547 ;
  assign y8166 = ~n22549 ;
  assign y8167 = ~n22550 ;
  assign y8168 = n22551 ;
  assign y8169 = ~n22554 ;
  assign y8170 = ~n22555 ;
  assign y8171 = n5886 ;
  assign y8172 = ~n22556 ;
  assign y8173 = ~n22558 ;
  assign y8174 = n22566 ;
  assign y8175 = ~1'b0 ;
  assign y8176 = ~1'b0 ;
  assign y8177 = ~n22568 ;
  assign y8178 = ~n22570 ;
  assign y8179 = ~n22573 ;
  assign y8180 = ~n22578 ;
  assign y8181 = ~n22580 ;
  assign y8182 = ~n12119 ;
  assign y8183 = ~n22581 ;
  assign y8184 = ~1'b0 ;
  assign y8185 = n22584 ;
  assign y8186 = ~n22588 ;
  assign y8187 = ~n22589 ;
  assign y8188 = n22592 ;
  assign y8189 = ~n22593 ;
  assign y8190 = n22594 ;
  assign y8191 = n22595 ;
  assign y8192 = n22598 ;
  assign y8193 = n22605 ;
  assign y8194 = 1'b0 ;
  assign y8195 = n3301 ;
  assign y8196 = ~n22606 ;
  assign y8197 = n22607 ;
  assign y8198 = ~n22608 ;
  assign y8199 = n22609 ;
  assign y8200 = n22610 ;
  assign y8201 = n22620 ;
  assign y8202 = ~1'b0 ;
  assign y8203 = ~1'b0 ;
  assign y8204 = ~n22621 ;
  assign y8205 = ~n22622 ;
  assign y8206 = ~n22624 ;
  assign y8207 = n22626 ;
  assign y8208 = ~1'b0 ;
  assign y8209 = n22628 ;
  assign y8210 = n22629 ;
  assign y8211 = n22630 ;
  assign y8212 = n1473 ;
  assign y8213 = n22632 ;
  assign y8214 = ~n22633 ;
  assign y8215 = n22635 ;
  assign y8216 = ~n22637 ;
  assign y8217 = ~1'b0 ;
  assign y8218 = ~1'b0 ;
  assign y8219 = ~1'b0 ;
  assign y8220 = n22639 ;
  assign y8221 = ~1'b0 ;
  assign y8222 = n22640 ;
  assign y8223 = ~n22641 ;
  assign y8224 = n22643 ;
  assign y8225 = ~n22647 ;
  assign y8226 = ~n22649 ;
  assign y8227 = n22653 ;
  assign y8228 = ~n22657 ;
  assign y8229 = 1'b0 ;
  assign y8230 = n22658 ;
  assign y8231 = ~n22659 ;
  assign y8232 = ~n22660 ;
  assign y8233 = n22662 ;
  assign y8234 = ~n22667 ;
  assign y8235 = n22669 ;
  assign y8236 = ~1'b0 ;
  assign y8237 = ~n22673 ;
  assign y8238 = ~n22674 ;
  assign y8239 = n22675 ;
  assign y8240 = ~n22676 ;
  assign y8241 = ~n22681 ;
  assign y8242 = n22682 ;
  assign y8243 = n22685 ;
  assign y8244 = ~n22692 ;
  assign y8245 = n22696 ;
  assign y8246 = n22699 ;
  assign y8247 = n22705 ;
  assign y8248 = n22707 ;
  assign y8249 = ~n22712 ;
  assign y8250 = ~n22714 ;
  assign y8251 = ~n22717 ;
  assign y8252 = ~n22718 ;
  assign y8253 = ~1'b0 ;
  assign y8254 = ~n610 ;
  assign y8255 = n22723 ;
  assign y8256 = n22727 ;
  assign y8257 = ~n22730 ;
  assign y8258 = ~n7006 ;
  assign y8259 = ~n22731 ;
  assign y8260 = ~n22734 ;
  assign y8261 = ~n22737 ;
  assign y8262 = ~1'b0 ;
  assign y8263 = ~n22740 ;
  assign y8264 = ~n22741 ;
  assign y8265 = n22742 ;
  assign y8266 = ~n22743 ;
  assign y8267 = ~n22751 ;
  assign y8268 = ~1'b0 ;
  assign y8269 = n22752 ;
  assign y8270 = ~n22757 ;
  assign y8271 = n22761 ;
  assign y8272 = n22767 ;
  assign y8273 = n22768 ;
  assign y8274 = ~n22770 ;
  assign y8275 = ~1'b0 ;
  assign y8276 = ~1'b0 ;
  assign y8277 = n22776 ;
  assign y8278 = ~n22777 ;
  assign y8279 = n22783 ;
  assign y8280 = n22786 ;
  assign y8281 = ~n22790 ;
  assign y8282 = n22791 ;
  assign y8283 = n22792 ;
  assign y8284 = ~n22798 ;
  assign y8285 = ~1'b0 ;
  assign y8286 = ~1'b0 ;
  assign y8287 = n22801 ;
  assign y8288 = ~n12501 ;
  assign y8289 = n22803 ;
  assign y8290 = n22808 ;
  assign y8291 = ~n22809 ;
  assign y8292 = n22813 ;
  assign y8293 = ~n22815 ;
  assign y8294 = ~n22816 ;
  assign y8295 = n22817 ;
  assign y8296 = n22818 ;
  assign y8297 = ~1'b0 ;
  assign y8298 = ~n22822 ;
  assign y8299 = ~1'b0 ;
  assign y8300 = n22824 ;
  assign y8301 = n22827 ;
  assign y8302 = ~n22828 ;
  assign y8303 = n22829 ;
  assign y8304 = ~n22830 ;
  assign y8305 = n22833 ;
  assign y8306 = n22835 ;
  assign y8307 = ~n22837 ;
  assign y8308 = ~1'b0 ;
  assign y8309 = ~n22839 ;
  assign y8310 = n22843 ;
  assign y8311 = ~n22847 ;
  assign y8312 = n22849 ;
  assign y8313 = n22852 ;
  assign y8314 = ~n22856 ;
  assign y8315 = n22857 ;
  assign y8316 = ~n22861 ;
  assign y8317 = ~n22869 ;
  assign y8318 = ~1'b0 ;
  assign y8319 = ~n22871 ;
  assign y8320 = ~n22874 ;
  assign y8321 = ~n22875 ;
  assign y8322 = ~n22880 ;
  assign y8323 = n22882 ;
  assign y8324 = n22883 ;
  assign y8325 = ~n22884 ;
  assign y8326 = ~n1314 ;
  assign y8327 = n22889 ;
  assign y8328 = n22892 ;
  assign y8329 = ~1'b0 ;
  assign y8330 = ~n22896 ;
  assign y8331 = ~1'b0 ;
  assign y8332 = ~n22897 ;
  assign y8333 = ~n22900 ;
  assign y8334 = ~n22904 ;
  assign y8335 = ~n22905 ;
  assign y8336 = ~n22906 ;
  assign y8337 = n22907 ;
  assign y8338 = n22909 ;
  assign y8339 = ~n22910 ;
  assign y8340 = 1'b0 ;
  assign y8341 = ~n22912 ;
  assign y8342 = ~n22913 ;
  assign y8343 = ~n22915 ;
  assign y8344 = n22916 ;
  assign y8345 = ~n22918 ;
  assign y8346 = n22920 ;
  assign y8347 = n22923 ;
  assign y8348 = ~n22929 ;
  assign y8349 = ~n22932 ;
  assign y8350 = n22934 ;
  assign y8351 = ~n22936 ;
  assign y8352 = n22937 ;
  assign y8353 = ~n22939 ;
  assign y8354 = n22941 ;
  assign y8355 = 1'b0 ;
  assign y8356 = ~1'b0 ;
  assign y8357 = n22942 ;
  assign y8358 = ~n22947 ;
  assign y8359 = n22948 ;
  assign y8360 = n22950 ;
  assign y8361 = ~n22954 ;
  assign y8362 = n22956 ;
  assign y8363 = n22957 ;
  assign y8364 = n22962 ;
  assign y8365 = ~n22963 ;
  assign y8366 = n22964 ;
  assign y8367 = ~1'b0 ;
  assign y8368 = n22966 ;
  assign y8369 = ~1'b0 ;
  assign y8370 = ~1'b0 ;
  assign y8371 = ~n22981 ;
  assign y8372 = ~n22985 ;
  assign y8373 = n22986 ;
  assign y8374 = ~n22987 ;
  assign y8375 = n22989 ;
  assign y8376 = ~1'b0 ;
  assign y8377 = n22990 ;
  assign y8378 = ~n22993 ;
  assign y8379 = n22997 ;
  assign y8380 = ~1'b0 ;
  assign y8381 = ~1'b0 ;
  assign y8382 = n23000 ;
  assign y8383 = ~n23007 ;
  assign y8384 = ~n23013 ;
  assign y8385 = ~n23014 ;
  assign y8386 = ~1'b0 ;
  assign y8387 = ~n23019 ;
  assign y8388 = 1'b0 ;
  assign y8389 = n23021 ;
  assign y8390 = ~n23023 ;
  assign y8391 = ~1'b0 ;
  assign y8392 = n23025 ;
  assign y8393 = n23026 ;
  assign y8394 = n23027 ;
  assign y8395 = n23031 ;
  assign y8396 = ~n23038 ;
  assign y8397 = n23040 ;
  assign y8398 = ~n23042 ;
  assign y8399 = ~1'b0 ;
  assign y8400 = ~n10065 ;
  assign y8401 = ~n23045 ;
  assign y8402 = n23047 ;
  assign y8403 = n23048 ;
  assign y8404 = ~1'b0 ;
  assign y8405 = n23049 ;
  assign y8406 = ~1'b0 ;
  assign y8407 = n23051 ;
  assign y8408 = ~n23052 ;
  assign y8409 = n23056 ;
  assign y8410 = ~n23061 ;
  assign y8411 = n23062 ;
  assign y8412 = ~n23066 ;
  assign y8413 = ~1'b0 ;
  assign y8414 = n23067 ;
  assign y8415 = ~n23069 ;
  assign y8416 = n23072 ;
  assign y8417 = n23073 ;
  assign y8418 = ~1'b0 ;
  assign y8419 = ~n23075 ;
  assign y8420 = n23079 ;
  assign y8421 = n23080 ;
  assign y8422 = n23082 ;
  assign y8423 = ~n23086 ;
  assign y8424 = ~n23088 ;
  assign y8425 = ~n13133 ;
  assign y8426 = ~n23091 ;
  assign y8427 = ~n23092 ;
  assign y8428 = ~n23093 ;
  assign y8429 = ~n23095 ;
  assign y8430 = ~n23097 ;
  assign y8431 = ~1'b0 ;
  assign y8432 = ~n23100 ;
  assign y8433 = n23102 ;
  assign y8434 = n18406 ;
  assign y8435 = n23103 ;
  assign y8436 = ~n23108 ;
  assign y8437 = ~n23110 ;
  assign y8438 = ~n23111 ;
  assign y8439 = ~1'b0 ;
  assign y8440 = n23113 ;
  assign y8441 = ~n23118 ;
  assign y8442 = ~n23121 ;
  assign y8443 = ~n23124 ;
  assign y8444 = ~1'b0 ;
  assign y8445 = ~n23126 ;
  assign y8446 = n23128 ;
  assign y8447 = ~1'b0 ;
  assign y8448 = n23129 ;
  assign y8449 = ~n23130 ;
  assign y8450 = ~n23142 ;
  assign y8451 = ~n5665 ;
  assign y8452 = n23143 ;
  assign y8453 = ~n23145 ;
  assign y8454 = ~n162 ;
  assign y8455 = ~n23147 ;
  assign y8456 = ~n23150 ;
  assign y8457 = ~1'b0 ;
  assign y8458 = ~n23151 ;
  assign y8459 = ~n23152 ;
  assign y8460 = n23155 ;
  assign y8461 = n23156 ;
  assign y8462 = n23158 ;
  assign y8463 = n23161 ;
  assign y8464 = ~1'b0 ;
  assign y8465 = ~n23163 ;
  assign y8466 = ~n23164 ;
  assign y8467 = ~1'b0 ;
  assign y8468 = ~n23166 ;
  assign y8469 = ~n23171 ;
  assign y8470 = ~1'b0 ;
  assign y8471 = n23172 ;
  assign y8472 = ~n23175 ;
  assign y8473 = ~n23179 ;
  assign y8474 = ~1'b0 ;
  assign y8475 = n23181 ;
  assign y8476 = ~n23187 ;
  assign y8477 = n23189 ;
  assign y8478 = ~n23190 ;
  assign y8479 = n23191 ;
  assign y8480 = ~1'b0 ;
  assign y8481 = n23195 ;
  assign y8482 = n23196 ;
  assign y8483 = ~n23199 ;
  assign y8484 = n23202 ;
  assign y8485 = n6288 ;
  assign y8486 = ~n23204 ;
  assign y8487 = ~n23206 ;
  assign y8488 = ~n23210 ;
  assign y8489 = n23212 ;
  assign y8490 = ~1'b0 ;
  assign y8491 = ~n20530 ;
  assign y8492 = ~n23218 ;
  assign y8493 = n23220 ;
  assign y8494 = ~1'b0 ;
  assign y8495 = ~1'b0 ;
  assign y8496 = n23221 ;
  assign y8497 = n1213 ;
  assign y8498 = n23224 ;
  assign y8499 = n23225 ;
  assign y8500 = n23229 ;
  assign y8501 = ~n19769 ;
  assign y8502 = n23231 ;
  assign y8503 = ~n3035 ;
  assign y8504 = n23233 ;
  assign y8505 = ~n23235 ;
  assign y8506 = ~n23236 ;
  assign y8507 = ~n23241 ;
  assign y8508 = ~n23245 ;
  assign y8509 = ~n23247 ;
  assign y8510 = ~1'b0 ;
  assign y8511 = ~n23248 ;
  assign y8512 = ~n23250 ;
  assign y8513 = n23254 ;
  assign y8514 = n23259 ;
  assign y8515 = n23262 ;
  assign y8516 = ~n23265 ;
  assign y8517 = ~n23267 ;
  assign y8518 = n14889 ;
  assign y8519 = ~n23270 ;
  assign y8520 = n23274 ;
  assign y8521 = n23277 ;
  assign y8522 = n23278 ;
  assign y8523 = n23287 ;
  assign y8524 = n23291 ;
  assign y8525 = ~n23296 ;
  assign y8526 = n23297 ;
  assign y8527 = ~1'b0 ;
  assign y8528 = ~1'b0 ;
  assign y8529 = n23298 ;
  assign y8530 = n23299 ;
  assign y8531 = ~n23300 ;
  assign y8532 = ~n23308 ;
  assign y8533 = ~1'b0 ;
  assign y8534 = n23310 ;
  assign y8535 = ~1'b0 ;
  assign y8536 = ~1'b0 ;
  assign y8537 = n23314 ;
  assign y8538 = ~n23318 ;
  assign y8539 = n23319 ;
  assign y8540 = n23320 ;
  assign y8541 = ~1'b0 ;
  assign y8542 = n23326 ;
  assign y8543 = n23328 ;
  assign y8544 = n23333 ;
  assign y8545 = ~1'b0 ;
  assign y8546 = ~n23334 ;
  assign y8547 = ~n23335 ;
  assign y8548 = n23337 ;
  assign y8549 = ~n23340 ;
  assign y8550 = ~1'b0 ;
  assign y8551 = ~n23341 ;
  assign y8552 = n23343 ;
  assign y8553 = ~n23346 ;
  assign y8554 = ~n23347 ;
  assign y8555 = ~n9245 ;
  assign y8556 = n23353 ;
  assign y8557 = n23354 ;
  assign y8558 = ~1'b0 ;
  assign y8559 = ~n23355 ;
  assign y8560 = ~1'b0 ;
  assign y8561 = ~n23359 ;
  assign y8562 = n23360 ;
  assign y8563 = n23361 ;
  assign y8564 = n23362 ;
  assign y8565 = n23364 ;
  assign y8566 = n23366 ;
  assign y8567 = ~1'b0 ;
  assign y8568 = ~1'b0 ;
  assign y8569 = n23368 ;
  assign y8570 = ~1'b0 ;
  assign y8571 = n23369 ;
  assign y8572 = ~n23370 ;
  assign y8573 = n23372 ;
  assign y8574 = ~n23379 ;
  assign y8575 = ~1'b0 ;
  assign y8576 = ~n23382 ;
  assign y8577 = ~n23385 ;
  assign y8578 = n23388 ;
  assign y8579 = ~n23392 ;
  assign y8580 = ~n23397 ;
  assign y8581 = n23400 ;
  assign y8582 = ~n23402 ;
  assign y8583 = ~n23403 ;
  assign y8584 = ~n23404 ;
  assign y8585 = ~n23406 ;
  assign y8586 = n23408 ;
  assign y8587 = n23412 ;
  assign y8588 = ~n23416 ;
  assign y8589 = n23419 ;
  assign y8590 = ~n23421 ;
  assign y8591 = n23427 ;
  assign y8592 = n23428 ;
  assign y8593 = ~n21349 ;
  assign y8594 = n23432 ;
  assign y8595 = n23437 ;
  assign y8596 = n23438 ;
  assign y8597 = ~1'b0 ;
  assign y8598 = ~1'b0 ;
  assign y8599 = n23443 ;
  assign y8600 = ~1'b0 ;
  assign y8601 = ~n23446 ;
  assign y8602 = ~n23453 ;
  assign y8603 = ~n23454 ;
  assign y8604 = n23456 ;
  assign y8605 = n23457 ;
  assign y8606 = n23459 ;
  assign y8607 = ~1'b0 ;
  assign y8608 = ~1'b0 ;
  assign y8609 = ~n23460 ;
  assign y8610 = ~1'b0 ;
  assign y8611 = n23462 ;
  assign y8612 = ~n23465 ;
  assign y8613 = n23470 ;
  assign y8614 = ~n23472 ;
  assign y8615 = n23479 ;
  assign y8616 = ~1'b0 ;
  assign y8617 = ~n23485 ;
  assign y8618 = ~n23487 ;
  assign y8619 = n23488 ;
  assign y8620 = n23489 ;
  assign y8621 = ~n11893 ;
  assign y8622 = ~n23492 ;
  assign y8623 = ~n23494 ;
  assign y8624 = 1'b0 ;
  assign y8625 = n23497 ;
  assign y8626 = n23498 ;
  assign y8627 = ~n8572 ;
  assign y8628 = n23502 ;
  assign y8629 = ~n23505 ;
  assign y8630 = n23509 ;
  assign y8631 = n8951 ;
  assign y8632 = ~n23511 ;
  assign y8633 = ~n23512 ;
  assign y8634 = ~n23515 ;
  assign y8635 = ~n23518 ;
  assign y8636 = n23521 ;
  assign y8637 = ~n5665 ;
  assign y8638 = n23530 ;
  assign y8639 = ~n23535 ;
  assign y8640 = ~1'b0 ;
  assign y8641 = n23542 ;
  assign y8642 = n5134 ;
  assign y8643 = ~n23543 ;
  assign y8644 = n23545 ;
  assign y8645 = ~1'b0 ;
  assign y8646 = ~1'b0 ;
  assign y8647 = n23547 ;
  assign y8648 = ~1'b0 ;
  assign y8649 = n23551 ;
  assign y8650 = ~n23560 ;
  assign y8651 = n23561 ;
  assign y8652 = ~n23564 ;
  assign y8653 = ~n23569 ;
  assign y8654 = ~n23570 ;
  assign y8655 = ~n23573 ;
  assign y8656 = ~1'b0 ;
  assign y8657 = ~1'b0 ;
  assign y8658 = ~1'b0 ;
  assign y8659 = n23574 ;
  assign y8660 = ~n23578 ;
  assign y8661 = ~n23579 ;
  assign y8662 = ~n23580 ;
  assign y8663 = n23581 ;
  assign y8664 = ~n23584 ;
  assign y8665 = n23588 ;
  assign y8666 = ~n23592 ;
  assign y8667 = ~1'b0 ;
  assign y8668 = n23593 ;
  assign y8669 = ~n23596 ;
  assign y8670 = ~n23597 ;
  assign y8671 = ~1'b0 ;
  assign y8672 = ~n23601 ;
  assign y8673 = ~n23602 ;
  assign y8674 = ~n23605 ;
  assign y8675 = ~n23606 ;
  assign y8676 = n23611 ;
  assign y8677 = ~n23612 ;
  assign y8678 = ~n23614 ;
  assign y8679 = ~1'b0 ;
  assign y8680 = ~n23617 ;
  assign y8681 = ~n23618 ;
  assign y8682 = n23623 ;
  assign y8683 = n23624 ;
  assign y8684 = n23625 ;
  assign y8685 = ~n23627 ;
  assign y8686 = n23629 ;
  assign y8687 = n23635 ;
  assign y8688 = n23636 ;
  assign y8689 = ~n23639 ;
  assign y8690 = ~n23640 ;
  assign y8691 = n23656 ;
  assign y8692 = ~n23657 ;
  assign y8693 = ~n23659 ;
  assign y8694 = ~n23661 ;
  assign y8695 = ~n23662 ;
  assign y8696 = ~1'b0 ;
  assign y8697 = ~n23664 ;
  assign y8698 = n23665 ;
  assign y8699 = n23666 ;
  assign y8700 = n23667 ;
  assign y8701 = n23669 ;
  assign y8702 = n23674 ;
  assign y8703 = 1'b0 ;
  assign y8704 = n23676 ;
  assign y8705 = ~n23679 ;
  assign y8706 = n23682 ;
  assign y8707 = n1647 ;
  assign y8708 = ~n20829 ;
  assign y8709 = n23687 ;
  assign y8710 = ~n23688 ;
  assign y8711 = ~n23690 ;
  assign y8712 = n23692 ;
  assign y8713 = n23696 ;
  assign y8714 = ~n23697 ;
  assign y8715 = ~n23698 ;
  assign y8716 = ~n23699 ;
  assign y8717 = ~n23701 ;
  assign y8718 = ~1'b0 ;
  assign y8719 = ~1'b0 ;
  assign y8720 = n23704 ;
  assign y8721 = ~1'b0 ;
  assign y8722 = n23709 ;
  assign y8723 = n23710 ;
  assign y8724 = n23711 ;
  assign y8725 = n23712 ;
  assign y8726 = n23717 ;
  assign y8727 = ~n23720 ;
  assign y8728 = ~n23723 ;
  assign y8729 = ~1'b0 ;
  assign y8730 = ~n23725 ;
  assign y8731 = ~1'b0 ;
  assign y8732 = ~1'b0 ;
  assign y8733 = n23733 ;
  assign y8734 = n23737 ;
  assign y8735 = ~n23738 ;
  assign y8736 = ~n23740 ;
  assign y8737 = ~1'b0 ;
  assign y8738 = ~1'b0 ;
  assign y8739 = n23473 ;
  assign y8740 = n4689 ;
  assign y8741 = n23742 ;
  assign y8742 = n23747 ;
  assign y8743 = n23750 ;
  assign y8744 = ~n23752 ;
  assign y8745 = ~1'b0 ;
  assign y8746 = ~n23753 ;
  assign y8747 = ~n23756 ;
  assign y8748 = ~1'b0 ;
  assign y8749 = ~n23760 ;
  assign y8750 = n23765 ;
  assign y8751 = ~n23766 ;
  assign y8752 = n23774 ;
  assign y8753 = ~n23775 ;
  assign y8754 = ~1'b0 ;
  assign y8755 = n23782 ;
  assign y8756 = n3626 ;
  assign y8757 = ~n8583 ;
  assign y8758 = n23783 ;
  assign y8759 = ~n23784 ;
  assign y8760 = ~1'b0 ;
  assign y8761 = ~1'b0 ;
  assign y8762 = n23788 ;
  assign y8763 = ~1'b0 ;
  assign y8764 = n23789 ;
  assign y8765 = n23790 ;
  assign y8766 = ~n23791 ;
  assign y8767 = ~n23795 ;
  assign y8768 = ~n23796 ;
  assign y8769 = ~n23801 ;
  assign y8770 = n23803 ;
  assign y8771 = n23805 ;
  assign y8772 = n23808 ;
  assign y8773 = ~1'b0 ;
  assign y8774 = ~n23811 ;
  assign y8775 = ~n23812 ;
  assign y8776 = n23813 ;
  assign y8777 = n23814 ;
  assign y8778 = ~1'b0 ;
  assign y8779 = ~n23816 ;
  assign y8780 = ~n23819 ;
  assign y8781 = n23826 ;
  assign y8782 = ~n21825 ;
  assign y8783 = n23830 ;
  assign y8784 = ~n23831 ;
  assign y8785 = ~n23841 ;
  assign y8786 = ~n23842 ;
  assign y8787 = n23845 ;
  assign y8788 = n23846 ;
  assign y8789 = ~1'b0 ;
  assign y8790 = n23848 ;
  assign y8791 = n23849 ;
  assign y8792 = n23852 ;
  assign y8793 = ~1'b0 ;
  assign y8794 = ~n23857 ;
  assign y8795 = ~1'b0 ;
  assign y8796 = ~n23861 ;
  assign y8797 = n23866 ;
  assign y8798 = ~n23867 ;
  assign y8799 = n23868 ;
  assign y8800 = ~n23876 ;
  assign y8801 = n23879 ;
  assign y8802 = ~n23881 ;
  assign y8803 = n23884 ;
  assign y8804 = n23889 ;
  assign y8805 = ~1'b0 ;
  assign y8806 = n10431 ;
  assign y8807 = n23891 ;
  assign y8808 = ~1'b0 ;
  assign y8809 = ~n23893 ;
  assign y8810 = n23897 ;
  assign y8811 = n23898 ;
  assign y8812 = ~n23899 ;
  assign y8813 = ~n23900 ;
  assign y8814 = ~n23901 ;
  assign y8815 = ~n23906 ;
  assign y8816 = n23908 ;
  assign y8817 = n23909 ;
  assign y8818 = ~n23910 ;
  assign y8819 = ~n23912 ;
  assign y8820 = ~n23913 ;
  assign y8821 = n23918 ;
  assign y8822 = ~n23919 ;
  assign y8823 = n23921 ;
  assign y8824 = n23923 ;
  assign y8825 = ~n23925 ;
  assign y8826 = ~n6279 ;
  assign y8827 = n23927 ;
  assign y8828 = n23929 ;
  assign y8829 = ~n23930 ;
  assign y8830 = ~n23934 ;
  assign y8831 = ~n23941 ;
  assign y8832 = ~n23943 ;
  assign y8833 = ~1'b0 ;
  assign y8834 = n23945 ;
  assign y8835 = n23946 ;
  assign y8836 = ~n23947 ;
  assign y8837 = ~n23949 ;
  assign y8838 = ~n23950 ;
  assign y8839 = ~n23951 ;
  assign y8840 = ~n23953 ;
  assign y8841 = n23957 ;
  assign y8842 = ~1'b0 ;
  assign y8843 = ~n23960 ;
  assign y8844 = ~n23964 ;
  assign y8845 = ~n23967 ;
  assign y8846 = n23968 ;
  assign y8847 = n23976 ;
  assign y8848 = ~n23978 ;
  assign y8849 = ~n23980 ;
  assign y8850 = ~1'b0 ;
  assign y8851 = ~n23984 ;
  assign y8852 = ~n23985 ;
  assign y8853 = n23991 ;
  assign y8854 = ~n23992 ;
  assign y8855 = ~n23998 ;
  assign y8856 = ~n24003 ;
  assign y8857 = ~n24007 ;
  assign y8858 = n24013 ;
  assign y8859 = ~n24018 ;
  assign y8860 = n24023 ;
  assign y8861 = n24026 ;
  assign y8862 = ~n24028 ;
  assign y8863 = ~n24030 ;
  assign y8864 = ~n24033 ;
  assign y8865 = n24034 ;
  assign y8866 = ~n24048 ;
  assign y8867 = ~n24050 ;
  assign y8868 = ~1'b0 ;
  assign y8869 = ~1'b0 ;
  assign y8870 = ~1'b0 ;
  assign y8871 = ~n24051 ;
  assign y8872 = ~n24055 ;
  assign y8873 = n24060 ;
  assign y8874 = ~n24063 ;
  assign y8875 = ~1'b0 ;
  assign y8876 = ~n24064 ;
  assign y8877 = n24066 ;
  assign y8878 = n24067 ;
  assign y8879 = n24070 ;
  assign y8880 = n24075 ;
  assign y8881 = n24076 ;
  assign y8882 = n24080 ;
  assign y8883 = ~n24081 ;
  assign y8884 = n24082 ;
  assign y8885 = n24084 ;
  assign y8886 = ~n24086 ;
  assign y8887 = n24087 ;
  assign y8888 = n24088 ;
  assign y8889 = ~n24092 ;
  assign y8890 = ~n24095 ;
  assign y8891 = n24097 ;
  assign y8892 = ~n24099 ;
  assign y8893 = n24107 ;
  assign y8894 = n24109 ;
  assign y8895 = n24111 ;
  assign y8896 = n24113 ;
  assign y8897 = ~n24114 ;
  assign y8898 = ~1'b0 ;
  assign y8899 = 1'b0 ;
  assign y8900 = ~1'b0 ;
  assign y8901 = n24116 ;
  assign y8902 = ~n24120 ;
  assign y8903 = n24123 ;
  assign y8904 = n24124 ;
  assign y8905 = n24125 ;
  assign y8906 = n24127 ;
  assign y8907 = ~n24129 ;
  assign y8908 = n24130 ;
  assign y8909 = ~n24132 ;
  assign y8910 = n24133 ;
  assign y8911 = ~n24136 ;
  assign y8912 = n24137 ;
  assign y8913 = n24144 ;
  assign y8914 = ~1'b0 ;
  assign y8915 = ~n24146 ;
  assign y8916 = n24149 ;
  assign y8917 = ~1'b0 ;
  assign y8918 = ~1'b0 ;
  assign y8919 = n24151 ;
  assign y8920 = n24156 ;
  assign y8921 = n24159 ;
  assign y8922 = n24160 ;
  assign y8923 = ~1'b0 ;
  assign y8924 = n24169 ;
  assign y8925 = ~1'b0 ;
  assign y8926 = ~n24170 ;
  assign y8927 = ~n24171 ;
  assign y8928 = n24175 ;
  assign y8929 = n24176 ;
  assign y8930 = ~1'b0 ;
  assign y8931 = ~1'b0 ;
  assign y8932 = n24178 ;
  assign y8933 = n24181 ;
  assign y8934 = n1271 ;
  assign y8935 = n24183 ;
  assign y8936 = n24184 ;
  assign y8937 = n24190 ;
  assign y8938 = ~n24191 ;
  assign y8939 = ~n24193 ;
  assign y8940 = n24201 ;
  assign y8941 = ~n24205 ;
  assign y8942 = ~n24207 ;
  assign y8943 = n24208 ;
  assign y8944 = ~n24212 ;
  assign y8945 = n24213 ;
  assign y8946 = ~n24216 ;
  assign y8947 = n24219 ;
  assign y8948 = ~n24222 ;
  assign y8949 = ~n24224 ;
  assign y8950 = ~1'b0 ;
  assign y8951 = ~n24229 ;
  assign y8952 = ~1'b0 ;
  assign y8953 = ~1'b0 ;
  assign y8954 = ~n24231 ;
  assign y8955 = ~n24232 ;
  assign y8956 = ~n24234 ;
  assign y8957 = ~n17576 ;
  assign y8958 = n24237 ;
  assign y8959 = ~1'b0 ;
  assign y8960 = ~n24242 ;
  assign y8961 = ~1'b0 ;
  assign y8962 = ~n24251 ;
  assign y8963 = n24252 ;
  assign y8964 = n24255 ;
  assign y8965 = ~n24259 ;
  assign y8966 = n24260 ;
  assign y8967 = ~n24263 ;
  assign y8968 = n24265 ;
  assign y8969 = ~n24268 ;
  assign y8970 = ~1'b0 ;
  assign y8971 = n24273 ;
  assign y8972 = n24275 ;
  assign y8973 = ~n24279 ;
  assign y8974 = ~n24280 ;
  assign y8975 = ~n3165 ;
  assign y8976 = ~n24283 ;
  assign y8977 = n24284 ;
  assign y8978 = ~n24285 ;
  assign y8979 = n24286 ;
  assign y8980 = ~n24291 ;
  assign y8981 = ~n24295 ;
  assign y8982 = n24298 ;
  assign y8983 = ~n24299 ;
  assign y8984 = ~n24301 ;
  assign y8985 = ~1'b0 ;
  assign y8986 = ~n24303 ;
  assign y8987 = n24304 ;
  assign y8988 = n24305 ;
  assign y8989 = n24312 ;
  assign y8990 = ~n24313 ;
  assign y8991 = n24317 ;
  assign y8992 = ~n24319 ;
  assign y8993 = ~n24320 ;
  assign y8994 = ~n24323 ;
  assign y8995 = ~n24324 ;
  assign y8996 = n24326 ;
  assign y8997 = ~n24329 ;
  assign y8998 = ~n24331 ;
  assign y8999 = n24332 ;
  assign y9000 = ~1'b0 ;
  assign y9001 = n24335 ;
  assign y9002 = ~n24336 ;
  assign y9003 = n24338 ;
  assign y9004 = n24342 ;
  assign y9005 = n24343 ;
  assign y9006 = ~n24349 ;
  assign y9007 = ~n24353 ;
  assign y9008 = n24355 ;
  assign y9009 = ~n24356 ;
  assign y9010 = ~n24357 ;
  assign y9011 = n24358 ;
  assign y9012 = ~1'b0 ;
  assign y9013 = n24362 ;
  assign y9014 = n24363 ;
  assign y9015 = ~n24364 ;
  assign y9016 = n24366 ;
  assign y9017 = n20315 ;
  assign y9018 = n24367 ;
  assign y9019 = ~1'b0 ;
  assign y9020 = ~1'b0 ;
  assign y9021 = ~n24371 ;
  assign y9022 = ~n24372 ;
  assign y9023 = n24380 ;
  assign y9024 = n24386 ;
  assign y9025 = ~n24387 ;
  assign y9026 = n24392 ;
  assign y9027 = ~n24394 ;
  assign y9028 = ~1'b0 ;
  assign y9029 = n24397 ;
  assign y9030 = ~1'b0 ;
  assign y9031 = ~1'b0 ;
  assign y9032 = ~n24400 ;
  assign y9033 = ~n24401 ;
  assign y9034 = ~n24406 ;
  assign y9035 = ~n24407 ;
  assign y9036 = n24411 ;
  assign y9037 = ~n24414 ;
  assign y9038 = n24419 ;
  assign y9039 = ~n24421 ;
  assign y9040 = ~n24425 ;
  assign y9041 = n24427 ;
  assign y9042 = ~n24430 ;
  assign y9043 = n24431 ;
  assign y9044 = ~n24432 ;
  assign y9045 = ~1'b0 ;
  assign y9046 = ~n24434 ;
  assign y9047 = ~1'b0 ;
  assign y9048 = n24435 ;
  assign y9049 = ~n24437 ;
  assign y9050 = n24440 ;
  assign y9051 = n12633 ;
  assign y9052 = ~1'b0 ;
  assign y9053 = n24441 ;
  assign y9054 = n24444 ;
  assign y9055 = n24448 ;
  assign y9056 = ~1'b0 ;
  assign y9057 = ~n24451 ;
  assign y9058 = ~1'b0 ;
  assign y9059 = n24454 ;
  assign y9060 = n24456 ;
  assign y9061 = n24458 ;
  assign y9062 = ~n24459 ;
  assign y9063 = n24462 ;
  assign y9064 = n24463 ;
  assign y9065 = n24465 ;
  assign y9066 = ~n24466 ;
  assign y9067 = n24469 ;
  assign y9068 = ~n24472 ;
  assign y9069 = ~n24476 ;
  assign y9070 = n24485 ;
  assign y9071 = n24487 ;
  assign y9072 = ~n24492 ;
  assign y9073 = n24494 ;
  assign y9074 = n24495 ;
  assign y9075 = n24496 ;
  assign y9076 = ~1'b0 ;
  assign y9077 = n24498 ;
  assign y9078 = ~1'b0 ;
  assign y9079 = ~n24502 ;
  assign y9080 = n14867 ;
  assign y9081 = n24503 ;
  assign y9082 = ~n24504 ;
  assign y9083 = n24506 ;
  assign y9084 = ~n24510 ;
  assign y9085 = n24520 ;
  assign y9086 = n24526 ;
  assign y9087 = ~n24530 ;
  assign y9088 = n24534 ;
  assign y9089 = ~n24538 ;
  assign y9090 = n24542 ;
  assign y9091 = n24544 ;
  assign y9092 = n24550 ;
  assign y9093 = ~n24552 ;
  assign y9094 = ~1'b0 ;
  assign y9095 = n24558 ;
  assign y9096 = n24559 ;
  assign y9097 = n24561 ;
  assign y9098 = ~n16021 ;
  assign y9099 = ~n24565 ;
  assign y9100 = n24568 ;
  assign y9101 = ~1'b0 ;
  assign y9102 = ~n24570 ;
  assign y9103 = n20098 ;
  assign y9104 = n24572 ;
  assign y9105 = n12350 ;
  assign y9106 = n24574 ;
  assign y9107 = ~n24577 ;
  assign y9108 = n24582 ;
  assign y9109 = ~1'b0 ;
  assign y9110 = ~n24584 ;
  assign y9111 = ~n24588 ;
  assign y9112 = n24590 ;
  assign y9113 = n24591 ;
  assign y9114 = ~n24595 ;
  assign y9115 = ~n24596 ;
  assign y9116 = n24598 ;
  assign y9117 = n24599 ;
  assign y9118 = ~n24601 ;
  assign y9119 = n24602 ;
  assign y9120 = ~n24603 ;
  assign y9121 = ~n24604 ;
  assign y9122 = ~n1175 ;
  assign y9123 = ~1'b0 ;
  assign y9124 = ~1'b0 ;
  assign y9125 = 1'b0 ;
  assign y9126 = ~1'b0 ;
  assign y9127 = ~1'b0 ;
  assign y9128 = n24606 ;
  assign y9129 = n24607 ;
  assign y9130 = ~n24618 ;
  assign y9131 = n24619 ;
  assign y9132 = n24622 ;
  assign y9133 = ~n24624 ;
  assign y9134 = ~1'b0 ;
  assign y9135 = n24627 ;
  assign y9136 = ~n24629 ;
  assign y9137 = n24630 ;
  assign y9138 = ~n24631 ;
  assign y9139 = ~n24636 ;
  assign y9140 = ~n24639 ;
  assign y9141 = ~n24645 ;
  assign y9142 = ~n24648 ;
  assign y9143 = ~1'b0 ;
  assign y9144 = n24650 ;
  assign y9145 = ~n24651 ;
  assign y9146 = n24653 ;
  assign y9147 = ~1'b0 ;
  assign y9148 = ~1'b0 ;
  assign y9149 = n24656 ;
  assign y9150 = n24657 ;
  assign y9151 = n24658 ;
  assign y9152 = ~n24663 ;
  assign y9153 = n24664 ;
  assign y9154 = n24665 ;
  assign y9155 = n24666 ;
  assign y9156 = n24667 ;
  assign y9157 = ~n24670 ;
  assign y9158 = n24672 ;
  assign y9159 = ~1'b0 ;
  assign y9160 = ~n24674 ;
  assign y9161 = ~n24677 ;
  assign y9162 = ~1'b0 ;
  assign y9163 = n24683 ;
  assign y9164 = ~1'b0 ;
  assign y9165 = n24687 ;
  assign y9166 = ~n24691 ;
  assign y9167 = ~n24692 ;
  assign y9168 = n24693 ;
  assign y9169 = ~n24695 ;
  assign y9170 = n24697 ;
  assign y9171 = n24698 ;
  assign y9172 = ~n24702 ;
  assign y9173 = n24703 ;
  assign y9174 = ~1'b0 ;
  assign y9175 = ~n24705 ;
  assign y9176 = ~1'b0 ;
  assign y9177 = ~n24706 ;
  assign y9178 = n24709 ;
  assign y9179 = ~n24710 ;
  assign y9180 = n24713 ;
  assign y9181 = ~1'b0 ;
  assign y9182 = ~n24718 ;
  assign y9183 = ~1'b0 ;
  assign y9184 = n24719 ;
  assign y9185 = n24728 ;
  assign y9186 = ~n24730 ;
  assign y9187 = ~1'b0 ;
  assign y9188 = ~1'b0 ;
  assign y9189 = ~n24733 ;
  assign y9190 = ~n24735 ;
  assign y9191 = ~n24736 ;
  assign y9192 = ~n24738 ;
  assign y9193 = n24740 ;
  assign y9194 = ~n8272 ;
  assign y9195 = n24741 ;
  assign y9196 = n24744 ;
  assign y9197 = n24746 ;
  assign y9198 = ~n24748 ;
  assign y9199 = n24753 ;
  assign y9200 = ~1'b0 ;
  assign y9201 = ~n24758 ;
  assign y9202 = ~n24760 ;
  assign y9203 = ~n24765 ;
  assign y9204 = ~n24766 ;
  assign y9205 = ~1'b0 ;
  assign y9206 = ~1'b0 ;
  assign y9207 = ~n24768 ;
  assign y9208 = ~1'b0 ;
  assign y9209 = ~n24770 ;
  assign y9210 = n24771 ;
  assign y9211 = n24772 ;
  assign y9212 = ~n24773 ;
  assign y9213 = ~n24776 ;
  assign y9214 = n24778 ;
  assign y9215 = ~n24779 ;
  assign y9216 = ~n24782 ;
  assign y9217 = ~n24784 ;
  assign y9218 = n24788 ;
  assign y9219 = ~1'b0 ;
  assign y9220 = ~n24791 ;
  assign y9221 = ~n24794 ;
  assign y9222 = n24795 ;
  assign y9223 = n24798 ;
  assign y9224 = ~1'b0 ;
  assign y9225 = n24800 ;
  assign y9226 = n24802 ;
  assign y9227 = ~n24805 ;
  assign y9228 = ~1'b0 ;
  assign y9229 = n24806 ;
  assign y9230 = ~n24812 ;
  assign y9231 = ~n1226 ;
  assign y9232 = n24815 ;
  assign y9233 = ~n24821 ;
  assign y9234 = ~1'b0 ;
  assign y9235 = ~1'b0 ;
  assign y9236 = ~n24825 ;
  assign y9237 = ~1'b0 ;
  assign y9238 = ~n10161 ;
  assign y9239 = n24827 ;
  assign y9240 = ~n24829 ;
  assign y9241 = ~n24831 ;
  assign y9242 = ~n24832 ;
  assign y9243 = ~1'b0 ;
  assign y9244 = ~n24833 ;
  assign y9245 = ~1'b0 ;
  assign y9246 = n24834 ;
  assign y9247 = ~n24836 ;
  assign y9248 = n24838 ;
  assign y9249 = ~n24845 ;
  assign y9250 = ~n24846 ;
  assign y9251 = 1'b0 ;
  assign y9252 = n24849 ;
  assign y9253 = ~1'b0 ;
  assign y9254 = ~n24851 ;
  assign y9255 = n24854 ;
  assign y9256 = ~1'b0 ;
  assign y9257 = ~n24855 ;
  assign y9258 = ~1'b0 ;
  assign y9259 = n24856 ;
  assign y9260 = ~n24857 ;
  assign y9261 = ~1'b0 ;
  assign y9262 = ~1'b0 ;
  assign y9263 = n24858 ;
  assign y9264 = ~1'b0 ;
  assign y9265 = n24860 ;
  assign y9266 = n24867 ;
  assign y9267 = n24872 ;
  assign y9268 = n24875 ;
  assign y9269 = n24877 ;
  assign y9270 = ~1'b0 ;
  assign y9271 = ~n24878 ;
  assign y9272 = ~1'b0 ;
  assign y9273 = ~n15300 ;
  assign y9274 = n24880 ;
  assign y9275 = n24882 ;
  assign y9276 = n24883 ;
  assign y9277 = n24886 ;
  assign y9278 = n24895 ;
  assign y9279 = ~n24896 ;
  assign y9280 = ~n24899 ;
  assign y9281 = ~n24900 ;
  assign y9282 = ~n24901 ;
  assign y9283 = ~n24904 ;
  assign y9284 = ~n24906 ;
  assign y9285 = ~n24908 ;
  assign y9286 = ~n24912 ;
  assign y9287 = n24916 ;
  assign y9288 = n24917 ;
  assign y9289 = ~n24919 ;
  assign y9290 = ~n24920 ;
  assign y9291 = n24921 ;
  assign y9292 = n24924 ;
  assign y9293 = ~n24928 ;
  assign y9294 = ~n24933 ;
  assign y9295 = ~1'b0 ;
  assign y9296 = ~1'b0 ;
  assign y9297 = n24934 ;
  assign y9298 = ~1'b0 ;
  assign y9299 = ~n24936 ;
  assign y9300 = n24938 ;
  assign y9301 = ~n24939 ;
  assign y9302 = n24940 ;
  assign y9303 = ~n24943 ;
  assign y9304 = n24945 ;
  assign y9305 = n24949 ;
  assign y9306 = n24950 ;
  assign y9307 = ~n24951 ;
  assign y9308 = n24953 ;
  assign y9309 = ~n24954 ;
  assign y9310 = ~n24960 ;
  assign y9311 = ~n24961 ;
  assign y9312 = ~n24962 ;
  assign y9313 = n24964 ;
  assign y9314 = ~1'b0 ;
  assign y9315 = ~n24970 ;
  assign y9316 = ~n24972 ;
  assign y9317 = n24974 ;
  assign y9318 = 1'b0 ;
  assign y9319 = ~1'b0 ;
  assign y9320 = n24975 ;
  assign y9321 = ~1'b0 ;
  assign y9322 = ~n24977 ;
  assign y9323 = ~n24982 ;
  assign y9324 = ~1'b0 ;
  assign y9325 = ~1'b0 ;
  assign y9326 = ~1'b0 ;
  assign y9327 = n24984 ;
  assign y9328 = n24987 ;
  assign y9329 = ~n24991 ;
  assign y9330 = n24992 ;
  assign y9331 = ~n24995 ;
  assign y9332 = ~n24997 ;
  assign y9333 = n25000 ;
  assign y9334 = ~1'b0 ;
  assign y9335 = n25003 ;
  assign y9336 = n25005 ;
  assign y9337 = n25012 ;
  assign y9338 = n25013 ;
  assign y9339 = ~n25014 ;
  assign y9340 = ~1'b0 ;
  assign y9341 = n25015 ;
  assign y9342 = ~1'b0 ;
  assign y9343 = ~n25020 ;
  assign y9344 = ~n25029 ;
  assign y9345 = ~n25032 ;
  assign y9346 = n25033 ;
  assign y9347 = n25034 ;
  assign y9348 = n25037 ;
  assign y9349 = ~1'b0 ;
  assign y9350 = ~1'b0 ;
  assign y9351 = n25038 ;
  assign y9352 = ~n25042 ;
  assign y9353 = n25044 ;
  assign y9354 = n25049 ;
  assign y9355 = ~n25051 ;
  assign y9356 = ~1'b0 ;
  assign y9357 = ~1'b0 ;
  assign y9358 = ~n25056 ;
  assign y9359 = n25058 ;
  assign y9360 = n25060 ;
  assign y9361 = ~n25065 ;
  assign y9362 = ~n25072 ;
  assign y9363 = n25075 ;
  assign y9364 = n25079 ;
  assign y9365 = ~n25082 ;
  assign y9366 = ~n25083 ;
  assign y9367 = n25088 ;
  assign y9368 = n25092 ;
  assign y9369 = ~n25094 ;
  assign y9370 = ~n25095 ;
  assign y9371 = ~n25096 ;
  assign y9372 = n25099 ;
  assign y9373 = ~n25100 ;
  assign y9374 = ~n25102 ;
  assign y9375 = ~1'b0 ;
  assign y9376 = n25106 ;
  assign y9377 = ~1'b0 ;
  assign y9378 = ~n25108 ;
  assign y9379 = n25109 ;
  assign y9380 = 1'b0 ;
  assign y9381 = ~n25110 ;
  assign y9382 = ~n25111 ;
  assign y9383 = ~n25112 ;
  assign y9384 = ~n25114 ;
  assign y9385 = ~1'b0 ;
  assign y9386 = n25116 ;
  assign y9387 = n25121 ;
  assign y9388 = n25124 ;
  assign y9389 = ~n25133 ;
  assign y9390 = n25135 ;
  assign y9391 = ~1'b0 ;
  assign y9392 = n25136 ;
  assign y9393 = ~n25138 ;
  assign y9394 = n25140 ;
  assign y9395 = ~n25141 ;
  assign y9396 = ~n25142 ;
  assign y9397 = 1'b0 ;
  assign y9398 = ~n25149 ;
  assign y9399 = ~n25152 ;
  assign y9400 = ~1'b0 ;
  assign y9401 = n25154 ;
  assign y9402 = ~n25156 ;
  assign y9403 = n25157 ;
  assign y9404 = n25159 ;
  assign y9405 = n25160 ;
  assign y9406 = ~n25162 ;
  assign y9407 = ~1'b0 ;
  assign y9408 = n25166 ;
  assign y9409 = ~n25170 ;
  assign y9410 = n25172 ;
  assign y9411 = ~n25176 ;
  assign y9412 = n25180 ;
  assign y9413 = n25184 ;
  assign y9414 = ~n25186 ;
  assign y9415 = n25189 ;
  assign y9416 = ~1'b0 ;
  assign y9417 = n25196 ;
  assign y9418 = ~1'b0 ;
  assign y9419 = ~1'b0 ;
  assign y9420 = ~n25197 ;
  assign y9421 = ~n25200 ;
  assign y9422 = n25201 ;
  assign y9423 = ~n25202 ;
  assign y9424 = ~1'b0 ;
  assign y9425 = ~n25203 ;
  assign y9426 = ~n1955 ;
  assign y9427 = ~n25204 ;
  assign y9428 = ~1'b0 ;
  assign y9429 = ~n12389 ;
  assign y9430 = n11242 ;
  assign y9431 = ~n25207 ;
  assign y9432 = n25208 ;
  assign y9433 = ~n25209 ;
  assign y9434 = ~1'b0 ;
  assign y9435 = ~1'b0 ;
  assign y9436 = ~1'b0 ;
  assign y9437 = ~1'b0 ;
  assign y9438 = n25211 ;
  assign y9439 = n25218 ;
  assign y9440 = n25220 ;
  assign y9441 = n25221 ;
  assign y9442 = n25222 ;
  assign y9443 = ~n25228 ;
  assign y9444 = ~1'b0 ;
  assign y9445 = ~1'b0 ;
  assign y9446 = ~1'b0 ;
  assign y9447 = ~n25229 ;
  assign y9448 = ~n25236 ;
  assign y9449 = ~n25237 ;
  assign y9450 = ~n25239 ;
  assign y9451 = n25241 ;
  assign y9452 = n25243 ;
  assign y9453 = ~1'b0 ;
  assign y9454 = n25245 ;
  assign y9455 = ~1'b0 ;
  assign y9456 = n25247 ;
  assign y9457 = n25259 ;
  assign y9458 = ~1'b0 ;
  assign y9459 = n25260 ;
  assign y9460 = ~n25273 ;
  assign y9461 = n25274 ;
  assign y9462 = n25281 ;
  assign y9463 = ~n25292 ;
  assign y9464 = n25295 ;
  assign y9465 = ~1'b0 ;
  assign y9466 = ~n25298 ;
  assign y9467 = ~n25301 ;
  assign y9468 = ~n25302 ;
  assign y9469 = n25305 ;
  assign y9470 = n1587 ;
  assign y9471 = n25307 ;
  assign y9472 = ~n25311 ;
  assign y9473 = ~n25314 ;
  assign y9474 = n25316 ;
  assign y9475 = ~n25318 ;
  assign y9476 = ~n25321 ;
  assign y9477 = n25323 ;
  assign y9478 = ~n21025 ;
  assign y9479 = n25324 ;
  assign y9480 = ~n25327 ;
  assign y9481 = ~n25330 ;
  assign y9482 = ~1'b0 ;
  assign y9483 = n25331 ;
  assign y9484 = ~1'b0 ;
  assign y9485 = n25333 ;
  assign y9486 = ~n25334 ;
  assign y9487 = ~n25340 ;
  assign y9488 = n25341 ;
  assign y9489 = ~n25342 ;
  assign y9490 = ~1'b0 ;
  assign y9491 = n25349 ;
  assign y9492 = ~n25351 ;
  assign y9493 = ~n25352 ;
  assign y9494 = n25353 ;
  assign y9495 = ~n25355 ;
  assign y9496 = n25357 ;
  assign y9497 = n25358 ;
  assign y9498 = n25359 ;
  assign y9499 = ~n25361 ;
  assign y9500 = ~n14591 ;
  assign y9501 = ~1'b0 ;
  assign y9502 = n25365 ;
  assign y9503 = ~1'b0 ;
  assign y9504 = n25369 ;
  assign y9505 = ~n25370 ;
  assign y9506 = n25371 ;
  assign y9507 = ~1'b0 ;
  assign y9508 = n25374 ;
  assign y9509 = n25378 ;
  assign y9510 = ~n25382 ;
  assign y9511 = ~n25384 ;
  assign y9512 = n25389 ;
  assign y9513 = n25390 ;
  assign y9514 = ~n25394 ;
  assign y9515 = ~n25395 ;
  assign y9516 = n25403 ;
  assign y9517 = ~n25404 ;
  assign y9518 = ~1'b0 ;
  assign y9519 = n25406 ;
  assign y9520 = ~n4000 ;
  assign y9521 = 1'b0 ;
  assign y9522 = ~n25409 ;
  assign y9523 = n25410 ;
  assign y9524 = n25413 ;
  assign y9525 = ~1'b0 ;
  assign y9526 = n25418 ;
  assign y9527 = ~n25419 ;
  assign y9528 = n25422 ;
  assign y9529 = n25424 ;
  assign y9530 = ~n25425 ;
  assign y9531 = ~1'b0 ;
  assign y9532 = ~n25429 ;
  assign y9533 = n25430 ;
  assign y9534 = ~1'b0 ;
  assign y9535 = n25432 ;
  assign y9536 = ~n25434 ;
  assign y9537 = ~n25436 ;
  assign y9538 = n25437 ;
  assign y9539 = ~n25439 ;
  assign y9540 = ~n25440 ;
  assign y9541 = ~1'b0 ;
  assign y9542 = ~1'b0 ;
  assign y9543 = n25443 ;
  assign y9544 = ~n25446 ;
  assign y9545 = ~n25449 ;
  assign y9546 = ~n25450 ;
  assign y9547 = ~n25451 ;
  assign y9548 = ~n25454 ;
  assign y9549 = ~n25455 ;
  assign y9550 = ~1'b0 ;
  assign y9551 = ~1'b0 ;
  assign y9552 = ~1'b0 ;
  assign y9553 = n25457 ;
  assign y9554 = ~1'b0 ;
  assign y9555 = n25459 ;
  assign y9556 = n25462 ;
  assign y9557 = ~n25465 ;
  assign y9558 = n9829 ;
  assign y9559 = ~n25466 ;
  assign y9560 = n25467 ;
  assign y9561 = n25475 ;
  assign y9562 = ~n25476 ;
  assign y9563 = n25478 ;
  assign y9564 = n25482 ;
  assign y9565 = ~n25491 ;
  assign y9566 = ~n25496 ;
  assign y9567 = n25497 ;
  assign y9568 = n25499 ;
  assign y9569 = n25501 ;
  assign y9570 = ~1'b0 ;
  assign y9571 = ~n25505 ;
  assign y9572 = ~1'b0 ;
  assign y9573 = ~1'b0 ;
  assign y9574 = ~1'b0 ;
  assign y9575 = ~n25506 ;
  assign y9576 = ~n25508 ;
  assign y9577 = ~n25509 ;
  assign y9578 = n25511 ;
  assign y9579 = ~n25512 ;
  assign y9580 = ~1'b0 ;
  assign y9581 = ~1'b0 ;
  assign y9582 = ~n25513 ;
  assign y9583 = ~1'b0 ;
  assign y9584 = ~1'b0 ;
  assign y9585 = n25515 ;
  assign y9586 = ~n25522 ;
  assign y9587 = ~n25523 ;
  assign y9588 = ~n25524 ;
  assign y9589 = ~n25529 ;
  assign y9590 = ~n25533 ;
  assign y9591 = ~1'b0 ;
  assign y9592 = n25539 ;
  assign y9593 = n25541 ;
  assign y9594 = ~1'b0 ;
  assign y9595 = n25544 ;
  assign y9596 = n25547 ;
  assign y9597 = n25548 ;
  assign y9598 = ~n25549 ;
  assign y9599 = n25553 ;
  assign y9600 = ~n25555 ;
  assign y9601 = n25559 ;
  assign y9602 = ~n25565 ;
  assign y9603 = ~n25566 ;
  assign y9604 = ~n25567 ;
  assign y9605 = ~n25569 ;
  assign y9606 = ~n25570 ;
  assign y9607 = ~n25571 ;
  assign y9608 = ~1'b0 ;
  assign y9609 = ~1'b0 ;
  assign y9610 = n25572 ;
  assign y9611 = ~n25575 ;
  assign y9612 = ~n25580 ;
  assign y9613 = n25581 ;
  assign y9614 = n25582 ;
  assign y9615 = n25584 ;
  assign y9616 = n25588 ;
  assign y9617 = ~n25591 ;
  assign y9618 = ~1'b0 ;
  assign y9619 = n25594 ;
  assign y9620 = ~1'b0 ;
  assign y9621 = ~1'b0 ;
  assign y9622 = n25600 ;
  assign y9623 = ~n25601 ;
  assign y9624 = ~n25614 ;
  assign y9625 = ~n25615 ;
  assign y9626 = n22080 ;
  assign y9627 = ~n25619 ;
  assign y9628 = n25623 ;
  assign y9629 = ~1'b0 ;
  assign y9630 = ~n25626 ;
  assign y9631 = ~n15256 ;
  assign y9632 = n25627 ;
  assign y9633 = ~n25629 ;
  assign y9634 = ~n25631 ;
  assign y9635 = ~n25633 ;
  assign y9636 = ~1'b0 ;
  assign y9637 = ~n25640 ;
  assign y9638 = ~n25644 ;
  assign y9639 = n25652 ;
  assign y9640 = ~n25653 ;
  assign y9641 = ~n25655 ;
  assign y9642 = ~n25656 ;
  assign y9643 = ~n25657 ;
  assign y9644 = ~n25658 ;
  assign y9645 = ~1'b0 ;
  assign y9646 = n25663 ;
  assign y9647 = n25667 ;
  assign y9648 = ~n25672 ;
  assign y9649 = ~1'b0 ;
  assign y9650 = ~n25674 ;
  assign y9651 = n25678 ;
  assign y9652 = ~n23084 ;
  assign y9653 = n25682 ;
  assign y9654 = n25683 ;
  assign y9655 = ~n25686 ;
  assign y9656 = n25687 ;
  assign y9657 = n25689 ;
  assign y9658 = n25690 ;
  assign y9659 = ~1'b0 ;
  assign y9660 = ~1'b0 ;
  assign y9661 = n25693 ;
  assign y9662 = ~n25695 ;
  assign y9663 = n25699 ;
  assign y9664 = ~n25703 ;
  assign y9665 = ~1'b0 ;
  assign y9666 = ~1'b0 ;
  assign y9667 = n25706 ;
  assign y9668 = n25710 ;
  assign y9669 = ~1'b0 ;
  assign y9670 = n25712 ;
  assign y9671 = n25713 ;
  assign y9672 = ~n25718 ;
  assign y9673 = ~n25719 ;
  assign y9674 = n25720 ;
  assign y9675 = ~1'b0 ;
  assign y9676 = ~n25721 ;
  assign y9677 = n9765 ;
  assign y9678 = n25722 ;
  assign y9679 = ~n25723 ;
  assign y9680 = ~n25730 ;
  assign y9681 = n25731 ;
  assign y9682 = ~n25734 ;
  assign y9683 = ~1'b0 ;
  assign y9684 = ~1'b0 ;
  assign y9685 = ~n25739 ;
  assign y9686 = ~n25741 ;
  assign y9687 = n25747 ;
  assign y9688 = ~n25750 ;
  assign y9689 = ~n25752 ;
  assign y9690 = n25756 ;
  assign y9691 = ~n25759 ;
  assign y9692 = n25761 ;
  assign y9693 = ~n25764 ;
  assign y9694 = n25767 ;
  assign y9695 = n25770 ;
  assign y9696 = ~1'b0 ;
  assign y9697 = ~n25774 ;
  assign y9698 = n25775 ;
  assign y9699 = ~n25777 ;
  assign y9700 = n25780 ;
  assign y9701 = ~n25781 ;
  assign y9702 = n25784 ;
  assign y9703 = ~1'b0 ;
  assign y9704 = ~1'b0 ;
  assign y9705 = ~n25789 ;
  assign y9706 = ~n25792 ;
  assign y9707 = ~n25798 ;
  assign y9708 = ~n25800 ;
  assign y9709 = n25801 ;
  assign y9710 = n2509 ;
  assign y9711 = n25803 ;
  assign y9712 = ~n25811 ;
  assign y9713 = ~n25814 ;
  assign y9714 = n25819 ;
  assign y9715 = ~1'b0 ;
  assign y9716 = ~n25821 ;
  assign y9717 = ~1'b0 ;
  assign y9718 = n1811 ;
  assign y9719 = n25823 ;
  assign y9720 = n25824 ;
  assign y9721 = ~n25825 ;
  assign y9722 = ~n25828 ;
  assign y9723 = n25829 ;
  assign y9724 = n25831 ;
  assign y9725 = ~n25838 ;
  assign y9726 = ~1'b0 ;
  assign y9727 = ~n25840 ;
  assign y9728 = ~1'b0 ;
  assign y9729 = ~n25841 ;
  assign y9730 = n25842 ;
  assign y9731 = ~n25843 ;
  assign y9732 = n25849 ;
  assign y9733 = n25850 ;
  assign y9734 = n25852 ;
  assign y9735 = n25853 ;
  assign y9736 = ~n25862 ;
  assign y9737 = ~1'b0 ;
  assign y9738 = ~1'b0 ;
  assign y9739 = ~n25865 ;
  assign y9740 = ~n25867 ;
  assign y9741 = ~n25868 ;
  assign y9742 = ~n25871 ;
  assign y9743 = ~1'b0 ;
  assign y9744 = n10434 ;
  assign y9745 = ~n25874 ;
  assign y9746 = n25877 ;
  assign y9747 = ~1'b0 ;
  assign y9748 = ~1'b0 ;
  assign y9749 = ~1'b0 ;
  assign y9750 = ~n25878 ;
  assign y9751 = ~n25879 ;
  assign y9752 = ~n25881 ;
  assign y9753 = n25885 ;
  assign y9754 = ~n25888 ;
  assign y9755 = ~n25891 ;
  assign y9756 = n3481 ;
  assign y9757 = n25896 ;
  assign y9758 = ~n25897 ;
  assign y9759 = n25898 ;
  assign y9760 = n25899 ;
  assign y9761 = n25904 ;
  assign y9762 = n25907 ;
  assign y9763 = ~n25911 ;
  assign y9764 = n25913 ;
  assign y9765 = ~1'b0 ;
  assign y9766 = n25918 ;
  assign y9767 = n25919 ;
  assign y9768 = n25922 ;
  assign y9769 = n25923 ;
  assign y9770 = ~n25926 ;
  assign y9771 = ~n25928 ;
  assign y9772 = ~1'b0 ;
  assign y9773 = ~n25929 ;
  assign y9774 = n25931 ;
  assign y9775 = n25935 ;
  assign y9776 = n25939 ;
  assign y9777 = n25942 ;
  assign y9778 = n25944 ;
  assign y9779 = ~n25946 ;
  assign y9780 = n25950 ;
  assign y9781 = ~1'b0 ;
  assign y9782 = ~1'b0 ;
  assign y9783 = n25954 ;
  assign y9784 = n6293 ;
  assign y9785 = ~n25956 ;
  assign y9786 = n25957 ;
  assign y9787 = n25959 ;
  assign y9788 = n25961 ;
  assign y9789 = n25968 ;
  assign y9790 = ~n25969 ;
  assign y9791 = n25971 ;
  assign y9792 = ~1'b0 ;
  assign y9793 = n25973 ;
  assign y9794 = ~n25974 ;
  assign y9795 = n25975 ;
  assign y9796 = n25977 ;
  assign y9797 = ~n25986 ;
  assign y9798 = ~n25989 ;
  assign y9799 = ~1'b0 ;
  assign y9800 = ~n25994 ;
  assign y9801 = ~1'b0 ;
  assign y9802 = ~n25995 ;
  assign y9803 = ~1'b0 ;
  assign y9804 = n25996 ;
  assign y9805 = n25997 ;
  assign y9806 = n25998 ;
  assign y9807 = n25999 ;
  assign y9808 = ~1'b0 ;
  assign y9809 = n26001 ;
  assign y9810 = ~n26003 ;
  assign y9811 = ~1'b0 ;
  assign y9812 = ~n26005 ;
  assign y9813 = ~n19945 ;
  assign y9814 = ~n26008 ;
  assign y9815 = ~n26009 ;
  assign y9816 = ~1'b0 ;
  assign y9817 = ~n10819 ;
  assign y9818 = ~1'b0 ;
  assign y9819 = n26011 ;
  assign y9820 = n26015 ;
  assign y9821 = ~1'b0 ;
  assign y9822 = ~n26021 ;
  assign y9823 = n26024 ;
  assign y9824 = ~1'b0 ;
  assign y9825 = n26030 ;
  assign y9826 = ~n26031 ;
  assign y9827 = ~1'b0 ;
  assign y9828 = ~1'b0 ;
  assign y9829 = n26033 ;
  assign y9830 = n26034 ;
  assign y9831 = n26035 ;
  assign y9832 = n26038 ;
  assign y9833 = n26040 ;
  assign y9834 = n26044 ;
  assign y9835 = n26046 ;
  assign y9836 = ~1'b0 ;
  assign y9837 = ~n26051 ;
  assign y9838 = ~n26062 ;
  assign y9839 = ~n26064 ;
  assign y9840 = n26065 ;
  assign y9841 = n26068 ;
  assign y9842 = ~n26070 ;
  assign y9843 = n26073 ;
  assign y9844 = n26074 ;
  assign y9845 = ~n26076 ;
  assign y9846 = ~1'b0 ;
  assign y9847 = ~n26078 ;
  assign y9848 = 1'b0 ;
  assign y9849 = ~n26081 ;
  assign y9850 = ~n26085 ;
  assign y9851 = n26088 ;
  assign y9852 = n26089 ;
  assign y9853 = n26090 ;
  assign y9854 = n26092 ;
  assign y9855 = n26093 ;
  assign y9856 = n26098 ;
  assign y9857 = n26099 ;
  assign y9858 = ~1'b0 ;
  assign y9859 = ~1'b0 ;
  assign y9860 = ~1'b0 ;
  assign y9861 = n26100 ;
  assign y9862 = n26101 ;
  assign y9863 = n26105 ;
  assign y9864 = n26106 ;
  assign y9865 = ~n26108 ;
  assign y9866 = ~n26111 ;
  assign y9867 = ~1'b0 ;
  assign y9868 = n26112 ;
  assign y9869 = ~n26113 ;
  assign y9870 = n26114 ;
  assign y9871 = ~1'b0 ;
  assign y9872 = ~n26115 ;
  assign y9873 = n26118 ;
  assign y9874 = ~n26125 ;
  assign y9875 = ~n26126 ;
  assign y9876 = ~1'b0 ;
  assign y9877 = ~n26127 ;
  assign y9878 = ~1'b0 ;
  assign y9879 = ~n26132 ;
  assign y9880 = ~1'b0 ;
  assign y9881 = ~n6366 ;
  assign y9882 = n26136 ;
  assign y9883 = n26138 ;
  assign y9884 = ~n26140 ;
  assign y9885 = ~1'b0 ;
  assign y9886 = ~n26142 ;
  assign y9887 = ~1'b0 ;
  assign y9888 = ~1'b0 ;
  assign y9889 = n26144 ;
  assign y9890 = ~n26147 ;
  assign y9891 = ~n26150 ;
  assign y9892 = ~n26151 ;
  assign y9893 = n26153 ;
  assign y9894 = ~1'b0 ;
  assign y9895 = n26157 ;
  assign y9896 = ~1'b0 ;
  assign y9897 = ~n26159 ;
  assign y9898 = n26162 ;
  assign y9899 = ~n26164 ;
  assign y9900 = ~n26170 ;
  assign y9901 = n26171 ;
  assign y9902 = ~n26176 ;
  assign y9903 = ~n26177 ;
  assign y9904 = ~n26181 ;
  assign y9905 = n26185 ;
  assign y9906 = ~n26187 ;
  assign y9907 = n26188 ;
  assign y9908 = ~n26189 ;
  assign y9909 = n26190 ;
  assign y9910 = ~n26194 ;
  assign y9911 = ~1'b0 ;
  assign y9912 = n26195 ;
  assign y9913 = n26197 ;
  assign y9914 = ~n26201 ;
  assign y9915 = ~n26202 ;
  assign y9916 = ~n26205 ;
  assign y9917 = ~1'b0 ;
  assign y9918 = ~n26207 ;
  assign y9919 = ~n26209 ;
  assign y9920 = n26212 ;
  assign y9921 = ~1'b0 ;
  assign y9922 = n26215 ;
  assign y9923 = n26219 ;
  assign y9924 = n26220 ;
  assign y9925 = n26225 ;
  assign y9926 = n26226 ;
  assign y9927 = ~n26228 ;
  assign y9928 = ~n26229 ;
  assign y9929 = ~1'b0 ;
  assign y9930 = n26231 ;
  assign y9931 = ~n26232 ;
  assign y9932 = n26235 ;
  assign y9933 = n26239 ;
  assign y9934 = n26242 ;
  assign y9935 = ~n26245 ;
  assign y9936 = ~1'b0 ;
  assign y9937 = ~n26246 ;
  assign y9938 = ~1'b0 ;
  assign y9939 = n26248 ;
  assign y9940 = n26250 ;
  assign y9941 = ~1'b0 ;
  assign y9942 = n26251 ;
  assign y9943 = n26253 ;
  assign y9944 = ~n26254 ;
  assign y9945 = ~n26256 ;
  assign y9946 = ~n26257 ;
  assign y9947 = ~n26260 ;
  assign y9948 = ~n26262 ;
  assign y9949 = ~n26264 ;
  assign y9950 = n26268 ;
  assign y9951 = ~1'b0 ;
  assign y9952 = n26270 ;
  assign y9953 = ~n26272 ;
  assign y9954 = n26273 ;
  assign y9955 = n26276 ;
  assign y9956 = ~n26282 ;
  assign y9957 = ~n26287 ;
  assign y9958 = ~n26291 ;
  assign y9959 = n26295 ;
  assign y9960 = n26296 ;
  assign y9961 = ~n26299 ;
  assign y9962 = n26302 ;
  assign y9963 = n26307 ;
  assign y9964 = ~n26309 ;
  assign y9965 = ~n26310 ;
  assign y9966 = n26317 ;
  assign y9967 = ~n26318 ;
  assign y9968 = ~n26327 ;
  assign y9969 = ~1'b0 ;
  assign y9970 = n26329 ;
  assign y9971 = ~n26333 ;
  assign y9972 = ~n26335 ;
  assign y9973 = ~n26336 ;
  assign y9974 = n26337 ;
  assign y9975 = n26340 ;
  assign y9976 = ~n26341 ;
  assign y9977 = ~n26345 ;
  assign y9978 = ~n26348 ;
  assign y9979 = ~n26350 ;
  assign y9980 = ~1'b0 ;
  assign y9981 = ~n26351 ;
  assign y9982 = ~n26352 ;
  assign y9983 = ~1'b0 ;
  assign y9984 = n26353 ;
  assign y9985 = n26355 ;
  assign y9986 = ~n26358 ;
  assign y9987 = ~1'b0 ;
  assign y9988 = ~n26360 ;
  assign y9989 = n26361 ;
  assign y9990 = ~n26363 ;
  assign y9991 = n26364 ;
  assign y9992 = n26366 ;
  assign y9993 = n26370 ;
  assign y9994 = n26374 ;
  assign y9995 = n26376 ;
  assign y9996 = ~n26379 ;
  assign y9997 = n26381 ;
  assign y9998 = ~1'b0 ;
  assign y9999 = ~n26385 ;
  assign y10000 = ~n26389 ;
  assign y10001 = ~n26393 ;
  assign y10002 = ~n26394 ;
  assign y10003 = n26395 ;
  assign y10004 = n1654 ;
  assign y10005 = ~n26398 ;
  assign y10006 = ~n26399 ;
  assign y10007 = ~n26401 ;
  assign y10008 = n26403 ;
  assign y10009 = n26404 ;
  assign y10010 = n26406 ;
  assign y10011 = ~n26409 ;
  assign y10012 = n26410 ;
  assign y10013 = n26412 ;
  assign y10014 = n26419 ;
  assign y10015 = ~n26421 ;
  assign y10016 = n26422 ;
  assign y10017 = n26424 ;
  assign y10018 = n26426 ;
  assign y10019 = ~n26428 ;
  assign y10020 = ~n26435 ;
  assign y10021 = ~n26439 ;
  assign y10022 = ~n26440 ;
  assign y10023 = ~n26441 ;
  assign y10024 = n26445 ;
  assign y10025 = n26448 ;
  assign y10026 = n26449 ;
  assign y10027 = ~1'b0 ;
  assign y10028 = n26451 ;
  assign y10029 = n26458 ;
  assign y10030 = n26462 ;
  assign y10031 = n4684 ;
  assign y10032 = ~n26465 ;
  assign y10033 = ~n26467 ;
  assign y10034 = n26468 ;
  assign y10035 = ~1'b0 ;
  assign y10036 = ~1'b0 ;
  assign y10037 = ~1'b0 ;
  assign y10038 = n26469 ;
  assign y10039 = ~1'b0 ;
  assign y10040 = n26477 ;
  assign y10041 = n26478 ;
  assign y10042 = n26484 ;
  assign y10043 = ~1'b0 ;
  assign y10044 = n26486 ;
  assign y10045 = n26487 ;
  assign y10046 = ~1'b0 ;
  assign y10047 = n26491 ;
  assign y10048 = ~n26492 ;
  assign y10049 = ~n26494 ;
  assign y10050 = ~n26497 ;
  assign y10051 = ~n16765 ;
  assign y10052 = ~n26502 ;
  assign y10053 = ~1'b0 ;
  assign y10054 = ~n26505 ;
  assign y10055 = ~1'b0 ;
  assign y10056 = ~1'b0 ;
  assign y10057 = ~n26508 ;
  assign y10058 = n26509 ;
  assign y10059 = n26514 ;
  assign y10060 = n26518 ;
  assign y10061 = ~n26519 ;
  assign y10062 = ~1'b0 ;
  assign y10063 = n26521 ;
  assign y10064 = ~1'b0 ;
  assign y10065 = ~1'b0 ;
  assign y10066 = ~n26526 ;
  assign y10067 = n26530 ;
  assign y10068 = n26533 ;
  assign y10069 = ~n26535 ;
  assign y10070 = n26540 ;
  assign y10071 = ~n26542 ;
  assign y10072 = ~n26546 ;
  assign y10073 = ~1'b0 ;
  assign y10074 = ~1'b0 ;
  assign y10075 = ~n26548 ;
  assign y10076 = ~n26550 ;
  assign y10077 = ~n26553 ;
  assign y10078 = n26555 ;
  assign y10079 = n26560 ;
  assign y10080 = ~n26563 ;
  assign y10081 = n26569 ;
  assign y10082 = ~n4714 ;
  assign y10083 = 1'b0 ;
  assign y10084 = ~1'b0 ;
  assign y10085 = ~1'b0 ;
  assign y10086 = n26570 ;
  assign y10087 = ~n26572 ;
  assign y10088 = ~n26575 ;
  assign y10089 = ~n26577 ;
  assign y10090 = ~n26580 ;
  assign y10091 = ~n26582 ;
  assign y10092 = ~n26587 ;
  assign y10093 = ~n26589 ;
  assign y10094 = n26591 ;
  assign y10095 = n26595 ;
  assign y10096 = n26596 ;
  assign y10097 = ~n26597 ;
  assign y10098 = n26601 ;
  assign y10099 = n26602 ;
  assign y10100 = n26603 ;
  assign y10101 = ~n26607 ;
  assign y10102 = ~n26609 ;
  assign y10103 = ~n26613 ;
  assign y10104 = ~1'b0 ;
  assign y10105 = ~1'b0 ;
  assign y10106 = n26616 ;
  assign y10107 = n26617 ;
  assign y10108 = ~n26619 ;
  assign y10109 = n26621 ;
  assign y10110 = ~1'b0 ;
  assign y10111 = ~n26623 ;
  assign y10112 = n26624 ;
  assign y10113 = n26625 ;
  assign y10114 = n26630 ;
  assign y10115 = ~n26632 ;
  assign y10116 = ~n26633 ;
  assign y10117 = ~n26634 ;
  assign y10118 = ~1'b0 ;
  assign y10119 = ~n26637 ;
  assign y10120 = ~1'b0 ;
  assign y10121 = ~1'b0 ;
  assign y10122 = ~n26642 ;
  assign y10123 = n26646 ;
  assign y10124 = ~n26651 ;
  assign y10125 = n26653 ;
  assign y10126 = n26654 ;
  assign y10127 = ~1'b0 ;
  assign y10128 = ~1'b0 ;
  assign y10129 = ~n26656 ;
  assign y10130 = n26658 ;
  assign y10131 = n26659 ;
  assign y10132 = ~n26661 ;
  assign y10133 = n26662 ;
  assign y10134 = ~n26663 ;
  assign y10135 = n26665 ;
  assign y10136 = n26668 ;
  assign y10137 = ~1'b0 ;
  assign y10138 = ~1'b0 ;
  assign y10139 = ~n3858 ;
  assign y10140 = ~n26669 ;
  assign y10141 = n26671 ;
  assign y10142 = ~n26673 ;
  assign y10143 = ~n26674 ;
  assign y10144 = ~n26677 ;
  assign y10145 = n26679 ;
  assign y10146 = ~n3706 ;
  assign y10147 = ~n26683 ;
  assign y10148 = ~1'b0 ;
  assign y10149 = n26686 ;
  assign y10150 = n26687 ;
  assign y10151 = n26688 ;
  assign y10152 = ~n26689 ;
  assign y10153 = n26695 ;
  assign y10154 = ~1'b0 ;
  assign y10155 = ~n26697 ;
  assign y10156 = n26701 ;
  assign y10157 = ~n26703 ;
  assign y10158 = ~n26704 ;
  assign y10159 = ~n3971 ;
  assign y10160 = n26707 ;
  assign y10161 = ~n26711 ;
  assign y10162 = ~n26713 ;
  assign y10163 = n26715 ;
  assign y10164 = n328 ;
  assign y10165 = ~1'b0 ;
  assign y10166 = n26717 ;
  assign y10167 = ~n26718 ;
  assign y10168 = n26725 ;
  assign y10169 = ~n26729 ;
  assign y10170 = ~1'b0 ;
  assign y10171 = ~n26731 ;
  assign y10172 = ~1'b0 ;
  assign y10173 = ~1'b0 ;
  assign y10174 = 1'b0 ;
  assign y10175 = ~n26733 ;
  assign y10176 = ~n26734 ;
  assign y10177 = ~n26738 ;
  assign y10178 = ~n26740 ;
  assign y10179 = ~n26741 ;
  assign y10180 = ~n26744 ;
  assign y10181 = ~n26747 ;
  assign y10182 = n26749 ;
  assign y10183 = n26753 ;
  assign y10184 = ~n26759 ;
  assign y10185 = ~n26761 ;
  assign y10186 = n26765 ;
  assign y10187 = 1'b0 ;
  assign y10188 = ~n26766 ;
  assign y10189 = n26767 ;
  assign y10190 = ~n26770 ;
  assign y10191 = ~1'b0 ;
  assign y10192 = n26774 ;
  assign y10193 = ~n26781 ;
  assign y10194 = n26784 ;
  assign y10195 = n26789 ;
  assign y10196 = ~1'b0 ;
  assign y10197 = ~n26791 ;
  assign y10198 = n26792 ;
  assign y10199 = n26797 ;
  assign y10200 = ~n26798 ;
  assign y10201 = ~n26802 ;
  assign y10202 = ~n26804 ;
  assign y10203 = n26807 ;
  assign y10204 = n26811 ;
  assign y10205 = ~n26813 ;
  assign y10206 = ~n26816 ;
  assign y10207 = n26820 ;
  assign y10208 = n26822 ;
  assign y10209 = n26826 ;
  assign y10210 = n23248 ;
  assign y10211 = ~n26831 ;
  assign y10212 = ~n26834 ;
  assign y10213 = ~1'b0 ;
  assign y10214 = ~n26840 ;
  assign y10215 = ~n26841 ;
  assign y10216 = n26842 ;
  assign y10217 = ~n26844 ;
  assign y10218 = ~1'b0 ;
  assign y10219 = 1'b0 ;
  assign y10220 = ~n26848 ;
  assign y10221 = ~1'b0 ;
  assign y10222 = ~1'b0 ;
  assign y10223 = n26850 ;
  assign y10224 = ~n26859 ;
  assign y10225 = n26861 ;
  assign y10226 = n26863 ;
  assign y10227 = ~n26864 ;
  assign y10228 = ~n17228 ;
  assign y10229 = n26865 ;
  assign y10230 = n26866 ;
  assign y10231 = ~n26867 ;
  assign y10232 = ~n26868 ;
  assign y10233 = ~n26871 ;
  assign y10234 = n26873 ;
  assign y10235 = n26878 ;
  assign y10236 = ~n26879 ;
  assign y10237 = n26882 ;
  assign y10238 = n26886 ;
  assign y10239 = n26888 ;
  assign y10240 = n26889 ;
  assign y10241 = ~1'b0 ;
  assign y10242 = ~n26890 ;
  assign y10243 = n26893 ;
  assign y10244 = ~n26896 ;
  assign y10245 = n26899 ;
  assign y10246 = n26903 ;
  assign y10247 = n26906 ;
  assign y10248 = ~1'b0 ;
  assign y10249 = ~n26913 ;
  assign y10250 = ~n26919 ;
  assign y10251 = ~n26921 ;
  assign y10252 = n26924 ;
  assign y10253 = ~n26926 ;
  assign y10254 = ~n26928 ;
  assign y10255 = n26931 ;
  assign y10256 = ~n26934 ;
  assign y10257 = 1'b0 ;
  assign y10258 = ~n26936 ;
  assign y10259 = ~n26938 ;
  assign y10260 = ~n26939 ;
  assign y10261 = ~n26943 ;
  assign y10262 = ~n26947 ;
  assign y10263 = n26955 ;
  assign y10264 = n26956 ;
  assign y10265 = n26959 ;
  assign y10266 = ~n26961 ;
  assign y10267 = n26962 ;
  assign y10268 = n26963 ;
  assign y10269 = ~1'b0 ;
  assign y10270 = n26966 ;
  assign y10271 = ~1'b0 ;
  assign y10272 = n26969 ;
  assign y10273 = ~n26970 ;
  assign y10274 = ~n26972 ;
  assign y10275 = ~n26973 ;
  assign y10276 = ~n6144 ;
  assign y10277 = ~n26976 ;
  assign y10278 = n26977 ;
  assign y10279 = n26980 ;
  assign y10280 = ~n26981 ;
  assign y10281 = ~n26982 ;
  assign y10282 = ~1'b0 ;
  assign y10283 = ~n26983 ;
  assign y10284 = ~n4971 ;
  assign y10285 = n26986 ;
  assign y10286 = ~n26990 ;
  assign y10287 = ~n26991 ;
  assign y10288 = n26993 ;
  assign y10289 = n26996 ;
  assign y10290 = ~1'b0 ;
  assign y10291 = n27001 ;
  assign y10292 = n27004 ;
  assign y10293 = ~n27006 ;
  assign y10294 = ~n27009 ;
  assign y10295 = ~n27010 ;
  assign y10296 = ~n27012 ;
  assign y10297 = ~n27014 ;
  assign y10298 = n27016 ;
  assign y10299 = ~n8217 ;
  assign y10300 = ~n27018 ;
  assign y10301 = ~1'b0 ;
  assign y10302 = ~n27022 ;
  assign y10303 = ~n27023 ;
  assign y10304 = ~n27024 ;
  assign y10305 = n27028 ;
  assign y10306 = ~n27030 ;
  assign y10307 = ~n27032 ;
  assign y10308 = ~1'b0 ;
  assign y10309 = ~n27034 ;
  assign y10310 = ~1'b0 ;
  assign y10311 = n27036 ;
  assign y10312 = ~n27039 ;
  assign y10313 = ~n27042 ;
  assign y10314 = n27047 ;
  assign y10315 = n27048 ;
  assign y10316 = n27049 ;
  assign y10317 = ~1'b0 ;
  assign y10318 = n27051 ;
  assign y10319 = ~n27057 ;
  assign y10320 = ~n27058 ;
  assign y10321 = ~1'b0 ;
  assign y10322 = ~1'b0 ;
  assign y10323 = ~n27059 ;
  assign y10324 = n27060 ;
  assign y10325 = ~n27061 ;
  assign y10326 = ~n27063 ;
  assign y10327 = ~n27069 ;
  assign y10328 = ~1'b0 ;
  assign y10329 = ~n27071 ;
  assign y10330 = ~n27075 ;
  assign y10331 = n27077 ;
  assign y10332 = n27078 ;
  assign y10333 = ~n27079 ;
  assign y10334 = n27083 ;
  assign y10335 = ~n27086 ;
  assign y10336 = ~n27088 ;
  assign y10337 = ~n27090 ;
  assign y10338 = n27097 ;
  assign y10339 = ~n27099 ;
  assign y10340 = ~n27103 ;
  assign y10341 = ~1'b0 ;
  assign y10342 = ~n27104 ;
  assign y10343 = ~n27108 ;
  assign y10344 = n27109 ;
  assign y10345 = ~n27115 ;
  assign y10346 = ~1'b0 ;
  assign y10347 = ~n27121 ;
  assign y10348 = n27123 ;
  assign y10349 = ~1'b0 ;
  assign y10350 = ~1'b0 ;
  assign y10351 = ~1'b0 ;
  assign y10352 = n27127 ;
  assign y10353 = ~n27128 ;
  assign y10354 = ~n27131 ;
  assign y10355 = ~1'b0 ;
  assign y10356 = ~n291 ;
  assign y10357 = ~n27136 ;
  assign y10358 = ~1'b0 ;
  assign y10359 = ~1'b0 ;
  assign y10360 = ~n27137 ;
  assign y10361 = n27139 ;
  assign y10362 = ~1'b0 ;
  assign y10363 = ~n8228 ;
  assign y10364 = ~n27140 ;
  assign y10365 = ~n27141 ;
  assign y10366 = n27146 ;
  assign y10367 = n27148 ;
  assign y10368 = n27151 ;
  assign y10369 = ~n27152 ;
  assign y10370 = ~n27153 ;
  assign y10371 = ~n27155 ;
  assign y10372 = ~n27156 ;
  assign y10373 = ~1'b0 ;
  assign y10374 = ~n27157 ;
  assign y10375 = ~n27159 ;
  assign y10376 = n27165 ;
  assign y10377 = n27170 ;
  assign y10378 = ~n27171 ;
  assign y10379 = ~n27174 ;
  assign y10380 = ~n27177 ;
  assign y10381 = ~1'b0 ;
  assign y10382 = n27179 ;
  assign y10383 = ~n27183 ;
  assign y10384 = n27184 ;
  assign y10385 = n27187 ;
  assign y10386 = n27190 ;
  assign y10387 = ~n27194 ;
  assign y10388 = ~1'b0 ;
  assign y10389 = ~1'b0 ;
  assign y10390 = ~1'b0 ;
  assign y10391 = ~1'b0 ;
  assign y10392 = ~n27196 ;
  assign y10393 = n27200 ;
  assign y10394 = ~n27202 ;
  assign y10395 = ~n27203 ;
  assign y10396 = n27205 ;
  assign y10397 = n27208 ;
  assign y10398 = n27210 ;
  assign y10399 = n27212 ;
  assign y10400 = ~n27214 ;
  assign y10401 = n27216 ;
  assign y10402 = ~1'b0 ;
  assign y10403 = ~1'b0 ;
  assign y10404 = n27220 ;
  assign y10405 = n27228 ;
  assign y10406 = n27230 ;
  assign y10407 = n27239 ;
  assign y10408 = ~n27240 ;
  assign y10409 = ~n27246 ;
  assign y10410 = ~n27250 ;
  assign y10411 = n27254 ;
  assign y10412 = n27257 ;
  assign y10413 = n27259 ;
  assign y10414 = ~n27261 ;
  assign y10415 = ~n27262 ;
  assign y10416 = n27264 ;
  assign y10417 = ~n27267 ;
  assign y10418 = ~n27268 ;
  assign y10419 = ~n27274 ;
  assign y10420 = n27275 ;
  assign y10421 = n27278 ;
  assign y10422 = ~1'b0 ;
  assign y10423 = ~1'b0 ;
  assign y10424 = ~1'b0 ;
  assign y10425 = n27279 ;
  assign y10426 = ~n27285 ;
  assign y10427 = ~n27289 ;
  assign y10428 = ~n27294 ;
  assign y10429 = ~n27295 ;
  assign y10430 = ~1'b0 ;
  assign y10431 = ~1'b0 ;
  assign y10432 = ~n27297 ;
  assign y10433 = ~n27302 ;
  assign y10434 = ~n27304 ;
  assign y10435 = ~n27307 ;
  assign y10436 = n27308 ;
  assign y10437 = n27311 ;
  assign y10438 = ~n27312 ;
  assign y10439 = ~n27318 ;
  assign y10440 = ~n27329 ;
  assign y10441 = ~1'b0 ;
  assign y10442 = n27330 ;
  assign y10443 = ~1'b0 ;
  assign y10444 = ~n27334 ;
  assign y10445 = ~n27347 ;
  assign y10446 = ~n27350 ;
  assign y10447 = n27352 ;
  assign y10448 = ~n27354 ;
  assign y10449 = ~n27359 ;
  assign y10450 = ~1'b0 ;
  assign y10451 = ~1'b0 ;
  assign y10452 = ~1'b0 ;
  assign y10453 = ~1'b0 ;
  assign y10454 = ~1'b0 ;
  assign y10455 = ~n27365 ;
  assign y10456 = n27366 ;
  assign y10457 = ~n27367 ;
  assign y10458 = ~n27369 ;
  assign y10459 = ~n27372 ;
  assign y10460 = n27376 ;
  assign y10461 = ~n27377 ;
  assign y10462 = n27379 ;
  assign y10463 = ~1'b0 ;
  assign y10464 = n27382 ;
  assign y10465 = n27385 ;
  assign y10466 = n27388 ;
  assign y10467 = ~n27391 ;
  assign y10468 = n27397 ;
  assign y10469 = n27398 ;
  assign y10470 = ~n27401 ;
  assign y10471 = ~1'b0 ;
  assign y10472 = ~n27404 ;
  assign y10473 = ~1'b0 ;
  assign y10474 = ~n27405 ;
  assign y10475 = ~1'b0 ;
  assign y10476 = ~1'b0 ;
  assign y10477 = ~n27406 ;
  assign y10478 = ~n27408 ;
  assign y10479 = n27410 ;
  assign y10480 = ~n27412 ;
  assign y10481 = n27414 ;
  assign y10482 = ~1'b0 ;
  assign y10483 = ~n27415 ;
  assign y10484 = n27416 ;
  assign y10485 = n27419 ;
  assign y10486 = ~n27421 ;
  assign y10487 = n27422 ;
  assign y10488 = n24536 ;
  assign y10489 = ~n27427 ;
  assign y10490 = n27431 ;
  assign y10491 = n27434 ;
  assign y10492 = ~1'b0 ;
  assign y10493 = ~1'b0 ;
  assign y10494 = ~n27441 ;
  assign y10495 = n27442 ;
  assign y10496 = ~n27443 ;
  assign y10497 = n27446 ;
  assign y10498 = n27448 ;
  assign y10499 = n27452 ;
  assign y10500 = n27454 ;
  assign y10501 = ~n27460 ;
  assign y10502 = n27462 ;
  assign y10503 = n27463 ;
  assign y10504 = ~n27465 ;
  assign y10505 = n27470 ;
  assign y10506 = ~n27473 ;
  assign y10507 = n27474 ;
  assign y10508 = n27477 ;
  assign y10509 = n27478 ;
  assign y10510 = n27481 ;
  assign y10511 = ~n27482 ;
  assign y10512 = n27485 ;
  assign y10513 = ~1'b0 ;
  assign y10514 = n27491 ;
  assign y10515 = n27494 ;
  assign y10516 = n27496 ;
  assign y10517 = ~n27502 ;
  assign y10518 = n27511 ;
  assign y10519 = ~n27515 ;
  assign y10520 = ~n27520 ;
  assign y10521 = n27525 ;
  assign y10522 = ~n27528 ;
  assign y10523 = ~1'b0 ;
  assign y10524 = ~n27529 ;
  assign y10525 = ~n27533 ;
  assign y10526 = ~n27535 ;
  assign y10527 = ~1'b0 ;
  assign y10528 = n27537 ;
  assign y10529 = n27540 ;
  assign y10530 = ~n27541 ;
  assign y10531 = ~n27544 ;
  assign y10532 = ~n27545 ;
  assign y10533 = ~n10026 ;
  assign y10534 = ~1'b0 ;
  assign y10535 = ~1'b0 ;
  assign y10536 = n27549 ;
  assign y10537 = ~1'b0 ;
  assign y10538 = ~1'b0 ;
  assign y10539 = ~n27552 ;
  assign y10540 = n27553 ;
  assign y10541 = n27554 ;
  assign y10542 = n27561 ;
  assign y10543 = ~n27564 ;
  assign y10544 = ~1'b0 ;
  assign y10545 = n27565 ;
  assign y10546 = n1212 ;
  assign y10547 = ~n27569 ;
  assign y10548 = ~1'b0 ;
  assign y10549 = ~n27570 ;
  assign y10550 = ~n27572 ;
  assign y10551 = n27573 ;
  assign y10552 = n27577 ;
  assign y10553 = ~n26786 ;
  assign y10554 = n27578 ;
  assign y10555 = n27580 ;
  assign y10556 = n27581 ;
  assign y10557 = n27583 ;
  assign y10558 = ~1'b0 ;
  assign y10559 = n27585 ;
  assign y10560 = ~n27587 ;
  assign y10561 = ~n27588 ;
  assign y10562 = ~n27590 ;
  assign y10563 = n27591 ;
  assign y10564 = ~n27593 ;
  assign y10565 = n14964 ;
  assign y10566 = ~n27597 ;
  assign y10567 = ~n27599 ;
  assign y10568 = n27601 ;
  assign y10569 = ~n27603 ;
  assign y10570 = ~n27604 ;
  assign y10571 = ~n27608 ;
  assign y10572 = ~n27609 ;
  assign y10573 = n27615 ;
  assign y10574 = ~n27617 ;
  assign y10575 = n27619 ;
  assign y10576 = ~1'b0 ;
  assign y10577 = n27622 ;
  assign y10578 = n27624 ;
  assign y10579 = ~n27629 ;
  assign y10580 = ~n27634 ;
  assign y10581 = n27635 ;
  assign y10582 = n27637 ;
  assign y10583 = n27638 ;
  assign y10584 = n165 ;
  assign y10585 = ~1'b0 ;
  assign y10586 = n27641 ;
  assign y10587 = ~1'b0 ;
  assign y10588 = ~n27643 ;
  assign y10589 = n27644 ;
  assign y10590 = ~n27645 ;
  assign y10591 = ~n27650 ;
  assign y10592 = n27651 ;
  assign y10593 = ~n27656 ;
  assign y10594 = ~1'b0 ;
  assign y10595 = n27657 ;
  assign y10596 = ~n27659 ;
  assign y10597 = ~n27662 ;
  assign y10598 = ~n27664 ;
  assign y10599 = n27665 ;
  assign y10600 = ~n27672 ;
  assign y10601 = n27673 ;
  assign y10602 = n27676 ;
  assign y10603 = ~n27677 ;
  assign y10604 = ~n27678 ;
  assign y10605 = ~1'b0 ;
  assign y10606 = n27681 ;
  assign y10607 = ~n27684 ;
  assign y10608 = n17677 ;
  assign y10609 = n27685 ;
  assign y10610 = ~n27686 ;
  assign y10611 = n27689 ;
  assign y10612 = ~n27691 ;
  assign y10613 = ~n27696 ;
  assign y10614 = ~n27700 ;
  assign y10615 = ~1'b0 ;
  assign y10616 = ~1'b0 ;
  assign y10617 = ~n27701 ;
  assign y10618 = n27704 ;
  assign y10619 = ~n27705 ;
  assign y10620 = ~n27707 ;
  assign y10621 = ~n27708 ;
  assign y10622 = n27712 ;
  assign y10623 = n27717 ;
  assign y10624 = n27720 ;
  assign y10625 = n27723 ;
  assign y10626 = n27728 ;
  assign y10627 = ~n27731 ;
  assign y10628 = ~n27732 ;
  assign y10629 = n27734 ;
  assign y10630 = ~n27736 ;
  assign y10631 = ~1'b0 ;
  assign y10632 = ~n27742 ;
  assign y10633 = n27743 ;
  assign y10634 = ~1'b0 ;
  assign y10635 = ~1'b0 ;
  assign y10636 = ~n27744 ;
  assign y10637 = ~n27745 ;
  assign y10638 = ~n27748 ;
  assign y10639 = n27749 ;
  assign y10640 = n27750 ;
  assign y10641 = ~1'b0 ;
  assign y10642 = ~1'b0 ;
  assign y10643 = ~n27753 ;
  assign y10644 = n27755 ;
  assign y10645 = ~n27758 ;
  assign y10646 = ~n27759 ;
  assign y10647 = ~n27763 ;
  assign y10648 = ~1'b0 ;
  assign y10649 = ~n27769 ;
  assign y10650 = ~1'b0 ;
  assign y10651 = ~1'b0 ;
  assign y10652 = ~n27771 ;
  assign y10653 = ~n27776 ;
  assign y10654 = ~1'b0 ;
  assign y10655 = n27777 ;
  assign y10656 = n27780 ;
  assign y10657 = n27781 ;
  assign y10658 = n27784 ;
  assign y10659 = ~n27785 ;
  assign y10660 = n27786 ;
  assign y10661 = ~n27788 ;
  assign y10662 = ~n27791 ;
  assign y10663 = ~1'b0 ;
  assign y10664 = ~1'b0 ;
  assign y10665 = ~1'b0 ;
  assign y10666 = ~1'b0 ;
  assign y10667 = ~n27797 ;
  assign y10668 = ~n27799 ;
  assign y10669 = n27800 ;
  assign y10670 = n27801 ;
  assign y10671 = ~n27802 ;
  assign y10672 = n27803 ;
  assign y10673 = n27804 ;
  assign y10674 = n27806 ;
  assign y10675 = ~1'b0 ;
  assign y10676 = n27809 ;
  assign y10677 = ~n27810 ;
  assign y10678 = n27811 ;
  assign y10679 = n27813 ;
  assign y10680 = n27815 ;
  assign y10681 = n27819 ;
  assign y10682 = n27821 ;
  assign y10683 = n27824 ;
  assign y10684 = ~1'b0 ;
  assign y10685 = n27827 ;
  assign y10686 = ~n27829 ;
  assign y10687 = n27831 ;
  assign y10688 = ~n27834 ;
  assign y10689 = ~n27835 ;
  assign y10690 = n27836 ;
  assign y10691 = ~n27837 ;
  assign y10692 = ~1'b0 ;
  assign y10693 = n27841 ;
  assign y10694 = ~n27844 ;
  assign y10695 = ~n27847 ;
  assign y10696 = ~1'b0 ;
  assign y10697 = ~n27850 ;
  assign y10698 = n27851 ;
  assign y10699 = n27854 ;
  assign y10700 = ~n27856 ;
  assign y10701 = ~n27859 ;
  assign y10702 = ~n27860 ;
  assign y10703 = ~n27862 ;
  assign y10704 = ~n27864 ;
  assign y10705 = n27867 ;
  assign y10706 = ~n27868 ;
  assign y10707 = n27873 ;
  assign y10708 = n27874 ;
  assign y10709 = ~n27876 ;
  assign y10710 = ~n27877 ;
  assign y10711 = ~n27879 ;
  assign y10712 = ~1'b0 ;
  assign y10713 = n27881 ;
  assign y10714 = ~1'b0 ;
  assign y10715 = n27882 ;
  assign y10716 = ~1'b0 ;
  assign y10717 = n27884 ;
  assign y10718 = ~n27886 ;
  assign y10719 = ~n27890 ;
  assign y10720 = n27891 ;
  assign y10721 = ~n27892 ;
  assign y10722 = n27896 ;
  assign y10723 = ~n27898 ;
  assign y10724 = n27902 ;
  assign y10725 = ~n27904 ;
  assign y10726 = ~1'b0 ;
  assign y10727 = n27906 ;
  assign y10728 = ~n27910 ;
  assign y10729 = ~n27913 ;
  assign y10730 = n27914 ;
  assign y10731 = ~1'b0 ;
  assign y10732 = n27917 ;
  assign y10733 = ~n27919 ;
  assign y10734 = ~n18644 ;
  assign y10735 = ~n27921 ;
  assign y10736 = ~1'b0 ;
  assign y10737 = n27930 ;
  assign y10738 = ~n27932 ;
  assign y10739 = ~n27935 ;
  assign y10740 = ~n27939 ;
  assign y10741 = ~n27941 ;
  assign y10742 = ~1'b0 ;
  assign y10743 = ~1'b0 ;
  assign y10744 = ~n27945 ;
  assign y10745 = 1'b0 ;
  assign y10746 = ~n27948 ;
  assign y10747 = ~1'b0 ;
  assign y10748 = ~n27950 ;
  assign y10749 = n27958 ;
  assign y10750 = ~n27963 ;
  assign y10751 = ~n27967 ;
  assign y10752 = ~1'b0 ;
  assign y10753 = n27972 ;
  assign y10754 = n27973 ;
  assign y10755 = ~1'b0 ;
  assign y10756 = n27977 ;
  assign y10757 = ~n27980 ;
  assign y10758 = n27982 ;
  assign y10759 = n27983 ;
  assign y10760 = n27989 ;
  assign y10761 = n27992 ;
  assign y10762 = ~n27993 ;
  assign y10763 = ~n27995 ;
  assign y10764 = ~n27998 ;
  assign y10765 = ~1'b0 ;
  assign y10766 = n27999 ;
  assign y10767 = n28000 ;
  assign y10768 = n28006 ;
  assign y10769 = n28007 ;
  assign y10770 = n28008 ;
  assign y10771 = n28010 ;
  assign y10772 = n28012 ;
  assign y10773 = n28013 ;
  assign y10774 = ~1'b0 ;
  assign y10775 = ~n28015 ;
  assign y10776 = n28016 ;
  assign y10777 = ~n28022 ;
  assign y10778 = ~n28024 ;
  assign y10779 = ~n1022 ;
  assign y10780 = n28025 ;
  assign y10781 = n28029 ;
  assign y10782 = ~n28030 ;
  assign y10783 = n28032 ;
  assign y10784 = n28034 ;
  assign y10785 = n28037 ;
  assign y10786 = n28042 ;
  assign y10787 = n28047 ;
  assign y10788 = n28050 ;
  assign y10789 = n22537 ;
  assign y10790 = ~n28051 ;
  assign y10791 = ~1'b0 ;
  assign y10792 = n28057 ;
  assign y10793 = ~n28062 ;
  assign y10794 = n28063 ;
  assign y10795 = ~n28067 ;
  assign y10796 = ~n28069 ;
  assign y10797 = n28070 ;
  assign y10798 = ~1'b0 ;
  assign y10799 = ~n28071 ;
  assign y10800 = ~1'b0 ;
  assign y10801 = ~n28077 ;
  assign y10802 = ~n28079 ;
  assign y10803 = ~n28083 ;
  assign y10804 = n28087 ;
  assign y10805 = ~n28088 ;
  assign y10806 = ~n28090 ;
  assign y10807 = n28093 ;
  assign y10808 = n28094 ;
  assign y10809 = n28095 ;
  assign y10810 = ~n26316 ;
  assign y10811 = n28096 ;
  assign y10812 = n28098 ;
  assign y10813 = n525 ;
  assign y10814 = n28100 ;
  assign y10815 = ~1'b0 ;
  assign y10816 = n28102 ;
  assign y10817 = ~n28104 ;
  assign y10818 = ~n28106 ;
  assign y10819 = ~n28109 ;
  assign y10820 = ~n28110 ;
  assign y10821 = n28113 ;
  assign y10822 = n28114 ;
  assign y10823 = ~n28119 ;
  assign y10824 = n28125 ;
  assign y10825 = n28127 ;
  assign y10826 = ~n28129 ;
  assign y10827 = ~1'b0 ;
  assign y10828 = ~n28131 ;
  assign y10829 = ~1'b0 ;
  assign y10830 = ~n28134 ;
  assign y10831 = ~n28138 ;
  assign y10832 = n28145 ;
  assign y10833 = ~n28147 ;
  assign y10834 = n28150 ;
  assign y10835 = n28154 ;
  assign y10836 = n28157 ;
  assign y10837 = n28162 ;
  assign y10838 = ~n28164 ;
  assign y10839 = ~n28168 ;
  assign y10840 = n28169 ;
  assign y10841 = n28170 ;
  assign y10842 = n28171 ;
  assign y10843 = n28172 ;
  assign y10844 = n28177 ;
  assign y10845 = n28178 ;
  assign y10846 = ~n28180 ;
  assign y10847 = ~n28181 ;
  assign y10848 = ~1'b0 ;
  assign y10849 = ~1'b0 ;
  assign y10850 = n28185 ;
  assign y10851 = n28188 ;
  assign y10852 = n28193 ;
  assign y10853 = ~n28194 ;
  assign y10854 = 1'b0 ;
  assign y10855 = n28195 ;
  assign y10856 = ~n28197 ;
  assign y10857 = ~n28201 ;
  assign y10858 = ~1'b0 ;
  assign y10859 = n28206 ;
  assign y10860 = ~n28208 ;
  assign y10861 = ~n28211 ;
  assign y10862 = ~n28218 ;
  assign y10863 = ~n28220 ;
  assign y10864 = n28221 ;
  assign y10865 = n28222 ;
  assign y10866 = ~1'b0 ;
  assign y10867 = n28225 ;
  assign y10868 = ~n28226 ;
  assign y10869 = ~n28238 ;
  assign y10870 = ~1'b0 ;
  assign y10871 = n28241 ;
  assign y10872 = n28244 ;
  assign y10873 = ~n28254 ;
  assign y10874 = n7157 ;
  assign y10875 = n28257 ;
  assign y10876 = n28259 ;
  assign y10877 = n28263 ;
  assign y10878 = ~n28267 ;
  assign y10879 = n28268 ;
  assign y10880 = n28270 ;
  assign y10881 = ~n28272 ;
  assign y10882 = ~n28273 ;
  assign y10883 = n28275 ;
  assign y10884 = n28279 ;
  assign y10885 = ~1'b0 ;
  assign y10886 = ~n28281 ;
  assign y10887 = ~n28285 ;
  assign y10888 = n28288 ;
  assign y10889 = ~n28291 ;
  assign y10890 = n28293 ;
  assign y10891 = ~1'b0 ;
  assign y10892 = ~n28299 ;
  assign y10893 = ~n28302 ;
  assign y10894 = ~n28303 ;
  assign y10895 = n28304 ;
  assign y10896 = ~n28305 ;
  assign y10897 = n28306 ;
  assign y10898 = n28308 ;
  assign y10899 = n28310 ;
  assign y10900 = ~1'b0 ;
  assign y10901 = ~1'b0 ;
  assign y10902 = n28311 ;
  assign y10903 = n28314 ;
  assign y10904 = ~n28317 ;
  assign y10905 = n28321 ;
  assign y10906 = ~n28323 ;
  assign y10907 = n28324 ;
  assign y10908 = ~n28327 ;
  assign y10909 = ~n28329 ;
  assign y10910 = ~n28330 ;
  assign y10911 = ~1'b0 ;
  assign y10912 = ~1'b0 ;
  assign y10913 = ~1'b0 ;
  assign y10914 = n28333 ;
  assign y10915 = n28334 ;
  assign y10916 = ~n28336 ;
  assign y10917 = n28342 ;
  assign y10918 = ~n28345 ;
  assign y10919 = ~1'b0 ;
  assign y10920 = ~n28349 ;
  assign y10921 = ~n28350 ;
  assign y10922 = ~n28352 ;
  assign y10923 = ~1'b0 ;
  assign y10924 = ~1'b0 ;
  assign y10925 = ~n28353 ;
  assign y10926 = n28359 ;
  assign y10927 = ~n28365 ;
  assign y10928 = n28367 ;
  assign y10929 = ~n28369 ;
  assign y10930 = n28371 ;
  assign y10931 = n28375 ;
  assign y10932 = ~1'b0 ;
  assign y10933 = ~1'b0 ;
  assign y10934 = ~n28376 ;
  assign y10935 = n28377 ;
  assign y10936 = ~n28389 ;
  assign y10937 = ~n28391 ;
  assign y10938 = n10853 ;
  assign y10939 = ~n28394 ;
  assign y10940 = ~n28395 ;
  assign y10941 = n28399 ;
  assign y10942 = n28401 ;
  assign y10943 = 1'b0 ;
  assign y10944 = n28407 ;
  assign y10945 = n28409 ;
  assign y10946 = ~n28410 ;
  assign y10947 = n28411 ;
  assign y10948 = ~n28414 ;
  assign y10949 = ~n28416 ;
  assign y10950 = n28417 ;
  assign y10951 = n28420 ;
  assign y10952 = ~1'b0 ;
  assign y10953 = ~1'b0 ;
  assign y10954 = ~n28429 ;
  assign y10955 = ~1'b0 ;
  assign y10956 = ~n28433 ;
  assign y10957 = n28434 ;
  assign y10958 = n28435 ;
  assign y10959 = n28437 ;
  assign y10960 = n28439 ;
  assign y10961 = ~n28445 ;
  assign y10962 = ~1'b0 ;
  assign y10963 = n28448 ;
  assign y10964 = n28450 ;
  assign y10965 = ~1'b0 ;
  assign y10966 = ~n28451 ;
  assign y10967 = ~n28453 ;
  assign y10968 = n28456 ;
  assign y10969 = ~n28460 ;
  assign y10970 = n28461 ;
  assign y10971 = ~n28462 ;
  assign y10972 = n28465 ;
  assign y10973 = ~1'b0 ;
  assign y10974 = ~n28466 ;
  assign y10975 = n28468 ;
  assign y10976 = ~n28470 ;
  assign y10977 = ~1'b0 ;
  assign y10978 = ~n28471 ;
  assign y10979 = ~n28476 ;
  assign y10980 = ~n28478 ;
  assign y10981 = ~n28483 ;
  assign y10982 = ~n28484 ;
  assign y10983 = n28488 ;
  assign y10984 = ~1'b0 ;
  assign y10985 = n28489 ;
  assign y10986 = n28491 ;
  assign y10987 = ~1'b0 ;
  assign y10988 = n28492 ;
  assign y10989 = n28493 ;
  assign y10990 = ~n28497 ;
  assign y10991 = ~n28498 ;
  assign y10992 = ~n28499 ;
  assign y10993 = n28500 ;
  assign y10994 = n28501 ;
  assign y10995 = n28504 ;
  assign y10996 = n28506 ;
  assign y10997 = ~1'b0 ;
  assign y10998 = n28509 ;
  assign y10999 = ~1'b0 ;
  assign y11000 = ~n28513 ;
  assign y11001 = ~n7421 ;
  assign y11002 = ~n28514 ;
  assign y11003 = n28516 ;
  assign y11004 = ~n28518 ;
  assign y11005 = ~n28519 ;
  assign y11006 = n28523 ;
  assign y11007 = ~n28525 ;
  assign y11008 = n28527 ;
  assign y11009 = ~n28530 ;
  assign y11010 = ~n28532 ;
  assign y11011 = n28538 ;
  assign y11012 = n28539 ;
  assign y11013 = n28542 ;
  assign y11014 = ~n28544 ;
  assign y11015 = n28546 ;
  assign y11016 = n28548 ;
  assign y11017 = ~n28552 ;
  assign y11018 = ~1'b0 ;
  assign y11019 = ~1'b0 ;
  assign y11020 = n28553 ;
  assign y11021 = n28555 ;
  assign y11022 = ~n28561 ;
  assign y11023 = ~n28563 ;
  assign y11024 = n28566 ;
  assign y11025 = ~n28567 ;
  assign y11026 = n28568 ;
  assign y11027 = n28569 ;
  assign y11028 = n9931 ;
  assign y11029 = ~n28571 ;
  assign y11030 = n28574 ;
  assign y11031 = ~n28577 ;
  assign y11032 = ~1'b0 ;
  assign y11033 = n28579 ;
  assign y11034 = n28586 ;
  assign y11035 = n28590 ;
  assign y11036 = ~n28591 ;
  assign y11037 = ~n28596 ;
  assign y11038 = ~n28602 ;
  assign y11039 = n28603 ;
  assign y11040 = ~n28606 ;
  assign y11041 = n28607 ;
  assign y11042 = ~n28608 ;
  assign y11043 = n28613 ;
  assign y11044 = n28615 ;
  assign y11045 = n28616 ;
  assign y11046 = ~n11687 ;
  assign y11047 = n28617 ;
  assign y11048 = n28618 ;
  assign y11049 = ~1'b0 ;
  assign y11050 = ~1'b0 ;
  assign y11051 = ~n28620 ;
  assign y11052 = n28624 ;
  assign y11053 = n28627 ;
  assign y11054 = n28629 ;
  assign y11055 = ~n28630 ;
  assign y11056 = ~n28631 ;
  assign y11057 = ~n28632 ;
  assign y11058 = n28634 ;
  assign y11059 = n28635 ;
  assign y11060 = n28636 ;
  assign y11061 = n28641 ;
  assign y11062 = ~n28643 ;
  assign y11063 = ~n28645 ;
  assign y11064 = n28650 ;
  assign y11065 = ~n28651 ;
  assign y11066 = ~n28653 ;
  assign y11067 = ~n28654 ;
  assign y11068 = n28657 ;
  assign y11069 = n28658 ;
  assign y11070 = ~n28665 ;
  assign y11071 = ~1'b0 ;
  assign y11072 = ~n28666 ;
  assign y11073 = ~n28667 ;
  assign y11074 = n28668 ;
  assign y11075 = ~n28673 ;
  assign y11076 = n28675 ;
  assign y11077 = n28676 ;
  assign y11078 = ~n28678 ;
  assign y11079 = ~1'b0 ;
  assign y11080 = n28679 ;
  assign y11081 = ~n28680 ;
  assign y11082 = ~n28683 ;
  assign y11083 = ~1'b0 ;
  assign y11084 = ~1'b0 ;
  assign y11085 = ~n28684 ;
  assign y11086 = ~n28686 ;
  assign y11087 = n4657 ;
  assign y11088 = ~n28687 ;
  assign y11089 = n28688 ;
  assign y11090 = ~n2761 ;
  assign y11091 = ~n28692 ;
  assign y11092 = ~n28694 ;
  assign y11093 = ~1'b0 ;
  assign y11094 = ~1'b0 ;
  assign y11095 = n28699 ;
  assign y11096 = ~n28700 ;
  assign y11097 = ~1'b0 ;
  assign y11098 = n28701 ;
  assign y11099 = n28707 ;
  assign y11100 = ~n28708 ;
  assign y11101 = n28709 ;
  assign y11102 = n28710 ;
  assign y11103 = n28713 ;
  assign y11104 = n17351 ;
  assign y11105 = ~1'b0 ;
  assign y11106 = n28715 ;
  assign y11107 = n28716 ;
  assign y11108 = n28719 ;
  assign y11109 = n28720 ;
  assign y11110 = n28721 ;
  assign y11111 = n28726 ;
  assign y11112 = n28729 ;
  assign y11113 = ~n28730 ;
  assign y11114 = n28734 ;
  assign y11115 = ~1'b0 ;
  assign y11116 = ~1'b0 ;
  assign y11117 = ~n28736 ;
  assign y11118 = n17475 ;
  assign y11119 = n28741 ;
  assign y11120 = ~n10817 ;
  assign y11121 = n7661 ;
  assign y11122 = n28743 ;
  assign y11123 = ~n28748 ;
  assign y11124 = ~n28753 ;
  assign y11125 = n28754 ;
  assign y11126 = n28756 ;
  assign y11127 = ~n28758 ;
  assign y11128 = ~n28761 ;
  assign y11129 = n28763 ;
  assign y11130 = ~n28764 ;
  assign y11131 = n28768 ;
  assign y11132 = n28769 ;
  assign y11133 = ~n28771 ;
  assign y11134 = n28775 ;
  assign y11135 = ~n28779 ;
  assign y11136 = n28780 ;
  assign y11137 = ~1'b0 ;
  assign y11138 = ~n28784 ;
  assign y11139 = ~n28785 ;
  assign y11140 = n28786 ;
  assign y11141 = n28787 ;
  assign y11142 = ~n28788 ;
  assign y11143 = ~n28789 ;
  assign y11144 = ~1'b0 ;
  assign y11145 = ~1'b0 ;
  assign y11146 = ~n28791 ;
  assign y11147 = ~1'b0 ;
  assign y11148 = ~n28794 ;
  assign y11149 = ~n28798 ;
  assign y11150 = n28800 ;
  assign y11151 = ~n28801 ;
  assign y11152 = ~n28803 ;
  assign y11153 = n28805 ;
  assign y11154 = n1511 ;
  assign y11155 = ~n28807 ;
  assign y11156 = ~1'b0 ;
  assign y11157 = n28808 ;
  assign y11158 = n28810 ;
  assign y11159 = n28811 ;
  assign y11160 = ~1'b0 ;
  assign y11161 = n28813 ;
  assign y11162 = ~n28815 ;
  assign y11163 = n28817 ;
  assign y11164 = ~n28821 ;
  assign y11165 = ~n12476 ;
  assign y11166 = ~n28825 ;
  assign y11167 = n28827 ;
  assign y11168 = ~1'b0 ;
  assign y11169 = ~n28830 ;
  assign y11170 = n28834 ;
  assign y11171 = n28835 ;
  assign y11172 = ~1'b0 ;
  assign y11173 = n28836 ;
  assign y11174 = n28840 ;
  assign y11175 = ~n28842 ;
  assign y11176 = ~1'b0 ;
  assign y11177 = n28844 ;
  assign y11178 = ~n28845 ;
  assign y11179 = ~1'b0 ;
  assign y11180 = n12203 ;
  assign y11181 = n28846 ;
  assign y11182 = n28849 ;
  assign y11183 = n28850 ;
  assign y11184 = 1'b0 ;
  assign y11185 = n28854 ;
  assign y11186 = ~1'b0 ;
  assign y11187 = 1'b0 ;
  assign y11188 = ~1'b0 ;
  assign y11189 = ~1'b0 ;
  assign y11190 = ~n28856 ;
  assign y11191 = n28857 ;
  assign y11192 = ~n28858 ;
  assign y11193 = ~n28862 ;
  assign y11194 = n28863 ;
  assign y11195 = ~n28864 ;
  assign y11196 = ~1'b0 ;
  assign y11197 = n28865 ;
  assign y11198 = ~n28870 ;
  assign y11199 = n28872 ;
  assign y11200 = ~1'b0 ;
  assign y11201 = ~1'b0 ;
  assign y11202 = n28873 ;
  assign y11203 = ~n28874 ;
  assign y11204 = ~n28875 ;
  assign y11205 = n28880 ;
  assign y11206 = ~1'b0 ;
  assign y11207 = ~n28882 ;
  assign y11208 = n28884 ;
  assign y11209 = ~1'b0 ;
  assign y11210 = ~1'b0 ;
  assign y11211 = n28892 ;
  assign y11212 = ~n28893 ;
  assign y11213 = ~n28894 ;
  assign y11214 = n15178 ;
  assign y11215 = ~n28897 ;
  assign y11216 = ~n28899 ;
  assign y11217 = ~1'b0 ;
  assign y11218 = ~n28901 ;
  assign y11219 = ~1'b0 ;
  assign y11220 = ~n28907 ;
  assign y11221 = n28908 ;
  assign y11222 = n28910 ;
  assign y11223 = n28911 ;
  assign y11224 = ~n28912 ;
  assign y11225 = ~n28913 ;
  assign y11226 = n28914 ;
  assign y11227 = n28915 ;
  assign y11228 = ~n28917 ;
  assign y11229 = n28921 ;
  assign y11230 = ~n28926 ;
  assign y11231 = n28928 ;
  assign y11232 = n28929 ;
  assign y11233 = ~n28930 ;
  assign y11234 = ~n28931 ;
  assign y11235 = ~n28934 ;
  assign y11236 = ~n28935 ;
  assign y11237 = ~n28936 ;
  assign y11238 = n28937 ;
  assign y11239 = n28943 ;
  assign y11240 = ~n28944 ;
  assign y11241 = n28945 ;
  assign y11242 = ~n28947 ;
  assign y11243 = n28951 ;
  assign y11244 = n28952 ;
  assign y11245 = ~n28953 ;
  assign y11246 = n28957 ;
  assign y11247 = ~n28966 ;
  assign y11248 = ~n28971 ;
  assign y11249 = ~n28973 ;
  assign y11250 = n28981 ;
  assign y11251 = n28982 ;
  assign y11252 = ~1'b0 ;
  assign y11253 = ~1'b0 ;
  assign y11254 = n28984 ;
  assign y11255 = ~n28988 ;
  assign y11256 = n28989 ;
  assign y11257 = ~n28991 ;
  assign y11258 = ~n28994 ;
  assign y11259 = ~n28997 ;
  assign y11260 = ~n29000 ;
  assign y11261 = n29003 ;
  assign y11262 = n29006 ;
  assign y11263 = ~n29011 ;
  assign y11264 = n24194 ;
  assign y11265 = n29013 ;
  assign y11266 = n29014 ;
  assign y11267 = ~n29015 ;
  assign y11268 = ~n29018 ;
  assign y11269 = n29021 ;
  assign y11270 = ~1'b0 ;
  assign y11271 = ~n29022 ;
  assign y11272 = n29024 ;
  assign y11273 = ~n29030 ;
  assign y11274 = ~n29031 ;
  assign y11275 = ~n29036 ;
  assign y11276 = ~n29038 ;
  assign y11277 = n29039 ;
  assign y11278 = ~n29041 ;
  assign y11279 = ~n29044 ;
  assign y11280 = n29046 ;
  assign y11281 = ~n29050 ;
  assign y11282 = ~n29051 ;
  assign y11283 = n29053 ;
  assign y11284 = n29056 ;
  assign y11285 = ~n29060 ;
  assign y11286 = ~1'b0 ;
  assign y11287 = ~n29073 ;
  assign y11288 = ~n29078 ;
  assign y11289 = ~n29080 ;
  assign y11290 = n29084 ;
  assign y11291 = ~n29087 ;
  assign y11292 = n29088 ;
  assign y11293 = n29090 ;
  assign y11294 = ~n29092 ;
  assign y11295 = ~n29095 ;
  assign y11296 = n5124 ;
  assign y11297 = n29100 ;
  assign y11298 = n29105 ;
  assign y11299 = ~n29106 ;
  assign y11300 = n29109 ;
  assign y11301 = ~n29111 ;
  assign y11302 = ~n29112 ;
  assign y11303 = n29113 ;
  assign y11304 = ~1'b0 ;
  assign y11305 = ~1'b0 ;
  assign y11306 = ~n29115 ;
  assign y11307 = n4802 ;
  assign y11308 = n29116 ;
  assign y11309 = n29117 ;
  assign y11310 = ~n29120 ;
  assign y11311 = ~n29121 ;
  assign y11312 = ~1'b0 ;
  assign y11313 = n29122 ;
  assign y11314 = ~1'b0 ;
  assign y11315 = ~n29127 ;
  assign y11316 = ~n29130 ;
  assign y11317 = ~1'b0 ;
  assign y11318 = ~n29132 ;
  assign y11319 = n29134 ;
  assign y11320 = ~n29137 ;
  assign y11321 = ~n29140 ;
  assign y11322 = n29141 ;
  assign y11323 = ~n29142 ;
  assign y11324 = ~n29146 ;
  assign y11325 = ~1'b0 ;
  assign y11326 = ~n29148 ;
  assign y11327 = ~1'b0 ;
  assign y11328 = ~n29150 ;
  assign y11329 = n29155 ;
  assign y11330 = n29156 ;
  assign y11331 = n29158 ;
  assign y11332 = ~n29160 ;
  assign y11333 = ~n29161 ;
  assign y11334 = ~1'b0 ;
  assign y11335 = ~n29163 ;
  assign y11336 = ~1'b0 ;
  assign y11337 = ~1'b0 ;
  assign y11338 = ~n29169 ;
  assign y11339 = ~n29171 ;
  assign y11340 = ~n29174 ;
  assign y11341 = n29175 ;
  assign y11342 = ~n29176 ;
  assign y11343 = ~n29184 ;
  assign y11344 = ~n29185 ;
  assign y11345 = ~1'b0 ;
  assign y11346 = ~1'b0 ;
  assign y11347 = ~n29187 ;
  assign y11348 = n29192 ;
  assign y11349 = ~1'b0 ;
  assign y11350 = ~1'b0 ;
  assign y11351 = n29193 ;
  assign y11352 = ~n24376 ;
  assign y11353 = ~n29194 ;
  assign y11354 = n29195 ;
  assign y11355 = ~n29197 ;
  assign y11356 = ~n29202 ;
  assign y11357 = n29204 ;
  assign y11358 = ~n29208 ;
  assign y11359 = n29210 ;
  assign y11360 = ~n29212 ;
  assign y11361 = n29214 ;
  assign y11362 = ~n29215 ;
  assign y11363 = n29219 ;
  assign y11364 = n4429 ;
  assign y11365 = ~n29220 ;
  assign y11366 = ~n29222 ;
  assign y11367 = ~1'b0 ;
  assign y11368 = n29224 ;
  assign y11369 = ~n29226 ;
  assign y11370 = ~1'b0 ;
  assign y11371 = ~1'b0 ;
  assign y11372 = ~n29229 ;
  assign y11373 = ~n29230 ;
  assign y11374 = n29234 ;
  assign y11375 = ~n29238 ;
  assign y11376 = n29244 ;
  assign y11377 = ~n29246 ;
  assign y11378 = ~1'b0 ;
  assign y11379 = ~n29253 ;
  assign y11380 = ~n29256 ;
  assign y11381 = n29257 ;
  assign y11382 = n29259 ;
  assign y11383 = n18779 ;
  assign y11384 = n29262 ;
  assign y11385 = n29267 ;
  assign y11386 = ~n29270 ;
  assign y11387 = ~n29271 ;
  assign y11388 = ~n29272 ;
  assign y11389 = ~n29274 ;
  assign y11390 = ~n29276 ;
  assign y11391 = ~1'b0 ;
  assign y11392 = ~1'b0 ;
  assign y11393 = n29277 ;
  assign y11394 = ~1'b0 ;
  assign y11395 = n29279 ;
  assign y11396 = n29281 ;
  assign y11397 = n29286 ;
  assign y11398 = ~n29288 ;
  assign y11399 = ~1'b0 ;
  assign y11400 = n29290 ;
  assign y11401 = ~n29291 ;
  assign y11402 = ~n29298 ;
  assign y11403 = n29301 ;
  assign y11404 = ~1'b0 ;
  assign y11405 = n29302 ;
  assign y11406 = ~n29303 ;
  assign y11407 = ~n29307 ;
  assign y11408 = n29308 ;
  assign y11409 = ~n29314 ;
  assign y11410 = ~n29315 ;
  assign y11411 = ~n29320 ;
  assign y11412 = ~n29321 ;
  assign y11413 = n29324 ;
  assign y11414 = ~n29326 ;
  assign y11415 = ~n29329 ;
  assign y11416 = ~n29331 ;
  assign y11417 = n29333 ;
  assign y11418 = ~n29334 ;
  assign y11419 = ~n29335 ;
  assign y11420 = ~n29337 ;
  assign y11421 = ~n29338 ;
  assign y11422 = ~n29340 ;
  assign y11423 = n29341 ;
  assign y11424 = ~n29343 ;
  assign y11425 = ~n29346 ;
  assign y11426 = n29347 ;
  assign y11427 = ~n29351 ;
  assign y11428 = ~n29357 ;
  assign y11429 = n29359 ;
  assign y11430 = ~1'b0 ;
  assign y11431 = n29364 ;
  assign y11432 = ~n29365 ;
  assign y11433 = ~1'b0 ;
  assign y11434 = ~1'b0 ;
  assign y11435 = ~n29370 ;
  assign y11436 = n29372 ;
  assign y11437 = n29373 ;
  assign y11438 = ~1'b0 ;
  assign y11439 = ~n29376 ;
  assign y11440 = n29378 ;
  assign y11441 = n29380 ;
  assign y11442 = n19751 ;
  assign y11443 = ~n29381 ;
  assign y11444 = ~1'b0 ;
  assign y11445 = n29382 ;
  assign y11446 = n29384 ;
  assign y11447 = ~1'b0 ;
  assign y11448 = ~n29390 ;
  assign y11449 = n29392 ;
  assign y11450 = ~n29394 ;
  assign y11451 = n29395 ;
  assign y11452 = ~n29396 ;
  assign y11453 = ~1'b0 ;
  assign y11454 = n29398 ;
  assign y11455 = ~1'b0 ;
  assign y11456 = ~n29402 ;
  assign y11457 = ~n29403 ;
  assign y11458 = n29405 ;
  assign y11459 = ~n29407 ;
  assign y11460 = n29408 ;
  assign y11461 = n29409 ;
  assign y11462 = n29410 ;
  assign y11463 = ~n29411 ;
  assign y11464 = n29413 ;
  assign y11465 = ~n29415 ;
  assign y11466 = n29416 ;
  assign y11467 = ~1'b0 ;
  assign y11468 = ~n29418 ;
  assign y11469 = ~1'b0 ;
  assign y11470 = ~n29419 ;
  assign y11471 = n29427 ;
  assign y11472 = ~n29428 ;
  assign y11473 = n29429 ;
  assign y11474 = n29431 ;
  assign y11475 = ~1'b0 ;
  assign y11476 = ~n4629 ;
  assign y11477 = ~n29433 ;
  assign y11478 = ~n29436 ;
  assign y11479 = n17000 ;
  assign y11480 = ~1'b0 ;
  assign y11481 = n29442 ;
  assign y11482 = n29446 ;
  assign y11483 = n29447 ;
  assign y11484 = ~n29448 ;
  assign y11485 = ~n29451 ;
  assign y11486 = ~1'b0 ;
  assign y11487 = n29452 ;
  assign y11488 = n29453 ;
  assign y11489 = n29456 ;
  assign y11490 = ~n29458 ;
  assign y11491 = ~n29463 ;
  assign y11492 = ~n29464 ;
  assign y11493 = ~n29465 ;
  assign y11494 = n6847 ;
  assign y11495 = n29466 ;
  assign y11496 = ~n29467 ;
  assign y11497 = ~n29469 ;
  assign y11498 = ~1'b0 ;
  assign y11499 = ~1'b0 ;
  assign y11500 = ~n29472 ;
  assign y11501 = ~1'b0 ;
  assign y11502 = n29474 ;
  assign y11503 = ~n29475 ;
  assign y11504 = ~n29477 ;
  assign y11505 = ~n29480 ;
  assign y11506 = n29488 ;
  assign y11507 = n29489 ;
  assign y11508 = ~1'b0 ;
  assign y11509 = ~n29494 ;
  assign y11510 = n29498 ;
  assign y11511 = ~1'b0 ;
  assign y11512 = n29503 ;
  assign y11513 = ~n29508 ;
  assign y11514 = ~n29510 ;
  assign y11515 = ~n29515 ;
  assign y11516 = ~n29517 ;
  assign y11517 = ~n29520 ;
  assign y11518 = ~n29524 ;
  assign y11519 = n29526 ;
  assign y11520 = n29528 ;
  assign y11521 = ~1'b0 ;
  assign y11522 = n29529 ;
  assign y11523 = ~n29531 ;
  assign y11524 = ~1'b0 ;
  assign y11525 = ~n29535 ;
  assign y11526 = n29537 ;
  assign y11527 = ~n11622 ;
  assign y11528 = n29540 ;
  assign y11529 = n29541 ;
  assign y11530 = ~1'b0 ;
  assign y11531 = n29543 ;
  assign y11532 = 1'b0 ;
  assign y11533 = ~n29545 ;
  assign y11534 = ~1'b0 ;
  assign y11535 = ~n29547 ;
  assign y11536 = n29550 ;
  assign y11537 = n29552 ;
  assign y11538 = ~n29555 ;
  assign y11539 = ~n29560 ;
  assign y11540 = ~n29561 ;
  assign y11541 = ~1'b0 ;
  assign y11542 = ~1'b0 ;
  assign y11543 = n29566 ;
  assign y11544 = n29567 ;
  assign y11545 = n27084 ;
  assign y11546 = n29569 ;
  assign y11547 = ~n29570 ;
  assign y11548 = ~n29573 ;
  assign y11549 = n29576 ;
  assign y11550 = n29578 ;
  assign y11551 = n29579 ;
  assign y11552 = n29580 ;
  assign y11553 = ~1'b0 ;
  assign y11554 = ~n29582 ;
  assign y11555 = ~n29584 ;
  assign y11556 = ~1'b0 ;
  assign y11557 = ~1'b0 ;
  assign y11558 = ~n29586 ;
  assign y11559 = n29588 ;
  assign y11560 = ~n29589 ;
  assign y11561 = ~n29590 ;
  assign y11562 = ~1'b0 ;
  assign y11563 = ~n29594 ;
  assign y11564 = 1'b0 ;
  assign y11565 = n19747 ;
  assign y11566 = ~n29598 ;
  assign y11567 = ~n29601 ;
  assign y11568 = n29602 ;
  assign y11569 = n29603 ;
  assign y11570 = ~n29604 ;
  assign y11571 = n29605 ;
  assign y11572 = n29607 ;
  assign y11573 = ~n29610 ;
  assign y11574 = ~1'b0 ;
  assign y11575 = ~n29614 ;
  assign y11576 = n29617 ;
  assign y11577 = ~1'b0 ;
  assign y11578 = ~1'b0 ;
  assign y11579 = ~1'b0 ;
  assign y11580 = ~n29618 ;
  assign y11581 = ~n29622 ;
  assign y11582 = n29626 ;
  assign y11583 = n29628 ;
  assign y11584 = ~n29630 ;
  assign y11585 = ~n29633 ;
  assign y11586 = ~n29636 ;
  assign y11587 = ~n29638 ;
  assign y11588 = n29642 ;
  assign y11589 = ~n29643 ;
  assign y11590 = n29644 ;
  assign y11591 = ~n29646 ;
  assign y11592 = ~n29649 ;
  assign y11593 = ~1'b0 ;
  assign y11594 = ~n29653 ;
  assign y11595 = ~1'b0 ;
  assign y11596 = n29655 ;
  assign y11597 = n29658 ;
  assign y11598 = n29660 ;
  assign y11599 = ~1'b0 ;
  assign y11600 = n29661 ;
  assign y11601 = ~n29665 ;
  assign y11602 = n29669 ;
  assign y11603 = ~1'b0 ;
  assign y11604 = n29671 ;
  assign y11605 = ~n29673 ;
  assign y11606 = ~1'b0 ;
  assign y11607 = ~n29678 ;
  assign y11608 = n1882 ;
  assign y11609 = n29679 ;
  assign y11610 = ~n29682 ;
  assign y11611 = ~n29683 ;
  assign y11612 = ~n29684 ;
  assign y11613 = n29687 ;
  assign y11614 = ~n29691 ;
  assign y11615 = n29692 ;
  assign y11616 = ~n29696 ;
  assign y11617 = n29700 ;
  assign y11618 = ~n29701 ;
  assign y11619 = ~1'b0 ;
  assign y11620 = ~1'b0 ;
  assign y11621 = n29702 ;
  assign y11622 = ~n29703 ;
  assign y11623 = ~n29705 ;
  assign y11624 = n29708 ;
  assign y11625 = n29709 ;
  assign y11626 = n29710 ;
  assign y11627 = n29711 ;
  assign y11628 = ~1'b0 ;
  assign y11629 = ~1'b0 ;
  assign y11630 = ~1'b0 ;
  assign y11631 = ~1'b0 ;
  assign y11632 = ~n29712 ;
  assign y11633 = 1'b0 ;
  assign y11634 = ~n29714 ;
  assign y11635 = ~n29715 ;
  assign y11636 = ~n29716 ;
  assign y11637 = ~n29722 ;
  assign y11638 = ~n29727 ;
  assign y11639 = ~1'b0 ;
  assign y11640 = ~n6659 ;
  assign y11641 = ~n29729 ;
  assign y11642 = n29730 ;
  assign y11643 = n29734 ;
  assign y11644 = n2896 ;
  assign y11645 = n29738 ;
  assign y11646 = n29739 ;
  assign y11647 = ~n29742 ;
  assign y11648 = ~1'b0 ;
  assign y11649 = ~n29743 ;
  assign y11650 = n29745 ;
  assign y11651 = ~n29749 ;
  assign y11652 = n29750 ;
  assign y11653 = ~n29752 ;
  assign y11654 = ~n29753 ;
  assign y11655 = ~n29756 ;
  assign y11656 = ~n29757 ;
  assign y11657 = n29760 ;
  assign y11658 = n29766 ;
  assign y11659 = ~1'b0 ;
  assign y11660 = n29770 ;
  assign y11661 = ~n29774 ;
  assign y11662 = ~n29779 ;
  assign y11663 = ~n29781 ;
  assign y11664 = ~1'b0 ;
endmodule
