module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 , y20242 , y20243 , y20244 , y20245 , y20246 , y20247 , y20248 , y20249 , y20250 , y20251 , y20252 , y20253 , y20254 , y20255 , y20256 , y20257 , y20258 , y20259 , y20260 , y20261 , y20262 , y20263 , y20264 , y20265 , y20266 , y20267 , y20268 , y20269 , y20270 , y20271 , y20272 , y20273 , y20274 , y20275 , y20276 , y20277 , y20278 , y20279 , y20280 , y20281 , y20282 , y20283 , y20284 , y20285 , y20286 , y20287 , y20288 , y20289 , y20290 , y20291 , y20292 , y20293 , y20294 , y20295 , y20296 , y20297 , y20298 , y20299 , y20300 , y20301 , y20302 , y20303 , y20304 , y20305 , y20306 , y20307 , y20308 , y20309 , y20310 , y20311 , y20312 , y20313 , y20314 , y20315 , y20316 , y20317 , y20318 , y20319 , y20320 , y20321 , y20322 , y20323 , y20324 , y20325 , y20326 , y20327 , y20328 , y20329 , y20330 , y20331 , y20332 , y20333 , y20334 , y20335 , y20336 , y20337 , y20338 , y20339 , y20340 , y20341 , y20342 , y20343 , y20344 , y20345 , y20346 , y20347 , y20348 , y20349 , y20350 , y20351 , y20352 , y20353 , y20354 , y20355 , y20356 , y20357 , y20358 , y20359 , y20360 , y20361 , y20362 , y20363 , y20364 , y20365 , y20366 , y20367 , y20368 , y20369 , y20370 , y20371 , y20372 , y20373 , y20374 , y20375 , y20376 , y20377 , y20378 , y20379 , y20380 , y20381 , y20382 , y20383 , y20384 , y20385 , y20386 , y20387 , y20388 , y20389 , y20390 , y20391 , y20392 , y20393 , y20394 , y20395 , y20396 , y20397 , y20398 , y20399 , y20400 , y20401 , y20402 , y20403 , y20404 , y20405 , y20406 , y20407 , y20408 , y20409 , y20410 , y20411 , y20412 , y20413 , y20414 , y20415 , y20416 , y20417 , y20418 , y20419 , y20420 , y20421 , y20422 , y20423 , y20424 , y20425 , y20426 , y20427 , y20428 , y20429 , y20430 , y20431 , y20432 , y20433 , y20434 , y20435 , y20436 , y20437 , y20438 , y20439 , y20440 , y20441 , y20442 , y20443 , y20444 , y20445 , y20446 , y20447 , y20448 , y20449 , y20450 , y20451 , y20452 , y20453 , y20454 , y20455 , y20456 , y20457 , y20458 , y20459 , y20460 , y20461 , y20462 , y20463 , y20464 , y20465 , y20466 , y20467 , y20468 , y20469 , y20470 , y20471 , y20472 , y20473 , y20474 , y20475 , y20476 , y20477 , y20478 , y20479 , y20480 , y20481 , y20482 , y20483 , y20484 , y20485 , y20486 , y20487 , y20488 , y20489 , y20490 , y20491 , y20492 , y20493 , y20494 , y20495 , y20496 , y20497 , y20498 , y20499 , y20500 , y20501 , y20502 , y20503 , y20504 , y20505 , y20506 , y20507 , y20508 , y20509 , y20510 , y20511 , y20512 , y20513 , y20514 , y20515 , y20516 , y20517 , y20518 , y20519 , y20520 , y20521 , y20522 , y20523 , y20524 , y20525 , y20526 , y20527 , y20528 , y20529 , y20530 , y20531 , y20532 , y20533 , y20534 , y20535 , y20536 , y20537 , y20538 , y20539 , y20540 , y20541 , y20542 , y20543 , y20544 , y20545 , y20546 , y20547 , y20548 , y20549 , y20550 , y20551 , y20552 , y20553 , y20554 , y20555 , y20556 , y20557 , y20558 , y20559 , y20560 , y20561 , y20562 , y20563 , y20564 , y20565 , y20566 , y20567 , y20568 , y20569 , y20570 , y20571 , y20572 , y20573 , y20574 , y20575 , y20576 , y20577 , y20578 , y20579 , y20580 , y20581 , y20582 , y20583 , y20584 , y20585 , y20586 , y20587 , y20588 , y20589 , y20590 , y20591 , y20592 , y20593 , y20594 , y20595 , y20596 , y20597 , y20598 , y20599 , y20600 , y20601 , y20602 , y20603 , y20604 , y20605 , y20606 , y20607 , y20608 , y20609 , y20610 , y20611 , y20612 , y20613 , y20614 , y20615 , y20616 , y20617 , y20618 , y20619 , y20620 , y20621 , y20622 , y20623 , y20624 , y20625 , y20626 , y20627 , y20628 , y20629 , y20630 , y20631 , y20632 , y20633 , y20634 , y20635 , y20636 , y20637 , y20638 , y20639 , y20640 , y20641 , y20642 , y20643 , y20644 , y20645 , y20646 , y20647 , y20648 , y20649 , y20650 , y20651 , y20652 , y20653 , y20654 , y20655 , y20656 , y20657 , y20658 , y20659 , y20660 , y20661 , y20662 , y20663 , y20664 , y20665 , y20666 , y20667 , y20668 , y20669 , y20670 , y20671 , y20672 , y20673 , y20674 , y20675 , y20676 , y20677 , y20678 , y20679 , y20680 , y20681 , y20682 , y20683 , y20684 , y20685 , y20686 , y20687 , y20688 , y20689 , y20690 , y20691 , y20692 , y20693 , y20694 , y20695 , y20696 , y20697 , y20698 , y20699 , y20700 , y20701 , y20702 , y20703 , y20704 , y20705 , y20706 , y20707 , y20708 , y20709 , y20710 , y20711 , y20712 , y20713 , y20714 , y20715 , y20716 , y20717 , y20718 , y20719 , y20720 , y20721 , y20722 , y20723 , y20724 , y20725 , y20726 , y20727 , y20728 , y20729 , y20730 , y20731 , y20732 , y20733 , y20734 , y20735 , y20736 , y20737 , y20738 , y20739 , y20740 , y20741 , y20742 , y20743 , y20744 , y20745 , y20746 , y20747 , y20748 , y20749 , y20750 , y20751 , y20752 , y20753 , y20754 , y20755 , y20756 , y20757 , y20758 , y20759 , y20760 , y20761 , y20762 , y20763 , y20764 , y20765 , y20766 , y20767 , y20768 , y20769 , y20770 , y20771 , y20772 , y20773 , y20774 , y20775 , y20776 , y20777 , y20778 , y20779 , y20780 , y20781 , y20782 , y20783 , y20784 , y20785 , y20786 , y20787 , y20788 , y20789 , y20790 , y20791 , y20792 , y20793 , y20794 , y20795 , y20796 , y20797 , y20798 , y20799 , y20800 , y20801 , y20802 , y20803 , y20804 , y20805 , y20806 , y20807 , y20808 , y20809 , y20810 , y20811 , y20812 , y20813 , y20814 , y20815 , y20816 , y20817 , y20818 , y20819 , y20820 , y20821 , y20822 , y20823 , y20824 , y20825 , y20826 , y20827 , y20828 , y20829 , y20830 , y20831 , y20832 , y20833 , y20834 , y20835 , y20836 , y20837 , y20838 , y20839 , y20840 , y20841 , y20842 , y20843 , y20844 , y20845 , y20846 , y20847 , y20848 , y20849 , y20850 , y20851 , y20852 , y20853 , y20854 , y20855 , y20856 , y20857 , y20858 , y20859 , y20860 , y20861 , y20862 , y20863 , y20864 , y20865 , y20866 , y20867 , y20868 , y20869 , y20870 , y20871 , y20872 , y20873 , y20874 , y20875 , y20876 , y20877 , y20878 , y20879 , y20880 , y20881 , y20882 , y20883 , y20884 , y20885 , y20886 , y20887 , y20888 , y20889 , y20890 , y20891 , y20892 , y20893 , y20894 , y20895 , y20896 , y20897 , y20898 , y20899 , y20900 , y20901 , y20902 , y20903 , y20904 , y20905 , y20906 , y20907 , y20908 , y20909 , y20910 , y20911 , y20912 , y20913 , y20914 , y20915 , y20916 , y20917 , y20918 , y20919 , y20920 , y20921 , y20922 , y20923 , y20924 , y20925 , y20926 , y20927 , y20928 , y20929 , y20930 , y20931 , y20932 , y20933 , y20934 , y20935 , y20936 , y20937 , y20938 , y20939 , y20940 , y20941 , y20942 , y20943 , y20944 , y20945 , y20946 , y20947 , y20948 , y20949 , y20950 , y20951 , y20952 , y20953 , y20954 , y20955 , y20956 , y20957 , y20958 , y20959 , y20960 , y20961 , y20962 , y20963 , y20964 , y20965 , y20966 , y20967 , y20968 , y20969 , y20970 , y20971 , y20972 , y20973 , y20974 , y20975 , y20976 , y20977 , y20978 , y20979 , y20980 , y20981 , y20982 , y20983 , y20984 , y20985 , y20986 , y20987 , y20988 , y20989 , y20990 , y20991 , y20992 , y20993 , y20994 , y20995 , y20996 , y20997 , y20998 , y20999 , y21000 , y21001 , y21002 , y21003 , y21004 , y21005 , y21006 , y21007 , y21008 , y21009 , y21010 , y21011 , y21012 , y21013 , y21014 , y21015 , y21016 , y21017 , y21018 , y21019 , y21020 , y21021 , y21022 , y21023 , y21024 , y21025 , y21026 , y21027 , y21028 , y21029 , y21030 , y21031 , y21032 , y21033 , y21034 , y21035 , y21036 , y21037 , y21038 , y21039 , y21040 , y21041 , y21042 , y21043 , y21044 , y21045 , y21046 , y21047 , y21048 , y21049 , y21050 , y21051 , y21052 , y21053 , y21054 , y21055 , y21056 , y21057 , y21058 , y21059 , y21060 , y21061 , y21062 , y21063 , y21064 , y21065 , y21066 , y21067 , y21068 , y21069 , y21070 , y21071 , y21072 , y21073 , y21074 , y21075 , y21076 , y21077 , y21078 , y21079 , y21080 , y21081 , y21082 , y21083 , y21084 , y21085 , y21086 , y21087 , y21088 , y21089 , y21090 , y21091 , y21092 , y21093 , y21094 , y21095 , y21096 , y21097 , y21098 , y21099 , y21100 , y21101 , y21102 , y21103 , y21104 , y21105 , y21106 , y21107 , y21108 , y21109 , y21110 , y21111 , y21112 , y21113 , y21114 , y21115 , y21116 , y21117 , y21118 , y21119 , y21120 , y21121 , y21122 , y21123 , y21124 , y21125 , y21126 , y21127 , y21128 , y21129 , y21130 , y21131 , y21132 , y21133 , y21134 , y21135 , y21136 , y21137 , y21138 , y21139 , y21140 , y21141 , y21142 , y21143 , y21144 , y21145 , y21146 , y21147 , y21148 , y21149 , y21150 , y21151 , y21152 , y21153 , y21154 , y21155 , y21156 , y21157 , y21158 , y21159 , y21160 , y21161 , y21162 , y21163 , y21164 , y21165 , y21166 , y21167 , y21168 , y21169 , y21170 , y21171 , y21172 , y21173 , y21174 , y21175 , y21176 , y21177 , y21178 , y21179 , y21180 , y21181 , y21182 , y21183 , y21184 , y21185 , y21186 , y21187 , y21188 , y21189 , y21190 , y21191 , y21192 , y21193 , y21194 , y21195 , y21196 , y21197 , y21198 , y21199 , y21200 , y21201 , y21202 , y21203 , y21204 , y21205 , y21206 , y21207 , y21208 , y21209 , y21210 , y21211 , y21212 , y21213 , y21214 , y21215 , y21216 , y21217 , y21218 , y21219 , y21220 , y21221 , y21222 , y21223 , y21224 , y21225 , y21226 , y21227 , y21228 , y21229 , y21230 , y21231 , y21232 , y21233 , y21234 , y21235 , y21236 , y21237 , y21238 , y21239 , y21240 , y21241 , y21242 , y21243 , y21244 , y21245 , y21246 , y21247 , y21248 , y21249 , y21250 , y21251 , y21252 , y21253 , y21254 , y21255 , y21256 , y21257 , y21258 , y21259 , y21260 , y21261 , y21262 , y21263 , y21264 , y21265 , y21266 , y21267 , y21268 , y21269 , y21270 , y21271 , y21272 , y21273 , y21274 , y21275 , y21276 , y21277 , y21278 , y21279 , y21280 , y21281 , y21282 , y21283 , y21284 , y21285 , y21286 , y21287 , y21288 , y21289 , y21290 , y21291 , y21292 , y21293 , y21294 , y21295 , y21296 , y21297 , y21298 , y21299 , y21300 , y21301 , y21302 , y21303 , y21304 , y21305 , y21306 , y21307 , y21308 , y21309 , y21310 , y21311 , y21312 , y21313 , y21314 , y21315 , y21316 , y21317 , y21318 , y21319 , y21320 , y21321 , y21322 , y21323 , y21324 , y21325 , y21326 , y21327 , y21328 , y21329 , y21330 , y21331 , y21332 , y21333 , y21334 , y21335 , y21336 , y21337 , y21338 , y21339 , y21340 , y21341 , y21342 , y21343 , y21344 , y21345 , y21346 , y21347 , y21348 , y21349 , y21350 , y21351 , y21352 , y21353 , y21354 , y21355 , y21356 , y21357 , y21358 , y21359 , y21360 , y21361 , y21362 , y21363 , y21364 , y21365 , y21366 , y21367 , y21368 , y21369 , y21370 , y21371 , y21372 , y21373 , y21374 , y21375 , y21376 , y21377 , y21378 , y21379 , y21380 , y21381 , y21382 , y21383 , y21384 , y21385 , y21386 , y21387 , y21388 , y21389 , y21390 , y21391 , y21392 , y21393 , y21394 , y21395 , y21396 , y21397 , y21398 , y21399 , y21400 , y21401 , y21402 , y21403 , y21404 , y21405 , y21406 , y21407 , y21408 , y21409 , y21410 , y21411 , y21412 , y21413 , y21414 , y21415 , y21416 , y21417 , y21418 , y21419 , y21420 , y21421 , y21422 , y21423 , y21424 , y21425 , y21426 , y21427 , y21428 , y21429 , y21430 , y21431 , y21432 , y21433 , y21434 , y21435 , y21436 , y21437 , y21438 , y21439 , y21440 , y21441 , y21442 , y21443 , y21444 , y21445 , y21446 , y21447 , y21448 , y21449 , y21450 , y21451 , y21452 , y21453 , y21454 , y21455 , y21456 , y21457 , y21458 , y21459 , y21460 , y21461 , y21462 , y21463 , y21464 , y21465 , y21466 , y21467 , y21468 , y21469 , y21470 , y21471 , y21472 , y21473 , y21474 , y21475 , y21476 , y21477 , y21478 , y21479 , y21480 , y21481 , y21482 , y21483 , y21484 , y21485 , y21486 , y21487 , y21488 , y21489 , y21490 , y21491 , y21492 , y21493 , y21494 , y21495 , y21496 , y21497 , y21498 , y21499 , y21500 , y21501 , y21502 , y21503 , y21504 , y21505 , y21506 , y21507 , y21508 , y21509 , y21510 , y21511 , y21512 , y21513 , y21514 , y21515 , y21516 , y21517 , y21518 , y21519 , y21520 , y21521 , y21522 , y21523 , y21524 , y21525 , y21526 , y21527 , y21528 , y21529 , y21530 , y21531 , y21532 , y21533 , y21534 , y21535 , y21536 , y21537 , y21538 , y21539 , y21540 , y21541 , y21542 , y21543 , y21544 , y21545 , y21546 , y21547 , y21548 , y21549 , y21550 , y21551 , y21552 , y21553 , y21554 , y21555 , y21556 , y21557 , y21558 , y21559 , y21560 , y21561 , y21562 , y21563 , y21564 , y21565 , y21566 , y21567 , y21568 , y21569 , y21570 , y21571 , y21572 , y21573 , y21574 , y21575 , y21576 , y21577 , y21578 , y21579 , y21580 , y21581 , y21582 , y21583 , y21584 , y21585 , y21586 , y21587 , y21588 , y21589 , y21590 , y21591 , y21592 , y21593 , y21594 , y21595 , y21596 , y21597 , y21598 , y21599 , y21600 , y21601 , y21602 , y21603 , y21604 , y21605 , y21606 , y21607 , y21608 , y21609 , y21610 , y21611 , y21612 , y21613 , y21614 , y21615 , y21616 , y21617 , y21618 , y21619 , y21620 , y21621 , y21622 , y21623 , y21624 , y21625 , y21626 , y21627 , y21628 , y21629 , y21630 , y21631 , y21632 , y21633 , y21634 , y21635 , y21636 , y21637 , y21638 , y21639 , y21640 , y21641 , y21642 , y21643 , y21644 , y21645 , y21646 , y21647 , y21648 , y21649 , y21650 , y21651 , y21652 , y21653 , y21654 , y21655 , y21656 , y21657 , y21658 , y21659 , y21660 , y21661 , y21662 , y21663 , y21664 , y21665 , y21666 , y21667 , y21668 , y21669 , y21670 , y21671 , y21672 , y21673 , y21674 , y21675 , y21676 , y21677 , y21678 , y21679 , y21680 , y21681 , y21682 , y21683 , y21684 , y21685 , y21686 , y21687 , y21688 , y21689 , y21690 , y21691 , y21692 , y21693 , y21694 , y21695 , y21696 , y21697 , y21698 , y21699 , y21700 , y21701 , y21702 , y21703 , y21704 , y21705 , y21706 , y21707 , y21708 , y21709 , y21710 , y21711 , y21712 , y21713 , y21714 , y21715 , y21716 , y21717 , y21718 , y21719 , y21720 , y21721 , y21722 , y21723 , y21724 , y21725 , y21726 , y21727 , y21728 , y21729 , y21730 , y21731 , y21732 , y21733 , y21734 , y21735 , y21736 , y21737 , y21738 , y21739 , y21740 , y21741 , y21742 , y21743 , y21744 , y21745 , y21746 , y21747 , y21748 , y21749 , y21750 , y21751 , y21752 , y21753 , y21754 , y21755 , y21756 , y21757 , y21758 , y21759 , y21760 , y21761 , y21762 , y21763 , y21764 , y21765 , y21766 , y21767 , y21768 , y21769 , y21770 , y21771 , y21772 , y21773 , y21774 , y21775 , y21776 , y21777 , y21778 , y21779 , y21780 , y21781 , y21782 , y21783 , y21784 , y21785 , y21786 , y21787 , y21788 , y21789 , y21790 , y21791 , y21792 , y21793 , y21794 , y21795 , y21796 , y21797 , y21798 , y21799 , y21800 , y21801 , y21802 , y21803 , y21804 , y21805 , y21806 , y21807 , y21808 , y21809 , y21810 , y21811 , y21812 , y21813 , y21814 , y21815 , y21816 , y21817 , y21818 , y21819 , y21820 , y21821 , y21822 , y21823 , y21824 , y21825 , y21826 , y21827 , y21828 , y21829 , y21830 , y21831 , y21832 , y21833 , y21834 , y21835 , y21836 , y21837 , y21838 , y21839 , y21840 , y21841 , y21842 , y21843 , y21844 , y21845 , y21846 , y21847 , y21848 , y21849 , y21850 , y21851 , y21852 , y21853 , y21854 , y21855 , y21856 , y21857 , y21858 , y21859 , y21860 , y21861 , y21862 , y21863 , y21864 , y21865 , y21866 , y21867 , y21868 , y21869 , y21870 , y21871 , y21872 , y21873 , y21874 , y21875 , y21876 , y21877 , y21878 , y21879 , y21880 , y21881 , y21882 , y21883 , y21884 , y21885 , y21886 , y21887 , y21888 , y21889 , y21890 , y21891 , y21892 , y21893 , y21894 , y21895 , y21896 , y21897 , y21898 , y21899 , y21900 , y21901 , y21902 , y21903 , y21904 , y21905 , y21906 , y21907 , y21908 , y21909 , y21910 , y21911 , y21912 , y21913 , y21914 , y21915 , y21916 , y21917 , y21918 , y21919 , y21920 , y21921 , y21922 , y21923 , y21924 , y21925 , y21926 , y21927 , y21928 , y21929 , y21930 , y21931 , y21932 , y21933 , y21934 , y21935 , y21936 , y21937 , y21938 , y21939 , y21940 , y21941 , y21942 , y21943 , y21944 , y21945 , y21946 , y21947 , y21948 , y21949 , y21950 , y21951 , y21952 , y21953 , y21954 , y21955 , y21956 , y21957 , y21958 , y21959 , y21960 , y21961 , y21962 , y21963 , y21964 , y21965 , y21966 , y21967 , y21968 , y21969 , y21970 , y21971 , y21972 , y21973 , y21974 , y21975 , y21976 , y21977 , y21978 , y21979 , y21980 , y21981 , y21982 , y21983 , y21984 , y21985 , y21986 , y21987 , y21988 , y21989 , y21990 , y21991 , y21992 , y21993 , y21994 , y21995 , y21996 , y21997 , y21998 , y21999 , y22000 , y22001 , y22002 , y22003 , y22004 , y22005 , y22006 , y22007 , y22008 , y22009 , y22010 , y22011 , y22012 , y22013 , y22014 , y22015 , y22016 , y22017 , y22018 , y22019 , y22020 , y22021 , y22022 , y22023 , y22024 , y22025 , y22026 , y22027 , y22028 , y22029 , y22030 , y22031 , y22032 , y22033 , y22034 , y22035 , y22036 , y22037 , y22038 , y22039 , y22040 , y22041 , y22042 , y22043 , y22044 , y22045 , y22046 , y22047 , y22048 , y22049 , y22050 , y22051 , y22052 , y22053 , y22054 , y22055 , y22056 , y22057 , y22058 , y22059 , y22060 , y22061 , y22062 , y22063 , y22064 , y22065 , y22066 , y22067 , y22068 , y22069 , y22070 , y22071 , y22072 , y22073 , y22074 , y22075 , y22076 , y22077 , y22078 , y22079 , y22080 , y22081 , y22082 , y22083 , y22084 , y22085 , y22086 , y22087 , y22088 , y22089 , y22090 , y22091 , y22092 , y22093 , y22094 , y22095 , y22096 , y22097 , y22098 , y22099 , y22100 , y22101 , y22102 , y22103 , y22104 , y22105 , y22106 , y22107 , y22108 , y22109 , y22110 , y22111 , y22112 , y22113 , y22114 , y22115 , y22116 , y22117 , y22118 , y22119 , y22120 , y22121 , y22122 , y22123 , y22124 , y22125 , y22126 , y22127 , y22128 , y22129 , y22130 , y22131 , y22132 , y22133 , y22134 , y22135 , y22136 , y22137 , y22138 , y22139 , y22140 , y22141 , y22142 , y22143 , y22144 , y22145 , y22146 , y22147 , y22148 , y22149 , y22150 , y22151 , y22152 , y22153 , y22154 , y22155 , y22156 , y22157 , y22158 , y22159 , y22160 , y22161 , y22162 , y22163 , y22164 , y22165 , y22166 , y22167 , y22168 , y22169 , y22170 , y22171 , y22172 , y22173 , y22174 , y22175 , y22176 , y22177 , y22178 , y22179 , y22180 , y22181 , y22182 , y22183 , y22184 , y22185 , y22186 , y22187 , y22188 , y22189 , y22190 , y22191 , y22192 , y22193 , y22194 , y22195 , y22196 , y22197 , y22198 , y22199 , y22200 , y22201 , y22202 , y22203 , y22204 , y22205 , y22206 , y22207 , y22208 , y22209 , y22210 , y22211 , y22212 , y22213 , y22214 , y22215 , y22216 , y22217 , y22218 , y22219 , y22220 , y22221 , y22222 , y22223 , y22224 , y22225 , y22226 , y22227 , y22228 , y22229 , y22230 , y22231 , y22232 , y22233 , y22234 , y22235 , y22236 , y22237 , y22238 , y22239 , y22240 , y22241 , y22242 , y22243 , y22244 , y22245 , y22246 , y22247 , y22248 , y22249 , y22250 , y22251 , y22252 , y22253 , y22254 , y22255 , y22256 , y22257 , y22258 , y22259 , y22260 , y22261 , y22262 , y22263 , y22264 , y22265 , y22266 , y22267 , y22268 , y22269 , y22270 , y22271 , y22272 , y22273 , y22274 , y22275 , y22276 , y22277 , y22278 , y22279 , y22280 , y22281 , y22282 , y22283 , y22284 , y22285 , y22286 , y22287 , y22288 , y22289 , y22290 , y22291 , y22292 , y22293 , y22294 , y22295 , y22296 , y22297 , y22298 , y22299 , y22300 , y22301 , y22302 , y22303 , y22304 , y22305 , y22306 , y22307 , y22308 , y22309 , y22310 , y22311 , y22312 , y22313 , y22314 , y22315 , y22316 , y22317 , y22318 , y22319 , y22320 , y22321 , y22322 , y22323 , y22324 , y22325 , y22326 , y22327 , y22328 , y22329 , y22330 , y22331 , y22332 , y22333 , y22334 , y22335 , y22336 , y22337 , y22338 , y22339 , y22340 , y22341 , y22342 , y22343 , y22344 , y22345 , y22346 , y22347 , y22348 , y22349 , y22350 , y22351 , y22352 , y22353 , y22354 , y22355 , y22356 , y22357 , y22358 , y22359 , y22360 , y22361 , y22362 , y22363 , y22364 , y22365 , y22366 , y22367 , y22368 , y22369 , y22370 , y22371 , y22372 , y22373 , y22374 , y22375 , y22376 , y22377 , y22378 , y22379 , y22380 , y22381 , y22382 , y22383 , y22384 , y22385 , y22386 , y22387 , y22388 , y22389 , y22390 , y22391 , y22392 , y22393 , y22394 , y22395 , y22396 , y22397 , y22398 , y22399 , y22400 , y22401 , y22402 , y22403 , y22404 , y22405 , y22406 , y22407 , y22408 , y22409 , y22410 , y22411 , y22412 , y22413 , y22414 , y22415 , y22416 , y22417 , y22418 , y22419 , y22420 , y22421 , y22422 , y22423 , y22424 , y22425 , y22426 , y22427 , y22428 , y22429 , y22430 , y22431 , y22432 , y22433 , y22434 , y22435 , y22436 , y22437 , y22438 , y22439 , y22440 , y22441 , y22442 , y22443 , y22444 , y22445 , y22446 , y22447 , y22448 , y22449 , y22450 , y22451 , y22452 , y22453 , y22454 , y22455 , y22456 , y22457 , y22458 , y22459 , y22460 , y22461 , y22462 , y22463 , y22464 , y22465 , y22466 , y22467 , y22468 , y22469 , y22470 , y22471 , y22472 , y22473 , y22474 , y22475 , y22476 , y22477 , y22478 , y22479 , y22480 , y22481 , y22482 , y22483 , y22484 , y22485 , y22486 , y22487 , y22488 , y22489 , y22490 , y22491 , y22492 , y22493 , y22494 , y22495 , y22496 , y22497 , y22498 , y22499 , y22500 , y22501 , y22502 , y22503 , y22504 , y22505 , y22506 , y22507 , y22508 , y22509 , y22510 , y22511 , y22512 , y22513 , y22514 , y22515 , y22516 , y22517 , y22518 , y22519 , y22520 , y22521 , y22522 , y22523 , y22524 , y22525 , y22526 , y22527 , y22528 , y22529 , y22530 , y22531 , y22532 , y22533 , y22534 , y22535 , y22536 , y22537 , y22538 , y22539 , y22540 , y22541 , y22542 , y22543 , y22544 , y22545 , y22546 , y22547 , y22548 , y22549 , y22550 , y22551 , y22552 , y22553 , y22554 , y22555 , y22556 , y22557 , y22558 , y22559 , y22560 , y22561 , y22562 , y22563 , y22564 , y22565 , y22566 , y22567 , y22568 , y22569 , y22570 , y22571 , y22572 , y22573 , y22574 , y22575 , y22576 , y22577 , y22578 , y22579 , y22580 , y22581 , y22582 , y22583 , y22584 , y22585 , y22586 , y22587 , y22588 , y22589 , y22590 , y22591 , y22592 , y22593 , y22594 , y22595 , y22596 , y22597 , y22598 , y22599 , y22600 , y22601 , y22602 , y22603 , y22604 , y22605 , y22606 , y22607 , y22608 , y22609 , y22610 , y22611 , y22612 , y22613 , y22614 , y22615 , y22616 , y22617 , y22618 , y22619 , y22620 , y22621 , y22622 , y22623 , y22624 , y22625 , y22626 , y22627 , y22628 , y22629 , y22630 , y22631 , y22632 , y22633 , y22634 , y22635 , y22636 , y22637 , y22638 , y22639 , y22640 , y22641 , y22642 , y22643 , y22644 , y22645 , y22646 , y22647 , y22648 , y22649 , y22650 , y22651 , y22652 , y22653 , y22654 , y22655 , y22656 , y22657 , y22658 , y22659 , y22660 , y22661 , y22662 , y22663 , y22664 , y22665 , y22666 , y22667 , y22668 , y22669 , y22670 , y22671 , y22672 , y22673 , y22674 , y22675 , y22676 , y22677 , y22678 , y22679 , y22680 , y22681 , y22682 , y22683 , y22684 , y22685 , y22686 , y22687 , y22688 , y22689 , y22690 , y22691 , y22692 , y22693 , y22694 , y22695 , y22696 , y22697 , y22698 , y22699 , y22700 , y22701 , y22702 , y22703 , y22704 , y22705 , y22706 , y22707 , y22708 , y22709 , y22710 , y22711 , y22712 , y22713 , y22714 , y22715 , y22716 , y22717 , y22718 , y22719 , y22720 , y22721 , y22722 , y22723 , y22724 , y22725 , y22726 , y22727 , y22728 , y22729 , y22730 , y22731 , y22732 , y22733 , y22734 , y22735 , y22736 , y22737 , y22738 , y22739 , y22740 , y22741 , y22742 , y22743 , y22744 , y22745 , y22746 , y22747 , y22748 , y22749 , y22750 , y22751 , y22752 , y22753 , y22754 , y22755 , y22756 , y22757 , y22758 , y22759 , y22760 , y22761 , y22762 , y22763 , y22764 , y22765 , y22766 , y22767 , y22768 , y22769 , y22770 , y22771 , y22772 , y22773 , y22774 , y22775 , y22776 , y22777 , y22778 , y22779 , y22780 , y22781 , y22782 , y22783 , y22784 , y22785 , y22786 , y22787 , y22788 , y22789 , y22790 , y22791 , y22792 , y22793 , y22794 , y22795 , y22796 , y22797 , y22798 , y22799 , y22800 , y22801 , y22802 , y22803 , y22804 , y22805 , y22806 , y22807 , y22808 , y22809 , y22810 , y22811 , y22812 , y22813 , y22814 , y22815 , y22816 , y22817 , y22818 , y22819 , y22820 , y22821 , y22822 , y22823 , y22824 , y22825 , y22826 , y22827 , y22828 , y22829 , y22830 , y22831 , y22832 , y22833 , y22834 , y22835 , y22836 , y22837 , y22838 , y22839 , y22840 , y22841 , y22842 , y22843 , y22844 , y22845 , y22846 , y22847 , y22848 , y22849 , y22850 , y22851 , y22852 , y22853 , y22854 , y22855 , y22856 , y22857 , y22858 , y22859 , y22860 , y22861 , y22862 , y22863 , y22864 , y22865 , y22866 , y22867 , y22868 , y22869 , y22870 , y22871 , y22872 , y22873 , y22874 , y22875 , y22876 , y22877 , y22878 , y22879 , y22880 , y22881 , y22882 , y22883 , y22884 , y22885 , y22886 , y22887 , y22888 , y22889 , y22890 , y22891 , y22892 , y22893 , y22894 , y22895 , y22896 , y22897 , y22898 , y22899 , y22900 , y22901 , y22902 , y22903 , y22904 , y22905 , y22906 , y22907 , y22908 , y22909 , y22910 , y22911 , y22912 , y22913 , y22914 , y22915 , y22916 , y22917 , y22918 , y22919 , y22920 , y22921 , y22922 , y22923 , y22924 , y22925 , y22926 , y22927 , y22928 , y22929 , y22930 , y22931 , y22932 , y22933 , y22934 , y22935 , y22936 , y22937 , y22938 , y22939 , y22940 , y22941 , y22942 , y22943 , y22944 , y22945 , y22946 , y22947 , y22948 , y22949 , y22950 , y22951 , y22952 , y22953 , y22954 , y22955 , y22956 , y22957 , y22958 , y22959 , y22960 , y22961 , y22962 , y22963 , y22964 , y22965 , y22966 , y22967 , y22968 , y22969 , y22970 , y22971 , y22972 , y22973 , y22974 , y22975 , y22976 , y22977 , y22978 , y22979 , y22980 , y22981 , y22982 , y22983 , y22984 , y22985 , y22986 , y22987 , y22988 , y22989 , y22990 , y22991 , y22992 , y22993 , y22994 , y22995 , y22996 , y22997 , y22998 , y22999 , y23000 , y23001 , y23002 , y23003 , y23004 , y23005 , y23006 , y23007 , y23008 , y23009 , y23010 , y23011 , y23012 , y23013 , y23014 , y23015 , y23016 , y23017 , y23018 , y23019 , y23020 , y23021 , y23022 , y23023 , y23024 , y23025 , y23026 , y23027 , y23028 , y23029 , y23030 , y23031 , y23032 , y23033 , y23034 , y23035 , y23036 , y23037 , y23038 , y23039 , y23040 , y23041 , y23042 , y23043 , y23044 , y23045 , y23046 , y23047 , y23048 , y23049 , y23050 , y23051 , y23052 , y23053 , y23054 , y23055 , y23056 , y23057 , y23058 , y23059 , y23060 , y23061 , y23062 , y23063 , y23064 , y23065 , y23066 , y23067 , y23068 , y23069 , y23070 , y23071 , y23072 , y23073 , y23074 , y23075 , y23076 , y23077 , y23078 , y23079 , y23080 , y23081 , y23082 , y23083 , y23084 , y23085 , y23086 , y23087 , y23088 , y23089 , y23090 , y23091 , y23092 , y23093 , y23094 , y23095 , y23096 , y23097 , y23098 , y23099 , y23100 , y23101 , y23102 , y23103 , y23104 , y23105 , y23106 , y23107 , y23108 , y23109 , y23110 , y23111 , y23112 , y23113 , y23114 , y23115 , y23116 , y23117 , y23118 , y23119 , y23120 , y23121 , y23122 , y23123 , y23124 , y23125 , y23126 , y23127 , y23128 , y23129 , y23130 , y23131 , y23132 , y23133 , y23134 , y23135 , y23136 , y23137 , y23138 , y23139 , y23140 , y23141 , y23142 , y23143 , y23144 , y23145 , y23146 , y23147 , y23148 , y23149 , y23150 , y23151 , y23152 , y23153 , y23154 , y23155 , y23156 , y23157 , y23158 , y23159 , y23160 , y23161 , y23162 , y23163 , y23164 , y23165 , y23166 , y23167 , y23168 , y23169 , y23170 , y23171 , y23172 , y23173 , y23174 , y23175 , y23176 , y23177 , y23178 , y23179 , y23180 , y23181 , y23182 , y23183 , y23184 , y23185 , y23186 , y23187 , y23188 , y23189 , y23190 , y23191 , y23192 , y23193 , y23194 , y23195 , y23196 , y23197 , y23198 , y23199 , y23200 , y23201 , y23202 , y23203 , y23204 , y23205 , y23206 , y23207 , y23208 , y23209 , y23210 , y23211 , y23212 , y23213 , y23214 , y23215 , y23216 , y23217 , y23218 , y23219 , y23220 , y23221 , y23222 , y23223 , y23224 , y23225 , y23226 , y23227 , y23228 , y23229 , y23230 , y23231 , y23232 , y23233 , y23234 , y23235 , y23236 , y23237 , y23238 , y23239 , y23240 , y23241 , y23242 , y23243 , y23244 , y23245 , y23246 , y23247 , y23248 , y23249 , y23250 , y23251 , y23252 , y23253 , y23254 , y23255 , y23256 , y23257 , y23258 , y23259 , y23260 , y23261 , y23262 , y23263 , y23264 , y23265 , y23266 , y23267 , y23268 , y23269 , y23270 , y23271 , y23272 , y23273 , y23274 , y23275 , y23276 , y23277 , y23278 , y23279 , y23280 , y23281 , y23282 , y23283 , y23284 , y23285 , y23286 , y23287 , y23288 , y23289 , y23290 , y23291 , y23292 , y23293 , y23294 , y23295 , y23296 , y23297 , y23298 , y23299 , y23300 , y23301 , y23302 , y23303 , y23304 , y23305 , y23306 , y23307 , y23308 , y23309 , y23310 , y23311 , y23312 , y23313 , y23314 , y23315 , y23316 , y23317 , y23318 , y23319 , y23320 , y23321 , y23322 , y23323 , y23324 , y23325 , y23326 , y23327 , y23328 , y23329 , y23330 , y23331 , y23332 , y23333 , y23334 , y23335 , y23336 , y23337 , y23338 , y23339 , y23340 , y23341 , y23342 , y23343 , y23344 , y23345 , y23346 , y23347 , y23348 , y23349 , y23350 , y23351 , y23352 , y23353 , y23354 , y23355 , y23356 , y23357 , y23358 , y23359 , y23360 , y23361 , y23362 , y23363 , y23364 , y23365 , y23366 , y23367 , y23368 , y23369 , y23370 , y23371 , y23372 , y23373 , y23374 , y23375 , y23376 , y23377 , y23378 , y23379 , y23380 , y23381 , y23382 , y23383 , y23384 , y23385 , y23386 , y23387 , y23388 , y23389 , y23390 , y23391 , y23392 , y23393 , y23394 , y23395 , y23396 , y23397 , y23398 , y23399 , y23400 , y23401 , y23402 , y23403 , y23404 , y23405 , y23406 , y23407 , y23408 , y23409 , y23410 , y23411 , y23412 , y23413 , y23414 , y23415 , y23416 , y23417 , y23418 , y23419 , y23420 , y23421 , y23422 , y23423 , y23424 , y23425 , y23426 , y23427 , y23428 , y23429 , y23430 , y23431 , y23432 , y23433 , y23434 , y23435 , y23436 , y23437 , y23438 , y23439 , y23440 , y23441 , y23442 , y23443 , y23444 , y23445 , y23446 , y23447 , y23448 , y23449 , y23450 , y23451 , y23452 , y23453 , y23454 , y23455 , y23456 , y23457 , y23458 , y23459 , y23460 , y23461 , y23462 , y23463 , y23464 , y23465 , y23466 , y23467 , y23468 , y23469 , y23470 , y23471 , y23472 , y23473 , y23474 , y23475 , y23476 , y23477 , y23478 , y23479 , y23480 , y23481 , y23482 , y23483 , y23484 , y23485 , y23486 , y23487 , y23488 , y23489 , y23490 , y23491 , y23492 , y23493 , y23494 , y23495 , y23496 , y23497 , y23498 , y23499 , y23500 , y23501 , y23502 , y23503 , y23504 , y23505 , y23506 , y23507 , y23508 , y23509 , y23510 , y23511 , y23512 , y23513 , y23514 , y23515 , y23516 , y23517 , y23518 , y23519 , y23520 , y23521 , y23522 , y23523 , y23524 , y23525 , y23526 , y23527 , y23528 , y23529 , y23530 , y23531 , y23532 , y23533 , y23534 , y23535 , y23536 , y23537 , y23538 , y23539 , y23540 , y23541 , y23542 , y23543 , y23544 , y23545 , y23546 , y23547 , y23548 , y23549 , y23550 , y23551 , y23552 , y23553 , y23554 , y23555 , y23556 , y23557 , y23558 , y23559 , y23560 , y23561 , y23562 , y23563 , y23564 , y23565 , y23566 , y23567 , y23568 , y23569 , y23570 , y23571 , y23572 , y23573 , y23574 , y23575 , y23576 , y23577 , y23578 , y23579 , y23580 , y23581 , y23582 , y23583 , y23584 , y23585 , y23586 , y23587 , y23588 , y23589 , y23590 , y23591 , y23592 , y23593 , y23594 , y23595 , y23596 , y23597 , y23598 , y23599 , y23600 , y23601 , y23602 , y23603 , y23604 , y23605 , y23606 , y23607 , y23608 , y23609 , y23610 , y23611 , y23612 , y23613 , y23614 , y23615 , y23616 , y23617 , y23618 , y23619 , y23620 , y23621 , y23622 , y23623 , y23624 , y23625 , y23626 , y23627 , y23628 , y23629 , y23630 , y23631 , y23632 , y23633 , y23634 , y23635 , y23636 , y23637 , y23638 , y23639 , y23640 , y23641 , y23642 , y23643 , y23644 , y23645 , y23646 , y23647 , y23648 , y23649 , y23650 , y23651 , y23652 , y23653 , y23654 , y23655 , y23656 , y23657 , y23658 , y23659 , y23660 , y23661 , y23662 , y23663 , y23664 , y23665 , y23666 , y23667 , y23668 , y23669 , y23670 , y23671 , y23672 , y23673 , y23674 , y23675 , y23676 , y23677 , y23678 , y23679 , y23680 , y23681 , y23682 , y23683 , y23684 , y23685 , y23686 , y23687 , y23688 , y23689 , y23690 , y23691 , y23692 , y23693 , y23694 , y23695 , y23696 , y23697 , y23698 , y23699 , y23700 , y23701 , y23702 , y23703 , y23704 , y23705 , y23706 , y23707 , y23708 , y23709 , y23710 , y23711 , y23712 , y23713 , y23714 , y23715 , y23716 , y23717 , y23718 , y23719 , y23720 , y23721 , y23722 , y23723 , y23724 , y23725 , y23726 , y23727 , y23728 , y23729 , y23730 , y23731 , y23732 , y23733 , y23734 , y23735 , y23736 , y23737 , y23738 , y23739 , y23740 , y23741 , y23742 , y23743 , y23744 , y23745 , y23746 , y23747 , y23748 , y23749 , y23750 , y23751 , y23752 , y23753 , y23754 , y23755 , y23756 , y23757 , y23758 , y23759 , y23760 , y23761 , y23762 , y23763 , y23764 , y23765 , y23766 , y23767 , y23768 , y23769 , y23770 , y23771 , y23772 , y23773 , y23774 , y23775 , y23776 , y23777 , y23778 , y23779 , y23780 , y23781 , y23782 , y23783 , y23784 , y23785 , y23786 , y23787 , y23788 , y23789 , y23790 , y23791 , y23792 , y23793 , y23794 , y23795 , y23796 , y23797 , y23798 , y23799 , y23800 , y23801 , y23802 , y23803 , y23804 , y23805 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 , y20242 , y20243 , y20244 , y20245 , y20246 , y20247 , y20248 , y20249 , y20250 , y20251 , y20252 , y20253 , y20254 , y20255 , y20256 , y20257 , y20258 , y20259 , y20260 , y20261 , y20262 , y20263 , y20264 , y20265 , y20266 , y20267 , y20268 , y20269 , y20270 , y20271 , y20272 , y20273 , y20274 , y20275 , y20276 , y20277 , y20278 , y20279 , y20280 , y20281 , y20282 , y20283 , y20284 , y20285 , y20286 , y20287 , y20288 , y20289 , y20290 , y20291 , y20292 , y20293 , y20294 , y20295 , y20296 , y20297 , y20298 , y20299 , y20300 , y20301 , y20302 , y20303 , y20304 , y20305 , y20306 , y20307 , y20308 , y20309 , y20310 , y20311 , y20312 , y20313 , y20314 , y20315 , y20316 , y20317 , y20318 , y20319 , y20320 , y20321 , y20322 , y20323 , y20324 , y20325 , y20326 , y20327 , y20328 , y20329 , y20330 , y20331 , y20332 , y20333 , y20334 , y20335 , y20336 , y20337 , y20338 , y20339 , y20340 , y20341 , y20342 , y20343 , y20344 , y20345 , y20346 , y20347 , y20348 , y20349 , y20350 , y20351 , y20352 , y20353 , y20354 , y20355 , y20356 , y20357 , y20358 , y20359 , y20360 , y20361 , y20362 , y20363 , y20364 , y20365 , y20366 , y20367 , y20368 , y20369 , y20370 , y20371 , y20372 , y20373 , y20374 , y20375 , y20376 , y20377 , y20378 , y20379 , y20380 , y20381 , y20382 , y20383 , y20384 , y20385 , y20386 , y20387 , y20388 , y20389 , y20390 , y20391 , y20392 , y20393 , y20394 , y20395 , y20396 , y20397 , y20398 , y20399 , y20400 , y20401 , y20402 , y20403 , y20404 , y20405 , y20406 , y20407 , y20408 , y20409 , y20410 , y20411 , y20412 , y20413 , y20414 , y20415 , y20416 , y20417 , y20418 , y20419 , y20420 , y20421 , y20422 , y20423 , y20424 , y20425 , y20426 , y20427 , y20428 , y20429 , y20430 , y20431 , y20432 , y20433 , y20434 , y20435 , y20436 , y20437 , y20438 , y20439 , y20440 , y20441 , y20442 , y20443 , y20444 , y20445 , y20446 , y20447 , y20448 , y20449 , y20450 , y20451 , y20452 , y20453 , y20454 , y20455 , y20456 , y20457 , y20458 , y20459 , y20460 , y20461 , y20462 , y20463 , y20464 , y20465 , y20466 , y20467 , y20468 , y20469 , y20470 , y20471 , y20472 , y20473 , y20474 , y20475 , y20476 , y20477 , y20478 , y20479 , y20480 , y20481 , y20482 , y20483 , y20484 , y20485 , y20486 , y20487 , y20488 , y20489 , y20490 , y20491 , y20492 , y20493 , y20494 , y20495 , y20496 , y20497 , y20498 , y20499 , y20500 , y20501 , y20502 , y20503 , y20504 , y20505 , y20506 , y20507 , y20508 , y20509 , y20510 , y20511 , y20512 , y20513 , y20514 , y20515 , y20516 , y20517 , y20518 , y20519 , y20520 , y20521 , y20522 , y20523 , y20524 , y20525 , y20526 , y20527 , y20528 , y20529 , y20530 , y20531 , y20532 , y20533 , y20534 , y20535 , y20536 , y20537 , y20538 , y20539 , y20540 , y20541 , y20542 , y20543 , y20544 , y20545 , y20546 , y20547 , y20548 , y20549 , y20550 , y20551 , y20552 , y20553 , y20554 , y20555 , y20556 , y20557 , y20558 , y20559 , y20560 , y20561 , y20562 , y20563 , y20564 , y20565 , y20566 , y20567 , y20568 , y20569 , y20570 , y20571 , y20572 , y20573 , y20574 , y20575 , y20576 , y20577 , y20578 , y20579 , y20580 , y20581 , y20582 , y20583 , y20584 , y20585 , y20586 , y20587 , y20588 , y20589 , y20590 , y20591 , y20592 , y20593 , y20594 , y20595 , y20596 , y20597 , y20598 , y20599 , y20600 , y20601 , y20602 , y20603 , y20604 , y20605 , y20606 , y20607 , y20608 , y20609 , y20610 , y20611 , y20612 , y20613 , y20614 , y20615 , y20616 , y20617 , y20618 , y20619 , y20620 , y20621 , y20622 , y20623 , y20624 , y20625 , y20626 , y20627 , y20628 , y20629 , y20630 , y20631 , y20632 , y20633 , y20634 , y20635 , y20636 , y20637 , y20638 , y20639 , y20640 , y20641 , y20642 , y20643 , y20644 , y20645 , y20646 , y20647 , y20648 , y20649 , y20650 , y20651 , y20652 , y20653 , y20654 , y20655 , y20656 , y20657 , y20658 , y20659 , y20660 , y20661 , y20662 , y20663 , y20664 , y20665 , y20666 , y20667 , y20668 , y20669 , y20670 , y20671 , y20672 , y20673 , y20674 , y20675 , y20676 , y20677 , y20678 , y20679 , y20680 , y20681 , y20682 , y20683 , y20684 , y20685 , y20686 , y20687 , y20688 , y20689 , y20690 , y20691 , y20692 , y20693 , y20694 , y20695 , y20696 , y20697 , y20698 , y20699 , y20700 , y20701 , y20702 , y20703 , y20704 , y20705 , y20706 , y20707 , y20708 , y20709 , y20710 , y20711 , y20712 , y20713 , y20714 , y20715 , y20716 , y20717 , y20718 , y20719 , y20720 , y20721 , y20722 , y20723 , y20724 , y20725 , y20726 , y20727 , y20728 , y20729 , y20730 , y20731 , y20732 , y20733 , y20734 , y20735 , y20736 , y20737 , y20738 , y20739 , y20740 , y20741 , y20742 , y20743 , y20744 , y20745 , y20746 , y20747 , y20748 , y20749 , y20750 , y20751 , y20752 , y20753 , y20754 , y20755 , y20756 , y20757 , y20758 , y20759 , y20760 , y20761 , y20762 , y20763 , y20764 , y20765 , y20766 , y20767 , y20768 , y20769 , y20770 , y20771 , y20772 , y20773 , y20774 , y20775 , y20776 , y20777 , y20778 , y20779 , y20780 , y20781 , y20782 , y20783 , y20784 , y20785 , y20786 , y20787 , y20788 , y20789 , y20790 , y20791 , y20792 , y20793 , y20794 , y20795 , y20796 , y20797 , y20798 , y20799 , y20800 , y20801 , y20802 , y20803 , y20804 , y20805 , y20806 , y20807 , y20808 , y20809 , y20810 , y20811 , y20812 , y20813 , y20814 , y20815 , y20816 , y20817 , y20818 , y20819 , y20820 , y20821 , y20822 , y20823 , y20824 , y20825 , y20826 , y20827 , y20828 , y20829 , y20830 , y20831 , y20832 , y20833 , y20834 , y20835 , y20836 , y20837 , y20838 , y20839 , y20840 , y20841 , y20842 , y20843 , y20844 , y20845 , y20846 , y20847 , y20848 , y20849 , y20850 , y20851 , y20852 , y20853 , y20854 , y20855 , y20856 , y20857 , y20858 , y20859 , y20860 , y20861 , y20862 , y20863 , y20864 , y20865 , y20866 , y20867 , y20868 , y20869 , y20870 , y20871 , y20872 , y20873 , y20874 , y20875 , y20876 , y20877 , y20878 , y20879 , y20880 , y20881 , y20882 , y20883 , y20884 , y20885 , y20886 , y20887 , y20888 , y20889 , y20890 , y20891 , y20892 , y20893 , y20894 , y20895 , y20896 , y20897 , y20898 , y20899 , y20900 , y20901 , y20902 , y20903 , y20904 , y20905 , y20906 , y20907 , y20908 , y20909 , y20910 , y20911 , y20912 , y20913 , y20914 , y20915 , y20916 , y20917 , y20918 , y20919 , y20920 , y20921 , y20922 , y20923 , y20924 , y20925 , y20926 , y20927 , y20928 , y20929 , y20930 , y20931 , y20932 , y20933 , y20934 , y20935 , y20936 , y20937 , y20938 , y20939 , y20940 , y20941 , y20942 , y20943 , y20944 , y20945 , y20946 , y20947 , y20948 , y20949 , y20950 , y20951 , y20952 , y20953 , y20954 , y20955 , y20956 , y20957 , y20958 , y20959 , y20960 , y20961 , y20962 , y20963 , y20964 , y20965 , y20966 , y20967 , y20968 , y20969 , y20970 , y20971 , y20972 , y20973 , y20974 , y20975 , y20976 , y20977 , y20978 , y20979 , y20980 , y20981 , y20982 , y20983 , y20984 , y20985 , y20986 , y20987 , y20988 , y20989 , y20990 , y20991 , y20992 , y20993 , y20994 , y20995 , y20996 , y20997 , y20998 , y20999 , y21000 , y21001 , y21002 , y21003 , y21004 , y21005 , y21006 , y21007 , y21008 , y21009 , y21010 , y21011 , y21012 , y21013 , y21014 , y21015 , y21016 , y21017 , y21018 , y21019 , y21020 , y21021 , y21022 , y21023 , y21024 , y21025 , y21026 , y21027 , y21028 , y21029 , y21030 , y21031 , y21032 , y21033 , y21034 , y21035 , y21036 , y21037 , y21038 , y21039 , y21040 , y21041 , y21042 , y21043 , y21044 , y21045 , y21046 , y21047 , y21048 , y21049 , y21050 , y21051 , y21052 , y21053 , y21054 , y21055 , y21056 , y21057 , y21058 , y21059 , y21060 , y21061 , y21062 , y21063 , y21064 , y21065 , y21066 , y21067 , y21068 , y21069 , y21070 , y21071 , y21072 , y21073 , y21074 , y21075 , y21076 , y21077 , y21078 , y21079 , y21080 , y21081 , y21082 , y21083 , y21084 , y21085 , y21086 , y21087 , y21088 , y21089 , y21090 , y21091 , y21092 , y21093 , y21094 , y21095 , y21096 , y21097 , y21098 , y21099 , y21100 , y21101 , y21102 , y21103 , y21104 , y21105 , y21106 , y21107 , y21108 , y21109 , y21110 , y21111 , y21112 , y21113 , y21114 , y21115 , y21116 , y21117 , y21118 , y21119 , y21120 , y21121 , y21122 , y21123 , y21124 , y21125 , y21126 , y21127 , y21128 , y21129 , y21130 , y21131 , y21132 , y21133 , y21134 , y21135 , y21136 , y21137 , y21138 , y21139 , y21140 , y21141 , y21142 , y21143 , y21144 , y21145 , y21146 , y21147 , y21148 , y21149 , y21150 , y21151 , y21152 , y21153 , y21154 , y21155 , y21156 , y21157 , y21158 , y21159 , y21160 , y21161 , y21162 , y21163 , y21164 , y21165 , y21166 , y21167 , y21168 , y21169 , y21170 , y21171 , y21172 , y21173 , y21174 , y21175 , y21176 , y21177 , y21178 , y21179 , y21180 , y21181 , y21182 , y21183 , y21184 , y21185 , y21186 , y21187 , y21188 , y21189 , y21190 , y21191 , y21192 , y21193 , y21194 , y21195 , y21196 , y21197 , y21198 , y21199 , y21200 , y21201 , y21202 , y21203 , y21204 , y21205 , y21206 , y21207 , y21208 , y21209 , y21210 , y21211 , y21212 , y21213 , y21214 , y21215 , y21216 , y21217 , y21218 , y21219 , y21220 , y21221 , y21222 , y21223 , y21224 , y21225 , y21226 , y21227 , y21228 , y21229 , y21230 , y21231 , y21232 , y21233 , y21234 , y21235 , y21236 , y21237 , y21238 , y21239 , y21240 , y21241 , y21242 , y21243 , y21244 , y21245 , y21246 , y21247 , y21248 , y21249 , y21250 , y21251 , y21252 , y21253 , y21254 , y21255 , y21256 , y21257 , y21258 , y21259 , y21260 , y21261 , y21262 , y21263 , y21264 , y21265 , y21266 , y21267 , y21268 , y21269 , y21270 , y21271 , y21272 , y21273 , y21274 , y21275 , y21276 , y21277 , y21278 , y21279 , y21280 , y21281 , y21282 , y21283 , y21284 , y21285 , y21286 , y21287 , y21288 , y21289 , y21290 , y21291 , y21292 , y21293 , y21294 , y21295 , y21296 , y21297 , y21298 , y21299 , y21300 , y21301 , y21302 , y21303 , y21304 , y21305 , y21306 , y21307 , y21308 , y21309 , y21310 , y21311 , y21312 , y21313 , y21314 , y21315 , y21316 , y21317 , y21318 , y21319 , y21320 , y21321 , y21322 , y21323 , y21324 , y21325 , y21326 , y21327 , y21328 , y21329 , y21330 , y21331 , y21332 , y21333 , y21334 , y21335 , y21336 , y21337 , y21338 , y21339 , y21340 , y21341 , y21342 , y21343 , y21344 , y21345 , y21346 , y21347 , y21348 , y21349 , y21350 , y21351 , y21352 , y21353 , y21354 , y21355 , y21356 , y21357 , y21358 , y21359 , y21360 , y21361 , y21362 , y21363 , y21364 , y21365 , y21366 , y21367 , y21368 , y21369 , y21370 , y21371 , y21372 , y21373 , y21374 , y21375 , y21376 , y21377 , y21378 , y21379 , y21380 , y21381 , y21382 , y21383 , y21384 , y21385 , y21386 , y21387 , y21388 , y21389 , y21390 , y21391 , y21392 , y21393 , y21394 , y21395 , y21396 , y21397 , y21398 , y21399 , y21400 , y21401 , y21402 , y21403 , y21404 , y21405 , y21406 , y21407 , y21408 , y21409 , y21410 , y21411 , y21412 , y21413 , y21414 , y21415 , y21416 , y21417 , y21418 , y21419 , y21420 , y21421 , y21422 , y21423 , y21424 , y21425 , y21426 , y21427 , y21428 , y21429 , y21430 , y21431 , y21432 , y21433 , y21434 , y21435 , y21436 , y21437 , y21438 , y21439 , y21440 , y21441 , y21442 , y21443 , y21444 , y21445 , y21446 , y21447 , y21448 , y21449 , y21450 , y21451 , y21452 , y21453 , y21454 , y21455 , y21456 , y21457 , y21458 , y21459 , y21460 , y21461 , y21462 , y21463 , y21464 , y21465 , y21466 , y21467 , y21468 , y21469 , y21470 , y21471 , y21472 , y21473 , y21474 , y21475 , y21476 , y21477 , y21478 , y21479 , y21480 , y21481 , y21482 , y21483 , y21484 , y21485 , y21486 , y21487 , y21488 , y21489 , y21490 , y21491 , y21492 , y21493 , y21494 , y21495 , y21496 , y21497 , y21498 , y21499 , y21500 , y21501 , y21502 , y21503 , y21504 , y21505 , y21506 , y21507 , y21508 , y21509 , y21510 , y21511 , y21512 , y21513 , y21514 , y21515 , y21516 , y21517 , y21518 , y21519 , y21520 , y21521 , y21522 , y21523 , y21524 , y21525 , y21526 , y21527 , y21528 , y21529 , y21530 , y21531 , y21532 , y21533 , y21534 , y21535 , y21536 , y21537 , y21538 , y21539 , y21540 , y21541 , y21542 , y21543 , y21544 , y21545 , y21546 , y21547 , y21548 , y21549 , y21550 , y21551 , y21552 , y21553 , y21554 , y21555 , y21556 , y21557 , y21558 , y21559 , y21560 , y21561 , y21562 , y21563 , y21564 , y21565 , y21566 , y21567 , y21568 , y21569 , y21570 , y21571 , y21572 , y21573 , y21574 , y21575 , y21576 , y21577 , y21578 , y21579 , y21580 , y21581 , y21582 , y21583 , y21584 , y21585 , y21586 , y21587 , y21588 , y21589 , y21590 , y21591 , y21592 , y21593 , y21594 , y21595 , y21596 , y21597 , y21598 , y21599 , y21600 , y21601 , y21602 , y21603 , y21604 , y21605 , y21606 , y21607 , y21608 , y21609 , y21610 , y21611 , y21612 , y21613 , y21614 , y21615 , y21616 , y21617 , y21618 , y21619 , y21620 , y21621 , y21622 , y21623 , y21624 , y21625 , y21626 , y21627 , y21628 , y21629 , y21630 , y21631 , y21632 , y21633 , y21634 , y21635 , y21636 , y21637 , y21638 , y21639 , y21640 , y21641 , y21642 , y21643 , y21644 , y21645 , y21646 , y21647 , y21648 , y21649 , y21650 , y21651 , y21652 , y21653 , y21654 , y21655 , y21656 , y21657 , y21658 , y21659 , y21660 , y21661 , y21662 , y21663 , y21664 , y21665 , y21666 , y21667 , y21668 , y21669 , y21670 , y21671 , y21672 , y21673 , y21674 , y21675 , y21676 , y21677 , y21678 , y21679 , y21680 , y21681 , y21682 , y21683 , y21684 , y21685 , y21686 , y21687 , y21688 , y21689 , y21690 , y21691 , y21692 , y21693 , y21694 , y21695 , y21696 , y21697 , y21698 , y21699 , y21700 , y21701 , y21702 , y21703 , y21704 , y21705 , y21706 , y21707 , y21708 , y21709 , y21710 , y21711 , y21712 , y21713 , y21714 , y21715 , y21716 , y21717 , y21718 , y21719 , y21720 , y21721 , y21722 , y21723 , y21724 , y21725 , y21726 , y21727 , y21728 , y21729 , y21730 , y21731 , y21732 , y21733 , y21734 , y21735 , y21736 , y21737 , y21738 , y21739 , y21740 , y21741 , y21742 , y21743 , y21744 , y21745 , y21746 , y21747 , y21748 , y21749 , y21750 , y21751 , y21752 , y21753 , y21754 , y21755 , y21756 , y21757 , y21758 , y21759 , y21760 , y21761 , y21762 , y21763 , y21764 , y21765 , y21766 , y21767 , y21768 , y21769 , y21770 , y21771 , y21772 , y21773 , y21774 , y21775 , y21776 , y21777 , y21778 , y21779 , y21780 , y21781 , y21782 , y21783 , y21784 , y21785 , y21786 , y21787 , y21788 , y21789 , y21790 , y21791 , y21792 , y21793 , y21794 , y21795 , y21796 , y21797 , y21798 , y21799 , y21800 , y21801 , y21802 , y21803 , y21804 , y21805 , y21806 , y21807 , y21808 , y21809 , y21810 , y21811 , y21812 , y21813 , y21814 , y21815 , y21816 , y21817 , y21818 , y21819 , y21820 , y21821 , y21822 , y21823 , y21824 , y21825 , y21826 , y21827 , y21828 , y21829 , y21830 , y21831 , y21832 , y21833 , y21834 , y21835 , y21836 , y21837 , y21838 , y21839 , y21840 , y21841 , y21842 , y21843 , y21844 , y21845 , y21846 , y21847 , y21848 , y21849 , y21850 , y21851 , y21852 , y21853 , y21854 , y21855 , y21856 , y21857 , y21858 , y21859 , y21860 , y21861 , y21862 , y21863 , y21864 , y21865 , y21866 , y21867 , y21868 , y21869 , y21870 , y21871 , y21872 , y21873 , y21874 , y21875 , y21876 , y21877 , y21878 , y21879 , y21880 , y21881 , y21882 , y21883 , y21884 , y21885 , y21886 , y21887 , y21888 , y21889 , y21890 , y21891 , y21892 , y21893 , y21894 , y21895 , y21896 , y21897 , y21898 , y21899 , y21900 , y21901 , y21902 , y21903 , y21904 , y21905 , y21906 , y21907 , y21908 , y21909 , y21910 , y21911 , y21912 , y21913 , y21914 , y21915 , y21916 , y21917 , y21918 , y21919 , y21920 , y21921 , y21922 , y21923 , y21924 , y21925 , y21926 , y21927 , y21928 , y21929 , y21930 , y21931 , y21932 , y21933 , y21934 , y21935 , y21936 , y21937 , y21938 , y21939 , y21940 , y21941 , y21942 , y21943 , y21944 , y21945 , y21946 , y21947 , y21948 , y21949 , y21950 , y21951 , y21952 , y21953 , y21954 , y21955 , y21956 , y21957 , y21958 , y21959 , y21960 , y21961 , y21962 , y21963 , y21964 , y21965 , y21966 , y21967 , y21968 , y21969 , y21970 , y21971 , y21972 , y21973 , y21974 , y21975 , y21976 , y21977 , y21978 , y21979 , y21980 , y21981 , y21982 , y21983 , y21984 , y21985 , y21986 , y21987 , y21988 , y21989 , y21990 , y21991 , y21992 , y21993 , y21994 , y21995 , y21996 , y21997 , y21998 , y21999 , y22000 , y22001 , y22002 , y22003 , y22004 , y22005 , y22006 , y22007 , y22008 , y22009 , y22010 , y22011 , y22012 , y22013 , y22014 , y22015 , y22016 , y22017 , y22018 , y22019 , y22020 , y22021 , y22022 , y22023 , y22024 , y22025 , y22026 , y22027 , y22028 , y22029 , y22030 , y22031 , y22032 , y22033 , y22034 , y22035 , y22036 , y22037 , y22038 , y22039 , y22040 , y22041 , y22042 , y22043 , y22044 , y22045 , y22046 , y22047 , y22048 , y22049 , y22050 , y22051 , y22052 , y22053 , y22054 , y22055 , y22056 , y22057 , y22058 , y22059 , y22060 , y22061 , y22062 , y22063 , y22064 , y22065 , y22066 , y22067 , y22068 , y22069 , y22070 , y22071 , y22072 , y22073 , y22074 , y22075 , y22076 , y22077 , y22078 , y22079 , y22080 , y22081 , y22082 , y22083 , y22084 , y22085 , y22086 , y22087 , y22088 , y22089 , y22090 , y22091 , y22092 , y22093 , y22094 , y22095 , y22096 , y22097 , y22098 , y22099 , y22100 , y22101 , y22102 , y22103 , y22104 , y22105 , y22106 , y22107 , y22108 , y22109 , y22110 , y22111 , y22112 , y22113 , y22114 , y22115 , y22116 , y22117 , y22118 , y22119 , y22120 , y22121 , y22122 , y22123 , y22124 , y22125 , y22126 , y22127 , y22128 , y22129 , y22130 , y22131 , y22132 , y22133 , y22134 , y22135 , y22136 , y22137 , y22138 , y22139 , y22140 , y22141 , y22142 , y22143 , y22144 , y22145 , y22146 , y22147 , y22148 , y22149 , y22150 , y22151 , y22152 , y22153 , y22154 , y22155 , y22156 , y22157 , y22158 , y22159 , y22160 , y22161 , y22162 , y22163 , y22164 , y22165 , y22166 , y22167 , y22168 , y22169 , y22170 , y22171 , y22172 , y22173 , y22174 , y22175 , y22176 , y22177 , y22178 , y22179 , y22180 , y22181 , y22182 , y22183 , y22184 , y22185 , y22186 , y22187 , y22188 , y22189 , y22190 , y22191 , y22192 , y22193 , y22194 , y22195 , y22196 , y22197 , y22198 , y22199 , y22200 , y22201 , y22202 , y22203 , y22204 , y22205 , y22206 , y22207 , y22208 , y22209 , y22210 , y22211 , y22212 , y22213 , y22214 , y22215 , y22216 , y22217 , y22218 , y22219 , y22220 , y22221 , y22222 , y22223 , y22224 , y22225 , y22226 , y22227 , y22228 , y22229 , y22230 , y22231 , y22232 , y22233 , y22234 , y22235 , y22236 , y22237 , y22238 , y22239 , y22240 , y22241 , y22242 , y22243 , y22244 , y22245 , y22246 , y22247 , y22248 , y22249 , y22250 , y22251 , y22252 , y22253 , y22254 , y22255 , y22256 , y22257 , y22258 , y22259 , y22260 , y22261 , y22262 , y22263 , y22264 , y22265 , y22266 , y22267 , y22268 , y22269 , y22270 , y22271 , y22272 , y22273 , y22274 , y22275 , y22276 , y22277 , y22278 , y22279 , y22280 , y22281 , y22282 , y22283 , y22284 , y22285 , y22286 , y22287 , y22288 , y22289 , y22290 , y22291 , y22292 , y22293 , y22294 , y22295 , y22296 , y22297 , y22298 , y22299 , y22300 , y22301 , y22302 , y22303 , y22304 , y22305 , y22306 , y22307 , y22308 , y22309 , y22310 , y22311 , y22312 , y22313 , y22314 , y22315 , y22316 , y22317 , y22318 , y22319 , y22320 , y22321 , y22322 , y22323 , y22324 , y22325 , y22326 , y22327 , y22328 , y22329 , y22330 , y22331 , y22332 , y22333 , y22334 , y22335 , y22336 , y22337 , y22338 , y22339 , y22340 , y22341 , y22342 , y22343 , y22344 , y22345 , y22346 , y22347 , y22348 , y22349 , y22350 , y22351 , y22352 , y22353 , y22354 , y22355 , y22356 , y22357 , y22358 , y22359 , y22360 , y22361 , y22362 , y22363 , y22364 , y22365 , y22366 , y22367 , y22368 , y22369 , y22370 , y22371 , y22372 , y22373 , y22374 , y22375 , y22376 , y22377 , y22378 , y22379 , y22380 , y22381 , y22382 , y22383 , y22384 , y22385 , y22386 , y22387 , y22388 , y22389 , y22390 , y22391 , y22392 , y22393 , y22394 , y22395 , y22396 , y22397 , y22398 , y22399 , y22400 , y22401 , y22402 , y22403 , y22404 , y22405 , y22406 , y22407 , y22408 , y22409 , y22410 , y22411 , y22412 , y22413 , y22414 , y22415 , y22416 , y22417 , y22418 , y22419 , y22420 , y22421 , y22422 , y22423 , y22424 , y22425 , y22426 , y22427 , y22428 , y22429 , y22430 , y22431 , y22432 , y22433 , y22434 , y22435 , y22436 , y22437 , y22438 , y22439 , y22440 , y22441 , y22442 , y22443 , y22444 , y22445 , y22446 , y22447 , y22448 , y22449 , y22450 , y22451 , y22452 , y22453 , y22454 , y22455 , y22456 , y22457 , y22458 , y22459 , y22460 , y22461 , y22462 , y22463 , y22464 , y22465 , y22466 , y22467 , y22468 , y22469 , y22470 , y22471 , y22472 , y22473 , y22474 , y22475 , y22476 , y22477 , y22478 , y22479 , y22480 , y22481 , y22482 , y22483 , y22484 , y22485 , y22486 , y22487 , y22488 , y22489 , y22490 , y22491 , y22492 , y22493 , y22494 , y22495 , y22496 , y22497 , y22498 , y22499 , y22500 , y22501 , y22502 , y22503 , y22504 , y22505 , y22506 , y22507 , y22508 , y22509 , y22510 , y22511 , y22512 , y22513 , y22514 , y22515 , y22516 , y22517 , y22518 , y22519 , y22520 , y22521 , y22522 , y22523 , y22524 , y22525 , y22526 , y22527 , y22528 , y22529 , y22530 , y22531 , y22532 , y22533 , y22534 , y22535 , y22536 , y22537 , y22538 , y22539 , y22540 , y22541 , y22542 , y22543 , y22544 , y22545 , y22546 , y22547 , y22548 , y22549 , y22550 , y22551 , y22552 , y22553 , y22554 , y22555 , y22556 , y22557 , y22558 , y22559 , y22560 , y22561 , y22562 , y22563 , y22564 , y22565 , y22566 , y22567 , y22568 , y22569 , y22570 , y22571 , y22572 , y22573 , y22574 , y22575 , y22576 , y22577 , y22578 , y22579 , y22580 , y22581 , y22582 , y22583 , y22584 , y22585 , y22586 , y22587 , y22588 , y22589 , y22590 , y22591 , y22592 , y22593 , y22594 , y22595 , y22596 , y22597 , y22598 , y22599 , y22600 , y22601 , y22602 , y22603 , y22604 , y22605 , y22606 , y22607 , y22608 , y22609 , y22610 , y22611 , y22612 , y22613 , y22614 , y22615 , y22616 , y22617 , y22618 , y22619 , y22620 , y22621 , y22622 , y22623 , y22624 , y22625 , y22626 , y22627 , y22628 , y22629 , y22630 , y22631 , y22632 , y22633 , y22634 , y22635 , y22636 , y22637 , y22638 , y22639 , y22640 , y22641 , y22642 , y22643 , y22644 , y22645 , y22646 , y22647 , y22648 , y22649 , y22650 , y22651 , y22652 , y22653 , y22654 , y22655 , y22656 , y22657 , y22658 , y22659 , y22660 , y22661 , y22662 , y22663 , y22664 , y22665 , y22666 , y22667 , y22668 , y22669 , y22670 , y22671 , y22672 , y22673 , y22674 , y22675 , y22676 , y22677 , y22678 , y22679 , y22680 , y22681 , y22682 , y22683 , y22684 , y22685 , y22686 , y22687 , y22688 , y22689 , y22690 , y22691 , y22692 , y22693 , y22694 , y22695 , y22696 , y22697 , y22698 , y22699 , y22700 , y22701 , y22702 , y22703 , y22704 , y22705 , y22706 , y22707 , y22708 , y22709 , y22710 , y22711 , y22712 , y22713 , y22714 , y22715 , y22716 , y22717 , y22718 , y22719 , y22720 , y22721 , y22722 , y22723 , y22724 , y22725 , y22726 , y22727 , y22728 , y22729 , y22730 , y22731 , y22732 , y22733 , y22734 , y22735 , y22736 , y22737 , y22738 , y22739 , y22740 , y22741 , y22742 , y22743 , y22744 , y22745 , y22746 , y22747 , y22748 , y22749 , y22750 , y22751 , y22752 , y22753 , y22754 , y22755 , y22756 , y22757 , y22758 , y22759 , y22760 , y22761 , y22762 , y22763 , y22764 , y22765 , y22766 , y22767 , y22768 , y22769 , y22770 , y22771 , y22772 , y22773 , y22774 , y22775 , y22776 , y22777 , y22778 , y22779 , y22780 , y22781 , y22782 , y22783 , y22784 , y22785 , y22786 , y22787 , y22788 , y22789 , y22790 , y22791 , y22792 , y22793 , y22794 , y22795 , y22796 , y22797 , y22798 , y22799 , y22800 , y22801 , y22802 , y22803 , y22804 , y22805 , y22806 , y22807 , y22808 , y22809 , y22810 , y22811 , y22812 , y22813 , y22814 , y22815 , y22816 , y22817 , y22818 , y22819 , y22820 , y22821 , y22822 , y22823 , y22824 , y22825 , y22826 , y22827 , y22828 , y22829 , y22830 , y22831 , y22832 , y22833 , y22834 , y22835 , y22836 , y22837 , y22838 , y22839 , y22840 , y22841 , y22842 , y22843 , y22844 , y22845 , y22846 , y22847 , y22848 , y22849 , y22850 , y22851 , y22852 , y22853 , y22854 , y22855 , y22856 , y22857 , y22858 , y22859 , y22860 , y22861 , y22862 , y22863 , y22864 , y22865 , y22866 , y22867 , y22868 , y22869 , y22870 , y22871 , y22872 , y22873 , y22874 , y22875 , y22876 , y22877 , y22878 , y22879 , y22880 , y22881 , y22882 , y22883 , y22884 , y22885 , y22886 , y22887 , y22888 , y22889 , y22890 , y22891 , y22892 , y22893 , y22894 , y22895 , y22896 , y22897 , y22898 , y22899 , y22900 , y22901 , y22902 , y22903 , y22904 , y22905 , y22906 , y22907 , y22908 , y22909 , y22910 , y22911 , y22912 , y22913 , y22914 , y22915 , y22916 , y22917 , y22918 , y22919 , y22920 , y22921 , y22922 , y22923 , y22924 , y22925 , y22926 , y22927 , y22928 , y22929 , y22930 , y22931 , y22932 , y22933 , y22934 , y22935 , y22936 , y22937 , y22938 , y22939 , y22940 , y22941 , y22942 , y22943 , y22944 , y22945 , y22946 , y22947 , y22948 , y22949 , y22950 , y22951 , y22952 , y22953 , y22954 , y22955 , y22956 , y22957 , y22958 , y22959 , y22960 , y22961 , y22962 , y22963 , y22964 , y22965 , y22966 , y22967 , y22968 , y22969 , y22970 , y22971 , y22972 , y22973 , y22974 , y22975 , y22976 , y22977 , y22978 , y22979 , y22980 , y22981 , y22982 , y22983 , y22984 , y22985 , y22986 , y22987 , y22988 , y22989 , y22990 , y22991 , y22992 , y22993 , y22994 , y22995 , y22996 , y22997 , y22998 , y22999 , y23000 , y23001 , y23002 , y23003 , y23004 , y23005 , y23006 , y23007 , y23008 , y23009 , y23010 , y23011 , y23012 , y23013 , y23014 , y23015 , y23016 , y23017 , y23018 , y23019 , y23020 , y23021 , y23022 , y23023 , y23024 , y23025 , y23026 , y23027 , y23028 , y23029 , y23030 , y23031 , y23032 , y23033 , y23034 , y23035 , y23036 , y23037 , y23038 , y23039 , y23040 , y23041 , y23042 , y23043 , y23044 , y23045 , y23046 , y23047 , y23048 , y23049 , y23050 , y23051 , y23052 , y23053 , y23054 , y23055 , y23056 , y23057 , y23058 , y23059 , y23060 , y23061 , y23062 , y23063 , y23064 , y23065 , y23066 , y23067 , y23068 , y23069 , y23070 , y23071 , y23072 , y23073 , y23074 , y23075 , y23076 , y23077 , y23078 , y23079 , y23080 , y23081 , y23082 , y23083 , y23084 , y23085 , y23086 , y23087 , y23088 , y23089 , y23090 , y23091 , y23092 , y23093 , y23094 , y23095 , y23096 , y23097 , y23098 , y23099 , y23100 , y23101 , y23102 , y23103 , y23104 , y23105 , y23106 , y23107 , y23108 , y23109 , y23110 , y23111 , y23112 , y23113 , y23114 , y23115 , y23116 , y23117 , y23118 , y23119 , y23120 , y23121 , y23122 , y23123 , y23124 , y23125 , y23126 , y23127 , y23128 , y23129 , y23130 , y23131 , y23132 , y23133 , y23134 , y23135 , y23136 , y23137 , y23138 , y23139 , y23140 , y23141 , y23142 , y23143 , y23144 , y23145 , y23146 , y23147 , y23148 , y23149 , y23150 , y23151 , y23152 , y23153 , y23154 , y23155 , y23156 , y23157 , y23158 , y23159 , y23160 , y23161 , y23162 , y23163 , y23164 , y23165 , y23166 , y23167 , y23168 , y23169 , y23170 , y23171 , y23172 , y23173 , y23174 , y23175 , y23176 , y23177 , y23178 , y23179 , y23180 , y23181 , y23182 , y23183 , y23184 , y23185 , y23186 , y23187 , y23188 , y23189 , y23190 , y23191 , y23192 , y23193 , y23194 , y23195 , y23196 , y23197 , y23198 , y23199 , y23200 , y23201 , y23202 , y23203 , y23204 , y23205 , y23206 , y23207 , y23208 , y23209 , y23210 , y23211 , y23212 , y23213 , y23214 , y23215 , y23216 , y23217 , y23218 , y23219 , y23220 , y23221 , y23222 , y23223 , y23224 , y23225 , y23226 , y23227 , y23228 , y23229 , y23230 , y23231 , y23232 , y23233 , y23234 , y23235 , y23236 , y23237 , y23238 , y23239 , y23240 , y23241 , y23242 , y23243 , y23244 , y23245 , y23246 , y23247 , y23248 , y23249 , y23250 , y23251 , y23252 , y23253 , y23254 , y23255 , y23256 , y23257 , y23258 , y23259 , y23260 , y23261 , y23262 , y23263 , y23264 , y23265 , y23266 , y23267 , y23268 , y23269 , y23270 , y23271 , y23272 , y23273 , y23274 , y23275 , y23276 , y23277 , y23278 , y23279 , y23280 , y23281 , y23282 , y23283 , y23284 , y23285 , y23286 , y23287 , y23288 , y23289 , y23290 , y23291 , y23292 , y23293 , y23294 , y23295 , y23296 , y23297 , y23298 , y23299 , y23300 , y23301 , y23302 , y23303 , y23304 , y23305 , y23306 , y23307 , y23308 , y23309 , y23310 , y23311 , y23312 , y23313 , y23314 , y23315 , y23316 , y23317 , y23318 , y23319 , y23320 , y23321 , y23322 , y23323 , y23324 , y23325 , y23326 , y23327 , y23328 , y23329 , y23330 , y23331 , y23332 , y23333 , y23334 , y23335 , y23336 , y23337 , y23338 , y23339 , y23340 , y23341 , y23342 , y23343 , y23344 , y23345 , y23346 , y23347 , y23348 , y23349 , y23350 , y23351 , y23352 , y23353 , y23354 , y23355 , y23356 , y23357 , y23358 , y23359 , y23360 , y23361 , y23362 , y23363 , y23364 , y23365 , y23366 , y23367 , y23368 , y23369 , y23370 , y23371 , y23372 , y23373 , y23374 , y23375 , y23376 , y23377 , y23378 , y23379 , y23380 , y23381 , y23382 , y23383 , y23384 , y23385 , y23386 , y23387 , y23388 , y23389 , y23390 , y23391 , y23392 , y23393 , y23394 , y23395 , y23396 , y23397 , y23398 , y23399 , y23400 , y23401 , y23402 , y23403 , y23404 , y23405 , y23406 , y23407 , y23408 , y23409 , y23410 , y23411 , y23412 , y23413 , y23414 , y23415 , y23416 , y23417 , y23418 , y23419 , y23420 , y23421 , y23422 , y23423 , y23424 , y23425 , y23426 , y23427 , y23428 , y23429 , y23430 , y23431 , y23432 , y23433 , y23434 , y23435 , y23436 , y23437 , y23438 , y23439 , y23440 , y23441 , y23442 , y23443 , y23444 , y23445 , y23446 , y23447 , y23448 , y23449 , y23450 , y23451 , y23452 , y23453 , y23454 , y23455 , y23456 , y23457 , y23458 , y23459 , y23460 , y23461 , y23462 , y23463 , y23464 , y23465 , y23466 , y23467 , y23468 , y23469 , y23470 , y23471 , y23472 , y23473 , y23474 , y23475 , y23476 , y23477 , y23478 , y23479 , y23480 , y23481 , y23482 , y23483 , y23484 , y23485 , y23486 , y23487 , y23488 , y23489 , y23490 , y23491 , y23492 , y23493 , y23494 , y23495 , y23496 , y23497 , y23498 , y23499 , y23500 , y23501 , y23502 , y23503 , y23504 , y23505 , y23506 , y23507 , y23508 , y23509 , y23510 , y23511 , y23512 , y23513 , y23514 , y23515 , y23516 , y23517 , y23518 , y23519 , y23520 , y23521 , y23522 , y23523 , y23524 , y23525 , y23526 , y23527 , y23528 , y23529 , y23530 , y23531 , y23532 , y23533 , y23534 , y23535 , y23536 , y23537 , y23538 , y23539 , y23540 , y23541 , y23542 , y23543 , y23544 , y23545 , y23546 , y23547 , y23548 , y23549 , y23550 , y23551 , y23552 , y23553 , y23554 , y23555 , y23556 , y23557 , y23558 , y23559 , y23560 , y23561 , y23562 , y23563 , y23564 , y23565 , y23566 , y23567 , y23568 , y23569 , y23570 , y23571 , y23572 , y23573 , y23574 , y23575 , y23576 , y23577 , y23578 , y23579 , y23580 , y23581 , y23582 , y23583 , y23584 , y23585 , y23586 , y23587 , y23588 , y23589 , y23590 , y23591 , y23592 , y23593 , y23594 , y23595 , y23596 , y23597 , y23598 , y23599 , y23600 , y23601 , y23602 , y23603 , y23604 , y23605 , y23606 , y23607 , y23608 , y23609 , y23610 , y23611 , y23612 , y23613 , y23614 , y23615 , y23616 , y23617 , y23618 , y23619 , y23620 , y23621 , y23622 , y23623 , y23624 , y23625 , y23626 , y23627 , y23628 , y23629 , y23630 , y23631 , y23632 , y23633 , y23634 , y23635 , y23636 , y23637 , y23638 , y23639 , y23640 , y23641 , y23642 , y23643 , y23644 , y23645 , y23646 , y23647 , y23648 , y23649 , y23650 , y23651 , y23652 , y23653 , y23654 , y23655 , y23656 , y23657 , y23658 , y23659 , y23660 , y23661 , y23662 , y23663 , y23664 , y23665 , y23666 , y23667 , y23668 , y23669 , y23670 , y23671 , y23672 , y23673 , y23674 , y23675 , y23676 , y23677 , y23678 , y23679 , y23680 , y23681 , y23682 , y23683 , y23684 , y23685 , y23686 , y23687 , y23688 , y23689 , y23690 , y23691 , y23692 , y23693 , y23694 , y23695 , y23696 , y23697 , y23698 , y23699 , y23700 , y23701 , y23702 , y23703 , y23704 , y23705 , y23706 , y23707 , y23708 , y23709 , y23710 , y23711 , y23712 , y23713 , y23714 , y23715 , y23716 , y23717 , y23718 , y23719 , y23720 , y23721 , y23722 , y23723 , y23724 , y23725 , y23726 , y23727 , y23728 , y23729 , y23730 , y23731 , y23732 , y23733 , y23734 , y23735 , y23736 , y23737 , y23738 , y23739 , y23740 , y23741 , y23742 , y23743 , y23744 , y23745 , y23746 , y23747 , y23748 , y23749 , y23750 , y23751 , y23752 , y23753 , y23754 , y23755 , y23756 , y23757 , y23758 , y23759 , y23760 , y23761 , y23762 , y23763 , y23764 , y23765 , y23766 , y23767 , y23768 , y23769 , y23770 , y23771 , y23772 , y23773 , y23774 , y23775 , y23776 , y23777 , y23778 , y23779 , y23780 , y23781 , y23782 , y23783 , y23784 , y23785 , y23786 , y23787 , y23788 , y23789 , y23790 , y23791 , y23792 , y23793 , y23794 , y23795 , y23796 , y23797 , y23798 , y23799 , y23800 , y23801 , y23802 , y23803 , y23804 , y23805 ;
  wire n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 ;
  assign n256 = x244 ^ x238 ^ x38 ;
  assign n257 = x186 & x227 ;
  assign n258 = ~x62 & n257 ;
  assign n259 = x211 ^ x191 ^ 1'b0 ;
  assign n260 = x221 & n259 ;
  assign n261 = n256 ^ x188 ^ 1'b0 ;
  assign n262 = x192 & ~n261 ;
  assign n263 = x221 ^ x112 ^ 1'b0 ;
  assign n264 = x169 ^ x132 ^ x44 ;
  assign n265 = n264 ^ n256 ^ 1'b0 ;
  assign n266 = x55 & n265 ;
  assign n267 = x82 & ~x205 ;
  assign n268 = x152 & x175 ;
  assign n269 = x58 & x64 ;
  assign n270 = ~x15 & n269 ;
  assign n271 = ( ~x42 & x184 ) | ( ~x42 & x229 ) | ( x184 & x229 ) ;
  assign n272 = x113 ^ x79 ^ 1'b0 ;
  assign n273 = x134 & x187 ;
  assign n274 = n273 ^ x246 ^ 1'b0 ;
  assign n275 = x3 & x151 ;
  assign n276 = ~x199 & n275 ;
  assign n277 = x133 & n276 ;
  assign n278 = x159 ^ x0 ^ 1'b0 ;
  assign n279 = x206 & n278 ;
  assign n280 = x76 & x210 ;
  assign n281 = ~x189 & n280 ;
  assign n282 = x78 & x180 ;
  assign n283 = n282 ^ n281 ^ 1'b0 ;
  assign n284 = x127 & x193 ;
  assign n285 = ~x201 & n284 ;
  assign n286 = x195 & x250 ;
  assign n287 = ~x169 & n286 ;
  assign n288 = n285 | n287 ;
  assign n289 = x96 | n288 ;
  assign n290 = x58 & x143 ;
  assign n291 = n290 ^ x83 ^ 1'b0 ;
  assign n292 = x81 ^ x58 ^ 1'b0 ;
  assign n293 = x34 & n292 ;
  assign n294 = ( x20 & x159 ) | ( x20 & ~n293 ) | ( x159 & ~n293 ) ;
  assign n295 = x198 & x221 ;
  assign n296 = n295 ^ x162 ^ 1'b0 ;
  assign n297 = x37 & x93 ;
  assign n298 = n297 ^ x90 ^ 1'b0 ;
  assign n299 = x38 & x142 ;
  assign n300 = n299 ^ x163 ^ 1'b0 ;
  assign n301 = n300 ^ x205 ^ 1'b0 ;
  assign n302 = x88 & ~n301 ;
  assign n304 = n266 ^ x164 ^ 1'b0 ;
  assign n305 = x44 & n304 ;
  assign n303 = x58 & x188 ;
  assign n306 = n305 ^ n303 ^ 1'b0 ;
  assign n307 = x118 & x144 ;
  assign n308 = ~x200 & n307 ;
  assign n309 = ( ~x90 & x190 ) | ( ~x90 & n308 ) | ( x190 & n308 ) ;
  assign n310 = n309 ^ x69 ^ x32 ;
  assign n311 = x18 & x130 ;
  assign n312 = ~x93 & n311 ;
  assign n313 = x45 & n260 ;
  assign n314 = n313 ^ x17 ^ 1'b0 ;
  assign n315 = ( x72 & ~x105 ) | ( x72 & n281 ) | ( ~x105 & n281 ) ;
  assign n316 = x131 & x140 ;
  assign n317 = ~n283 & n316 ;
  assign n318 = ( x55 & x82 ) | ( x55 & ~x240 ) | ( x82 & ~x240 ) ;
  assign n319 = x1 & n318 ;
  assign n320 = n319 ^ x240 ^ 1'b0 ;
  assign n326 = x86 & n305 ;
  assign n327 = n326 ^ x248 ^ 1'b0 ;
  assign n325 = ( ~x80 & x113 ) | ( ~x80 & x204 ) | ( x113 & x204 ) ;
  assign n328 = n327 ^ n325 ^ 1'b0 ;
  assign n321 = x146 & x213 ;
  assign n322 = n321 ^ n272 ^ 1'b0 ;
  assign n323 = ( x126 & x190 ) | ( x126 & n322 ) | ( x190 & n322 ) ;
  assign n324 = x9 & n323 ;
  assign n329 = n328 ^ n324 ^ 1'b0 ;
  assign n330 = x235 & ~n300 ;
  assign n331 = n330 ^ x241 ^ 1'b0 ;
  assign n332 = ( x161 & ~n263 ) | ( x161 & n331 ) | ( ~n263 & n331 ) ;
  assign n333 = x232 ^ x213 ^ x199 ;
  assign n334 = n333 ^ x169 ^ 1'b0 ;
  assign n335 = n305 ^ x224 ^ x120 ;
  assign n336 = n335 ^ x162 ^ x100 ;
  assign n337 = x32 & x107 ;
  assign n338 = n337 ^ x39 ^ 1'b0 ;
  assign n339 = x205 & x206 ;
  assign n340 = ~x71 & n339 ;
  assign n341 = x83 & x138 ;
  assign n342 = n341 ^ x64 ^ 1'b0 ;
  assign n343 = x178 & ~n342 ;
  assign n344 = n343 ^ x74 ^ 1'b0 ;
  assign n345 = x33 & x58 ;
  assign n346 = ~x101 & n345 ;
  assign n347 = n274 | n306 ;
  assign n348 = n346 | n347 ;
  assign n349 = x220 ^ x151 ^ x0 ;
  assign n350 = x134 ^ x104 ^ 1'b0 ;
  assign n351 = x97 & n350 ;
  assign n352 = x228 ^ x92 ^ 1'b0 ;
  assign n353 = x121 & n352 ;
  assign n354 = n353 ^ n276 ^ 1'b0 ;
  assign n355 = x35 & ~n354 ;
  assign n356 = x253 ^ x165 ^ 1'b0 ;
  assign n357 = x121 & n356 ;
  assign n358 = n357 ^ n260 ^ 1'b0 ;
  assign n359 = ~n277 & n358 ;
  assign n360 = x41 & x155 ;
  assign n361 = ~x217 & n360 ;
  assign n362 = x167 & n266 ;
  assign n363 = n362 ^ x138 ^ 1'b0 ;
  assign n364 = n363 ^ n271 ^ 1'b0 ;
  assign n365 = x222 ^ x121 ^ x23 ;
  assign n366 = ( x126 & x206 ) | ( x126 & n365 ) | ( x206 & n365 ) ;
  assign n367 = x184 ^ x148 ^ 1'b0 ;
  assign n368 = x18 & x197 ;
  assign n369 = n368 ^ x186 ^ 1'b0 ;
  assign n370 = x250 ^ x203 ^ x78 ;
  assign n371 = x66 & n266 ;
  assign n372 = n371 ^ x14 ^ 1'b0 ;
  assign n373 = x20 & x132 ;
  assign n374 = ~x166 & n373 ;
  assign n375 = x117 | n374 ;
  assign n376 = n372 | n375 ;
  assign n377 = x211 ^ x47 ^ 1'b0 ;
  assign n378 = x173 & n377 ;
  assign n379 = x146 ^ x104 ^ 1'b0 ;
  assign n380 = x40 & n379 ;
  assign n381 = x91 & ~n327 ;
  assign n382 = n381 ^ x1 ^ 1'b0 ;
  assign n383 = n380 & ~n382 ;
  assign n384 = ~x115 & n383 ;
  assign n385 = n384 ^ n266 ^ x178 ;
  assign n386 = n277 ^ x201 ^ 1'b0 ;
  assign n387 = n385 & ~n386 ;
  assign n388 = x187 & n263 ;
  assign n389 = n388 ^ n310 ^ 1'b0 ;
  assign n390 = x246 ^ x160 ^ 1'b0 ;
  assign n391 = x149 & n390 ;
  assign n393 = n256 ^ x73 ^ 1'b0 ;
  assign n392 = x220 & ~n296 ;
  assign n394 = n393 ^ n392 ^ 1'b0 ;
  assign n395 = n391 & n394 ;
  assign n396 = x56 & x171 ;
  assign n397 = ~x181 & n396 ;
  assign n398 = n308 ^ x174 ^ 1'b0 ;
  assign n399 = n335 | n398 ;
  assign n400 = ( x46 & ~x130 ) | ( x46 & x171 ) | ( ~x130 & x171 ) ;
  assign n401 = n400 ^ x69 ^ 1'b0 ;
  assign n402 = ~n327 & n401 ;
  assign n403 = n402 ^ x241 ^ 1'b0 ;
  assign n404 = x241 & n403 ;
  assign n405 = n404 ^ x61 ^ 1'b0 ;
  assign n406 = x203 & n405 ;
  assign n407 = n394 ^ x172 ^ 1'b0 ;
  assign n408 = x155 ^ x67 ^ 1'b0 ;
  assign n409 = n407 & n408 ;
  assign n410 = x49 & x69 ;
  assign n411 = ~x130 & n410 ;
  assign n412 = x46 & x188 ;
  assign n413 = ~x116 & n412 ;
  assign n414 = n370 | n413 ;
  assign n415 = n380 | n414 ;
  assign n416 = n325 ^ x22 ^ 1'b0 ;
  assign n417 = ~x71 & n416 ;
  assign n418 = x5 & x225 ;
  assign n419 = ~x121 & n418 ;
  assign n420 = ~x146 & x222 ;
  assign n421 = x145 & ~x206 ;
  assign n422 = n415 & n421 ;
  assign n423 = n422 ^ x92 ^ 1'b0 ;
  assign n424 = ( x80 & ~x109 ) | ( x80 & x207 ) | ( ~x109 & x207 ) ;
  assign n425 = n277 ^ x224 ^ x65 ;
  assign n426 = ( x67 & n296 ) | ( x67 & ~n425 ) | ( n296 & ~n425 ) ;
  assign n427 = x19 & x156 ;
  assign n428 = n427 ^ n300 ^ 1'b0 ;
  assign n429 = n385 & n428 ;
  assign n430 = ~x214 & n429 ;
  assign n431 = n430 ^ x176 ^ 1'b0 ;
  assign n432 = x105 ^ x11 ^ 1'b0 ;
  assign n433 = n432 ^ n425 ^ 1'b0 ;
  assign n434 = x25 & x161 ;
  assign n435 = n434 ^ x61 ^ 1'b0 ;
  assign n436 = x111 & n435 ;
  assign n437 = n436 ^ n402 ^ x196 ;
  assign n439 = x74 & x84 ;
  assign n440 = ~x163 & n439 ;
  assign n441 = x29 & ~n440 ;
  assign n442 = ~x192 & n441 ;
  assign n443 = x154 & ~n442 ;
  assign n444 = n315 & n443 ;
  assign n438 = x104 & x239 ;
  assign n445 = n444 ^ n438 ^ 1'b0 ;
  assign n446 = x238 ^ x9 ^ 1'b0 ;
  assign n448 = x246 ^ x195 ^ x181 ;
  assign n447 = x119 & n400 ;
  assign n449 = n448 ^ n447 ^ 1'b0 ;
  assign n450 = x41 & ~x96 ;
  assign n451 = n450 ^ x199 ^ 1'b0 ;
  assign n452 = x30 & n451 ;
  assign n453 = n452 ^ n312 ^ 1'b0 ;
  assign n456 = x56 & x217 ;
  assign n457 = n456 ^ x98 ^ 1'b0 ;
  assign n454 = x181 & ~n440 ;
  assign n455 = ~x238 & n454 ;
  assign n458 = n457 ^ n455 ^ n306 ;
  assign n459 = n458 ^ x184 ^ 1'b0 ;
  assign n460 = x42 & x217 ;
  assign n461 = n460 ^ n387 ^ 1'b0 ;
  assign n462 = x143 & n256 ;
  assign n463 = x54 & ~n462 ;
  assign n464 = n463 ^ x71 ^ 1'b0 ;
  assign n465 = x66 & x166 ;
  assign n466 = ~x188 & n465 ;
  assign n467 = ~n464 & n466 ;
  assign n468 = x220 & n467 ;
  assign n469 = n344 & n468 ;
  assign n470 = n270 ^ x20 ^ 1'b0 ;
  assign n471 = x121 & ~n470 ;
  assign n472 = x137 & n471 ;
  assign n473 = n472 ^ x217 ^ 1'b0 ;
  assign n474 = x228 & ~n473 ;
  assign n475 = ~x118 & n474 ;
  assign n476 = n267 ^ x21 ^ 1'b0 ;
  assign n477 = x110 & ~n476 ;
  assign n478 = x222 & x232 ;
  assign n479 = ~x138 & n478 ;
  assign n480 = x134 & ~n479 ;
  assign n481 = ~x52 & n480 ;
  assign n482 = n477 & ~n481 ;
  assign n483 = n482 ^ x85 ^ 1'b0 ;
  assign n484 = x206 & ~n440 ;
  assign n485 = n484 ^ x216 ^ 1'b0 ;
  assign n486 = x142 & n485 ;
  assign n487 = n276 ^ x209 ^ 1'b0 ;
  assign n488 = x121 & ~n487 ;
  assign n489 = ~n320 & n488 ;
  assign n490 = ~n486 & n489 ;
  assign n491 = x117 & n479 ;
  assign n492 = x130 & ~x158 ;
  assign n493 = x86 & n492 ;
  assign n494 = n493 ^ x233 ^ 1'b0 ;
  assign n499 = x198 & ~n457 ;
  assign n500 = n499 ^ x173 ^ 1'b0 ;
  assign n501 = x19 & n382 ;
  assign n502 = n501 ^ x190 ^ 1'b0 ;
  assign n503 = ~n500 & n502 ;
  assign n496 = n294 & ~n416 ;
  assign n495 = x91 & x104 ;
  assign n497 = n496 ^ n495 ^ 1'b0 ;
  assign n498 = ( n271 & n300 ) | ( n271 & n497 ) | ( n300 & n497 ) ;
  assign n504 = n503 ^ n498 ^ 1'b0 ;
  assign n505 = n483 | n504 ;
  assign n506 = x178 & x195 ;
  assign n507 = ~x20 & n506 ;
  assign n508 = x0 & x3 ;
  assign n509 = n508 ^ x254 ^ 1'b0 ;
  assign n510 = ~n507 & n509 ;
  assign n511 = x243 ^ x88 ^ x20 ;
  assign n512 = x172 & ~n267 ;
  assign n513 = n512 ^ x45 ^ 1'b0 ;
  assign n514 = n513 ^ n430 ^ 1'b0 ;
  assign n515 = x62 & x125 ;
  assign n516 = ~x155 & n515 ;
  assign n517 = x192 & ~n516 ;
  assign n518 = ~n328 & n517 ;
  assign n519 = n518 ^ x108 ^ 1'b0 ;
  assign n520 = n346 | n519 ;
  assign n521 = x1 & ~n256 ;
  assign n522 = ~n323 & n521 ;
  assign n523 = n306 ^ n268 ^ x3 ;
  assign n524 = x250 ^ x208 ^ 1'b0 ;
  assign n525 = x15 & n524 ;
  assign n526 = x54 & x174 ;
  assign n527 = ~n525 & n526 ;
  assign n528 = n527 ^ x90 ^ 1'b0 ;
  assign n529 = x2 & ~n528 ;
  assign n530 = n527 | n529 ;
  assign n531 = x82 ^ x78 ^ 1'b0 ;
  assign n532 = x254 & n531 ;
  assign n533 = n532 ^ n451 ^ 1'b0 ;
  assign n534 = x45 & n533 ;
  assign n535 = x118 & ~n294 ;
  assign n536 = x38 & x175 ;
  assign n537 = n536 ^ n264 ^ 1'b0 ;
  assign n538 = x231 & ~n309 ;
  assign n539 = n538 ^ x14 ^ 1'b0 ;
  assign n540 = ( ~x38 & x119 ) | ( ~x38 & x135 ) | ( x119 & x135 ) ;
  assign n541 = x33 & n540 ;
  assign n542 = n320 & n541 ;
  assign n543 = x169 & ~n542 ;
  assign n544 = n543 ^ x4 ^ 1'b0 ;
  assign n545 = ~n539 & n544 ;
  assign n546 = n353 ^ x137 ^ 1'b0 ;
  assign n547 = n433 & n546 ;
  assign n548 = n518 ^ n488 ^ 1'b0 ;
  assign n549 = x106 & x181 ;
  assign n550 = ~x173 & n549 ;
  assign n551 = x153 & ~n455 ;
  assign n552 = n550 & n551 ;
  assign n553 = x229 ^ x70 ^ 1'b0 ;
  assign n554 = x84 & n553 ;
  assign n555 = n291 & n554 ;
  assign n556 = x140 ^ x30 ^ 1'b0 ;
  assign n557 = n556 ^ n464 ^ 1'b0 ;
  assign n558 = x213 & ~n557 ;
  assign n559 = x4 & x95 ;
  assign n560 = ~x180 & n559 ;
  assign n561 = n402 ^ x36 ^ 1'b0 ;
  assign n562 = x195 & n561 ;
  assign n563 = ~n560 & n562 ;
  assign n564 = n563 ^ x153 ^ 1'b0 ;
  assign n565 = n357 ^ x115 ^ 1'b0 ;
  assign n566 = x59 & n565 ;
  assign n567 = n566 ^ x194 ^ x153 ;
  assign n568 = n567 ^ x154 ^ 1'b0 ;
  assign n569 = x211 & ~n568 ;
  assign n570 = x10 & n387 ;
  assign n571 = ~n569 & n570 ;
  assign n572 = x85 & ~n571 ;
  assign n573 = x82 & x164 ;
  assign n574 = n296 & n573 ;
  assign n575 = x173 ^ x127 ^ 1'b0 ;
  assign n576 = ~n555 & n575 ;
  assign n577 = n384 & n576 ;
  assign n578 = x35 ^ x12 ^ 1'b0 ;
  assign n579 = x190 & n578 ;
  assign n580 = ( x86 & n333 ) | ( x86 & n579 ) | ( n333 & n579 ) ;
  assign n581 = x225 | n411 ;
  assign n582 = ~n382 & n581 ;
  assign n583 = n582 ^ x133 ^ 1'b0 ;
  assign n584 = x79 & n503 ;
  assign n585 = ~x167 & n584 ;
  assign n586 = n369 | n585 ;
  assign n587 = n583 & ~n586 ;
  assign n588 = x4 & x8 ;
  assign n589 = n588 ^ x135 ^ 1'b0 ;
  assign n590 = x71 ^ x43 ^ 1'b0 ;
  assign n591 = x152 & n590 ;
  assign n592 = x253 & n591 ;
  assign n594 = x210 & ~n317 ;
  assign n595 = n370 & n594 ;
  assign n593 = ( x80 & x149 ) | ( x80 & n327 ) | ( x149 & n327 ) ;
  assign n596 = n595 ^ n593 ^ 1'b0 ;
  assign n597 = ( x98 & ~x193 ) | ( x98 & n433 ) | ( ~x193 & n433 ) ;
  assign n600 = x178 & x196 ;
  assign n601 = ~x118 & n600 ;
  assign n602 = x163 & ~n601 ;
  assign n603 = n602 ^ n260 ^ 1'b0 ;
  assign n598 = x114 & x168 ;
  assign n599 = ~x230 & n598 ;
  assign n604 = n603 ^ n599 ^ 1'b0 ;
  assign n605 = x173 & x218 ;
  assign n606 = ~n604 & n605 ;
  assign n610 = x58 & ~n327 ;
  assign n611 = n610 ^ x194 ^ 1'b0 ;
  assign n612 = n611 ^ x78 ^ 1'b0 ;
  assign n613 = n310 & ~n612 ;
  assign n607 = x46 & x62 ;
  assign n608 = n607 ^ x112 ^ 1'b0 ;
  assign n609 = n283 & ~n608 ;
  assign n614 = n613 ^ n609 ^ 1'b0 ;
  assign n615 = n289 ^ x91 ^ x34 ;
  assign n616 = n615 ^ x73 ^ 1'b0 ;
  assign n617 = n492 & ~n616 ;
  assign n618 = ~n614 & n617 ;
  assign n621 = ( ~x97 & x123 ) | ( ~x97 & n351 ) | ( x123 & n351 ) ;
  assign n619 = ~x159 & n451 ;
  assign n620 = x120 & ~n619 ;
  assign n622 = n621 ^ n620 ^ 1'b0 ;
  assign n623 = x75 & x212 ;
  assign n624 = ~x76 & n623 ;
  assign n625 = ( ~x73 & n293 ) | ( ~x73 & n415 ) | ( n293 & n415 ) ;
  assign n626 = x190 & x243 ;
  assign n627 = n626 ^ n597 ^ 1'b0 ;
  assign n628 = x212 | n507 ;
  assign n629 = n440 & n628 ;
  assign n632 = n436 ^ n347 ^ x196 ;
  assign n630 = x13 & x29 ;
  assign n631 = n630 ^ n615 ^ 1'b0 ;
  assign n633 = n632 ^ n631 ^ 1'b0 ;
  assign n634 = ~n629 & n633 ;
  assign n635 = n424 & ~n540 ;
  assign n636 = ~n348 & n366 ;
  assign n637 = n635 & n636 ;
  assign n638 = ~x9 & n400 ;
  assign n639 = x118 & x191 ;
  assign n640 = n639 ^ n428 ^ 1'b0 ;
  assign n641 = x0 & ~n640 ;
  assign n642 = ~x95 & n641 ;
  assign n643 = n642 ^ n614 ^ n424 ;
  assign n644 = x20 & x254 ;
  assign n645 = n644 ^ x187 ^ 1'b0 ;
  assign n646 = n488 ^ x24 ^ 1'b0 ;
  assign n647 = ~n442 & n646 ;
  assign n648 = n539 ^ x132 ^ 1'b0 ;
  assign n649 = x114 & ~n648 ;
  assign n650 = n613 & n649 ;
  assign n651 = ~n647 & n650 ;
  assign n652 = n349 | n507 ;
  assign n653 = n444 & ~n652 ;
  assign n654 = n589 | n653 ;
  assign n655 = n315 & ~n654 ;
  assign n656 = x134 & x212 ;
  assign n657 = ~x168 & n656 ;
  assign n658 = n657 ^ n497 ^ 1'b0 ;
  assign n659 = x125 & n658 ;
  assign n660 = ~n419 & n632 ;
  assign n661 = n660 ^ x157 ^ 1'b0 ;
  assign n662 = n338 | n661 ;
  assign n663 = x120 | n662 ;
  assign n664 = x246 & ~n426 ;
  assign n665 = n611 & n664 ;
  assign n666 = ( x109 & x237 ) | ( x109 & n665 ) | ( x237 & n665 ) ;
  assign n667 = x171 & n260 ;
  assign n668 = ~n477 & n667 ;
  assign n670 = x102 ^ x21 ^ 1'b0 ;
  assign n671 = x87 & n670 ;
  assign n669 = x13 & x246 ;
  assign n672 = n671 ^ n669 ^ 1'b0 ;
  assign n673 = ~n589 & n672 ;
  assign n674 = x41 & x138 ;
  assign n675 = n674 ^ x99 ^ 1'b0 ;
  assign n676 = x213 & ~n333 ;
  assign n677 = n676 ^ n653 ^ 1'b0 ;
  assign n678 = n677 ^ n380 ^ 1'b0 ;
  assign n679 = n675 | n678 ;
  assign n680 = ( x92 & x231 ) | ( x92 & n450 ) | ( x231 & n450 ) ;
  assign n690 = ~n298 & n318 ;
  assign n691 = n690 ^ n268 ^ 1'b0 ;
  assign n692 = n442 ^ n320 ^ 1'b0 ;
  assign n693 = n692 ^ x239 ^ 1'b0 ;
  assign n694 = n466 | n693 ;
  assign n695 = n694 ^ n272 ^ 1'b0 ;
  assign n696 = x241 & ~n300 ;
  assign n697 = ~x92 & n696 ;
  assign n698 = x60 & ~n697 ;
  assign n699 = n695 & n698 ;
  assign n700 = n691 | n699 ;
  assign n701 = x208 | n700 ;
  assign n681 = x76 & x168 ;
  assign n682 = n681 ^ n271 ^ 1'b0 ;
  assign n683 = x10 & x94 ;
  assign n684 = ~x228 & n683 ;
  assign n685 = n391 & ~n684 ;
  assign n686 = n685 ^ n448 ^ 1'b0 ;
  assign n687 = n498 ^ n323 ^ 1'b0 ;
  assign n688 = n686 & ~n687 ;
  assign n689 = ~n682 & n688 ;
  assign n702 = n701 ^ n689 ^ 1'b0 ;
  assign n703 = n680 & n702 ;
  assign n704 = x243 & ~n661 ;
  assign n705 = n704 ^ x236 ^ 1'b0 ;
  assign n706 = n264 ^ x193 ^ 1'b0 ;
  assign n707 = x41 & ~n706 ;
  assign n708 = n407 ^ n365 ^ x44 ;
  assign n709 = ~x18 & n708 ;
  assign n710 = ( x249 & n413 ) | ( x249 & n475 ) | ( n413 & n475 ) ;
  assign n711 = x213 ^ x144 ^ x107 ;
  assign n712 = n569 ^ x91 ^ 1'b0 ;
  assign n713 = ~n711 & n712 ;
  assign n714 = x9 & ~n707 ;
  assign n715 = x56 & n380 ;
  assign n716 = ~x13 & n715 ;
  assign n717 = n716 ^ x173 ^ 1'b0 ;
  assign n718 = x131 & ~n717 ;
  assign n719 = ( n446 & n530 ) | ( n446 & n621 ) | ( n530 & n621 ) ;
  assign n720 = n719 ^ x1 ^ 1'b0 ;
  assign n721 = x6 & x250 ;
  assign n722 = n721 ^ n442 ^ 1'b0 ;
  assign n723 = ( n331 & ~n387 ) | ( n331 & n722 ) | ( ~n387 & n722 ) ;
  assign n724 = ~x207 & x225 ;
  assign n725 = n415 & ~n724 ;
  assign n726 = x116 & x159 ;
  assign n727 = ~n488 & n726 ;
  assign n728 = n727 ^ x138 ^ x85 ;
  assign n729 = n666 & ~n728 ;
  assign n730 = x118 & n272 ;
  assign n731 = n730 ^ n431 ^ 1'b0 ;
  assign n732 = n731 ^ n618 ^ 1'b0 ;
  assign n733 = ( x21 & ~x254 ) | ( x21 & n603 ) | ( ~x254 & n603 ) ;
  assign n734 = x55 & ~n733 ;
  assign n735 = n734 ^ n334 ^ 1'b0 ;
  assign n736 = n613 ^ n281 ^ 1'b0 ;
  assign n737 = x164 & ~n736 ;
  assign n738 = ~x46 & x153 ;
  assign n739 = n256 & ~n738 ;
  assign n740 = x157 & ~n615 ;
  assign n741 = n663 ^ n433 ^ 1'b0 ;
  assign n742 = n740 & n741 ;
  assign n743 = x227 & ~n374 ;
  assign n744 = n507 & n743 ;
  assign n745 = n315 | n682 ;
  assign n746 = n744 & ~n745 ;
  assign n747 = n746 ^ n500 ^ 1'b0 ;
  assign n748 = x3 & x73 ;
  assign n749 = n748 ^ n413 ^ 1'b0 ;
  assign n750 = x102 & n749 ;
  assign n751 = n750 ^ x14 ^ 1'b0 ;
  assign n752 = x97 & n437 ;
  assign n753 = x254 & ~n752 ;
  assign n754 = n753 ^ x232 ^ 1'b0 ;
  assign n755 = x227 & ~n707 ;
  assign n756 = x38 & x104 ;
  assign n757 = n756 ^ n585 ^ x197 ;
  assign n758 = x235 ^ x47 ^ 1'b0 ;
  assign n759 = n496 & n758 ;
  assign n760 = n296 ^ x254 ^ 1'b0 ;
  assign n761 = n327 | n760 ;
  assign n762 = n761 ^ n752 ^ 1'b0 ;
  assign n763 = n759 & n762 ;
  assign n764 = x28 & ~n446 ;
  assign n765 = n764 ^ x221 ^ x157 ;
  assign n766 = n550 ^ n518 ^ x180 ;
  assign n767 = ( x11 & x162 ) | ( x11 & n766 ) | ( x162 & n766 ) ;
  assign n768 = x149 & n767 ;
  assign n769 = n768 ^ n585 ^ 1'b0 ;
  assign n770 = x231 & ~n274 ;
  assign n771 = n483 & n770 ;
  assign n772 = n771 ^ n492 ^ 1'b0 ;
  assign n783 = n277 | n281 ;
  assign n784 = x41 | n783 ;
  assign n785 = ~n624 & n784 ;
  assign n786 = n785 ^ n618 ^ 1'b0 ;
  assign n773 = x175 & ~n448 ;
  assign n774 = ~x153 & n773 ;
  assign n775 = x43 & x53 ;
  assign n776 = ~x58 & n775 ;
  assign n777 = x15 & ~n776 ;
  assign n778 = ~x230 & n777 ;
  assign n779 = ( x34 & ~x171 ) | ( x34 & n778 ) | ( ~x171 & n778 ) ;
  assign n780 = n779 ^ x200 ^ 1'b0 ;
  assign n781 = n780 ^ n281 ^ 1'b0 ;
  assign n782 = ~n774 & n781 ;
  assign n787 = n786 ^ n782 ^ 1'b0 ;
  assign n788 = n448 ^ x225 ^ 1'b0 ;
  assign n789 = x118 & ~n788 ;
  assign n790 = n789 ^ n406 ^ 1'b0 ;
  assign n791 = n728 & ~n790 ;
  assign n792 = n791 ^ x99 ^ 1'b0 ;
  assign n794 = n509 ^ x187 ^ 1'b0 ;
  assign n795 = x244 ^ x113 ^ 1'b0 ;
  assign n796 = n794 & n795 ;
  assign n793 = x221 & n272 ;
  assign n797 = n796 ^ n793 ^ 1'b0 ;
  assign n803 = x0 & x26 ;
  assign n804 = n803 ^ x61 ^ 1'b0 ;
  assign n805 = n342 ^ x134 ^ 1'b0 ;
  assign n806 = x11 & ~n805 ;
  assign n807 = ( ~x26 & n804 ) | ( ~x26 & n806 ) | ( n804 & n806 ) ;
  assign n798 = x253 & n543 ;
  assign n799 = ~x0 & n798 ;
  assign n800 = x166 & ~n799 ;
  assign n801 = n317 & n800 ;
  assign n802 = x99 & ~n801 ;
  assign n808 = n807 ^ n802 ^ 1'b0 ;
  assign n809 = ( x29 & x202 ) | ( x29 & ~n416 ) | ( x202 & ~n416 ) ;
  assign n810 = n759 & ~n809 ;
  assign n811 = x148 & ~n491 ;
  assign n812 = ~x37 & n811 ;
  assign n813 = ( ~x155 & x231 ) | ( ~x155 & n411 ) | ( x231 & n411 ) ;
  assign n814 = x196 & ~n794 ;
  assign n815 = n814 ^ x205 ^ 1'b0 ;
  assign n816 = n393 ^ x12 ^ 1'b0 ;
  assign n817 = x235 & ~n816 ;
  assign n818 = x214 & n817 ;
  assign n819 = n818 ^ x33 ^ 1'b0 ;
  assign n820 = n296 | n819 ;
  assign n821 = x112 | n820 ;
  assign n822 = x208 & x253 ;
  assign n823 = ~x250 & n822 ;
  assign n824 = x86 & ~n823 ;
  assign n825 = n363 & n824 ;
  assign n826 = ~n738 & n825 ;
  assign n827 = x108 & n732 ;
  assign n828 = n466 & n827 ;
  assign n829 = n374 ^ x123 ^ 1'b0 ;
  assign n830 = x99 & n829 ;
  assign n833 = x39 & x131 ;
  assign n834 = ~x50 & n833 ;
  assign n835 = ~n585 & n834 ;
  assign n831 = n287 ^ x56 ^ 1'b0 ;
  assign n832 = x110 & n831 ;
  assign n836 = n835 ^ n832 ^ 1'b0 ;
  assign n837 = n631 ^ x188 ^ 1'b0 ;
  assign n838 = x190 & n837 ;
  assign n839 = n838 ^ x191 ^ 1'b0 ;
  assign n840 = x252 ^ x146 ^ x46 ;
  assign n841 = x104 & x188 ;
  assign n842 = n841 ^ x169 ^ 1'b0 ;
  assign n843 = n479 | n842 ;
  assign n844 = n843 ^ x167 ^ 1'b0 ;
  assign n845 = n844 ^ x228 ^ 1'b0 ;
  assign n848 = n440 ^ x216 ^ x47 ;
  assign n846 = n632 ^ x68 ^ 1'b0 ;
  assign n847 = n510 & n846 ;
  assign n849 = n848 ^ n847 ^ 1'b0 ;
  assign n850 = n845 & n849 ;
  assign n851 = ( x233 & n840 ) | ( x233 & ~n850 ) | ( n840 & ~n850 ) ;
  assign n852 = x121 & ~n665 ;
  assign n853 = x184 & n852 ;
  assign n854 = x33 & ~n676 ;
  assign n855 = ~n491 & n854 ;
  assign n856 = n853 & n855 ;
  assign n857 = n834 | n856 ;
  assign n858 = n475 & ~n857 ;
  assign n859 = x58 ^ x5 ^ 1'b0 ;
  assign n860 = n540 & n859 ;
  assign n861 = n860 ^ n789 ^ 1'b0 ;
  assign n862 = x225 & n861 ;
  assign n863 = n516 ^ n310 ^ 1'b0 ;
  assign n864 = n353 & n845 ;
  assign n865 = n329 & n864 ;
  assign n866 = n865 ^ n663 ^ 1'b0 ;
  assign n867 = n679 | n866 ;
  assign n868 = n867 ^ n831 ^ 1'b0 ;
  assign n869 = n703 & ~n868 ;
  assign n870 = x91 & n869 ;
  assign n871 = ~x122 & n870 ;
  assign n872 = x77 & ~x245 ;
  assign n873 = n552 | n872 ;
  assign n874 = n873 ^ n814 ^ 1'b0 ;
  assign n875 = ( ~x69 & n310 ) | ( ~x69 & n477 ) | ( n310 & n477 ) ;
  assign n876 = n579 & ~n875 ;
  assign n877 = n305 ^ x80 ^ 1'b0 ;
  assign n878 = n389 | n446 ;
  assign n879 = n878 ^ n332 ^ 1'b0 ;
  assign n880 = ( x31 & ~x142 ) | ( x31 & n854 ) | ( ~x142 & n854 ) ;
  assign n881 = ~n347 & n880 ;
  assign n882 = ~n271 & n881 ;
  assign n883 = n742 ^ x7 ^ 1'b0 ;
  assign n884 = ~n731 & n757 ;
  assign n885 = ~n703 & n884 ;
  assign n886 = n883 | n885 ;
  assign n887 = x50 & n395 ;
  assign n888 = ~x214 & n887 ;
  assign n889 = n772 ^ x246 ^ x75 ;
  assign n890 = n889 ^ n720 ^ 1'b0 ;
  assign n891 = x84 ^ x45 ^ 1'b0 ;
  assign n892 = x58 & x224 ;
  assign n893 = ~x135 & n892 ;
  assign n894 = x222 | n893 ;
  assign n895 = x119 & x129 ;
  assign n896 = n895 ^ n677 ^ 1'b0 ;
  assign n897 = ~n671 & n896 ;
  assign n898 = x211 & ~n335 ;
  assign n899 = ~x36 & n898 ;
  assign n902 = x3 & x83 ;
  assign n903 = n902 ^ n477 ^ 1'b0 ;
  assign n900 = n455 ^ x158 ^ x9 ;
  assign n901 = ~n893 & n900 ;
  assign n904 = n903 ^ n901 ^ 1'b0 ;
  assign n905 = x216 & ~n431 ;
  assign n906 = ( n899 & n904 ) | ( n899 & n905 ) | ( n904 & n905 ) ;
  assign n907 = ( x44 & ~x93 ) | ( x44 & x110 ) | ( ~x93 & x110 ) ;
  assign n908 = n399 ^ x39 ^ 1'b0 ;
  assign n909 = n907 | n908 ;
  assign n910 = n308 ^ x33 ^ 1'b0 ;
  assign n911 = n566 & ~n910 ;
  assign n912 = x194 & x212 ;
  assign n913 = n912 ^ x57 ^ 1'b0 ;
  assign n914 = n911 & n913 ;
  assign n915 = n809 ^ n440 ^ 1'b0 ;
  assign n916 = ( x42 & x103 ) | ( x42 & ~x190 ) | ( x103 & ~x190 ) ;
  assign n917 = n553 ^ n281 ^ x31 ;
  assign n918 = x60 & n917 ;
  assign n919 = n461 & n918 ;
  assign n920 = ( n389 & n860 ) | ( n389 & ~n919 ) | ( n860 & ~n919 ) ;
  assign n921 = ( n854 & ~n916 ) | ( n854 & n920 ) | ( ~n916 & n920 ) ;
  assign n922 = ~x48 & x94 ;
  assign n923 = x226 ^ x28 ^ x6 ;
  assign n924 = n923 ^ x146 ^ 1'b0 ;
  assign n925 = ~n922 & n924 ;
  assign n927 = ~x8 & x95 ;
  assign n926 = x193 & ~n880 ;
  assign n928 = n927 ^ n926 ^ 1'b0 ;
  assign n929 = n928 ^ x98 ^ 1'b0 ;
  assign n930 = ~n830 & n929 ;
  assign n931 = n516 ^ x31 ^ 1'b0 ;
  assign n932 = n535 & n931 ;
  assign n933 = ~x213 & n806 ;
  assign n934 = n692 ^ x187 ^ 1'b0 ;
  assign n935 = x87 & ~n934 ;
  assign n936 = n935 ^ x88 ^ 1'b0 ;
  assign n937 = n933 & n936 ;
  assign n940 = n260 ^ x69 ^ 1'b0 ;
  assign n938 = x191 & n518 ;
  assign n939 = x85 & ~n938 ;
  assign n941 = n940 ^ n939 ^ 1'b0 ;
  assign n942 = x128 & x240 ;
  assign n943 = n942 ^ x218 ^ 1'b0 ;
  assign n944 = x22 & n899 ;
  assign n945 = n943 | n944 ;
  assign n946 = x51 | n945 ;
  assign n947 = n433 & ~n677 ;
  assign n948 = ~n262 & n947 ;
  assign n949 = n789 | n948 ;
  assign n950 = n375 & n914 ;
  assign n951 = n950 ^ n338 ^ 1'b0 ;
  assign n952 = ~n364 & n688 ;
  assign n953 = n952 ^ x32 ^ 1'b0 ;
  assign n954 = n871 ^ n518 ^ 1'b0 ;
  assign n955 = x214 & ~n595 ;
  assign n956 = n335 & n955 ;
  assign n957 = n956 ^ x99 ^ 1'b0 ;
  assign n958 = ~n867 & n957 ;
  assign n959 = n679 & n831 ;
  assign n960 = n617 ^ n425 ^ 1'b0 ;
  assign n961 = x19 & n960 ;
  assign n962 = x83 & n961 ;
  assign n963 = ~x155 & n962 ;
  assign n964 = n963 ^ n839 ^ n389 ;
  assign n965 = x168 & ~n320 ;
  assign n966 = n965 ^ n599 ^ 1'b0 ;
  assign n967 = ~n812 & n966 ;
  assign n968 = n967 ^ n258 ^ 1'b0 ;
  assign n969 = x33 & n657 ;
  assign n970 = x101 & ~n334 ;
  assign n971 = n705 & ~n778 ;
  assign n972 = x59 & ~n277 ;
  assign n973 = n972 ^ n525 ^ 1'b0 ;
  assign n974 = x10 & ~n813 ;
  assign n975 = n974 ^ n830 ^ 1'b0 ;
  assign n976 = ~n973 & n975 ;
  assign n977 = ~n769 & n976 ;
  assign n978 = n911 ^ n725 ^ 1'b0 ;
  assign n979 = x11 & x237 ;
  assign n980 = ~n449 & n979 ;
  assign n981 = n980 ^ n913 ^ 1'b0 ;
  assign n982 = ~n535 & n981 ;
  assign n983 = x61 & ~x206 ;
  assign n984 = x43 | n983 ;
  assign n985 = ( ~n281 & n903 ) | ( ~n281 & n984 ) | ( n903 & n984 ) ;
  assign n986 = n985 ^ n875 ^ 1'b0 ;
  assign n987 = n349 | n562 ;
  assign n988 = n842 ^ x82 ^ 1'b0 ;
  assign n989 = x170 ^ x71 ^ 1'b0 ;
  assign n990 = x253 & n989 ;
  assign n991 = ~n733 & n990 ;
  assign n992 = n966 ^ x63 ^ 1'b0 ;
  assign n993 = n449 ^ n375 ^ x119 ;
  assign n994 = n790 | n993 ;
  assign n995 = x46 & ~n453 ;
  assign n996 = n391 ^ n294 ^ x95 ;
  assign n997 = ( x213 & ~n817 ) | ( x213 & n996 ) | ( ~n817 & n996 ) ;
  assign n998 = n479 | n963 ;
  assign n1000 = n511 ^ n417 ^ 1'b0 ;
  assign n1001 = x123 & ~n1000 ;
  assign n999 = x232 & n666 ;
  assign n1002 = n1001 ^ n999 ^ 1'b0 ;
  assign n1003 = x16 & ~n1002 ;
  assign n1004 = ~x64 & n1003 ;
  assign n1010 = n776 ^ x144 ^ 1'b0 ;
  assign n1005 = n631 ^ x139 ^ 1'b0 ;
  assign n1006 = n351 & n1005 ;
  assign n1007 = x119 ^ x89 ^ 1'b0 ;
  assign n1008 = x220 & n1007 ;
  assign n1009 = n1006 & n1008 ;
  assign n1011 = n1010 ^ n1009 ^ 1'b0 ;
  assign n1012 = n862 & n1011 ;
  assign n1013 = n1012 ^ n305 ^ 1'b0 ;
  assign n1014 = n1013 ^ n562 ^ n364 ;
  assign n1019 = x53 & n779 ;
  assign n1020 = n1019 ^ x215 ^ x121 ;
  assign n1015 = n518 ^ x181 ^ 1'b0 ;
  assign n1016 = n518 | n1015 ;
  assign n1017 = n789 & n1016 ;
  assign n1018 = ( n854 & ~n893 ) | ( n854 & n1017 ) | ( ~n893 & n1017 ) ;
  assign n1021 = n1020 ^ n1018 ^ n449 ;
  assign n1022 = x129 & ~n761 ;
  assign n1023 = n1022 ^ x177 ^ 1'b0 ;
  assign n1024 = x134 ^ x66 ^ 1'b0 ;
  assign n1025 = ~n473 & n1024 ;
  assign n1026 = n567 ^ n431 ^ 1'b0 ;
  assign n1027 = n434 & ~n1026 ;
  assign n1029 = n888 ^ n327 ^ 1'b0 ;
  assign n1030 = x231 & n1029 ;
  assign n1028 = n333 ^ x153 ^ x146 ;
  assign n1031 = n1030 ^ n1028 ^ 1'b0 ;
  assign n1032 = x209 & n1031 ;
  assign n1033 = n1027 & n1032 ;
  assign n1034 = ~x181 & n1033 ;
  assign n1035 = n975 & ~n1034 ;
  assign n1036 = n1035 ^ x199 ^ 1'b0 ;
  assign n1037 = n340 ^ x144 ^ x33 ;
  assign n1038 = n430 ^ n399 ^ 1'b0 ;
  assign n1039 = n425 & n1038 ;
  assign n1041 = n440 | n776 ;
  assign n1042 = x44 | n1041 ;
  assign n1040 = ~n574 & n911 ;
  assign n1043 = n1042 ^ n1040 ^ 1'b0 ;
  assign n1044 = n450 | n1043 ;
  assign n1045 = n1039 | n1044 ;
  assign n1046 = x47 & x80 ;
  assign n1047 = ~x232 & n1046 ;
  assign n1048 = n1047 ^ x229 ^ x62 ;
  assign n1049 = n1048 ^ n900 ^ 1'b0 ;
  assign n1050 = n840 | n1049 ;
  assign n1051 = n437 & ~n1050 ;
  assign n1052 = ~n365 & n417 ;
  assign n1053 = n1052 ^ x229 ^ 1'b0 ;
  assign n1054 = n689 ^ x16 ^ 1'b0 ;
  assign n1055 = ~n624 & n1054 ;
  assign n1056 = ~n661 & n1055 ;
  assign n1057 = n1053 & n1056 ;
  assign n1058 = x226 & ~n1057 ;
  assign n1059 = n574 & n1058 ;
  assign n1060 = n289 | n300 ;
  assign n1061 = ~n587 & n1060 ;
  assign n1062 = n1061 ^ x68 ^ 1'b0 ;
  assign n1069 = x24 & ~n375 ;
  assign n1063 = n613 ^ n318 ^ 1'b0 ;
  assign n1064 = x125 & n1063 ;
  assign n1065 = n494 ^ x16 ^ 1'b0 ;
  assign n1066 = x187 & ~n1065 ;
  assign n1067 = n1066 ^ x103 ^ 1'b0 ;
  assign n1068 = n1064 & ~n1067 ;
  assign n1070 = n1069 ^ n1068 ^ 1'b0 ;
  assign n1071 = x135 | n1062 ;
  assign n1072 = n378 & n794 ;
  assign n1073 = n1072 ^ x119 ^ 1'b0 ;
  assign n1074 = x148 & ~n1073 ;
  assign n1075 = n1074 ^ x55 ^ 1'b0 ;
  assign n1076 = n733 ^ x46 ^ 1'b0 ;
  assign n1077 = x39 & ~n1076 ;
  assign n1078 = n1077 ^ n809 ^ 1'b0 ;
  assign n1079 = n276 | n1064 ;
  assign n1082 = n927 ^ x250 ^ 1'b0 ;
  assign n1083 = x163 & ~n1082 ;
  assign n1084 = n1083 ^ n312 ^ 1'b0 ;
  assign n1085 = n355 & ~n1084 ;
  assign n1080 = x110 & ~x207 ;
  assign n1081 = ~n767 & n1080 ;
  assign n1086 = n1085 ^ n1081 ^ 1'b0 ;
  assign n1087 = n1079 | n1086 ;
  assign n1088 = n1087 ^ x44 ^ 1'b0 ;
  assign n1089 = ~x150 & x229 ;
  assign n1090 = x204 & n1089 ;
  assign n1091 = n1090 ^ n423 ^ 1'b0 ;
  assign n1092 = n437 | n1025 ;
  assign n1093 = n298 | n740 ;
  assign n1094 = x249 ^ x168 ^ x47 ;
  assign n1095 = n393 & ~n1094 ;
  assign n1096 = n1095 ^ n446 ^ 1'b0 ;
  assign n1097 = x24 | n865 ;
  assign n1098 = n1097 ^ n535 ^ 1'b0 ;
  assign n1099 = n1080 ^ n473 ^ 1'b0 ;
  assign n1100 = x175 & ~n613 ;
  assign n1101 = n1100 ^ n672 ^ x230 ;
  assign n1102 = n779 | n1049 ;
  assign n1103 = n1102 ^ n421 ^ 1'b0 ;
  assign n1104 = n1103 ^ n988 ^ 1'b0 ;
  assign n1105 = n1101 | n1104 ;
  assign n1106 = n430 ^ x56 ^ 1'b0 ;
  assign n1107 = x80 & ~n1106 ;
  assign n1108 = ~n382 & n931 ;
  assign n1109 = n1108 ^ x122 ^ 1'b0 ;
  assign n1110 = n1109 ^ x215 ^ 1'b0 ;
  assign n1111 = n1107 & ~n1110 ;
  assign n1112 = n1111 ^ n417 ^ 1'b0 ;
  assign n1113 = x107 & x244 ;
  assign n1114 = ~n1112 & n1113 ;
  assign n1115 = x158 & n266 ;
  assign n1116 = n274 & n1115 ;
  assign n1117 = n778 ^ x118 ^ 1'b0 ;
  assign n1118 = x17 & ~n1117 ;
  assign n1119 = ( ~x163 & n540 ) | ( ~x163 & n842 ) | ( n540 & n842 ) ;
  assign n1120 = n1118 & n1119 ;
  assign n1121 = n1120 ^ n713 ^ n694 ;
  assign n1122 = n903 ^ n897 ^ 1'b0 ;
  assign n1123 = n1121 & n1122 ;
  assign n1124 = n787 ^ n485 ^ n306 ;
  assign n1125 = n270 ^ x173 ^ 1'b0 ;
  assign n1128 = n550 ^ n312 ^ 1'b0 ;
  assign n1129 = n591 & n1128 ;
  assign n1126 = ( n283 & ~n380 ) | ( n283 & n425 ) | ( ~n380 & n425 ) ;
  assign n1127 = ~n300 & n1126 ;
  assign n1130 = n1129 ^ n1127 ^ 1'b0 ;
  assign n1131 = n661 ^ n455 ^ 1'b0 ;
  assign n1132 = x199 & n1131 ;
  assign n1133 = n314 | n1132 ;
  assign n1134 = n790 ^ n500 ^ 1'b0 ;
  assign n1135 = x180 & ~n932 ;
  assign n1136 = x89 & n415 ;
  assign n1137 = n1136 ^ n503 ^ 1'b0 ;
  assign n1138 = n1010 | n1080 ;
  assign n1139 = ~n1137 & n1138 ;
  assign n1140 = n1139 ^ n1039 ^ 1'b0 ;
  assign n1147 = n394 ^ x154 ^ x92 ;
  assign n1148 = ( n407 & ~n694 ) | ( n407 & n1147 ) | ( ~n694 & n1147 ) ;
  assign n1141 = x175 ^ x101 ^ 1'b0 ;
  assign n1142 = x2 & n1141 ;
  assign n1143 = n1142 ^ x243 ^ 1'b0 ;
  assign n1144 = n540 & n1143 ;
  assign n1145 = ~n317 & n1144 ;
  assign n1146 = ~x199 & n1145 ;
  assign n1149 = n1148 ^ n1146 ^ 1'b0 ;
  assign n1150 = x113 ^ x61 ^ 1'b0 ;
  assign n1151 = ~n457 & n1150 ;
  assign n1152 = ( x112 & n1049 ) | ( x112 & ~n1151 ) | ( n1049 & ~n1151 ) ;
  assign n1153 = ( n395 & ~n763 ) | ( n395 & n1152 ) | ( ~n763 & n1152 ) ;
  assign n1154 = x78 | n778 ;
  assign n1155 = n1154 ^ n907 ^ 1'b0 ;
  assign n1156 = n262 & n1155 ;
  assign n1157 = n1156 ^ n542 ^ x55 ;
  assign n1158 = ~n969 & n1157 ;
  assign n1159 = n1158 ^ x186 ^ 1'b0 ;
  assign n1160 = n738 ^ n634 ^ 1'b0 ;
  assign n1161 = ( ~x130 & x167 ) | ( ~x130 & n1160 ) | ( x167 & n1160 ) ;
  assign n1162 = ~n374 & n1161 ;
  assign n1163 = ~x254 & n1162 ;
  assign n1164 = n555 ^ x195 ^ 1'b0 ;
  assign n1165 = n618 | n1164 ;
  assign n1166 = n1097 & ~n1165 ;
  assign n1167 = n1166 ^ n975 ^ 1'b0 ;
  assign n1168 = n562 & n1167 ;
  assign n1169 = x122 & ~n778 ;
  assign n1170 = x118 & x249 ;
  assign n1171 = n1169 & n1170 ;
  assign n1172 = n1171 ^ n713 ^ 1'b0 ;
  assign n1173 = n1172 ^ n907 ^ 1'b0 ;
  assign n1174 = x48 & ~n1173 ;
  assign n1175 = ~x104 & n796 ;
  assign n1176 = n713 ^ n374 ^ 1'b0 ;
  assign n1177 = n784 ^ x244 ^ x95 ;
  assign n1178 = x17 & ~x139 ;
  assign n1179 = x159 & ~n1178 ;
  assign n1180 = n1179 ^ n1109 ^ 1'b0 ;
  assign n1181 = x145 ^ x73 ^ 1'b0 ;
  assign n1182 = n1180 & n1181 ;
  assign n1183 = x241 & n799 ;
  assign n1184 = n1183 ^ x164 ^ 1'b0 ;
  assign n1185 = n810 | n1184 ;
  assign n1186 = n1185 ^ n1103 ^ 1'b0 ;
  assign n1188 = ~n513 & n1064 ;
  assign n1189 = n1188 ^ n896 ^ 1'b0 ;
  assign n1187 = ~n287 & n1042 ;
  assign n1190 = n1189 ^ n1187 ^ 1'b0 ;
  assign n1191 = x87 & x102 ;
  assign n1192 = ~x54 & n1191 ;
  assign n1193 = n619 & n1089 ;
  assign n1194 = n294 & ~n1193 ;
  assign n1195 = n1194 ^ n871 ^ 1'b0 ;
  assign n1196 = n611 ^ x87 ^ 1'b0 ;
  assign n1197 = n1195 & n1196 ;
  assign n1198 = ~x168 & x205 ;
  assign n1199 = ( x235 & n448 ) | ( x235 & n1198 ) | ( n448 & n1198 ) ;
  assign n1202 = x23 & ~n614 ;
  assign n1203 = n1202 ^ n1064 ^ 1'b0 ;
  assign n1200 = ( x38 & ~x236 ) | ( x38 & n455 ) | ( ~x236 & n455 ) ;
  assign n1201 = n828 | n1200 ;
  assign n1204 = n1203 ^ n1201 ^ 1'b0 ;
  assign n1205 = n794 & ~n830 ;
  assign n1206 = ~x141 & n1205 ;
  assign n1207 = x184 & ~n497 ;
  assign n1208 = n1207 ^ x124 ^ 1'b0 ;
  assign n1209 = n774 ^ n477 ^ 1'b0 ;
  assign n1210 = n1208 | n1209 ;
  assign n1211 = n1210 ^ x222 ^ 1'b0 ;
  assign n1212 = n556 & ~n1211 ;
  assign n1213 = n1212 ^ n500 ^ 1'b0 ;
  assign n1214 = ~n333 & n553 ;
  assign n1215 = ~n540 & n1214 ;
  assign n1216 = n1215 ^ n867 ^ 1'b0 ;
  assign n1217 = ~n692 & n1216 ;
  assign n1218 = x177 & ~n752 ;
  assign n1219 = ~x146 & n1218 ;
  assign n1220 = ( ~x251 & n624 ) | ( ~x251 & n1126 ) | ( n624 & n1126 ) ;
  assign n1221 = ( x10 & ~n1219 ) | ( x10 & n1220 ) | ( ~n1219 & n1220 ) ;
  assign n1222 = x193 & n1221 ;
  assign n1223 = n1222 ^ n716 ^ 1'b0 ;
  assign n1224 = x101 & x198 ;
  assign n1225 = ~n380 & n1224 ;
  assign n1226 = ~n496 & n925 ;
  assign n1227 = n1225 & n1226 ;
  assign n1228 = n1161 ^ n689 ^ 1'b0 ;
  assign n1229 = n1228 ^ n618 ^ 1'b0 ;
  assign n1230 = x187 & ~n1229 ;
  assign n1231 = n442 ^ n293 ^ 1'b0 ;
  assign n1236 = n425 & ~n1137 ;
  assign n1237 = ~n680 & n1236 ;
  assign n1232 = n844 ^ x191 ^ x87 ;
  assign n1233 = x97 & n632 ;
  assign n1234 = n1233 ^ n461 ^ 1'b0 ;
  assign n1235 = ~n1232 & n1234 ;
  assign n1238 = n1237 ^ n1235 ^ 1'b0 ;
  assign n1239 = n628 ^ x205 ^ 1'b0 ;
  assign n1240 = x153 & n1239 ;
  assign n1241 = ~n308 & n357 ;
  assign n1242 = ~x41 & n1241 ;
  assign n1243 = x241 & ~n349 ;
  assign n1244 = ~x153 & n1243 ;
  assign n1245 = ( n1240 & ~n1242 ) | ( n1240 & n1244 ) | ( ~n1242 & n1244 ) ;
  assign n1246 = n272 ^ x1 ^ 1'b0 ;
  assign n1247 = ~n457 & n1246 ;
  assign n1248 = n1247 ^ x237 ^ 1'b0 ;
  assign n1249 = ~n457 & n1248 ;
  assign n1250 = n1118 ^ n449 ^ 1'b0 ;
  assign n1251 = n603 | n1250 ;
  assign n1252 = n1251 ^ n260 ^ 1'b0 ;
  assign n1253 = x108 & ~n829 ;
  assign n1254 = n1253 ^ n804 ^ 1'b0 ;
  assign n1255 = ~n707 & n1254 ;
  assign n1257 = ~n424 & n917 ;
  assign n1256 = n883 | n1200 ;
  assign n1258 = n1257 ^ n1256 ^ 1'b0 ;
  assign n1259 = x32 & n1258 ;
  assign n1260 = n840 | n1259 ;
  assign n1261 = n1260 ^ n314 ^ 1'b0 ;
  assign n1262 = n958 ^ n530 ^ 1'b0 ;
  assign n1263 = x141 & x144 ;
  assign n1264 = ~x190 & n1263 ;
  assign n1265 = n946 & n1264 ;
  assign n1266 = n285 | n595 ;
  assign n1267 = n1265 & ~n1266 ;
  assign n1268 = x29 & n302 ;
  assign n1269 = n1268 ^ n1264 ^ 1'b0 ;
  assign n1270 = ~n711 & n1269 ;
  assign n1271 = n1242 & n1270 ;
  assign n1272 = x206 & ~n1156 ;
  assign n1273 = ~x107 & x187 ;
  assign n1274 = x118 | n643 ;
  assign n1275 = ~n1273 & n1274 ;
  assign n1276 = ~n1272 & n1275 ;
  assign n1277 = n839 & n985 ;
  assign n1278 = n1277 ^ n677 ^ 1'b0 ;
  assign n1279 = n1051 ^ n1027 ^ 1'b0 ;
  assign n1280 = n613 & ~n643 ;
  assign n1281 = n1280 ^ x54 ^ 1'b0 ;
  assign n1282 = x121 & ~n479 ;
  assign n1283 = n317 & n1282 ;
  assign n1284 = n1281 | n1283 ;
  assign n1285 = n395 & ~n997 ;
  assign n1286 = ~x134 & n1285 ;
  assign n1287 = n1286 ^ n604 ^ 1'b0 ;
  assign n1288 = n751 | n1287 ;
  assign n1289 = x187 & ~n695 ;
  assign n1290 = n1289 ^ n863 ^ 1'b0 ;
  assign n1292 = ( x106 & n338 ) | ( x106 & n498 ) | ( n338 & n498 ) ;
  assign n1291 = n367 & ~n819 ;
  assign n1293 = n1292 ^ n1291 ^ 1'b0 ;
  assign n1294 = n710 | n1293 ;
  assign n1295 = ( n459 & ~n613 ) | ( n459 & n906 ) | ( ~n613 & n906 ) ;
  assign n1296 = n404 ^ x244 ^ 1'b0 ;
  assign n1297 = n1295 & n1296 ;
  assign n1298 = ( ~n287 & n430 ) | ( ~n287 & n1297 ) | ( n430 & n1297 ) ;
  assign n1299 = ~n692 & n1186 ;
  assign n1300 = n1299 ^ n638 ^ 1'b0 ;
  assign n1301 = n1211 ^ n724 ^ n638 ;
  assign n1302 = n1023 | n1051 ;
  assign n1303 = n1302 ^ n1125 ^ 1'b0 ;
  assign n1304 = x182 & ~n1126 ;
  assign n1305 = x137 & ~n863 ;
  assign n1306 = n738 & n1305 ;
  assign n1307 = ~n963 & n1306 ;
  assign n1308 = n801 | n1307 ;
  assign n1309 = n1304 & ~n1308 ;
  assign n1310 = n331 | n1309 ;
  assign n1311 = x58 | n1310 ;
  assign n1312 = x217 & ~n963 ;
  assign n1313 = n1312 ^ n1309 ^ n262 ;
  assign n1314 = n359 & n686 ;
  assign n1315 = n1314 ^ n1135 ^ 1'b0 ;
  assign n1316 = n1313 & n1315 ;
  assign n1317 = ~n477 & n1186 ;
  assign n1318 = x127 & n914 ;
  assign n1319 = ~n276 & n1156 ;
  assign n1320 = ~n657 & n970 ;
  assign n1321 = ~x27 & n1320 ;
  assign n1322 = n1321 ^ n1315 ^ n888 ;
  assign n1323 = x227 & x232 ;
  assign n1324 = ~x136 & n1323 ;
  assign n1325 = n491 | n1324 ;
  assign n1326 = n835 & ~n1325 ;
  assign n1327 = n302 & ~n481 ;
  assign n1328 = ~x137 & n1327 ;
  assign n1329 = n1328 ^ n661 ^ 1'b0 ;
  assign n1330 = ~n677 & n1329 ;
  assign n1331 = n579 & n1330 ;
  assign n1332 = n1326 & n1331 ;
  assign n1333 = n883 ^ x122 ^ 1'b0 ;
  assign n1334 = n675 ^ x146 ^ 1'b0 ;
  assign n1335 = x163 & ~n1334 ;
  assign n1336 = ( ~x208 & n491 ) | ( ~x208 & n705 ) | ( n491 & n705 ) ;
  assign n1337 = n1336 ^ n1185 ^ 1'b0 ;
  assign n1338 = n1335 & n1337 ;
  assign n1339 = x16 & x220 ;
  assign n1340 = n1114 & n1339 ;
  assign n1343 = x147 & n473 ;
  assign n1341 = n318 & ~n333 ;
  assign n1342 = n1341 ^ n1190 ^ 1'b0 ;
  assign n1344 = n1343 ^ n1342 ^ x102 ;
  assign n1345 = n580 ^ n459 ^ 1'b0 ;
  assign n1346 = n1345 ^ n1290 ^ 1'b0 ;
  assign n1347 = n413 & ~n709 ;
  assign n1348 = n637 | n1347 ;
  assign n1349 = n338 & ~n1348 ;
  assign n1350 = x84 & n387 ;
  assign n1351 = n804 & n1350 ;
  assign n1352 = n1351 ^ n953 ^ x153 ;
  assign n1353 = n789 & n941 ;
  assign n1354 = n1328 | n1353 ;
  assign n1355 = n1099 ^ n724 ^ 1'b0 ;
  assign n1356 = x115 & ~n1355 ;
  assign n1357 = n888 ^ n875 ^ 1'b0 ;
  assign n1358 = n1356 & ~n1357 ;
  assign n1359 = ~n766 & n806 ;
  assign n1360 = ~n279 & n1359 ;
  assign n1361 = n1360 ^ n1094 ^ 1'b0 ;
  assign n1362 = n498 & n663 ;
  assign n1363 = n647 & n742 ;
  assign n1364 = ~n428 & n1363 ;
  assign n1365 = n964 ^ n778 ^ n302 ;
  assign n1366 = n1176 & ~n1365 ;
  assign n1367 = n376 ^ x186 ^ 1'b0 ;
  assign n1368 = n1258 & n1367 ;
  assign n1369 = ~n659 & n729 ;
  assign n1370 = n956 ^ n711 ^ 1'b0 ;
  assign n1371 = x247 & n1370 ;
  assign n1372 = n794 ^ n498 ^ 1'b0 ;
  assign n1373 = n1371 & ~n1372 ;
  assign n1374 = ( ~n739 & n1100 ) | ( ~n739 & n1373 ) | ( n1100 & n1373 ) ;
  assign n1375 = x81 & ~n464 ;
  assign n1376 = n1375 ^ n732 ^ 1'b0 ;
  assign n1377 = n738 & ~n1376 ;
  assign n1378 = n1374 & n1377 ;
  assign n1379 = n271 & ~n430 ;
  assign n1380 = x125 & x148 ;
  assign n1381 = n309 & n1380 ;
  assign n1382 = x203 & n1381 ;
  assign n1383 = x191 & ~n1382 ;
  assign n1384 = n496 ^ x180 ^ 1'b0 ;
  assign n1385 = n1159 ^ n893 ^ 1'b0 ;
  assign n1386 = ( n464 & n492 ) | ( n464 & n872 ) | ( n492 & n872 ) ;
  assign n1387 = x57 | n1386 ;
  assign n1388 = n949 ^ n369 ^ 1'b0 ;
  assign n1389 = n1176 ^ n618 ^ 1'b0 ;
  assign n1390 = x137 & x248 ;
  assign n1391 = ~x243 & n1390 ;
  assign n1392 = x42 | n1391 ;
  assign n1393 = ( n789 & n925 ) | ( n789 & n1250 ) | ( n925 & n1250 ) ;
  assign n1394 = n1125 ^ x11 ^ 1'b0 ;
  assign n1395 = n1393 & ~n1394 ;
  assign n1396 = n671 & ~n1051 ;
  assign n1397 = n571 & n1396 ;
  assign n1398 = n1397 ^ x172 ^ 1'b0 ;
  assign n1399 = x181 & x234 ;
  assign n1400 = n1398 & n1399 ;
  assign n1401 = x140 & ~n635 ;
  assign n1402 = ~n794 & n1401 ;
  assign n1403 = n543 & ~n1013 ;
  assign n1404 = n1403 ^ n987 ^ 1'b0 ;
  assign n1405 = n1099 ^ n703 ^ 1'b0 ;
  assign n1406 = n1313 & ~n1398 ;
  assign n1408 = x102 & n525 ;
  assign n1409 = ~x170 & n1408 ;
  assign n1407 = x231 & n532 ;
  assign n1410 = n1409 ^ n1407 ^ 1'b0 ;
  assign n1411 = ( ~x70 & n498 ) | ( ~x70 & n1410 ) | ( n498 & n1410 ) ;
  assign n1412 = x98 ^ x48 ^ 1'b0 ;
  assign n1413 = ~n1411 & n1412 ;
  assign n1414 = n1142 & n1371 ;
  assign n1415 = n1414 ^ x121 ^ 1'b0 ;
  assign n1416 = n1415 ^ n1011 ^ 1'b0 ;
  assign n1417 = n501 ^ n399 ^ 1'b0 ;
  assign n1418 = ~n507 & n1417 ;
  assign n1419 = n1418 ^ x45 ^ 1'b0 ;
  assign n1420 = ( n446 & ~n1382 ) | ( n446 & n1419 ) | ( ~n1382 & n1419 ) ;
  assign n1421 = n569 & ~n1420 ;
  assign n1422 = ~n1416 & n1421 ;
  assign n1423 = n796 ^ n627 ^ 1'b0 ;
  assign n1424 = n601 | n889 ;
  assign n1425 = n1424 ^ n1123 ^ 1'b0 ;
  assign n1426 = n1307 | n1425 ;
  assign n1427 = n1423 & ~n1426 ;
  assign n1428 = ~x150 & n1427 ;
  assign n1429 = x50 & x106 ;
  assign n1430 = n606 & n1429 ;
  assign n1431 = x252 & ~n1430 ;
  assign n1432 = n1431 ^ n1048 ^ 1'b0 ;
  assign n1433 = n575 & ~n1203 ;
  assign n1434 = n1433 ^ n714 ^ 1'b0 ;
  assign n1435 = n518 & ~n1434 ;
  assign n1436 = x0 & ~n1002 ;
  assign n1437 = ~x115 & n1436 ;
  assign n1438 = n389 | n1437 ;
  assign n1439 = n1067 & ~n1438 ;
  assign n1440 = n1437 ^ n1213 ^ 1'b0 ;
  assign n1441 = n1409 ^ x185 ^ 1'b0 ;
  assign n1442 = ( x41 & n893 ) | ( x41 & n916 ) | ( n893 & n916 ) ;
  assign n1443 = ( x124 & ~x189 ) | ( x124 & n761 ) | ( ~x189 & n761 ) ;
  assign n1444 = x165 & ~n314 ;
  assign n1445 = n1443 & n1444 ;
  assign n1446 = n1144 & ~n1445 ;
  assign n1447 = n1446 ^ x191 ^ 1'b0 ;
  assign n1448 = n1442 & ~n1447 ;
  assign n1449 = ~n1441 & n1448 ;
  assign n1450 = n755 & ~n1147 ;
  assign n1451 = ( x54 & ~n567 ) | ( x54 & n1450 ) | ( ~n567 & n1450 ) ;
  assign n1452 = ~n1449 & n1451 ;
  assign n1453 = n1452 ^ n714 ^ 1'b0 ;
  assign n1454 = x103 & n535 ;
  assign n1455 = n1453 & n1454 ;
  assign n1456 = n1455 ^ n744 ^ 1'b0 ;
  assign n1457 = n260 | n1288 ;
  assign n1458 = ~n891 & n1376 ;
  assign n1461 = n911 & n917 ;
  assign n1462 = n1461 ^ n264 ^ 1'b0 ;
  assign n1459 = n1060 ^ n819 ^ 1'b0 ;
  assign n1460 = n1379 & n1459 ;
  assign n1463 = n1462 ^ n1460 ^ 1'b0 ;
  assign n1464 = x124 & ~n1049 ;
  assign n1465 = n1464 ^ x221 ^ 1'b0 ;
  assign n1466 = x59 & ~x183 ;
  assign n1467 = n916 ^ n739 ^ 1'b0 ;
  assign n1468 = n1051 ^ n363 ^ 1'b0 ;
  assign n1469 = n1208 | n1468 ;
  assign n1470 = n1469 ^ x194 ^ 1'b0 ;
  assign n1471 = n1140 ^ x12 ^ 1'b0 ;
  assign n1472 = n1203 ^ n1028 ^ 1'b0 ;
  assign n1473 = n1471 | n1472 ;
  assign n1474 = ( x82 & n977 ) | ( x82 & n1467 ) | ( n977 & n1467 ) ;
  assign n1475 = n1219 ^ n1129 ^ 1'b0 ;
  assign n1476 = x25 & x230 ;
  assign n1477 = n642 & n1476 ;
  assign n1478 = n1100 & ~n1477 ;
  assign n1479 = ~n419 & n534 ;
  assign n1480 = n1479 ^ n984 ^ 1'b0 ;
  assign n1481 = n361 & n471 ;
  assign n1483 = x248 & ~n1381 ;
  assign n1484 = n1483 ^ n957 ^ 1'b0 ;
  assign n1485 = n1081 ^ x132 ^ 1'b0 ;
  assign n1486 = n1484 & ~n1485 ;
  assign n1482 = n1083 ^ x207 ^ x31 ;
  assign n1487 = n1486 ^ n1482 ^ n448 ;
  assign n1488 = n1023 | n1244 ;
  assign n1489 = n1487 & ~n1488 ;
  assign n1490 = n413 ^ x208 ^ 1'b0 ;
  assign n1491 = n1490 ^ n908 ^ 1'b0 ;
  assign n1492 = n796 & n1491 ;
  assign n1501 = ( x4 & ~x60 ) | ( x4 & x208 ) | ( ~x60 & x208 ) ;
  assign n1502 = x172 & n1501 ;
  assign n1503 = n1502 ^ n503 ^ 1'b0 ;
  assign n1496 = n349 ^ x181 ^ 1'b0 ;
  assign n1497 = n1496 ^ n615 ^ n402 ;
  assign n1498 = x137 & n1497 ;
  assign n1499 = ~n1089 & n1498 ;
  assign n1494 = n668 ^ n256 ^ 1'b0 ;
  assign n1493 = n1165 | n1450 ;
  assign n1495 = n1494 ^ n1493 ^ 1'b0 ;
  assign n1500 = n1499 ^ n1495 ^ 1'b0 ;
  assign n1504 = n1503 ^ n1500 ^ 1'b0 ;
  assign n1505 = n369 & ~n1398 ;
  assign n1506 = n694 & n1231 ;
  assign n1507 = n893 ^ n545 ^ 1'b0 ;
  assign n1508 = n821 & ~n1507 ;
  assign n1509 = n1508 ^ n1252 ^ 1'b0 ;
  assign n1510 = n1509 ^ x236 ^ 1'b0 ;
  assign n1511 = n713 ^ n294 ^ 1'b0 ;
  assign n1512 = ~n329 & n1511 ;
  assign n1513 = ( ~x41 & n854 ) | ( ~x41 & n1512 ) | ( n854 & n1512 ) ;
  assign n1516 = n666 ^ n340 ^ 1'b0 ;
  assign n1514 = ( x56 & ~x221 ) | ( x56 & n455 ) | ( ~x221 & n455 ) ;
  assign n1515 = n1410 & ~n1514 ;
  assign n1517 = n1516 ^ n1515 ^ 1'b0 ;
  assign n1518 = ~n306 & n1293 ;
  assign n1519 = n1518 ^ n749 ^ 1'b0 ;
  assign n1520 = n1303 ^ n1290 ^ 1'b0 ;
  assign n1521 = n679 | n1520 ;
  assign n1522 = n1521 ^ n780 ^ 1'b0 ;
  assign n1523 = ( x252 & ~n260 ) | ( x252 & n1129 ) | ( ~n260 & n1129 ) ;
  assign n1524 = ~n399 & n1523 ;
  assign n1525 = n1524 ^ x141 ^ 1'b0 ;
  assign n1526 = x55 & ~n1525 ;
  assign n1527 = ~x178 & n1526 ;
  assign n1528 = n1522 & n1527 ;
  assign n1529 = x88 & n688 ;
  assign n1530 = ~n604 & n1529 ;
  assign n1531 = n464 | n1530 ;
  assign n1532 = n1531 ^ n577 ^ 1'b0 ;
  assign n1533 = n1532 ^ n445 ^ 1'b0 ;
  assign n1534 = n402 & ~n1533 ;
  assign n1535 = n464 | n1534 ;
  assign n1536 = n1535 ^ x88 ^ 1'b0 ;
  assign n1537 = n421 & ~n711 ;
  assign n1538 = ~n1254 & n1537 ;
  assign n1539 = x16 & n1538 ;
  assign n1540 = n372 | n1539 ;
  assign n1541 = n701 | n1540 ;
  assign n1542 = n1366 & n1541 ;
  assign n1543 = n1542 ^ n853 ^ 1'b0 ;
  assign n1544 = n1409 ^ n1064 ^ 1'b0 ;
  assign n1545 = n794 ^ n510 ^ x104 ;
  assign n1546 = n1247 & ~n1545 ;
  assign n1547 = ~x155 & n1546 ;
  assign n1548 = n651 ^ n466 ^ 1'b0 ;
  assign n1549 = ~n550 & n1083 ;
  assign n1550 = n1549 ^ n1254 ^ 1'b0 ;
  assign n1551 = ~x46 & x158 ;
  assign n1552 = x173 | n1551 ;
  assign n1553 = n1552 ^ n1195 ^ 1'b0 ;
  assign n1560 = n679 ^ n513 ^ 1'b0 ;
  assign n1561 = ~n611 & n1560 ;
  assign n1554 = x64 | n725 ;
  assign n1555 = ~n314 & n659 ;
  assign n1556 = ~x221 & n1555 ;
  assign n1557 = ~n298 & n1556 ;
  assign n1558 = n1557 ^ x88 ^ 1'b0 ;
  assign n1559 = ~n1554 & n1558 ;
  assign n1562 = n1561 ^ n1559 ^ 1'b0 ;
  assign n1563 = n266 & ~n603 ;
  assign n1564 = n1028 ^ n808 ^ 1'b0 ;
  assign n1565 = x19 & n1564 ;
  assign n1566 = ( x118 & n1554 ) | ( x118 & ~n1565 ) | ( n1554 & ~n1565 ) ;
  assign n1567 = n1566 ^ n1085 ^ 1'b0 ;
  assign n1568 = x217 & ~n1567 ;
  assign n1569 = n1332 & n1453 ;
  assign n1570 = n1048 ^ n496 ^ 1'b0 ;
  assign n1571 = x7 & n1570 ;
  assign n1572 = n530 ^ n511 ^ 1'b0 ;
  assign n1573 = n1571 & ~n1572 ;
  assign n1574 = x185 & ~n738 ;
  assign n1575 = ~n749 & n1574 ;
  assign n1576 = x73 & x243 ;
  assign n1577 = n1576 ^ x10 ^ 1'b0 ;
  assign n1578 = x78 & ~n1577 ;
  assign n1579 = n996 & n1578 ;
  assign n1580 = n488 ^ x223 ^ 1'b0 ;
  assign n1581 = x236 & n1580 ;
  assign n1582 = n860 & n1581 ;
  assign n1583 = n1579 & n1582 ;
  assign n1584 = n893 | n1583 ;
  assign n1585 = n1584 ^ x141 ^ 1'b0 ;
  assign n1586 = n1585 ^ n464 ^ 1'b0 ;
  assign n1587 = n542 ^ x221 ^ 1'b0 ;
  assign n1588 = n1182 & ~n1587 ;
  assign n1589 = n778 ^ n680 ^ 1'b0 ;
  assign n1590 = n1049 & n1589 ;
  assign n1591 = n659 | n1590 ;
  assign n1592 = ( ~x71 & n1156 ) | ( ~x71 & n1324 ) | ( n1156 & n1324 ) ;
  assign n1593 = n619 | n911 ;
  assign n1594 = x63 & ~n957 ;
  assign n1595 = n1593 & n1594 ;
  assign n1596 = n1595 ^ n488 ^ 1'b0 ;
  assign n1597 = n332 | n893 ;
  assign n1598 = n1597 ^ x214 ^ 1'b0 ;
  assign n1599 = n1170 & n1598 ;
  assign n1600 = n1599 ^ n1065 ^ 1'b0 ;
  assign n1601 = x48 & n366 ;
  assign n1602 = ~x111 & n1601 ;
  assign n1603 = ( x222 & ~n789 ) | ( x222 & n1602 ) | ( ~n789 & n1602 ) ;
  assign n1604 = x204 & n1330 ;
  assign n1605 = n1603 & n1604 ;
  assign n1606 = n809 ^ n661 ^ x151 ;
  assign n1607 = n1606 ^ x80 ^ 1'b0 ;
  assign n1608 = ~n1605 & n1607 ;
  assign n1609 = x68 & x139 ;
  assign n1610 = n1609 ^ n479 ^ 1'b0 ;
  assign n1611 = ~n1417 & n1610 ;
  assign n1612 = ( n353 & ~n599 ) | ( n353 & n807 ) | ( ~n599 & n807 ) ;
  assign n1613 = n1279 ^ n543 ^ x57 ;
  assign n1614 = ~n363 & n1042 ;
  assign n1615 = ~n520 & n1614 ;
  assign n1616 = ~n1345 & n1510 ;
  assign n1617 = n1616 ^ x120 ^ 1'b0 ;
  assign n1619 = n1138 ^ n966 ^ 1'b0 ;
  assign n1618 = n845 & n984 ;
  assign n1620 = n1619 ^ n1618 ^ 1'b0 ;
  assign n1621 = x228 & n1356 ;
  assign n1622 = ~n1620 & n1621 ;
  assign n1623 = x182 ^ x121 ^ 1'b0 ;
  assign n1624 = n1623 ^ n1037 ^ 1'b0 ;
  assign n1626 = n374 | n553 ;
  assign n1625 = n679 | n1306 ;
  assign n1627 = n1626 ^ n1625 ^ 1'b0 ;
  assign n1628 = x206 & ~n1627 ;
  assign n1629 = n764 ^ n638 ^ 1'b0 ;
  assign n1630 = n1424 | n1629 ;
  assign n1631 = x90 & x184 ;
  assign n1632 = n1631 ^ n1417 ^ 1'b0 ;
  assign n1633 = n1632 ^ n534 ^ n498 ;
  assign n1634 = n357 | n1633 ;
  assign n1635 = x214 & n769 ;
  assign n1636 = x18 & ~x212 ;
  assign n1637 = n1636 ^ n631 ^ 1'b0 ;
  assign n1638 = x42 & ~n1637 ;
  assign n1639 = n1385 ^ n671 ^ 1'b0 ;
  assign n1640 = ~n779 & n877 ;
  assign n1641 = n1640 ^ x203 ^ 1'b0 ;
  assign n1642 = x221 & ~n514 ;
  assign n1643 = n1642 ^ n1264 ^ 1'b0 ;
  assign n1644 = n1643 ^ n477 ^ 1'b0 ;
  assign n1645 = ~n1304 & n1644 ;
  assign n1650 = n604 & ~n1119 ;
  assign n1651 = ~x86 & n1650 ;
  assign n1649 = n692 ^ x132 ^ 1'b0 ;
  assign n1652 = n1651 ^ n1649 ^ 1'b0 ;
  assign n1653 = ~n397 & n1652 ;
  assign n1646 = x157 & ~n309 ;
  assign n1647 = n1646 ^ x215 ^ 1'b0 ;
  assign n1648 = x133 & n1647 ;
  assign n1654 = n1653 ^ n1648 ^ n1288 ;
  assign n1655 = x227 & ~n813 ;
  assign n1656 = n1655 ^ x196 ^ 1'b0 ;
  assign n1657 = ~x135 & n425 ;
  assign n1658 = n1254 ^ x191 ^ 1'b0 ;
  assign n1659 = ~n792 & n1658 ;
  assign n1660 = n1441 & n1659 ;
  assign n1661 = n1660 ^ x150 ^ 1'b0 ;
  assign n1662 = ~n1657 & n1661 ;
  assign n1663 = x180 & ~n1328 ;
  assign n1664 = n645 & n1663 ;
  assign n1665 = n1664 ^ n1495 ^ n372 ;
  assign n1666 = x122 & x139 ;
  assign n1667 = ~x227 & n1666 ;
  assign n1668 = n949 ^ x90 ^ 1'b0 ;
  assign n1669 = ~n1667 & n1668 ;
  assign n1670 = n336 & n1367 ;
  assign n1671 = n1670 ^ x198 ^ 1'b0 ;
  assign n1672 = n545 & ~n1671 ;
  assign n1673 = x133 & ~n908 ;
  assign n1674 = n1069 & n1673 ;
  assign n1675 = x228 & ~n1674 ;
  assign n1676 = ~n862 & n1675 ;
  assign n1677 = n599 | n1676 ;
  assign n1678 = n1677 ^ x127 ^ 1'b0 ;
  assign n1679 = n1678 ^ n1417 ^ 1'b0 ;
  assign n1680 = ~n1530 & n1679 ;
  assign n1681 = n376 | n933 ;
  assign n1682 = x181 & n1681 ;
  assign n1683 = n1037 ^ n787 ^ 1'b0 ;
  assign n1684 = n1371 & ~n1683 ;
  assign n1685 = n890 & ~n891 ;
  assign n1686 = ~x4 & n1685 ;
  assign n1687 = n1686 ^ n842 ^ 1'b0 ;
  assign n1688 = n1684 & n1687 ;
  assign n1689 = ~x235 & n305 ;
  assign n1690 = n1689 ^ n808 ^ n642 ;
  assign n1691 = n1635 ^ n1369 ^ 1'b0 ;
  assign n1692 = n907 & n1691 ;
  assign n1693 = n591 & n1692 ;
  assign n1694 = ~n1092 & n1693 ;
  assign n1695 = n731 ^ x136 ^ 1'b0 ;
  assign n1696 = n904 | n1695 ;
  assign n1697 = n525 & ~n1602 ;
  assign n1698 = n1098 & n1697 ;
  assign n1699 = n1698 ^ n1563 ^ 1'b0 ;
  assign n1700 = n359 & ~n1130 ;
  assign n1701 = n1700 ^ n1581 ^ 1'b0 ;
  assign n1703 = n421 & ~n823 ;
  assign n1704 = n334 & n1703 ;
  assign n1705 = x95 & n1664 ;
  assign n1706 = n1705 ^ n894 ^ 1'b0 ;
  assign n1707 = n1704 | n1706 ;
  assign n1708 = n1300 & n1707 ;
  assign n1702 = x125 & x230 ;
  assign n1709 = n1708 ^ n1702 ^ 1'b0 ;
  assign n1710 = n963 ^ n840 ^ n264 ;
  assign n1711 = ( x61 & n651 ) | ( x61 & n1254 ) | ( n651 & n1254 ) ;
  assign n1712 = n1711 ^ n613 ^ x69 ;
  assign n1713 = ~n466 & n1269 ;
  assign n1714 = n727 & n1713 ;
  assign n1715 = n606 | n1714 ;
  assign n1716 = n1715 ^ n540 ^ 1'b0 ;
  assign n1717 = ~n1712 & n1716 ;
  assign n1718 = ~n1710 & n1717 ;
  assign n1720 = n993 ^ n353 ^ n314 ;
  assign n1719 = x95 & x96 ;
  assign n1721 = n1720 ^ n1719 ^ 1'b0 ;
  assign n1722 = n431 ^ x6 ^ 1'b0 ;
  assign n1723 = ~n1172 & n1722 ;
  assign n1724 = ~n1208 & n1723 ;
  assign n1725 = ~n990 & n1724 ;
  assign n1726 = ( x148 & n946 ) | ( x148 & n1725 ) | ( n946 & n1725 ) ;
  assign n1727 = n1217 | n1345 ;
  assign n1728 = x24 & ~x242 ;
  assign n1729 = n1034 & ~n1728 ;
  assign n1730 = n1190 & n1626 ;
  assign n1731 = ~n893 & n1474 ;
  assign n1732 = x52 & x108 ;
  assign n1733 = ~x219 & n1732 ;
  assign n1734 = x174 ^ x108 ^ 1'b0 ;
  assign n1735 = ~n1120 & n1734 ;
  assign n1736 = ( n682 & n1649 ) | ( n682 & n1735 ) | ( n1649 & n1735 ) ;
  assign n1737 = ( ~n479 & n893 ) | ( ~n479 & n1577 ) | ( n893 & n1577 ) ;
  assign n1738 = n1225 & ~n1737 ;
  assign n1739 = n1172 ^ n1069 ^ 1'b0 ;
  assign n1740 = n1738 & ~n1739 ;
  assign n1741 = ~n1456 & n1740 ;
  assign n1742 = n931 & n953 ;
  assign n1743 = x107 & n394 ;
  assign n1744 = n1743 ^ n325 ^ 1'b0 ;
  assign n1745 = n1322 ^ x253 ^ 1'b0 ;
  assign n1746 = ~n665 & n1745 ;
  assign n1747 = n1230 ^ n953 ^ 1'b0 ;
  assign n1748 = n1623 & ~n1747 ;
  assign n1749 = n877 ^ n682 ^ 1'b0 ;
  assign n1752 = ~x17 & x187 ;
  assign n1750 = n491 | n558 ;
  assign n1751 = x231 & ~n1750 ;
  assign n1753 = n1752 ^ n1751 ^ 1'b0 ;
  assign n1754 = n409 & ~n433 ;
  assign n1755 = n1754 ^ n882 ^ 1'b0 ;
  assign n1756 = ~n1362 & n1755 ;
  assign n1757 = ( n589 & ~n603 ) | ( n589 & n1726 ) | ( ~n603 & n1726 ) ;
  assign n1758 = n949 ^ n334 ^ 1'b0 ;
  assign n1759 = x12 & n1758 ;
  assign n1760 = n1105 ^ n355 ^ 1'b0 ;
  assign n1761 = x12 & x213 ;
  assign n1762 = ~n271 & n1761 ;
  assign n1763 = ( ~x150 & x170 ) | ( ~x150 & n1343 ) | ( x170 & n1343 ) ;
  assign n1764 = x251 & ~n599 ;
  assign n1765 = n1764 ^ n619 ^ 1'b0 ;
  assign n1766 = n1765 ^ n419 ^ n413 ;
  assign n1767 = n727 | n1766 ;
  assign n1768 = n1763 | n1767 ;
  assign n1769 = n1768 ^ n529 ^ 1'b0 ;
  assign n1770 = n907 & n1769 ;
  assign n1771 = ~n1762 & n1770 ;
  assign n1772 = n1771 ^ n671 ^ 1'b0 ;
  assign n1773 = n682 | n1671 ;
  assign n1774 = x107 | n1773 ;
  assign n1775 = x48 & ~n1774 ;
  assign n1776 = n391 & n1775 ;
  assign n1777 = n1776 ^ n1465 ^ 1'b0 ;
  assign n1778 = x236 & ~n872 ;
  assign n1779 = x115 & ~n1778 ;
  assign n1780 = n1779 ^ x211 ^ 1'b0 ;
  assign n1781 = x146 & ~n819 ;
  assign n1782 = ~n808 & n1781 ;
  assign n1783 = n1468 | n1782 ;
  assign n1784 = n1783 ^ n920 ^ 1'b0 ;
  assign n1788 = x97 & x116 ;
  assign n1785 = x3 & ~n880 ;
  assign n1786 = n1785 ^ n1132 ^ 1'b0 ;
  assign n1787 = x223 & ~n1786 ;
  assign n1789 = n1788 ^ n1787 ^ 1'b0 ;
  assign n1790 = x182 & ~n908 ;
  assign n1791 = n1200 & n1790 ;
  assign n1792 = n672 ^ n367 ^ 1'b0 ;
  assign n1793 = n1784 & n1792 ;
  assign n1794 = n804 | n1100 ;
  assign n1795 = n1410 | n1794 ;
  assign n1796 = n556 & n1795 ;
  assign n1797 = n1667 ^ n1603 ^ 1'b0 ;
  assign n1798 = x160 & ~n1797 ;
  assign n1799 = x179 & n457 ;
  assign n1800 = n1045 & n1799 ;
  assign n1801 = n419 & n1800 ;
  assign n1803 = n1345 ^ n900 ^ x80 ;
  assign n1804 = n737 & ~n1803 ;
  assign n1802 = n1632 ^ x218 ^ 1'b0 ;
  assign n1805 = n1804 ^ n1802 ^ 1'b0 ;
  assign n1806 = n604 ^ x221 ^ 1'b0 ;
  assign n1807 = ~n1805 & n1806 ;
  assign n1808 = x91 & ~n462 ;
  assign n1809 = ~n1001 & n1808 ;
  assign n1810 = x174 | n1016 ;
  assign n1811 = x104 & ~n603 ;
  assign n1812 = ~x231 & n1811 ;
  assign n1813 = n772 & ~n959 ;
  assign n1814 = ~n1812 & n1813 ;
  assign n1816 = n848 ^ n281 ^ 1'b0 ;
  assign n1817 = n419 | n1816 ;
  assign n1818 = n1817 ^ n747 ^ 1'b0 ;
  assign n1819 = x250 & ~n1818 ;
  assign n1815 = ( x6 & n1160 ) | ( x6 & ~n1445 ) | ( n1160 & ~n1445 ) ;
  assign n1820 = n1819 ^ n1815 ^ x88 ;
  assign n1821 = n763 ^ n462 ^ 1'b0 ;
  assign n1822 = x27 & ~n1821 ;
  assign n1823 = n548 ^ x11 ^ 1'b0 ;
  assign n1824 = n1651 | n1823 ;
  assign n1825 = n615 | n1824 ;
  assign n1826 = n695 & ~n1825 ;
  assign n1827 = x44 & n351 ;
  assign n1828 = n1827 ^ n331 ^ 1'b0 ;
  assign n1830 = ~x141 & n917 ;
  assign n1829 = n1307 ^ x4 ^ 1'b0 ;
  assign n1831 = n1830 ^ n1829 ^ 1'b0 ;
  assign n1832 = n1828 & n1831 ;
  assign n1833 = ( x172 & ~n537 ) | ( x172 & n1042 ) | ( ~n537 & n1042 ) ;
  assign n1834 = x181 & ~n511 ;
  assign n1835 = n498 & n1834 ;
  assign n1836 = x125 & ~n1835 ;
  assign n1837 = n1836 ^ x143 ^ 1'b0 ;
  assign n1838 = n1837 ^ n882 ^ n327 ;
  assign n1839 = n1838 ^ n992 ^ 1'b0 ;
  assign n1840 = n1839 ^ x171 ^ 1'b0 ;
  assign n1841 = n1833 & n1840 ;
  assign n1842 = n1193 ^ n1169 ^ 1'b0 ;
  assign n1843 = n1841 & ~n1842 ;
  assign n1844 = n1777 ^ x182 ^ 1'b0 ;
  assign n1845 = n889 ^ n440 ^ 1'b0 ;
  assign n1846 = n1473 ^ n389 ^ 1'b0 ;
  assign n1847 = ~n771 & n1534 ;
  assign n1848 = n1847 ^ x163 ^ 1'b0 ;
  assign n1849 = n1674 ^ n778 ^ 1'b0 ;
  assign n1850 = x6 & n1849 ;
  assign n1851 = n764 ^ x254 ^ 1'b0 ;
  assign n1852 = n511 ^ x169 ^ 1'b0 ;
  assign n1853 = n1851 | n1852 ;
  assign n1854 = n1602 & ~n1853 ;
  assign n1855 = n464 ^ x183 ^ 1'b0 ;
  assign n1856 = n448 | n1855 ;
  assign n1857 = ~n1219 & n1856 ;
  assign n1858 = ~n1854 & n1857 ;
  assign n1859 = n1850 & n1858 ;
  assign n1860 = n1105 ^ n637 ^ 1'b0 ;
  assign n1861 = n1859 & n1860 ;
  assign n1862 = n1478 ^ n1148 ^ 1'b0 ;
  assign n1863 = ~n891 & n1148 ;
  assign n1864 = n430 & n1863 ;
  assign n1865 = n860 & ~n1864 ;
  assign n1866 = n1865 ^ n314 ^ 1'b0 ;
  assign n1867 = n1433 ^ n810 ^ x94 ;
  assign n1868 = n1153 | n1867 ;
  assign n1869 = n1868 ^ n1835 ^ 1'b0 ;
  assign n1870 = ~n953 & n1869 ;
  assign n1871 = n625 ^ n593 ^ 1'b0 ;
  assign n1872 = n1148 & ~n1641 ;
  assign n1873 = n1871 & n1872 ;
  assign n1874 = n577 ^ n516 ^ 1'b0 ;
  assign n1875 = n1874 ^ n1157 ^ 1'b0 ;
  assign n1876 = n1409 ^ n1089 ^ 1'b0 ;
  assign n1877 = n1116 | n1876 ;
  assign n1878 = n558 & n1374 ;
  assign n1879 = n387 | n1869 ;
  assign n1880 = n1269 ^ x125 ^ 1'b0 ;
  assign n1881 = n708 & n713 ;
  assign n1882 = ~n1880 & n1881 ;
  assign n1883 = x132 & ~n994 ;
  assign n1884 = n1882 & n1883 ;
  assign n1885 = n1884 ^ n1698 ^ n1261 ;
  assign n1886 = n774 | n1057 ;
  assign n1887 = n486 | n1886 ;
  assign n1888 = n1887 ^ n863 ^ 1'b0 ;
  assign n1889 = n581 & ~n1888 ;
  assign n1890 = ( x184 & ~n477 ) | ( x184 & n1614 ) | ( ~n477 & n1614 ) ;
  assign n1891 = n1195 & ~n1890 ;
  assign n1892 = n1627 ^ n604 ^ 1'b0 ;
  assign n1893 = n1064 & n1892 ;
  assign n1894 = x53 | n1250 ;
  assign n1895 = n1628 | n1664 ;
  assign n1896 = n1895 ^ x80 ^ 1'b0 ;
  assign n1897 = n431 & ~n1084 ;
  assign n1898 = ~n325 & n1897 ;
  assign n1899 = ( x22 & n579 ) | ( x22 & n1539 ) | ( n579 & n1539 ) ;
  assign n1900 = n1899 ^ x202 ^ 1'b0 ;
  assign n1901 = x132 ^ x115 ^ 1'b0 ;
  assign n1908 = n1595 | n1762 ;
  assign n1909 = n1908 ^ n323 ^ 1'b0 ;
  assign n1902 = ~n329 & n613 ;
  assign n1903 = n1902 ^ n1649 ^ 1'b0 ;
  assign n1904 = n404 & ~n823 ;
  assign n1905 = ~n1343 & n1904 ;
  assign n1906 = n1905 ^ n1558 ^ 1'b0 ;
  assign n1907 = n1903 & n1906 ;
  assign n1910 = n1909 ^ n1907 ^ 1'b0 ;
  assign n1911 = n1910 ^ n318 ^ 1'b0 ;
  assign n1912 = n624 ^ x130 ^ 1'b0 ;
  assign n1913 = n581 | n1912 ;
  assign n1914 = n1913 ^ x32 ^ 1'b0 ;
  assign n1915 = x228 & n1548 ;
  assign n1916 = n1914 & n1915 ;
  assign n1917 = ~n729 & n1916 ;
  assign n1918 = x148 & ~n347 ;
  assign n1919 = n1918 ^ n787 ^ 1'b0 ;
  assign n1920 = n1919 ^ n1342 ^ 1'b0 ;
  assign n1921 = n1682 & ~n1920 ;
  assign n1922 = n1312 ^ n1011 ^ 1'b0 ;
  assign n1923 = n1922 ^ n963 ^ 1'b0 ;
  assign n1924 = x210 & ~n1923 ;
  assign n1925 = ~x39 & n1924 ;
  assign n1926 = n1921 & n1925 ;
  assign n1927 = n838 & n1126 ;
  assign n1928 = n1927 ^ x254 ^ 1'b0 ;
  assign n1929 = n276 & ~n1928 ;
  assign n1930 = n727 | n1443 ;
  assign n1931 = n1930 ^ n372 ^ 1'b0 ;
  assign n1932 = n1042 | n1931 ;
  assign n1933 = n1932 ^ n272 ^ 1'b0 ;
  assign n1934 = n1345 ^ x51 ^ 1'b0 ;
  assign n1935 = n1048 & ~n1934 ;
  assign n1936 = ~n406 & n1935 ;
  assign n1942 = n1903 ^ n874 ^ 1'b0 ;
  assign n1943 = n1880 & ~n1942 ;
  assign n1937 = n1144 ^ n794 ^ 1'b0 ;
  assign n1938 = x225 & n1178 ;
  assign n1939 = n1938 ^ n1850 ^ 1'b0 ;
  assign n1940 = n1937 | n1939 ;
  assign n1941 = n491 | n1940 ;
  assign n1944 = n1943 ^ n1941 ^ 1'b0 ;
  assign n1945 = n1042 ^ x180 ^ 1'b0 ;
  assign n1946 = n1945 ^ n1622 ^ 1'b0 ;
  assign n1947 = n1851 & n1946 ;
  assign n1948 = n1538 ^ x248 ^ 1'b0 ;
  assign n1949 = x21 & ~n571 ;
  assign n1950 = n1378 & n1949 ;
  assign n1951 = x94 & ~n334 ;
  assign n1952 = n682 & n1951 ;
  assign n1953 = n547 | n1952 ;
  assign n1954 = n1369 & ~n1953 ;
  assign n1962 = ( n789 & n810 ) | ( n789 & ~n1443 ) | ( n810 & ~n1443 ) ;
  assign n1963 = n949 ^ x176 ^ 1'b0 ;
  assign n1964 = ( ~n1126 & n1962 ) | ( ~n1126 & n1963 ) | ( n1962 & n1963 ) ;
  assign n1959 = ~n668 & n1610 ;
  assign n1960 = ~n933 & n1959 ;
  assign n1955 = n1786 ^ n869 ^ 1'b0 ;
  assign n1956 = x72 & ~n1955 ;
  assign n1957 = n742 ^ x85 ^ 1'b0 ;
  assign n1958 = n1956 & n1957 ;
  assign n1961 = n1960 ^ n1958 ^ 1'b0 ;
  assign n1965 = n1964 ^ n1961 ^ n357 ;
  assign n1966 = n1893 ^ n723 ^ 1'b0 ;
  assign n1967 = ~n651 & n966 ;
  assign n1968 = n1967 ^ x129 ^ 1'b0 ;
  assign n1969 = ~x98 & n375 ;
  assign n1970 = n1969 ^ n520 ^ 1'b0 ;
  assign n1971 = ~n1968 & n1970 ;
  assign n1972 = n467 & n737 ;
  assign n1973 = ~n409 & n1972 ;
  assign n1974 = x117 & ~n314 ;
  assign n1975 = n1974 ^ n382 ^ 1'b0 ;
  assign n1976 = n1975 ^ x44 ^ 1'b0 ;
  assign n1977 = x17 & n1976 ;
  assign n1978 = n1977 ^ n722 ^ 1'b0 ;
  assign n1979 = ~n1973 & n1978 ;
  assign n1980 = n1979 ^ n1975 ^ 1'b0 ;
  assign n1981 = ~n935 & n982 ;
  assign n1982 = ( x100 & n1352 ) | ( x100 & ~n1981 ) | ( n1352 & ~n1981 ) ;
  assign n1983 = n1982 ^ n473 ^ x6 ;
  assign n1984 = ~n440 & n891 ;
  assign n1985 = n1984 ^ x175 ^ 1'b0 ;
  assign n1986 = n1008 ^ n970 ^ 1'b0 ;
  assign n1988 = n315 | n882 ;
  assign n1989 = n1988 ^ x72 ^ 1'b0 ;
  assign n1987 = x93 & n1129 ;
  assign n1990 = n1989 ^ n1987 ^ 1'b0 ;
  assign n1991 = ~n312 & n1975 ;
  assign n1992 = ~x232 & n1991 ;
  assign n1993 = n1245 & ~n1992 ;
  assign n1994 = n880 & n1146 ;
  assign n1995 = ( ~n668 & n1993 ) | ( ~n668 & n1994 ) | ( n1993 & n1994 ) ;
  assign n1996 = x33 & x60 ;
  assign n1997 = n1996 ^ x96 ^ 1'b0 ;
  assign n1998 = n1606 & n1997 ;
  assign n1999 = n1962 ^ n689 ^ 1'b0 ;
  assign n2000 = n973 | n1999 ;
  assign n2001 = n1514 & ~n2000 ;
  assign n2002 = n1341 | n1729 ;
  assign n2003 = n2002 ^ n1950 ^ 1'b0 ;
  assign n2004 = n1589 ^ n724 ^ 1'b0 ;
  assign n2005 = n896 ^ x206 ^ 1'b0 ;
  assign n2006 = n2004 & n2005 ;
  assign n2007 = n799 & n1144 ;
  assign n2012 = x149 & ~n1445 ;
  assign n2013 = ~n1711 & n2012 ;
  assign n2008 = n718 & n751 ;
  assign n2009 = n708 & n2008 ;
  assign n2010 = n2009 ^ n1124 ^ 1'b0 ;
  assign n2011 = n1913 & n2010 ;
  assign n2014 = n2013 ^ n2011 ^ 1'b0 ;
  assign n2015 = n444 ^ n402 ^ 1'b0 ;
  assign n2016 = n387 ^ x18 ^ 1'b0 ;
  assign n2017 = x200 & n2016 ;
  assign n2018 = n475 & n2017 ;
  assign n2019 = x47 & x143 ;
  assign n2020 = n2019 ^ x118 ^ 1'b0 ;
  assign n2021 = x123 & ~n2020 ;
  assign n2022 = n1577 & n2021 ;
  assign n2023 = n1495 & n2022 ;
  assign n2024 = n1725 | n2023 ;
  assign n2027 = n545 ^ x40 ^ x35 ;
  assign n2028 = n1577 ^ x202 ^ 1'b0 ;
  assign n2029 = n2027 | n2028 ;
  assign n2025 = x96 & n1606 ;
  assign n2026 = n552 & n2025 ;
  assign n2030 = n2029 ^ n2026 ^ 1'b0 ;
  assign n2036 = x102 ^ x44 ^ 1'b0 ;
  assign n2037 = x26 & n2036 ;
  assign n2038 = n1085 & n2037 ;
  assign n2039 = n2038 ^ x166 ^ 1'b0 ;
  assign n2040 = ( n957 & n1433 ) | ( n957 & ~n2039 ) | ( n1433 & ~n2039 ) ;
  assign n2031 = n1453 & ~n1960 ;
  assign n2032 = n2031 ^ n1011 ^ 1'b0 ;
  assign n2033 = n776 | n2032 ;
  assign n2034 = n2033 ^ n651 ^ 1'b0 ;
  assign n2035 = n2034 ^ n1527 ^ 1'b0 ;
  assign n2041 = n2040 ^ n2035 ^ 1'b0 ;
  assign n2042 = n1966 ^ n1153 ^ 1'b0 ;
  assign n2043 = x180 & ~n2042 ;
  assign n2044 = x129 & n1045 ;
  assign n2045 = n2044 ^ n1867 ^ 1'b0 ;
  assign n2046 = x192 & x193 ;
  assign n2047 = n1051 & n2046 ;
  assign n2048 = n1662 & ~n2047 ;
  assign n2049 = x131 & n1723 ;
  assign n2050 = ( x124 & ~n1989 ) | ( x124 & n2049 ) | ( ~n1989 & n2049 ) ;
  assign n2051 = n937 ^ n365 ^ 1'b0 ;
  assign n2052 = ~n1575 & n2051 ;
  assign n2053 = n2052 ^ n283 ^ 1'b0 ;
  assign n2054 = n1474 & n1662 ;
  assign n2055 = x129 | n1219 ;
  assign n2056 = n287 & n492 ;
  assign n2057 = n2055 & n2056 ;
  assign n2058 = ~n2016 & n2057 ;
  assign n2059 = n511 | n635 ;
  assign n2060 = n1766 & ~n2059 ;
  assign n2061 = n2060 ^ n1288 ^ 1'b0 ;
  assign n2062 = n380 | n2061 ;
  assign n2063 = ~n577 & n819 ;
  assign n2064 = n2063 ^ n1579 ^ 1'b0 ;
  assign n2065 = n839 | n1647 ;
  assign n2066 = n943 | n1426 ;
  assign n2067 = n366 | n2066 ;
  assign n2068 = n1981 ^ n1963 ^ 1'b0 ;
  assign n2069 = n2067 & ~n2068 ;
  assign n2070 = x94 & ~x200 ;
  assign n2071 = n1456 & n1975 ;
  assign n2072 = n2071 ^ n659 ^ 1'b0 ;
  assign n2073 = n899 ^ x76 ^ 1'b0 ;
  assign n2074 = n632 & n2073 ;
  assign n2075 = n2074 ^ n1373 ^ 1'b0 ;
  assign n2076 = n1134 & n2075 ;
  assign n2077 = ~x218 & n2076 ;
  assign n2078 = n1583 | n2077 ;
  assign n2080 = n1505 ^ n1149 ^ x163 ;
  assign n2079 = x20 & ~n274 ;
  assign n2081 = n2080 ^ n2079 ^ 1'b0 ;
  assign n2082 = n984 & n2081 ;
  assign n2083 = n283 & ~n682 ;
  assign n2084 = x88 & ~n716 ;
  assign n2085 = n980 & n2084 ;
  assign n2086 = n916 ^ x113 ^ 1'b0 ;
  assign n2087 = n2086 ^ n835 ^ 1'b0 ;
  assign n2088 = ~n462 & n2087 ;
  assign n2089 = n2088 ^ n1665 ^ 1'b0 ;
  assign n2090 = n2089 ^ x178 ^ 1'b0 ;
  assign n2091 = ~n2085 & n2090 ;
  assign n2092 = n1064 ^ n957 ^ x115 ;
  assign n2093 = n2092 ^ n1900 ^ n1172 ;
  assign n2094 = n1912 ^ x6 ^ 1'b0 ;
  assign n2095 = n919 | n2094 ;
  assign n2096 = n1876 ^ x163 ^ 1'b0 ;
  assign n2097 = n2096 ^ n571 ^ 1'b0 ;
  assign n2098 = n2095 & ~n2097 ;
  assign n2099 = ~n500 & n746 ;
  assign n2100 = x84 & ~n2099 ;
  assign n2101 = ~n1615 & n2100 ;
  assign n2102 = n359 & n558 ;
  assign n2103 = ~x176 & n1643 ;
  assign n2104 = n1919 ^ n444 ^ x154 ;
  assign n2105 = ~n331 & n2104 ;
  assign n2106 = n589 ^ n312 ^ 1'b0 ;
  assign n2107 = n2106 ^ n1986 ^ n1349 ;
  assign n2108 = x134 | n1019 ;
  assign n2109 = n2108 ^ x25 ^ 1'b0 ;
  assign n2110 = n937 & n2109 ;
  assign n2111 = x17 & ~n346 ;
  assign n2112 = ~n1160 & n2111 ;
  assign n2113 = n725 ^ x12 ^ 1'b0 ;
  assign n2114 = x154 | n1081 ;
  assign n2115 = n267 | n1998 ;
  assign n2116 = n2115 ^ n395 ^ 1'b0 ;
  assign n2117 = x109 ^ x21 ^ 1'b0 ;
  assign n2118 = n1345 ^ n755 ^ 1'b0 ;
  assign n2119 = n2117 & n2118 ;
  assign n2120 = n2119 ^ x229 ^ 1'b0 ;
  assign n2121 = n1345 ^ n281 ^ 1'b0 ;
  assign n2122 = n2120 | n2121 ;
  assign n2123 = n2122 ^ n1107 ^ 1'b0 ;
  assign n2132 = n1782 ^ n970 ^ 1'b0 ;
  assign n2133 = n1606 & ~n2132 ;
  assign n2130 = n1307 ^ x185 ^ x3 ;
  assign n2124 = x130 & n1089 ;
  assign n2125 = n879 & n2124 ;
  assign n2126 = n1011 & ~n2125 ;
  assign n2127 = n274 & n2126 ;
  assign n2128 = n1297 & ~n1495 ;
  assign n2129 = ~n2127 & n2128 ;
  assign n2131 = n2130 ^ n2129 ^ 1'b0 ;
  assign n2134 = n2133 ^ n2131 ^ 1'b0 ;
  assign n2135 = n1354 | n2134 ;
  assign n2136 = x225 & ~n2135 ;
  assign n2137 = n2136 ^ n1909 ^ 1'b0 ;
  assign n2138 = n699 ^ n575 ^ 1'b0 ;
  assign n2139 = n542 | n2138 ;
  assign n2140 = n2139 ^ x27 ^ 1'b0 ;
  assign n2141 = n395 | n2140 ;
  assign n2142 = n359 & n932 ;
  assign n2143 = ( n530 & n986 ) | ( n530 & n1447 ) | ( n986 & n1447 ) ;
  assign n2144 = n1913 ^ n1797 ^ n1193 ;
  assign n2145 = x16 & ~n2144 ;
  assign n2146 = n2145 ^ n809 ^ 1'b0 ;
  assign n2147 = n862 & ~n1279 ;
  assign n2148 = n2147 ^ n461 ^ 1'b0 ;
  assign n2149 = n826 & ~n2148 ;
  assign n2152 = x106 & n1815 ;
  assign n2153 = n1690 & n2152 ;
  assign n2150 = n1632 ^ n986 ^ n589 ;
  assign n2151 = ~n1864 & n2150 ;
  assign n2154 = n2153 ^ n2151 ^ 1'b0 ;
  assign n2155 = n1756 & n2154 ;
  assign n2156 = n1328 ^ n592 ^ 1'b0 ;
  assign n2157 = n838 & ~n2156 ;
  assign n2158 = ~x116 & n1174 ;
  assign n2159 = n2157 | n2158 ;
  assign n2160 = x95 & ~n505 ;
  assign n2161 = ~n1765 & n2160 ;
  assign n2162 = n1180 & n2161 ;
  assign n2163 = n2162 ^ n943 ^ 1'b0 ;
  assign n2164 = n2163 ^ n1850 ^ 1'b0 ;
  assign n2165 = ~x223 & n1513 ;
  assign n2166 = n389 | n2165 ;
  assign n2167 = n1338 | n2166 ;
  assign n2168 = n322 | n627 ;
  assign n2169 = n643 & ~n2168 ;
  assign n2170 = ( x232 & ~n434 ) | ( x232 & n2169 ) | ( ~n434 & n2169 ) ;
  assign n2171 = x228 | n2170 ;
  assign n2172 = n1680 ^ n1272 ^ 1'b0 ;
  assign n2174 = x250 & ~n1788 ;
  assign n2175 = n1417 & n2174 ;
  assign n2176 = ~n293 & n2175 ;
  assign n2177 = x175 | n2176 ;
  assign n2173 = n825 | n880 ;
  assign n2178 = n2177 ^ n2173 ^ 1'b0 ;
  assign n2179 = n771 ^ n705 ^ 1'b0 ;
  assign n2180 = n1111 & ~n2179 ;
  assign n2181 = n2180 ^ x26 ^ 1'b0 ;
  assign n2182 = ~n574 & n2181 ;
  assign n2183 = n2182 ^ n1803 ^ 1'b0 ;
  assign n2184 = n2183 ^ n789 ^ 1'b0 ;
  assign n2186 = x88 & n1129 ;
  assign n2187 = n2186 ^ n1094 ^ 1'b0 ;
  assign n2188 = n1059 & n1170 ;
  assign n2189 = x32 & ~n2188 ;
  assign n2190 = ( n1249 & ~n2187 ) | ( n1249 & n2189 ) | ( ~n2187 & n2189 ) ;
  assign n2185 = n281 | n627 ;
  assign n2191 = n2190 ^ n2185 ^ 1'b0 ;
  assign n2192 = n1424 ^ n996 ^ 1'b0 ;
  assign n2193 = n737 & ~n2192 ;
  assign n2194 = x144 ^ x83 ^ 1'b0 ;
  assign n2195 = n387 & ~n2194 ;
  assign n2196 = n853 & n2195 ;
  assign n2197 = n925 & ~n2196 ;
  assign n2198 = n2197 ^ n2034 ^ 1'b0 ;
  assign n2199 = n1377 ^ n789 ^ 1'b0 ;
  assign n2200 = n2099 ^ n1391 ^ 1'b0 ;
  assign n2201 = ~n776 & n1523 ;
  assign n2202 = ~n794 & n2201 ;
  assign n2203 = n1347 & ~n2202 ;
  assign n2208 = ( x10 & ~x117 ) | ( x10 & x207 ) | ( ~x117 & x207 ) ;
  assign n2209 = n2208 ^ n831 ^ n675 ;
  assign n2210 = n831 & ~n1193 ;
  assign n2211 = n357 & n2210 ;
  assign n2212 = n402 & n2211 ;
  assign n2213 = n2209 & n2212 ;
  assign n2204 = ( ~x176 & n492 ) | ( ~x176 & n966 ) | ( n492 & n966 ) ;
  assign n2205 = n614 ^ n369 ^ 1'b0 ;
  assign n2206 = n806 & n2205 ;
  assign n2207 = n2204 & n2206 ;
  assign n2214 = n2213 ^ n2207 ^ 1'b0 ;
  assign n2215 = n312 | n1929 ;
  assign n2216 = x162 | n1961 ;
  assign n2217 = x214 & ~n312 ;
  assign n2218 = ~x158 & n2217 ;
  assign n2219 = n2218 ^ n801 ^ 1'b0 ;
  assign n2220 = n2172 & n2219 ;
  assign n2221 = n1381 & n2220 ;
  assign n2222 = n2208 ^ n766 ^ 1'b0 ;
  assign n2223 = n442 | n2222 ;
  assign n2224 = n424 & ~n2223 ;
  assign n2225 = n920 & n1312 ;
  assign n2226 = n1027 & n1405 ;
  assign n2227 = n1647 ^ x166 ^ 1'b0 ;
  assign n2228 = x31 & n466 ;
  assign n2229 = x108 ^ x94 ^ x3 ;
  assign n2230 = n2229 ^ n466 ^ n333 ;
  assign n2231 = n1893 & ~n2230 ;
  assign n2232 = ~n587 & n1014 ;
  assign n2233 = x75 & n2232 ;
  assign n2234 = n2233 ^ x198 ^ 1'b0 ;
  assign n2235 = n2234 ^ n1278 ^ 1'b0 ;
  assign n2236 = x247 & ~n2235 ;
  assign n2237 = ~x30 & n2236 ;
  assign n2238 = ~x195 & n1833 ;
  assign n2239 = n2238 ^ n500 ^ 1'b0 ;
  assign n2240 = x190 & n2239 ;
  assign n2241 = n402 & n2240 ;
  assign n2242 = ~n1956 & n2241 ;
  assign n2243 = n1397 & n1716 ;
  assign n2244 = n291 & n1723 ;
  assign n2245 = n1613 & ~n1882 ;
  assign n2246 = x206 ^ x125 ^ x102 ;
  assign n2247 = n2246 ^ n1219 ^ 1'b0 ;
  assign n2248 = n2247 ^ n635 ^ 1'b0 ;
  assign n2249 = n1428 & ~n2248 ;
  assign n2250 = n733 ^ x218 ^ 1'b0 ;
  assign n2251 = x171 & n2232 ;
  assign n2252 = n603 & n2251 ;
  assign n2253 = n732 & ~n2252 ;
  assign n2254 = ~n789 & n2253 ;
  assign n2255 = n2250 & ~n2254 ;
  assign n2256 = n1060 & n2255 ;
  assign n2257 = n1998 ^ n1215 ^ 1'b0 ;
  assign n2258 = n464 & n1622 ;
  assign n2259 = n2242 ^ n1926 ^ x252 ;
  assign n2260 = ( n406 & n842 ) | ( n406 & n1931 ) | ( n842 & n1931 ) ;
  assign n2261 = n2260 ^ n1539 ^ 1'b0 ;
  assign n2262 = x247 & n2261 ;
  assign n2263 = n2262 ^ n1039 ^ 1'b0 ;
  assign n2264 = n1477 ^ n466 ^ x60 ;
  assign n2265 = n1189 & ~n2218 ;
  assign n2267 = n1963 ^ n1182 ^ x112 ;
  assign n2266 = ~n1378 & n1945 ;
  assign n2268 = n2267 ^ n2266 ^ 1'b0 ;
  assign n2269 = x143 & n1124 ;
  assign n2270 = ~n2229 & n2269 ;
  assign n2271 = n411 & n2270 ;
  assign n2272 = n2039 ^ n1619 ^ 1'b0 ;
  assign n2273 = n2271 | n2272 ;
  assign n2274 = n2273 ^ n1148 ^ 1'b0 ;
  assign n2275 = n2274 ^ x251 ^ 1'b0 ;
  assign n2276 = ( x107 & x250 ) | ( x107 & n1037 ) | ( x250 & n1037 ) ;
  assign n2277 = n1786 ^ n1592 ^ 1'b0 ;
  assign n2278 = n395 & n518 ;
  assign n2279 = n1695 & n2278 ;
  assign n2280 = x165 & n732 ;
  assign n2281 = n2280 ^ n925 ^ 1'b0 ;
  assign n2282 = n697 | n2073 ;
  assign n2283 = ( ~n415 & n581 ) | ( ~n415 & n2282 ) | ( n581 & n2282 ) ;
  assign n2284 = x132 & n694 ;
  assign n2285 = ~n444 & n2284 ;
  assign n2286 = ~x0 & n2285 ;
  assign n2287 = x136 & n385 ;
  assign n2288 = n847 & n2287 ;
  assign n2289 = ~n1788 & n2288 ;
  assign n2290 = x247 & ~n411 ;
  assign n2291 = ~n1170 & n2290 ;
  assign n2292 = n2291 ^ n1351 ^ 1'b0 ;
  assign n2293 = x189 & n2292 ;
  assign n2294 = x232 & n891 ;
  assign n2295 = n1635 & n2294 ;
  assign n2296 = ~n2293 & n2295 ;
  assign n2297 = n1651 ^ n970 ^ 1'b0 ;
  assign n2298 = n2296 | n2297 ;
  assign n2299 = n466 | n2298 ;
  assign n2300 = n325 & ~n941 ;
  assign n2301 = ~x65 & n2300 ;
  assign n2302 = n1950 ^ n1577 ^ 1'b0 ;
  assign n2303 = n268 & n707 ;
  assign n2304 = n765 & n2303 ;
  assign n2307 = n281 ^ x234 ^ x73 ;
  assign n2305 = n1599 ^ x150 ^ 1'b0 ;
  assign n2306 = n2305 ^ n1552 ^ n722 ;
  assign n2308 = n2307 ^ n2306 ^ 1'b0 ;
  assign n2309 = ( n2282 & n2304 ) | ( n2282 & n2308 ) | ( n2304 & n2308 ) ;
  assign n2310 = n1467 | n2194 ;
  assign n2311 = ~n1306 & n1932 ;
  assign n2312 = n579 & ~n764 ;
  assign n2313 = n1356 ^ x72 ^ 1'b0 ;
  assign n2314 = ~n481 & n2313 ;
  assign n2315 = n2312 & n2314 ;
  assign n2316 = n2311 & n2315 ;
  assign n2317 = n2133 ^ n1002 ^ n914 ;
  assign n2318 = n1746 ^ n1338 ^ 1'b0 ;
  assign n2319 = n325 & n2318 ;
  assign n2320 = ( x67 & n651 ) | ( x67 & n2319 ) | ( n651 & n2319 ) ;
  assign n2321 = n1639 ^ x149 ^ 1'b0 ;
  assign n2322 = n2161 | n2321 ;
  assign n2323 = n1002 | n1775 ;
  assign n2324 = x181 & n2120 ;
  assign n2325 = n2324 ^ n1193 ^ 1'b0 ;
  assign n2326 = n1379 & n1494 ;
  assign n2327 = n1583 ^ n742 ^ 1'b0 ;
  assign n2328 = n2326 & ~n2327 ;
  assign n2329 = n863 & n1333 ;
  assign n2330 = n819 & n2329 ;
  assign n2331 = n274 ^ x58 ^ 1'b0 ;
  assign n2332 = n2331 ^ n769 ^ 1'b0 ;
  assign n2333 = n2332 ^ n1341 ^ 1'b0 ;
  assign n2334 = n1240 & ~n2333 ;
  assign n2335 = n2334 ^ n1718 ^ 1'b0 ;
  assign n2338 = n376 | n442 ;
  assign n2339 = n2338 ^ n1174 ^ 1'b0 ;
  assign n2340 = n1496 & ~n2339 ;
  assign n2336 = n627 | n699 ;
  assign n2337 = n2336 ^ n2218 ^ 1'b0 ;
  assign n2341 = n2340 ^ n2337 ^ 1'b0 ;
  assign n2342 = x39 & x184 ;
  assign n2343 = ~n2341 & n2342 ;
  assign n2344 = x162 & n262 ;
  assign n2345 = n2344 ^ n904 ^ 1'b0 ;
  assign n2346 = n883 | n1232 ;
  assign n2347 = n759 | n2346 ;
  assign n2348 = ~n677 & n986 ;
  assign n2349 = n485 | n1132 ;
  assign n2350 = n1862 & n2349 ;
  assign n2351 = n2272 & n2350 ;
  assign n2352 = n399 | n1912 ;
  assign n2353 = n2352 ^ x175 ^ 1'b0 ;
  assign n2354 = n1385 & n1413 ;
  assign n2355 = ( n466 & n2353 ) | ( n466 & n2354 ) | ( n2353 & n2354 ) ;
  assign n2356 = n863 | n1249 ;
  assign n2357 = n799 & ~n2356 ;
  assign n2358 = n2070 ^ n932 ^ 1'b0 ;
  assign n2359 = x26 & x119 ;
  assign n2360 = n2359 ^ n1728 ^ 1'b0 ;
  assign n2361 = ~n1416 & n2360 ;
  assign n2362 = n738 & ~n2361 ;
  assign n2364 = x186 & n749 ;
  assign n2365 = n2364 ^ x231 ^ 1'b0 ;
  assign n2363 = ~n611 & n2048 ;
  assign n2366 = n2365 ^ n2363 ^ 1'b0 ;
  assign n2367 = n2282 & ~n2366 ;
  assign n2368 = x76 & n479 ;
  assign n2369 = n2367 ^ n2307 ^ 1'b0 ;
  assign n2370 = n1124 ^ x178 ^ 1'b0 ;
  assign n2371 = n1219 ^ n982 ^ 1'b0 ;
  assign n2372 = ~x77 & n2015 ;
  assign n2373 = n1254 & n1459 ;
  assign n2374 = n1016 & n2373 ;
  assign n2375 = n2011 ^ x169 ^ 1'b0 ;
  assign n2376 = n2135 ^ n1680 ^ 1'b0 ;
  assign n2377 = n262 & ~n1780 ;
  assign n2378 = n2377 ^ n479 ^ 1'b0 ;
  assign n2379 = n1462 ^ x149 ^ 1'b0 ;
  assign n2380 = x187 & n2379 ;
  assign n2381 = x90 & ~n1704 ;
  assign n2382 = ~x254 & n2381 ;
  assign n2383 = x40 & n455 ;
  assign n2384 = n874 | n2383 ;
  assign n2385 = n2384 ^ n397 ^ 1'b0 ;
  assign n2386 = n2382 | n2385 ;
  assign n2387 = n2386 ^ n1167 ^ 1'b0 ;
  assign n2388 = ~n423 & n1121 ;
  assign n2389 = n640 & n2388 ;
  assign n2390 = x251 ^ x172 ^ 1'b0 ;
  assign n2391 = n1723 & ~n2390 ;
  assign n2392 = n2391 ^ x186 ^ 1'b0 ;
  assign n2393 = x115 & ~n2392 ;
  assign n2394 = n1539 & n2393 ;
  assign n2395 = ( ~x107 & n1078 ) | ( ~x107 & n2394 ) | ( n1078 & n2394 ) ;
  assign n2396 = n328 & ~n1204 ;
  assign n2397 = n1176 & n2396 ;
  assign n2398 = n2020 | n2226 ;
  assign n2399 = n2397 & ~n2398 ;
  assign n2400 = n1725 ^ n1259 ^ n1064 ;
  assign n2401 = x195 | n1190 ;
  assign n2402 = n1720 | n1838 ;
  assign n2403 = n530 | n668 ;
  assign n2404 = n2402 & n2403 ;
  assign n2405 = n1605 ^ x14 ^ 1'b0 ;
  assign n2406 = n1990 | n2405 ;
  assign n2407 = ~x199 & n1245 ;
  assign n2408 = x216 & n1577 ;
  assign n2409 = x44 ^ x38 ^ 1'b0 ;
  assign n2410 = n2409 ^ x204 ^ 1'b0 ;
  assign n2411 = n591 | n2410 ;
  assign n2412 = n1915 ^ x40 ^ 1'b0 ;
  assign n2413 = n355 & n2412 ;
  assign n2414 = x150 & n558 ;
  assign n2415 = n671 & ~n1496 ;
  assign n2416 = n2415 ^ n389 ^ x10 ;
  assign n2417 = n2414 & n2416 ;
  assign n2418 = ~n2413 & n2417 ;
  assign n2419 = n1332 ^ n1276 ^ 1'b0 ;
  assign n2420 = n415 & n2419 ;
  assign n2421 = ~n879 & n1366 ;
  assign n2422 = ~n1091 & n2421 ;
  assign n2423 = x132 & n318 ;
  assign n2424 = n270 & n2423 ;
  assign n2425 = n2424 ^ n1170 ^ 1'b0 ;
  assign n2426 = n1496 & ~n2425 ;
  assign n2427 = n799 | n1402 ;
  assign n2428 = x103 | n2427 ;
  assign n2429 = x169 & ~n527 ;
  assign n2430 = ~x230 & n2429 ;
  assign n2431 = x127 & n2430 ;
  assign n2432 = n1671 & ~n2431 ;
  assign n2433 = ~n2428 & n2432 ;
  assign n2434 = n1525 ^ x212 ^ 1'b0 ;
  assign n2435 = n1451 & n2434 ;
  assign n2436 = n2435 ^ x133 ^ 1'b0 ;
  assign n2437 = n2436 ^ n1636 ^ 1'b0 ;
  assign n2438 = n1964 & n2437 ;
  assign n2439 = n613 ^ x180 ^ 1'b0 ;
  assign n2440 = n891 & ~n2418 ;
  assign n2441 = n2440 ^ n2114 ^ 1'b0 ;
  assign n2442 = x161 ^ x0 ^ 1'b0 ;
  assign n2443 = n739 ^ x118 ^ 1'b0 ;
  assign n2444 = n695 ^ n661 ^ 1'b0 ;
  assign n2445 = n1148 & n2444 ;
  assign n2446 = ( n2442 & n2443 ) | ( n2442 & ~n2445 ) | ( n2443 & ~n2445 ) ;
  assign n2447 = x146 & ~n1409 ;
  assign n2448 = n1333 | n2447 ;
  assign n2449 = n932 ^ n817 ^ 1'b0 ;
  assign n2450 = n2448 | n2449 ;
  assign n2451 = n2450 ^ n1221 ^ 1'b0 ;
  assign n2452 = n851 | n2451 ;
  assign n2453 = n455 ^ x154 ^ 1'b0 ;
  assign n2454 = n1269 & ~n1397 ;
  assign n2455 = n2365 & n2454 ;
  assign n2456 = ~n765 & n2455 ;
  assign n2457 = n1112 & ~n1167 ;
  assign n2458 = n627 & n2457 ;
  assign n2459 = x233 & n749 ;
  assign n2460 = n2459 ^ n1295 ^ 1'b0 ;
  assign n2461 = n1034 ^ x81 ^ 1'b0 ;
  assign n2462 = n1581 & ~n2461 ;
  assign n2463 = n796 & ~n2462 ;
  assign n2464 = n1208 ^ n591 ^ n277 ;
  assign n2465 = n2464 ^ n688 ^ 1'b0 ;
  assign n2466 = n640 ^ x48 ^ 1'b0 ;
  assign n2467 = ~n1768 & n2466 ;
  assign n2468 = n2269 | n2467 ;
  assign n2476 = n1067 | n1855 ;
  assign n2469 = n921 ^ n399 ^ 1'b0 ;
  assign n2470 = x7 & ~n1762 ;
  assign n2471 = n1602 & n2470 ;
  assign n2472 = n2471 ^ n532 ^ 1'b0 ;
  assign n2473 = n1265 ^ n271 ^ 1'b0 ;
  assign n2474 = ( n993 & n2472 ) | ( n993 & ~n2473 ) | ( n2472 & ~n2473 ) ;
  assign n2475 = n2469 | n2474 ;
  assign n2477 = n2476 ^ n2475 ^ 1'b0 ;
  assign n2478 = n2214 ^ n1137 ^ 1'b0 ;
  assign n2479 = n2326 & ~n2478 ;
  assign n2480 = n2445 ^ n344 ^ 1'b0 ;
  assign n2481 = n1548 & ~n2480 ;
  assign n2482 = ( ~n322 & n732 ) | ( ~n322 & n840 ) | ( n732 & n840 ) ;
  assign n2483 = n938 ^ n281 ^ 1'b0 ;
  assign n2484 = x176 & n2483 ;
  assign n2485 = n1711 & n2484 ;
  assign n2486 = x166 ^ x1 ^ 1'b0 ;
  assign n2487 = n1977 & n2486 ;
  assign n2488 = n875 & n2487 ;
  assign n2489 = n1780 & n2488 ;
  assign n2490 = x42 & ~n322 ;
  assign n2491 = n2490 ^ n1614 ^ 1'b0 ;
  assign n2492 = n2491 ^ n361 ^ 1'b0 ;
  assign n2493 = ~x63 & n671 ;
  assign n2494 = ~n1998 & n2493 ;
  assign n2495 = n890 & ~n1593 ;
  assign n2496 = n1447 & n2495 ;
  assign n2497 = n1779 ^ n1487 ^ 1'b0 ;
  assign n2498 = n2497 ^ n613 ^ 1'b0 ;
  assign n2499 = n2496 | n2498 ;
  assign n2500 = x241 ^ x93 ^ 1'b0 ;
  assign n2501 = x109 & x130 ;
  assign n2502 = n2501 ^ n509 ^ 1'b0 ;
  assign n2503 = n634 ^ n543 ^ 1'b0 ;
  assign n2504 = n2016 & n2503 ;
  assign n2505 = n1083 & n2504 ;
  assign n2506 = ~n781 & n2505 ;
  assign n2507 = ( ~n462 & n1501 ) | ( ~n462 & n1876 ) | ( n1501 & n1876 ) ;
  assign n2508 = n2507 ^ x125 ^ 1'b0 ;
  assign n2509 = ~x89 & n471 ;
  assign n2510 = n1776 ^ x228 ^ 1'b0 ;
  assign n2511 = ~n2509 & n2510 ;
  assign n2512 = x156 & ~n699 ;
  assign n2513 = ~n1395 & n2512 ;
  assign n2514 = ~n430 & n1937 ;
  assign n2515 = x207 ^ x162 ^ 1'b0 ;
  assign n2516 = ~n2306 & n2515 ;
  assign n2517 = ~n2514 & n2516 ;
  assign n2518 = ~n1856 & n2517 ;
  assign n2519 = n2513 | n2518 ;
  assign n2520 = n2519 ^ n1335 ^ 1'b0 ;
  assign n2521 = n2099 ^ n691 ^ 1'b0 ;
  assign n2522 = n1599 & ~n1867 ;
  assign n2523 = n2096 & n2522 ;
  assign n2524 = n1208 | n2523 ;
  assign n2525 = n2227 | n2524 ;
  assign n2526 = ~x71 & n1682 ;
  assign n2530 = n340 & n2174 ;
  assign n2527 = n1440 | n1923 ;
  assign n2528 = n1219 & ~n2527 ;
  assign n2529 = ~n809 & n2528 ;
  assign n2531 = n2530 ^ n2529 ^ n1395 ;
  assign n2532 = n1593 & n2056 ;
  assign n2534 = n1151 ^ n631 ^ 1'b0 ;
  assign n2533 = ( n778 & ~n1307 ) | ( n778 & n1393 ) | ( ~n1307 & n1393 ) ;
  assign n2535 = n2534 ^ n2533 ^ n765 ;
  assign n2536 = ~n1509 & n2535 ;
  assign n2537 = n2536 ^ n2430 ^ 1'b0 ;
  assign n2538 = x34 | n1912 ;
  assign n2539 = n1721 & n2538 ;
  assign n2540 = n2539 ^ n1382 ^ 1'b0 ;
  assign n2541 = n2540 ^ n1986 ^ 1'b0 ;
  assign n2542 = n1001 ^ n430 ^ x196 ;
  assign n2543 = n935 ^ n426 ^ 1'b0 ;
  assign n2544 = n2542 & ~n2543 ;
  assign n2545 = n2244 ^ n2114 ^ n1870 ;
  assign n2554 = n2210 ^ n274 ^ 1'b0 ;
  assign n2555 = n2554 ^ n2020 ^ 1'b0 ;
  assign n2556 = ~n1286 & n2555 ;
  assign n2546 = n1494 ^ n1016 ^ 1'b0 ;
  assign n2547 = n2072 | n2546 ;
  assign n2548 = x113 & ~n281 ;
  assign n2549 = ~n302 & n2548 ;
  assign n2550 = n2549 ^ n1678 ^ n1571 ;
  assign n2551 = n2550 ^ n1075 ^ 1'b0 ;
  assign n2552 = n731 | n2551 ;
  assign n2553 = n2547 | n2552 ;
  assign n2557 = n2556 ^ n2553 ^ 1'b0 ;
  assign n2560 = ~n491 & n571 ;
  assign n2561 = n1453 & ~n1544 ;
  assign n2562 = n2560 & n2561 ;
  assign n2558 = x35 & n2340 ;
  assign n2559 = n2558 ^ n903 ^ 1'b0 ;
  assign n2563 = n2562 ^ n2559 ^ 1'b0 ;
  assign n2564 = x16 & ~n2563 ;
  assign n2565 = x14 & ~n1447 ;
  assign n2566 = n1397 & n2565 ;
  assign n2567 = n876 | n2566 ;
  assign n2568 = n2567 ^ n2216 ^ n389 ;
  assign n2569 = n922 | n1180 ;
  assign n2570 = n2569 ^ n1973 ^ 1'b0 ;
  assign n2571 = n2018 ^ n1049 ^ 1'b0 ;
  assign n2572 = n2571 ^ n1989 ^ 1'b0 ;
  assign n2573 = x61 & ~n840 ;
  assign n2574 = ~n911 & n2573 ;
  assign n2576 = n737 & ~n920 ;
  assign n2575 = n893 | n1324 ;
  assign n2577 = n2576 ^ n2575 ^ 1'b0 ;
  assign n2578 = n701 & n2577 ;
  assign n2579 = n2574 & n2578 ;
  assign n2580 = x189 & n823 ;
  assign n2581 = n400 ^ x37 ^ 1'b0 ;
  assign n2582 = n1133 & n2581 ;
  assign n2583 = x41 & ~n1099 ;
  assign n2584 = ~n2582 & n2583 ;
  assign n2585 = n2584 ^ n847 ^ 1'b0 ;
  assign n2586 = n2501 | n2585 ;
  assign n2587 = n1948 & ~n2586 ;
  assign n2588 = n1349 ^ x173 ^ 1'b0 ;
  assign n2589 = n532 & ~n2588 ;
  assign n2590 = ( n1317 & n1541 ) | ( n1317 & n2589 ) | ( n1541 & n2589 ) ;
  assign n2592 = n543 & ~n1073 ;
  assign n2591 = n672 | n1698 ;
  assign n2593 = n2592 ^ n2591 ^ 1'b0 ;
  assign n2594 = n2593 ^ n1091 ^ x122 ;
  assign n2595 = n2594 ^ n1710 ^ n957 ;
  assign n2596 = n2595 ^ n1589 ^ n705 ;
  assign n2597 = n844 & ~n959 ;
  assign n2598 = ~x164 & n2597 ;
  assign n2599 = n2596 & ~n2598 ;
  assign n2600 = n2265 & n2599 ;
  assign n2601 = x138 & n471 ;
  assign n2602 = ~x139 & n2601 ;
  assign n2603 = x77 & ~n2602 ;
  assign n2604 = ~n1118 & n2603 ;
  assign n2605 = n2604 ^ n2139 ^ 1'b0 ;
  assign n2606 = n1213 & n2605 ;
  assign n2607 = n2492 ^ n1228 ^ 1'b0 ;
  assign n2608 = n448 | n2607 ;
  assign n2609 = x56 & ~n2368 ;
  assign n2610 = n2372 ^ n1273 ^ 1'b0 ;
  assign n2611 = n327 | n2610 ;
  assign n2612 = n579 & ~n883 ;
  assign n2613 = n964 & n2612 ;
  assign n2614 = n1589 | n2613 ;
  assign n2615 = n2466 ^ x167 ^ 1'b0 ;
  assign n2616 = ~n2614 & n2615 ;
  assign n2617 = n2611 & n2616 ;
  assign n2618 = n1501 & ~n1536 ;
  assign n2619 = n688 & ~n2618 ;
  assign n2620 = n1633 & n2619 ;
  assign n2621 = x155 & ~n691 ;
  assign n2622 = n2621 ^ n334 ^ 1'b0 ;
  assign n2623 = n977 | n2622 ;
  assign n2624 = ( n1151 & n1813 ) | ( n1151 & ~n2623 ) | ( n1813 & ~n2623 ) ;
  assign n2625 = x6 & x89 ;
  assign n2626 = x139 & n2625 ;
  assign n2627 = n2626 ^ n2007 ^ 1'b0 ;
  assign n2628 = n757 & ~n2627 ;
  assign n2629 = n2628 ^ n792 ^ 1'b0 ;
  assign n2630 = n2629 ^ n2550 ^ 1'b0 ;
  assign n2631 = ~n2351 & n2630 ;
  assign n2632 = n444 | n1303 ;
  assign n2633 = n2632 ^ n462 ^ 1'b0 ;
  assign n2634 = n668 | n1477 ;
  assign n2635 = n2056 & ~n2338 ;
  assign n2636 = n2635 ^ n291 ^ 1'b0 ;
  assign n2637 = x202 & n518 ;
  assign n2638 = ~n1799 & n2637 ;
  assign n2639 = x88 & ~n2638 ;
  assign n2640 = n2639 ^ n518 ^ 1'b0 ;
  assign n2641 = ~x67 & n2640 ;
  assign n2642 = n2641 ^ n1519 ^ 1'b0 ;
  assign n2643 = n1151 & ~n2642 ;
  assign n2644 = n817 & n2643 ;
  assign n2645 = ~n382 & n591 ;
  assign n2646 = ~x168 & n2645 ;
  assign n2647 = n510 & ~n2646 ;
  assign n2648 = n2647 ^ n1365 ^ 1'b0 ;
  assign n2649 = x252 & ~n2648 ;
  assign n2650 = n2468 & n2649 ;
  assign n2651 = ~n2644 & n2650 ;
  assign n2652 = n483 | n943 ;
  assign n2653 = n1903 | n2652 ;
  assign n2654 = ( n825 & n1678 ) | ( n825 & n2653 ) | ( n1678 & n2653 ) ;
  assign n2655 = n781 & ~n1065 ;
  assign n2656 = n1591 & n1734 ;
  assign n2657 = n1676 & n2656 ;
  assign n2658 = n2655 & ~n2657 ;
  assign n2659 = n1657 & n2658 ;
  assign n2660 = x211 & ~n657 ;
  assign n2661 = n2660 ^ x172 ^ 1'b0 ;
  assign n2662 = x43 & ~n1075 ;
  assign n2663 = n2662 ^ x152 ^ 1'b0 ;
  assign n2664 = n1598 & ~n2663 ;
  assign n2665 = ~n1223 & n2664 ;
  assign n2666 = n1556 ^ x117 ^ 1'b0 ;
  assign n2667 = n2666 ^ n1369 ^ 1'b0 ;
  assign n2668 = x60 & n2667 ;
  assign n2669 = n1585 & n1678 ;
  assign n2670 = ~x59 & n2669 ;
  assign n2671 = n2670 ^ x56 ^ 1'b0 ;
  assign n2672 = n1600 & ~n2671 ;
  assign n2673 = n1782 ^ n1081 ^ 1'b0 ;
  assign n2674 = n2672 & n2673 ;
  assign n2675 = n2244 | n2674 ;
  assign n2676 = n877 ^ n604 ^ 1'b0 ;
  assign n2677 = x12 & n2676 ;
  assign n2678 = n1217 & ~n1238 ;
  assign n2679 = n1828 & ~n2678 ;
  assign n2680 = n604 & n2679 ;
  assign n2681 = ~n2677 & n2680 ;
  assign n2683 = n992 ^ n797 ^ 1'b0 ;
  assign n2684 = n1341 & n2683 ;
  assign n2682 = x157 & n2420 ;
  assign n2685 = n2684 ^ n2682 ^ n2289 ;
  assign n2686 = n948 ^ n943 ^ n876 ;
  assign n2687 = ~n756 & n1919 ;
  assign n2688 = x226 & ~n838 ;
  assign n2689 = n1294 & ~n2501 ;
  assign n2690 = n583 ^ x185 ^ 1'b0 ;
  assign n2691 = n2689 & ~n2690 ;
  assign n2692 = x164 & n464 ;
  assign n2693 = n2692 ^ n995 ^ 1'b0 ;
  assign n2694 = n2693 ^ n580 ^ 1'b0 ;
  assign n2695 = n2691 & n2694 ;
  assign n2696 = n2688 & n2695 ;
  assign n2697 = n1228 | n2696 ;
  assign n2698 = n1931 ^ x218 ^ 1'b0 ;
  assign n2699 = x203 & n2698 ;
  assign n2700 = x126 & ~n317 ;
  assign n2701 = ~x179 & n2700 ;
  assign n2702 = n826 | n2701 ;
  assign n2703 = n2702 ^ n2496 ^ 1'b0 ;
  assign n2704 = ~x80 & n1796 ;
  assign n2705 = n1433 & ~n2704 ;
  assign n2706 = n572 & ~n671 ;
  assign n2707 = n1730 & n2706 ;
  assign n2708 = n2707 ^ n2696 ^ 1'b0 ;
  assign n2709 = n1923 ^ n1796 ^ 1'b0 ;
  assign n2710 = n1062 | n2709 ;
  assign n2711 = n1262 & n2710 ;
  assign n2712 = x42 & n1581 ;
  assign n2713 = n2712 ^ n727 ^ 1'b0 ;
  assign n2714 = n980 | n2713 ;
  assign n2715 = x202 & n2714 ;
  assign n2716 = n498 ^ n437 ^ 1'b0 ;
  assign n2717 = n850 & ~n1116 ;
  assign n2718 = n2717 ^ n2018 ^ 1'b0 ;
  assign n2719 = n2718 ^ n1739 ^ 1'b0 ;
  assign n2720 = n2643 ^ x107 ^ 1'b0 ;
  assign n2721 = ~n1639 & n2720 ;
  assign n2734 = n1060 ^ n618 ^ 1'b0 ;
  assign n2735 = n784 & n2734 ;
  assign n2736 = n1085 & ~n2735 ;
  assign n2737 = ~n1067 & n2736 ;
  assign n2738 = n2737 ^ n694 ^ 1'b0 ;
  assign n2728 = n270 | n680 ;
  assign n2729 = n2728 ^ n2337 ^ 1'b0 ;
  assign n2730 = n2472 | n2729 ;
  assign n2731 = n2730 ^ n1871 ^ 1'b0 ;
  assign n2732 = n1672 & n2731 ;
  assign n2725 = n564 | n1968 ;
  assign n2722 = n1943 ^ x228 ^ 1'b0 ;
  assign n2723 = n666 & n890 ;
  assign n2724 = ~n2722 & n2723 ;
  assign n2726 = n2725 ^ n2724 ^ n1223 ;
  assign n2727 = n2154 & ~n2726 ;
  assign n2733 = n2732 ^ n2727 ^ 1'b0 ;
  assign n2739 = n2738 ^ n2733 ^ 1'b0 ;
  assign n2740 = ~x113 & n2468 ;
  assign n2744 = x27 & n1501 ;
  assign n2745 = n340 & n2744 ;
  assign n2741 = n1100 & ~n2034 ;
  assign n2742 = n2250 & ~n2741 ;
  assign n2743 = ~x31 & n2742 ;
  assign n2746 = n2745 ^ n2743 ^ 1'b0 ;
  assign n2747 = n825 ^ x188 ^ 1'b0 ;
  assign n2748 = n2747 ^ x155 ^ 1'b0 ;
  assign n2749 = ~n1817 & n2748 ;
  assign n2750 = n2749 ^ n1242 ^ 1'b0 ;
  assign n2751 = x227 & ~n927 ;
  assign n2752 = n2751 ^ n671 ^ 1'b0 ;
  assign n2753 = x34 & ~n1404 ;
  assign n2754 = ~n1659 & n2753 ;
  assign n2755 = ( n2365 & n2752 ) | ( n2365 & ~n2754 ) | ( n2752 & ~n2754 ) ;
  assign n2756 = n1993 ^ n699 ^ 1'b0 ;
  assign n2757 = ~n2585 & n2694 ;
  assign n2758 = n2757 ^ n1915 ^ 1'b0 ;
  assign n2759 = x92 & n2758 ;
  assign n2760 = n2759 ^ n1151 ^ 1'b0 ;
  assign n2761 = ~n1667 & n2760 ;
  assign n2762 = n560 ^ x29 ^ 1'b0 ;
  assign n2763 = n1439 | n2762 ;
  assign n2764 = ~x75 & n1126 ;
  assign n2765 = ( x31 & ~n1528 ) | ( x31 & n1674 ) | ( ~n1528 & n1674 ) ;
  assign n2766 = x111 & ~n1583 ;
  assign n2767 = n2766 ^ n755 ^ 1'b0 ;
  assign n2768 = n1309 ^ x33 ^ 1'b0 ;
  assign n2769 = n2337 | n2768 ;
  assign n2770 = n314 | n432 ;
  assign n2771 = n2534 ^ n1788 ^ 1'b0 ;
  assign n2772 = ~n2770 & n2771 ;
  assign n2773 = n2772 ^ n1099 ^ 1'b0 ;
  assign n2774 = ~n2769 & n2773 ;
  assign n2775 = n1557 ^ x213 ^ 1'b0 ;
  assign n2776 = n2775 ^ n1575 ^ 1'b0 ;
  assign n2777 = ~n1227 & n2358 ;
  assign n2778 = n2777 ^ n621 ^ 1'b0 ;
  assign n2779 = n1779 ^ n535 ^ 1'b0 ;
  assign n2780 = n1598 & n1737 ;
  assign n2781 = n684 & n2780 ;
  assign n2782 = n1086 | n1701 ;
  assign n2783 = n2782 ^ n1020 ^ 1'b0 ;
  assign n2784 = x57 & ~n2491 ;
  assign n2785 = n2784 ^ n1156 ^ 1'b0 ;
  assign n2786 = x232 & ~n1447 ;
  assign n2787 = n2785 & n2786 ;
  assign n2788 = n2787 ^ n2224 ^ n790 ;
  assign n2789 = n1846 ^ x189 ^ 1'b0 ;
  assign n2790 = ~n958 & n1565 ;
  assign n2791 = n2335 & ~n2790 ;
  assign n2792 = ~n325 & n2791 ;
  assign n2793 = n1167 & ~n2072 ;
  assign n2794 = ~n1064 & n2793 ;
  assign n2795 = n2794 ^ n1023 ^ 1'b0 ;
  assign n2796 = n514 | n776 ;
  assign n2797 = n2735 ^ n710 ^ n592 ;
  assign n2798 = n315 ^ x128 ^ 1'b0 ;
  assign n2799 = n272 ^ x63 ^ 1'b0 ;
  assign n2800 = n444 | n1973 ;
  assign n2801 = n2800 ^ x212 ^ 1'b0 ;
  assign n2802 = ~n423 & n1300 ;
  assign n2803 = n1405 & n2802 ;
  assign n2804 = n2095 | n2803 ;
  assign n2805 = n604 ^ n466 ^ x54 ;
  assign n2806 = n891 ^ n458 ^ 1'b0 ;
  assign n2807 = x241 & ~n2806 ;
  assign n2808 = n1011 & n2807 ;
  assign n2809 = ~n2805 & n2808 ;
  assign n2810 = ( n327 & ~n1882 ) | ( n327 & n2809 ) | ( ~n1882 & n2809 ) ;
  assign n2811 = n2666 | n2810 ;
  assign n2812 = n2811 ^ n2114 ^ 1'b0 ;
  assign n2813 = ( n298 & n2804 ) | ( n298 & n2812 ) | ( n2804 & n2812 ) ;
  assign n2814 = n2801 & ~n2813 ;
  assign n2815 = n2814 ^ n2556 ^ 1'b0 ;
  assign n2816 = ~n1739 & n2170 ;
  assign n2817 = n713 & ~n2816 ;
  assign n2818 = n458 & ~n1185 ;
  assign n2819 = n2818 ^ n814 ^ 1'b0 ;
  assign n2820 = n880 | n2370 ;
  assign n2821 = n2819 | n2820 ;
  assign n2822 = n1167 | n1273 ;
  assign n2823 = n2822 ^ n391 ^ 1'b0 ;
  assign n2824 = ~n1986 & n2823 ;
  assign n2825 = ~n1356 & n2824 ;
  assign n2826 = n2825 ^ n571 ^ 1'b0 ;
  assign n2827 = ~n2711 & n2826 ;
  assign n2828 = n668 & ~n2027 ;
  assign n2829 = n2039 ^ n475 ^ 1'b0 ;
  assign n2830 = n2828 & ~n2829 ;
  assign n2831 = n705 ^ n638 ^ x207 ;
  assign n2832 = x95 & ~n2831 ;
  assign n2833 = ~n2830 & n2832 ;
  assign n2834 = ~n697 & n1144 ;
  assign n2835 = ~n838 & n2834 ;
  assign n2836 = n1170 & ~n2835 ;
  assign n2837 = n2836 ^ x145 ^ 1'b0 ;
  assign n2838 = n2837 ^ x26 ^ 1'b0 ;
  assign n2839 = n2833 | n2838 ;
  assign n2840 = x62 & ~x159 ;
  assign n2841 = n1475 & ~n2840 ;
  assign n2842 = n272 & ~n2841 ;
  assign n2843 = ~n1500 & n2842 ;
  assign n2844 = ~n1021 & n1048 ;
  assign n2846 = n529 | n1183 ;
  assign n2845 = n2622 ^ x101 ^ 1'b0 ;
  assign n2847 = n2846 ^ n2845 ^ 1'b0 ;
  assign n2848 = n2844 | n2847 ;
  assign n2849 = n293 & ~n2848 ;
  assign n2850 = n1917 & n2849 ;
  assign n2851 = n2293 ^ n1757 ^ 1'b0 ;
  assign n2852 = n1490 & n2851 ;
  assign n2853 = ~x106 & x181 ;
  assign n2854 = n1712 | n2853 ;
  assign n2855 = n2852 | n2854 ;
  assign n2856 = ~n1779 & n2123 ;
  assign n2857 = n1627 ^ n347 ^ 1'b0 ;
  assign n2858 = n2324 & n2857 ;
  assign n2859 = n1328 ^ x168 ^ 1'b0 ;
  assign n2860 = n2706 ^ n434 ^ 1'b0 ;
  assign n2861 = x250 & n2860 ;
  assign n2862 = n449 & ~n2122 ;
  assign n2863 = n2862 ^ n1267 ^ 1'b0 ;
  assign n2864 = n2863 ^ n872 ^ 1'b0 ;
  assign n2865 = n2861 & ~n2864 ;
  assign n2866 = n2865 ^ n1297 ^ 1'b0 ;
  assign n2867 = ~n1638 & n2866 ;
  assign n2872 = x3 | n1376 ;
  assign n2871 = n1094 ^ n722 ^ 1'b0 ;
  assign n2868 = n1737 ^ x79 ^ 1'b0 ;
  assign n2869 = x174 & ~n348 ;
  assign n2870 = n2868 & n2869 ;
  assign n2873 = n2872 ^ n2871 ^ n2870 ;
  assign n2874 = x214 ^ x68 ^ 1'b0 ;
  assign n2875 = n794 & n2874 ;
  assign n2876 = ~n963 & n1217 ;
  assign n2877 = n2876 ^ n2123 ^ 1'b0 ;
  assign n2884 = n314 | n2409 ;
  assign n2878 = n1501 & ~n1589 ;
  assign n2879 = n2878 ^ n2469 ^ 1'b0 ;
  assign n2880 = n860 & n1971 ;
  assign n2881 = n2880 ^ n404 ^ 1'b0 ;
  assign n2882 = n2879 & ~n2881 ;
  assign n2883 = n2771 & n2882 ;
  assign n2885 = n2884 ^ n2883 ^ n2240 ;
  assign n2886 = n2507 ^ n1565 ^ 1'b0 ;
  assign n2887 = ~n485 & n2886 ;
  assign n2888 = n1244 ^ n925 ^ 1'b0 ;
  assign n2889 = n1172 | n2888 ;
  assign n2890 = n969 | n1610 ;
  assign n2891 = n686 & n2890 ;
  assign n2892 = n580 ^ n353 ^ 1'b0 ;
  assign n2893 = x30 & n2892 ;
  assign n2894 = ~n879 & n931 ;
  assign n2895 = ~n2893 & n2894 ;
  assign n2896 = n2283 ^ n842 ^ 1'b0 ;
  assign n2897 = n1328 ^ x196 ^ 1'b0 ;
  assign n2898 = x176 | n2804 ;
  assign n2899 = n342 | n450 ;
  assign n2900 = n2899 ^ n666 ^ 1'b0 ;
  assign n2901 = x179 & n880 ;
  assign n2902 = n2901 ^ n287 ^ 1'b0 ;
  assign n2903 = n2900 & n2902 ;
  assign n2904 = n415 & ~n2903 ;
  assign n2905 = n2904 ^ n1741 ^ n1011 ;
  assign n2906 = n2681 ^ n1176 ^ 1'b0 ;
  assign n2907 = ~n1491 & n2906 ;
  assign n2908 = x36 & n2907 ;
  assign n2909 = n2908 ^ n1993 ^ 1'b0 ;
  assign n2914 = ~n511 & n729 ;
  assign n2915 = n2914 ^ n957 ^ 1'b0 ;
  assign n2911 = ( n569 & n1786 ) | ( n569 & ~n2823 ) | ( n1786 & ~n2823 ) ;
  assign n2910 = ~n1101 & n2187 ;
  assign n2912 = n2911 ^ n2910 ^ 1'b0 ;
  assign n2913 = n2779 & n2912 ;
  assign n2916 = n2915 ^ n2913 ^ 1'b0 ;
  assign n2917 = n2104 ^ n497 ^ 1'b0 ;
  assign n2918 = x39 & ~n2917 ;
  assign n2919 = n2918 ^ n1484 ^ x185 ;
  assign n2920 = ~n1960 & n2121 ;
  assign n2921 = n937 ^ n593 ^ 1'b0 ;
  assign n2922 = n2230 & n2921 ;
  assign n2923 = n973 | n1167 ;
  assign n2924 = n2922 | n2923 ;
  assign n2925 = ( ~x118 & n1126 ) | ( ~x118 & n2080 ) | ( n1126 & n2080 ) ;
  assign n2926 = ( x238 & ~n1217 ) | ( x238 & n2925 ) | ( ~n1217 & n2925 ) ;
  assign n2927 = ( x29 & ~x230 ) | ( x29 & n1853 ) | ( ~x230 & n1853 ) ;
  assign n2928 = x63 & ~n2927 ;
  assign n2929 = n1550 ^ n1064 ^ 1'b0 ;
  assign n2930 = n1466 & ~n2929 ;
  assign n2931 = n2928 & ~n2930 ;
  assign n2932 = n2931 ^ n2330 ^ 1'b0 ;
  assign n2933 = n2037 & ~n2932 ;
  assign n2934 = n2518 ^ n856 ^ x3 ;
  assign n2935 = x189 & ~n334 ;
  assign n2936 = ( x4 & n992 ) | ( x4 & n2935 ) | ( n992 & n2935 ) ;
  assign n2937 = n2501 | n2936 ;
  assign n2938 = x73 & x245 ;
  assign n2939 = n2785 & n2938 ;
  assign n2940 = n2113 ^ n1416 ^ 1'b0 ;
  assign n2941 = n2497 | n2633 ;
  assign n2942 = n1388 | n2941 ;
  assign n2943 = x115 & n618 ;
  assign n2944 = ~n1819 & n2943 ;
  assign n2945 = n2408 & n2944 ;
  assign n2946 = n1297 ^ n1099 ^ n891 ;
  assign n2947 = x2 & n875 ;
  assign n2948 = ~n353 & n2947 ;
  assign n2956 = ~x33 & x188 ;
  assign n2949 = n1288 ^ x135 ^ 1'b0 ;
  assign n2953 = x84 & ~n987 ;
  assign n2950 = n466 & ~n1154 ;
  assign n2951 = x86 & n2950 ;
  assign n2952 = n317 | n2951 ;
  assign n2954 = n2953 ^ n2952 ^ 1'b0 ;
  assign n2955 = n2949 & ~n2954 ;
  assign n2957 = n2956 ^ n2955 ^ 1'b0 ;
  assign n2958 = n1463 ^ x72 ^ 1'b0 ;
  assign n2959 = n1581 & n2055 ;
  assign n2960 = n1997 & ~n2267 ;
  assign n2965 = x165 & x235 ;
  assign n2966 = n1208 & n2965 ;
  assign n2961 = n490 | n649 ;
  assign n2962 = n466 ^ x128 ^ 1'b0 ;
  assign n2963 = n2961 | n2962 ;
  assign n2964 = n2963 ^ n1445 ^ 1'b0 ;
  assign n2967 = n2966 ^ n2964 ^ 1'b0 ;
  assign n2968 = n2706 ^ n2061 ^ n1592 ;
  assign n2969 = n663 & ~n2968 ;
  assign n2970 = n2967 & n2969 ;
  assign n2971 = n1832 & ~n2970 ;
  assign n2972 = n256 & n2971 ;
  assign n2973 = n1753 & n2712 ;
  assign n2974 = n2973 ^ n938 ^ 1'b0 ;
  assign n2975 = n2972 & n2974 ;
  assign n2976 = x139 | n2265 ;
  assign n2977 = n2976 ^ n2403 ^ 1'b0 ;
  assign n2978 = ~n2975 & n2977 ;
  assign n2979 = x184 | n1539 ;
  assign n2980 = n809 & ~n2979 ;
  assign n2981 = ~n542 & n1887 ;
  assign n2982 = ~n2187 & n2981 ;
  assign n2983 = n1328 | n1838 ;
  assign n2984 = ( n569 & ~n1709 ) | ( n569 & n2983 ) | ( ~n1709 & n2983 ) ;
  assign n2985 = n2984 ^ n931 ^ 1'b0 ;
  assign n2986 = ~n2982 & n2985 ;
  assign n2987 = ~n1426 & n1645 ;
  assign n2988 = n1198 & n2987 ;
  assign n2989 = ~n1272 & n2414 ;
  assign n2990 = n2989 ^ n1793 ^ 1'b0 ;
  assign n2991 = n2990 ^ n2247 ^ 1'b0 ;
  assign n2992 = n1681 & ~n2991 ;
  assign n2993 = n915 & ~n1784 ;
  assign n2994 = n1415 | n2993 ;
  assign n2995 = n2994 ^ n2828 ^ 1'b0 ;
  assign n2996 = n547 ^ x167 ^ 1'b0 ;
  assign n2997 = ~n1733 & n2996 ;
  assign n2998 = n2571 ^ n436 ^ 1'b0 ;
  assign n2999 = n1423 & n2998 ;
  assign n3000 = ( n1051 & n2997 ) | ( n1051 & ~n2999 ) | ( n2997 & ~n2999 ) ;
  assign n3001 = ~n481 & n1433 ;
  assign n3002 = ~n2161 & n3001 ;
  assign n3003 = n1069 & n3002 ;
  assign n3004 = x5 & ~n1482 ;
  assign n3005 = n3003 & n3004 ;
  assign n3006 = n2493 ^ n1251 ^ 1'b0 ;
  assign n3007 = n2911 | n3006 ;
  assign n3008 = n325 & n890 ;
  assign n3009 = n3007 & n3008 ;
  assign n3010 = n385 & ~n922 ;
  assign n3011 = ~n2123 & n3010 ;
  assign n3012 = n707 | n1910 ;
  assign n3013 = n716 | n1651 ;
  assign n3014 = n2051 | n3013 ;
  assign n3015 = n2961 ^ x184 ^ 1'b0 ;
  assign n3016 = n560 | n3015 ;
  assign n3017 = n2135 | n3016 ;
  assign n3018 = x97 | n3017 ;
  assign n3019 = n3018 ^ n2243 ^ 1'b0 ;
  assign n3020 = n3019 ^ n2963 ^ 1'b0 ;
  assign n3021 = n3014 & n3020 ;
  assign n3022 = n500 & n2326 ;
  assign n3023 = n1161 | n3022 ;
  assign n3024 = n2414 ^ n891 ^ 1'b0 ;
  assign n3025 = ~n865 & n3024 ;
  assign n3026 = n399 | n2951 ;
  assign n3027 = n3026 ^ n1422 ^ 1'b0 ;
  assign n3028 = n3027 ^ n320 ^ 1'b0 ;
  assign n3033 = x19 & n453 ;
  assign n3034 = n3033 ^ x72 ^ 1'b0 ;
  assign n3035 = ~n695 & n3034 ;
  assign n3029 = n2692 ^ n2382 ^ 1'b0 ;
  assign n3030 = n810 | n3029 ;
  assign n3031 = x253 & ~n1882 ;
  assign n3032 = n3030 & n3031 ;
  assign n3036 = n3035 ^ n3032 ^ n1065 ;
  assign n3037 = x53 & n2010 ;
  assign n3038 = ~n611 & n1227 ;
  assign n3039 = n847 & ~n3038 ;
  assign n3040 = n2893 | n3039 ;
  assign n3041 = n1639 | n2809 ;
  assign n3049 = x226 & n2596 ;
  assign n3042 = n2638 ^ n498 ^ n385 ;
  assign n3043 = n367 & ~n3042 ;
  assign n3044 = n3043 ^ n1230 ^ 1'b0 ;
  assign n3045 = ~n1193 & n3044 ;
  assign n3046 = n3045 ^ n1118 ^ n647 ;
  assign n3047 = n1381 ^ x76 ^ 1'b0 ;
  assign n3048 = n3046 & ~n3047 ;
  assign n3050 = n3049 ^ n3048 ^ 1'b0 ;
  assign n3051 = x75 & ~n1999 ;
  assign n3052 = n3051 ^ x185 ^ 1'b0 ;
  assign n3053 = x76 & ~n393 ;
  assign n3054 = n3053 ^ n404 ^ 1'b0 ;
  assign n3055 = n550 & ~n1321 ;
  assign n3056 = n3055 ^ n2341 ^ 1'b0 ;
  assign n3057 = n3054 | n3056 ;
  assign n3059 = n291 ^ x164 ^ 1'b0 ;
  assign n3058 = n1165 | n1240 ;
  assign n3060 = n3059 ^ n3058 ^ n746 ;
  assign n3061 = n3060 ^ n1494 ^ 1'b0 ;
  assign n3062 = n2674 & ~n3061 ;
  assign n3063 = x230 & ~n2281 ;
  assign n3064 = n3063 ^ n851 ^ 1'b0 ;
  assign n3065 = ~n1326 & n2206 ;
  assign n3066 = ~n3064 & n3065 ;
  assign n3067 = ~x175 & n1579 ;
  assign n3068 = n2037 ^ n959 ^ 1'b0 ;
  assign n3069 = n2710 | n3068 ;
  assign n3070 = n3069 ^ n1707 ^ 1'b0 ;
  assign n3072 = n1120 ^ x240 ^ 1'b0 ;
  assign n3073 = ~n1701 & n3072 ;
  assign n3071 = x80 & ~n638 ;
  assign n3074 = n3073 ^ n3071 ^ 1'b0 ;
  assign n3077 = n1208 ^ n1100 ^ 1'b0 ;
  assign n3075 = n1016 ^ n375 ^ 1'b0 ;
  assign n3076 = ( n2016 & ~n2069 ) | ( n2016 & n3075 ) | ( ~n2069 & n3075 ) ;
  assign n3078 = n3077 ^ n3076 ^ 1'b0 ;
  assign n3079 = n2397 ^ n529 ^ 1'b0 ;
  assign n3080 = n2077 | n3079 ;
  assign n3084 = x247 & ~n716 ;
  assign n3085 = ~n353 & n3084 ;
  assign n3086 = n871 & ~n3085 ;
  assign n3081 = n376 | n977 ;
  assign n3082 = n3081 ^ n564 ^ 1'b0 ;
  assign n3083 = x115 & ~n3082 ;
  assign n3087 = n3086 ^ n3083 ^ 1'b0 ;
  assign n3088 = n3087 ^ n1725 ^ 1'b0 ;
  assign n3089 = n916 & n2305 ;
  assign n3090 = n349 & n3089 ;
  assign n3091 = n490 | n1514 ;
  assign n3092 = n1714 ^ n300 ^ 1'b0 ;
  assign n3093 = n2211 & ~n3092 ;
  assign n3094 = n3093 ^ n338 ^ 1'b0 ;
  assign n3095 = n853 | n2029 ;
  assign n3096 = n3094 | n3095 ;
  assign n3097 = n862 & n3096 ;
  assign n3098 = n3097 ^ n695 ^ 1'b0 ;
  assign n3099 = n3098 ^ n1969 ^ n1850 ;
  assign n3100 = n619 & n3099 ;
  assign n3101 = ~x107 & n391 ;
  assign n3102 = n444 & n3101 ;
  assign n3103 = n1092 & ~n2260 ;
  assign n3104 = n1707 & n3103 ;
  assign n3105 = x241 & n513 ;
  assign n3106 = n3105 ^ x135 ^ 1'b0 ;
  assign n3114 = n759 & ~n951 ;
  assign n3112 = x239 & n1245 ;
  assign n3113 = ~n518 & n3112 ;
  assign n3108 = n1714 & ~n1952 ;
  assign n3109 = ( n1358 & ~n2016 ) | ( n1358 & n3108 ) | ( ~n2016 & n3108 ) ;
  assign n3107 = ~x175 & n453 ;
  assign n3110 = n3109 ^ n3107 ^ 1'b0 ;
  assign n3111 = n3110 ^ n359 ^ x100 ;
  assign n3115 = n3114 ^ n3113 ^ n3111 ;
  assign n3116 = x120 & ~n1312 ;
  assign n3117 = n1237 & n2375 ;
  assign n3118 = ( x93 & n774 ) | ( x93 & ~n1958 ) | ( n774 & ~n1958 ) ;
  assign n3119 = n1489 ^ n1317 ^ 1'b0 ;
  assign n3124 = n397 ^ n264 ^ x214 ;
  assign n3125 = n3124 ^ x71 ^ 1'b0 ;
  assign n3126 = n417 & ~n3125 ;
  assign n3120 = n3085 ^ n1649 ^ 1'b0 ;
  assign n3121 = x125 & n3120 ;
  assign n3122 = n3121 ^ n2569 ^ x34 ;
  assign n3123 = n1689 & n3122 ;
  assign n3127 = n3126 ^ n3123 ^ 1'b0 ;
  assign n3128 = n617 & n931 ;
  assign n3129 = n3128 ^ n534 ^ 1'b0 ;
  assign n3130 = n3129 ^ x49 ^ 1'b0 ;
  assign n3131 = n289 & ~n3130 ;
  assign n3136 = ~n285 & n2445 ;
  assign n3137 = n3136 ^ n937 ^ 1'b0 ;
  assign n3132 = n903 | n1973 ;
  assign n3133 = n461 & ~n3132 ;
  assign n3134 = ~n1126 & n1862 ;
  assign n3135 = n3133 | n3134 ;
  assign n3138 = n3137 ^ n3135 ^ 1'b0 ;
  assign n3139 = n2893 ^ n560 ^ n430 ;
  assign n3140 = n937 & n3139 ;
  assign n3141 = n1051 ^ x82 ^ 1'b0 ;
  assign n3142 = n2200 & ~n3141 ;
  assign n3143 = n1539 ^ n1424 ^ 1'b0 ;
  assign n3144 = ~n2523 & n3143 ;
  assign n3145 = n444 ^ x158 ^ 1'b0 ;
  assign n3146 = x137 ^ x14 ^ 1'b0 ;
  assign n3147 = n1071 ^ x176 ^ 1'b0 ;
  assign n3148 = n3147 ^ n534 ^ 1'b0 ;
  assign n3149 = n1659 & ~n3148 ;
  assign n3150 = ( n3145 & n3146 ) | ( n3145 & n3149 ) | ( n3146 & n3149 ) ;
  assign n3151 = n1541 ^ n1330 ^ 1'b0 ;
  assign n3152 = n1257 & ~n3151 ;
  assign n3153 = n3152 ^ n333 ^ 1'b0 ;
  assign n3154 = n3150 & ~n3153 ;
  assign n3155 = n2297 ^ n2237 ^ 1'b0 ;
  assign n3156 = n1671 ^ n1364 ^ 1'b0 ;
  assign n3157 = n1475 & ~n3156 ;
  assign n3158 = n1157 & n3157 ;
  assign n3159 = n1272 ^ n1203 ^ 1'b0 ;
  assign n3161 = ~x30 & n402 ;
  assign n3160 = n491 & ~n657 ;
  assign n3162 = n3161 ^ n3160 ^ 1'b0 ;
  assign n3163 = n451 & ~n3162 ;
  assign n3166 = x155 | n744 ;
  assign n3167 = ~n1779 & n3166 ;
  assign n3168 = n1211 & n3167 ;
  assign n3164 = x48 & n1059 ;
  assign n3165 = ( n2353 & ~n2466 ) | ( n2353 & n3164 ) | ( ~n2466 & n3164 ) ;
  assign n3169 = n3168 ^ n3165 ^ 1'b0 ;
  assign n3170 = n560 | n835 ;
  assign n3171 = n3170 ^ n684 ^ 1'b0 ;
  assign n3172 = n3171 ^ n737 ^ 1'b0 ;
  assign n3173 = n831 ^ x195 ^ 1'b0 ;
  assign n3174 = ~n1286 & n3173 ;
  assign n3175 = ~n1360 & n3174 ;
  assign n3176 = ~n1481 & n3175 ;
  assign n3182 = n1762 ^ x146 ^ 1'b0 ;
  assign n3177 = ( ~x29 & n334 ) | ( ~x29 & n1977 ) | ( n334 & n1977 ) ;
  assign n3178 = n1001 & n3177 ;
  assign n3179 = ( n1793 & n2448 ) | ( n1793 & n3178 ) | ( n2448 & n3178 ) ;
  assign n3180 = n975 | n3179 ;
  assign n3181 = n2675 & ~n3180 ;
  assign n3183 = n3182 ^ n3181 ^ 1'b0 ;
  assign n3184 = n1705 & n3183 ;
  assign n3188 = ~n550 & n2949 ;
  assign n3189 = n3188 ^ n919 ^ 1'b0 ;
  assign n3190 = ~n3075 & n3189 ;
  assign n3185 = n2267 ^ n842 ^ 1'b0 ;
  assign n3186 = n738 | n3185 ;
  assign n3187 = n3184 | n3186 ;
  assign n3191 = n3190 ^ n3187 ^ 1'b0 ;
  assign n3192 = n2927 ^ n1958 ^ 1'b0 ;
  assign n3193 = n940 & n3192 ;
  assign n3194 = n1885 & n3193 ;
  assign n3195 = n3194 ^ n835 ^ 1'b0 ;
  assign n3196 = n599 & ~n927 ;
  assign n3197 = ~n285 & n3196 ;
  assign n3198 = n1351 | n2741 ;
  assign n3199 = ~n1741 & n2521 ;
  assign n3201 = n2577 ^ n1368 ^ 1'b0 ;
  assign n3200 = x247 & ~n2065 ;
  assign n3202 = n3201 ^ n3200 ^ 1'b0 ;
  assign n3203 = n1259 ^ n601 ^ 1'b0 ;
  assign n3204 = n3203 ^ n1283 ^ 1'b0 ;
  assign n3205 = n3164 | n3204 ;
  assign n3206 = n1812 & n1896 ;
  assign n3207 = ~n446 & n894 ;
  assign n3208 = ~n2726 & n3207 ;
  assign n3209 = ~n1459 & n3208 ;
  assign n3210 = n2618 ^ n340 ^ 1'b0 ;
  assign n3211 = n2243 ^ n1369 ^ 1'b0 ;
  assign n3212 = x37 & n1344 ;
  assign n3213 = n1192 & n3212 ;
  assign n3214 = x128 | n3213 ;
  assign n3215 = n3214 ^ n372 ^ 1'b0 ;
  assign n3216 = n1534 ^ n1198 ^ 1'b0 ;
  assign n3217 = ( n1247 & n3215 ) | ( n1247 & n3216 ) | ( n3215 & n3216 ) ;
  assign n3218 = n815 | n2113 ;
  assign n3220 = x22 & ~n983 ;
  assign n3221 = ~n2533 & n3220 ;
  assign n3219 = n1813 & n2779 ;
  assign n3222 = n3221 ^ n3219 ^ 1'b0 ;
  assign n3223 = ( x62 & ~x228 ) | ( x62 & n434 ) | ( ~x228 & n434 ) ;
  assign n3224 = x58 & x176 ;
  assign n3225 = n897 & n3224 ;
  assign n3226 = n3225 ^ n1369 ^ 1'b0 ;
  assign n3227 = n3223 & n3226 ;
  assign n3228 = ~n424 & n3227 ;
  assign n3229 = n3114 | n3228 ;
  assign n3230 = n1544 & ~n3229 ;
  assign n3231 = n3230 ^ n2204 ^ 1'b0 ;
  assign n3232 = n2332 ^ n1254 ^ 1'b0 ;
  assign n3233 = n3179 ^ n547 ^ 1'b0 ;
  assign n3234 = n3174 ^ n325 ^ 1'b0 ;
  assign n3235 = n1495 & ~n2640 ;
  assign n3236 = n1711 & n1893 ;
  assign n3237 = n3236 ^ n431 ^ 1'b0 ;
  assign n3238 = n3237 ^ n2008 ^ n1333 ;
  assign n3239 = n569 ^ n271 ^ 1'b0 ;
  assign n3240 = ~n809 & n3239 ;
  assign n3241 = n932 ^ n359 ^ 1'b0 ;
  assign n3242 = n1867 | n3241 ;
  assign n3243 = x249 | n3242 ;
  assign n3244 = n627 | n2681 ;
  assign n3245 = n1684 | n3244 ;
  assign n3246 = n2544 ^ x29 ^ 1'b0 ;
  assign n3250 = n1523 ^ n415 ^ 1'b0 ;
  assign n3247 = n2846 ^ x110 ^ 1'b0 ;
  assign n3248 = ~n1200 & n3247 ;
  assign n3249 = ( ~n1369 & n1393 ) | ( ~n1369 & n3248 ) | ( n1393 & n3248 ) ;
  assign n3251 = n3250 ^ n3249 ^ n2072 ;
  assign n3252 = n2513 ^ n1931 ^ 1'b0 ;
  assign n3253 = n1462 & ~n3252 ;
  assign n3254 = n3253 ^ n2733 ^ 1'b0 ;
  assign n3255 = n1480 | n3254 ;
  assign n3256 = n3255 ^ n1689 ^ 1'b0 ;
  assign n3257 = n1463 | n1866 ;
  assign n3258 = ( n293 & n1116 ) | ( n293 & ~n3257 ) | ( n1116 & ~n3257 ) ;
  assign n3259 = n2045 | n3258 ;
  assign n3260 = n3259 ^ n1450 ^ 1'b0 ;
  assign n3261 = n1132 & ~n1948 ;
  assign n3262 = ~n634 & n3261 ;
  assign n3263 = ~n3260 & n3262 ;
  assign n3264 = n1943 ^ n856 ^ 1'b0 ;
  assign n3265 = n635 & ~n1837 ;
  assign n3266 = x29 & ~n3265 ;
  assign n3267 = ( x107 & ~n2260 ) | ( x107 & n2314 ) | ( ~n2260 & n2314 ) ;
  assign n3268 = n1114 | n2967 ;
  assign n3269 = n3131 | n3268 ;
  assign n3270 = n1231 ^ n676 ^ 1'b0 ;
  assign n3271 = n847 & n3270 ;
  assign n3272 = n3271 ^ n1528 ^ 1'b0 ;
  assign n3273 = n1475 | n3272 ;
  assign n3274 = n3273 ^ n3049 ^ 1'b0 ;
  assign n3275 = ( n2334 & ~n2445 ) | ( n2334 & n3058 ) | ( ~n2445 & n3058 ) ;
  assign n3276 = n789 & n1599 ;
  assign n3277 = n3276 ^ n1138 ^ 1'b0 ;
  assign n3278 = n1802 & n2936 ;
  assign n3279 = n3277 & n3278 ;
  assign n3280 = x98 & ~n711 ;
  assign n3281 = n3280 ^ n908 ^ 1'b0 ;
  assign n3282 = x24 & n2764 ;
  assign n3283 = n518 & n3282 ;
  assign n3284 = n1788 | n3283 ;
  assign n3290 = x162 & n891 ;
  assign n3287 = n507 & ~n589 ;
  assign n3285 = ~n535 & n2208 ;
  assign n3286 = n461 & n3285 ;
  assign n3288 = n3287 ^ n3286 ^ n2085 ;
  assign n3289 = n1368 | n3288 ;
  assign n3291 = n3290 ^ n3289 ^ 1'b0 ;
  assign n3296 = x121 & n765 ;
  assign n3292 = x130 & n2086 ;
  assign n3293 = n3292 ^ x77 ^ 1'b0 ;
  assign n3294 = n2840 ^ n488 ^ 1'b0 ;
  assign n3295 = ~n3293 & n3294 ;
  assign n3297 = n3296 ^ n3295 ^ 1'b0 ;
  assign n3298 = x195 & n509 ;
  assign n3299 = n763 & n2542 ;
  assign n3300 = ~n831 & n3299 ;
  assign n3301 = n2127 ^ n617 ^ 1'b0 ;
  assign n3302 = n3300 | n3301 ;
  assign n3303 = n2640 & ~n3302 ;
  assign n3304 = n3298 & n3303 ;
  assign n3305 = n2582 ^ n1134 ^ 1'b0 ;
  assign n3306 = ~n2455 & n3305 ;
  assign n3307 = n3306 ^ n3064 ^ 1'b0 ;
  assign n3308 = n537 | n3307 ;
  assign n3309 = n2550 ^ n2494 ^ 1'b0 ;
  assign n3310 = n1416 & n3309 ;
  assign n3311 = n3310 ^ n1861 ^ 1'b0 ;
  assign n3312 = n2221 ^ n2191 ^ x147 ;
  assign n3313 = x156 & n3186 ;
  assign n3314 = n988 | n2884 ;
  assign n3315 = n1332 & ~n3314 ;
  assign n3316 = ( ~n809 & n1657 ) | ( ~n809 & n1788 ) | ( n1657 & n1788 ) ;
  assign n3317 = n2967 ^ n516 ^ 1'b0 ;
  assign n3318 = n1844 | n3317 ;
  assign n3319 = n3316 & ~n3318 ;
  assign n3320 = n2219 & ~n2831 ;
  assign n3321 = n3082 & n3320 ;
  assign n3322 = n983 | n2297 ;
  assign n3323 = n3322 ^ n1979 ^ 1'b0 ;
  assign n3324 = ~n694 & n3323 ;
  assign n3325 = ~n2858 & n3324 ;
  assign n3326 = n2030 ^ n1437 ^ 1'b0 ;
  assign n3327 = ( ~n434 & n1435 ) | ( ~n434 & n3326 ) | ( n1435 & n3326 ) ;
  assign n3330 = n1107 & ~n3161 ;
  assign n3331 = n3330 ^ n1326 ^ 1'b0 ;
  assign n3328 = n1822 ^ n1590 ^ 1'b0 ;
  assign n3329 = n3328 ^ n2780 ^ 1'b0 ;
  assign n3332 = n3331 ^ n3329 ^ n890 ;
  assign n3333 = n831 | n1386 ;
  assign n3334 = n433 & ~n922 ;
  assign n3335 = n3334 ^ x171 ^ 1'b0 ;
  assign n3336 = n1217 ^ n1053 ^ 1'b0 ;
  assign n3337 = n1495 & ~n3336 ;
  assign n3338 = n2756 | n3337 ;
  assign n3339 = n1037 | n3338 ;
  assign n3340 = x236 | n2020 ;
  assign n3341 = n328 & ~n1130 ;
  assign n3342 = n3341 ^ n3335 ^ 1'b0 ;
  assign n3343 = ~n2934 & n3342 ;
  assign n3344 = n1680 & n3343 ;
  assign n3348 = x192 & n1519 ;
  assign n3345 = n1550 ^ x64 ^ 1'b0 ;
  assign n3346 = n1981 | n3345 ;
  assign n3347 = n2533 & ~n3346 ;
  assign n3349 = n3348 ^ n3347 ^ 1'b0 ;
  assign n3350 = n958 & ~n3234 ;
  assign n3351 = ~n3349 & n3350 ;
  assign n3352 = n1336 & ~n3351 ;
  assign n3353 = n1384 ^ n334 ^ x37 ;
  assign n3354 = n1504 | n2829 ;
  assign n3355 = n3353 | n3354 ;
  assign n3356 = n266 & ~n677 ;
  assign n3357 = n413 & n3356 ;
  assign n3358 = x159 & ~n969 ;
  assign n3359 = ~n1295 & n3358 ;
  assign n3360 = n3359 ^ n2140 ^ 1'b0 ;
  assign n3361 = n3357 | n3360 ;
  assign n3362 = n3355 | n3361 ;
  assign n3366 = x245 & n2015 ;
  assign n3367 = ~x248 & n3366 ;
  assign n3363 = n1272 ^ x45 ^ 1'b0 ;
  assign n3364 = ~n1178 & n3363 ;
  assign n3365 = x238 & n3364 ;
  assign n3368 = n3367 ^ n3365 ^ 1'b0 ;
  assign n3369 = n3362 & n3368 ;
  assign n3370 = n3369 ^ n3234 ^ 1'b0 ;
  assign n3371 = ~x192 & n1500 ;
  assign n3372 = n1620 ^ n977 ^ 1'b0 ;
  assign n3373 = n752 | n2868 ;
  assign n3374 = n752 & ~n3373 ;
  assign n3375 = n1312 | n3374 ;
  assign n3376 = n542 | n547 ;
  assign n3377 = n3376 ^ n1151 ^ 1'b0 ;
  assign n3378 = n3377 ^ n3012 ^ n309 ;
  assign n3379 = n1463 ^ n921 ^ 1'b0 ;
  assign n3380 = ~n1752 & n3379 ;
  assign n3381 = x247 | n1630 ;
  assign n3382 = n3381 ^ n1501 ^ 1'b0 ;
  assign n3383 = n3382 ^ n613 ^ 1'b0 ;
  assign n3384 = n378 & ~n1569 ;
  assign n3385 = ~n1735 & n3384 ;
  assign n3386 = n986 & ~n3385 ;
  assign n3387 = n2016 ^ x198 ^ 1'b0 ;
  assign n3388 = x251 & n3387 ;
  assign n3389 = n2502 | n3388 ;
  assign n3390 = n880 | n1711 ;
  assign n3391 = n2015 | n3390 ;
  assign n3392 = n3391 ^ n2375 ^ 1'b0 ;
  assign n3393 = n3150 & ~n3392 ;
  assign n3394 = n1695 ^ n969 ^ 1'b0 ;
  assign n3395 = ~n1376 & n3394 ;
  assign n3396 = n3123 & n3395 ;
  assign n3397 = ( n2056 & ~n2276 ) | ( n2056 & n3207 ) | ( ~n2276 & n3207 ) ;
  assign n3398 = n3397 ^ x82 ^ 1'b0 ;
  assign n3399 = n1230 & n3398 ;
  assign n3400 = n527 | n1657 ;
  assign n3401 = ~n946 & n2117 ;
  assign n3402 = ~n430 & n1581 ;
  assign n3403 = n3402 ^ x238 ^ 1'b0 ;
  assign n3404 = x50 & ~n2279 ;
  assign n3405 = ( n3401 & ~n3403 ) | ( n3401 & n3404 ) | ( ~n3403 & n3404 ) ;
  assign n3406 = n1195 & ~n1674 ;
  assign n3407 = n3406 ^ n351 ^ 1'b0 ;
  assign n3408 = x200 & n3407 ;
  assign n3409 = n3405 & ~n3408 ;
  assign n3410 = n333 & n3409 ;
  assign n3411 = n1770 & n2433 ;
  assign n3412 = n3411 ^ n406 ^ 1'b0 ;
  assign n3415 = n3287 ^ n909 ^ n407 ;
  assign n3416 = n3415 ^ n1841 ^ x121 ;
  assign n3413 = ~x172 & n1880 ;
  assign n3414 = n1010 | n3413 ;
  assign n3417 = n3416 ^ n3414 ^ 1'b0 ;
  assign n3420 = ~x204 & n915 ;
  assign n3421 = ~n2884 & n3420 ;
  assign n3422 = n1983 & n3421 ;
  assign n3423 = n3422 ^ n2477 ^ 1'b0 ;
  assign n3418 = ~x195 & n2697 ;
  assign n3419 = n3418 ^ x13 ^ 1'b0 ;
  assign n3424 = n3423 ^ n3419 ^ 1'b0 ;
  assign n3425 = n413 ^ x232 ^ 1'b0 ;
  assign n3426 = ~n2265 & n3425 ;
  assign n3427 = n3426 ^ n3396 ^ 1'b0 ;
  assign n3428 = n828 ^ x42 ^ 1'b0 ;
  assign n3429 = n366 & ~n3428 ;
  assign n3430 = n3171 ^ n2891 ^ 1'b0 ;
  assign n3431 = ~n3328 & n3430 ;
  assign n3432 = n1654 & n3431 ;
  assign n3433 = n2738 & ~n3109 ;
  assign n3434 = n2900 ^ n1361 ^ 1'b0 ;
  assign n3435 = n3433 & ~n3434 ;
  assign n3436 = n1610 & ~n2594 ;
  assign n3437 = ~x181 & n3436 ;
  assign n3438 = n3329 & ~n3437 ;
  assign n3439 = ~n2312 & n3438 ;
  assign n3440 = n2827 | n3348 ;
  assign n3441 = n1968 ^ n642 ^ 1'b0 ;
  assign n3442 = ~n285 & n3441 ;
  assign n3443 = n2895 ^ n1550 ^ 1'b0 ;
  assign n3444 = ~n1177 & n3443 ;
  assign n3445 = n2465 ^ n445 ^ 1'b0 ;
  assign n3446 = n3444 & n3445 ;
  assign n3447 = n1247 ^ n1043 ^ n917 ;
  assign n3448 = ~n1147 & n3447 ;
  assign n3449 = n3448 ^ x223 ^ 1'b0 ;
  assign n3450 = ( n395 & n1593 ) | ( n395 & n3449 ) | ( n1593 & n3449 ) ;
  assign n3451 = n2549 ^ n1633 ^ 1'b0 ;
  assign n3452 = n3451 ^ n1754 ^ 1'b0 ;
  assign n3453 = n1456 & n3452 ;
  assign n3454 = ~x26 & n3453 ;
  assign n3455 = ~n3450 & n3454 ;
  assign n3456 = n1674 | n3455 ;
  assign n3457 = n3456 ^ n1744 ^ 1'b0 ;
  assign n3458 = n1352 & ~n1381 ;
  assign n3459 = n3458 ^ n1435 ^ 1'b0 ;
  assign n3460 = ~x175 & n3459 ;
  assign n3461 = n380 & ~n577 ;
  assign n3462 = ( ~x35 & x40 ) | ( ~x35 & n1471 ) | ( x40 & n1471 ) ;
  assign n3463 = n2219 ^ n325 ^ 1'b0 ;
  assign n3464 = ~n3462 & n3463 ;
  assign n3465 = n466 & n2239 ;
  assign n3466 = n3465 ^ n983 ^ 1'b0 ;
  assign n3467 = n3464 & ~n3466 ;
  assign n3468 = ( n2452 & n3388 ) | ( n2452 & n3467 ) | ( n3388 & n3467 ) ;
  assign n3469 = ~n264 & n1887 ;
  assign n3470 = n3469 ^ x148 ^ 1'b0 ;
  assign n3471 = x76 & ~n419 ;
  assign n3472 = n3471 ^ n1070 ^ 1'b0 ;
  assign n3473 = n1114 | n1288 ;
  assign n3474 = n3473 ^ n322 ^ 1'b0 ;
  assign n3475 = n3474 ^ n466 ^ 1'b0 ;
  assign n3476 = n2420 & ~n3475 ;
  assign n3477 = n2853 & n3476 ;
  assign n3478 = ( ~n3470 & n3472 ) | ( ~n3470 & n3477 ) | ( n3472 & n3477 ) ;
  assign n3479 = n2196 ^ n1844 ^ 1'b0 ;
  assign n3480 = ~n1354 & n3479 ;
  assign n3481 = n2165 & n3480 ;
  assign n3482 = x247 & ~n1219 ;
  assign n3483 = n1667 & n3482 ;
  assign n3484 = n1315 | n3483 ;
  assign n3485 = n1097 | n3484 ;
  assign n3486 = n3485 ^ n1088 ^ 1'b0 ;
  assign n3487 = n1938 ^ n1558 ^ 1'b0 ;
  assign n3488 = n3396 & ~n3487 ;
  assign n3489 = n1815 & ~n2142 ;
  assign n3490 = n3489 ^ n425 ^ 1'b0 ;
  assign n3492 = n2137 ^ n799 ^ 1'b0 ;
  assign n3493 = ~n2796 & n3492 ;
  assign n3494 = n1669 & n2304 ;
  assign n3495 = n3003 | n3494 ;
  assign n3496 = n3493 | n3495 ;
  assign n3491 = n968 ^ n614 ^ n416 ;
  assign n3497 = n3496 ^ n3491 ^ 1'b0 ;
  assign n3498 = ~n1547 & n3497 ;
  assign n3499 = ( ~n697 & n858 ) | ( ~n697 & n1828 ) | ( n858 & n1828 ) ;
  assign n3500 = n980 & n2722 ;
  assign n3501 = n3499 & ~n3500 ;
  assign n3502 = ~n445 & n3501 ;
  assign n3503 = n3463 ^ n2775 ^ 1'b0 ;
  assign n3504 = n2929 & ~n3503 ;
  assign n3505 = n1830 | n2464 ;
  assign n3506 = ( x75 & n665 ) | ( x75 & n3505 ) | ( n665 & n3505 ) ;
  assign n3507 = ~n710 & n3506 ;
  assign n3508 = ~x193 & n3507 ;
  assign n3509 = n1917 ^ n1828 ^ 1'b0 ;
  assign n3510 = n3509 ^ n2410 ^ 1'b0 ;
  assign n3511 = ~n1183 & n3510 ;
  assign n3512 = n2154 & n3511 ;
  assign n3513 = n1758 & n3512 ;
  assign n3514 = n2508 ^ x82 ^ 1'b0 ;
  assign n3516 = n466 & n532 ;
  assign n3517 = n3516 ^ n3248 ^ 1'b0 ;
  assign n3515 = n1876 | n3272 ;
  assign n3518 = n3517 ^ n3515 ^ 1'b0 ;
  assign n3519 = n1089 & n1829 ;
  assign n3520 = n3519 ^ n1710 ^ 1'b0 ;
  assign n3521 = n3451 ^ x89 ^ 1'b0 ;
  assign n3522 = n1426 | n3521 ;
  assign n3523 = n668 | n3522 ;
  assign n3524 = n2164 ^ x160 ^ 1'b0 ;
  assign n3525 = n3523 & n3524 ;
  assign n3526 = ~n1172 & n3525 ;
  assign n3527 = n3520 & n3526 ;
  assign n3528 = n264 ^ x131 ^ 1'b0 ;
  assign n3529 = n2953 | n3528 ;
  assign n3530 = x201 | n3529 ;
  assign n3531 = n1636 | n2281 ;
  assign n3532 = n3530 | n3531 ;
  assign n3533 = n2509 | n3529 ;
  assign n3534 = n3533 ^ n2920 ^ 1'b0 ;
  assign n3535 = ~n920 & n2768 ;
  assign n3536 = n2936 ^ n1935 ^ 1'b0 ;
  assign n3537 = n3536 ^ n3225 ^ 1'b0 ;
  assign n3538 = n1373 & ~n1603 ;
  assign n3539 = ~n1295 & n3538 ;
  assign n3540 = n3419 | n3539 ;
  assign n3541 = n3540 ^ n2299 ^ 1'b0 ;
  assign n3542 = n2926 ^ n2198 ^ 1'b0 ;
  assign n3546 = ~n867 & n963 ;
  assign n3544 = x95 | n2223 ;
  assign n3543 = n3165 ^ n2704 ^ 1'b0 ;
  assign n3545 = n3544 ^ n3543 ^ 1'b0 ;
  assign n3547 = n3546 ^ n3545 ^ n407 ;
  assign n3548 = n689 & ~n2085 ;
  assign n3549 = ~n1124 & n3548 ;
  assign n3550 = n1807 ^ n1550 ^ 1'b0 ;
  assign n3551 = ~n3549 & n3550 ;
  assign n3552 = n2865 ^ n1736 ^ n585 ;
  assign n3553 = x247 & ~n3552 ;
  assign n3554 = ~n3551 & n3553 ;
  assign n3555 = ~n676 & n2119 ;
  assign n3556 = n2907 ^ x48 ^ 1'b0 ;
  assign n3557 = ~n3555 & n3556 ;
  assign n3558 = n3557 ^ n3288 ^ 1'b0 ;
  assign n3559 = n628 & ~n1999 ;
  assign n3560 = n3559 ^ x25 ^ 1'b0 ;
  assign n3561 = n1364 | n2974 ;
  assign n3562 = n1328 | n3359 ;
  assign n3563 = n3562 ^ n893 ^ 1'b0 ;
  assign n3564 = x113 & ~n2594 ;
  assign n3565 = n2823 ^ n1938 ^ 1'b0 ;
  assign n3567 = ( ~x229 & x235 ) | ( ~x229 & n274 ) | ( x235 & n274 ) ;
  assign n3566 = x238 & ~n469 ;
  assign n3568 = n3567 ^ n3566 ^ 1'b0 ;
  assign n3569 = n720 | n3568 ;
  assign n3570 = ~n1149 & n3569 ;
  assign n3571 = n3177 & n3570 ;
  assign n3572 = n2210 & n2240 ;
  assign n3573 = ~n1586 & n3572 ;
  assign n3574 = n1356 & n2925 ;
  assign n3575 = ~n264 & n3207 ;
  assign n3576 = n3575 ^ n1347 ^ 1'b0 ;
  assign n3580 = n888 | n3293 ;
  assign n3581 = n3580 ^ n302 ^ 1'b0 ;
  assign n3577 = n1632 ^ n1585 ^ x151 ;
  assign n3578 = ~n1489 & n3577 ;
  assign n3579 = ~n3450 & n3578 ;
  assign n3582 = n3581 ^ n3579 ^ n834 ;
  assign n3583 = n3582 ^ n752 ^ 1'b0 ;
  assign n3584 = ~n1147 & n3583 ;
  assign n3585 = n3293 ^ n997 ^ 1'b0 ;
  assign n3586 = n2008 & n3585 ;
  assign n3587 = x87 & n3586 ;
  assign n3588 = n479 & n3587 ;
  assign n3589 = n3588 ^ n1219 ^ 1'b0 ;
  assign n3590 = n3589 ^ n2424 ^ n466 ;
  assign n3591 = n854 | n1185 ;
  assign n3592 = n3147 & ~n3591 ;
  assign n3593 = n635 & n2110 ;
  assign n3594 = n3593 ^ n436 ^ 1'b0 ;
  assign n3595 = n2043 ^ n1619 ^ 1'b0 ;
  assign n3596 = n353 & n3595 ;
  assign n3601 = n1049 ^ n632 ^ x16 ;
  assign n3602 = n387 & n739 ;
  assign n3603 = ~n854 & n3602 ;
  assign n3604 = n3601 & ~n3603 ;
  assign n3597 = x149 & ~n751 ;
  assign n3598 = n3597 ^ n1501 ^ 1'b0 ;
  assign n3599 = n3598 ^ x33 ^ 1'b0 ;
  assign n3600 = n2034 & n3599 ;
  assign n3605 = n3604 ^ n3600 ^ 1'b0 ;
  assign n3606 = ~n1649 & n3605 ;
  assign n3607 = n1081 & ~n2316 ;
  assign n3608 = ~n865 & n3607 ;
  assign n3609 = n2576 ^ n908 ^ 1'b0 ;
  assign n3610 = n1838 & ~n3609 ;
  assign n3611 = n3610 ^ n889 ^ 1'b0 ;
  assign n3615 = ~n3151 & n3250 ;
  assign n3612 = x234 & ~n1938 ;
  assign n3613 = n2967 & n3612 ;
  assign n3614 = ( x177 & ~n3059 ) | ( x177 & n3613 ) | ( ~n3059 & n3613 ) ;
  assign n3616 = n3615 ^ n3614 ^ 1'b0 ;
  assign n3617 = n2661 ^ n2634 ^ 1'b0 ;
  assign n3618 = n671 & n3157 ;
  assign n3619 = n3618 ^ n640 ^ 1'b0 ;
  assign n3620 = ~n258 & n2866 ;
  assign n3621 = ~n2988 & n3620 ;
  assign n3622 = ~n2117 & n3621 ;
  assign n3623 = n1297 ^ n1288 ^ 1'b0 ;
  assign n3624 = n842 & ~n3623 ;
  assign n3625 = ~n716 & n1341 ;
  assign n3626 = n3625 ^ x174 ^ 1'b0 ;
  assign n3627 = n2494 ^ n710 ^ 1'b0 ;
  assign n3628 = x80 & n1116 ;
  assign n3629 = n2835 ^ n1735 ^ 1'b0 ;
  assign n3630 = n3629 ^ n1725 ^ 1'b0 ;
  assign n3631 = n2192 & ~n3630 ;
  assign n3632 = n2679 ^ n1945 ^ 1'b0 ;
  assign n3633 = x75 & n3632 ;
  assign n3634 = n428 & ~n1647 ;
  assign n3635 = ~n2927 & n3007 ;
  assign n3636 = n3634 & ~n3635 ;
  assign n3637 = ~n3633 & n3636 ;
  assign n3638 = n2268 & n2360 ;
  assign n3639 = n3637 & n3638 ;
  assign n3640 = ( ~n1527 & n2745 ) | ( ~n1527 & n2787 ) | ( n2745 & n2787 ) ;
  assign n3641 = n2604 & ~n3640 ;
  assign n3642 = n1779 | n3572 ;
  assign n3643 = n3642 ^ n991 ^ 1'b0 ;
  assign n3644 = n1342 ^ x73 ^ 1'b0 ;
  assign n3645 = ~n516 & n3644 ;
  assign n3646 = n1175 ^ x16 ^ 1'b0 ;
  assign n3647 = n3646 ^ n523 ^ 1'b0 ;
  assign n3648 = ( n477 & n3645 ) | ( n477 & ~n3647 ) | ( n3645 & ~n3647 ) ;
  assign n3649 = n3648 ^ n2974 ^ 1'b0 ;
  assign n3650 = n3109 ^ n1378 ^ x93 ;
  assign n3651 = n2328 & ~n3650 ;
  assign n3652 = n1294 & ~n3403 ;
  assign n3653 = n3652 ^ n1696 ^ 1'b0 ;
  assign n3654 = n2623 | n3653 ;
  assign n3655 = n3298 ^ n1382 ^ 1'b0 ;
  assign n3656 = n615 | n3655 ;
  assign n3657 = n1553 | n3054 ;
  assign n3658 = x158 ^ x97 ^ 1'b0 ;
  assign n3659 = ~n943 & n3658 ;
  assign n3660 = n1919 & ~n3258 ;
  assign n3661 = n3660 ^ n1361 ^ 1'b0 ;
  assign n3662 = n3659 & n3661 ;
  assign n3663 = n3657 & n3662 ;
  assign n3664 = n957 ^ x111 ^ 1'b0 ;
  assign n3665 = ~n3663 & n3664 ;
  assign n3666 = ( x199 & n1170 ) | ( x199 & ~n1803 ) | ( n1170 & ~n1803 ) ;
  assign n3667 = x143 & ~n1453 ;
  assign n3668 = n2770 & ~n3667 ;
  assign n3669 = n267 | n1203 ;
  assign n3670 = n3669 ^ n332 ^ 1'b0 ;
  assign n3671 = ( x240 & ~n747 ) | ( x240 & n3670 ) | ( ~n747 & n3670 ) ;
  assign n3672 = n1400 ^ n975 ^ x127 ;
  assign n3673 = n3672 ^ n2077 ^ 1'b0 ;
  assign n3674 = ( ~n1506 & n2396 ) | ( ~n1506 & n3673 ) | ( n2396 & n3673 ) ;
  assign n3675 = n3671 | n3674 ;
  assign n3676 = n3675 ^ n2351 ^ 1'b0 ;
  assign n3677 = n2484 ^ n825 ^ 1'b0 ;
  assign n3679 = n2646 ^ n1279 ^ n677 ;
  assign n3680 = n3679 ^ n1250 ^ 1'b0 ;
  assign n3678 = ~n838 & n2596 ;
  assign n3681 = n3680 ^ n3678 ^ 1'b0 ;
  assign n3682 = x7 & ~n3681 ;
  assign n3683 = n3682 ^ n3615 ^ 1'b0 ;
  assign n3684 = ( n2376 & n3677 ) | ( n2376 & ~n3683 ) | ( n3677 & ~n3683 ) ;
  assign n3685 = x63 & n2841 ;
  assign n3686 = n1528 ^ n548 ^ 1'b0 ;
  assign n3687 = n784 & n3364 ;
  assign n3688 = n3686 & n3687 ;
  assign n3689 = n1608 ^ n627 ^ 1'b0 ;
  assign n3690 = n1583 ^ n1081 ^ n699 ;
  assign n3691 = n3689 & n3690 ;
  assign n3692 = n3691 ^ n1875 ^ 1'b0 ;
  assign n3693 = n3688 | n3692 ;
  assign n3694 = ( n2956 & n3685 ) | ( n2956 & ~n3693 ) | ( n3685 & ~n3693 ) ;
  assign n3695 = n3694 ^ n475 ^ 1'b0 ;
  assign n3696 = n1965 & ~n2345 ;
  assign n3697 = x36 & ~n1992 ;
  assign n3698 = n3696 & n3697 ;
  assign n3701 = ( n1037 & ~n1151 ) | ( n1037 & n2577 ) | ( ~n1151 & n2577 ) ;
  assign n3702 = n437 & n3701 ;
  assign n3699 = n1360 ^ x112 ^ 1'b0 ;
  assign n3700 = n2102 & ~n3699 ;
  assign n3703 = n3702 ^ n3700 ^ 1'b0 ;
  assign n3704 = n3703 ^ n2489 ^ n752 ;
  assign n3705 = ( n3305 & n3455 ) | ( n3305 & ~n3704 ) | ( n3455 & ~n3704 ) ;
  assign n3706 = x188 & n353 ;
  assign n3707 = ~n2108 & n3706 ;
  assign n3708 = n2816 | n3594 ;
  assign n3709 = n3708 ^ n511 ^ 1'b0 ;
  assign n3710 = n3648 ^ n514 ^ 1'b0 ;
  assign n3711 = n1513 & ~n3419 ;
  assign n3712 = ~n2936 & n3711 ;
  assign n3714 = ~n673 & n747 ;
  assign n3715 = n1276 ^ n1130 ^ 1'b0 ;
  assign n3716 = n3714 & n3715 ;
  assign n3713 = n2644 & n3154 ;
  assign n3717 = n3716 ^ n3713 ^ 1'b0 ;
  assign n3718 = ~n382 & n1508 ;
  assign n3719 = n3718 ^ x67 ^ 1'b0 ;
  assign n3720 = n2879 ^ n2237 ^ 1'b0 ;
  assign n3721 = n3719 | n3720 ;
  assign n3722 = n842 & ~n3685 ;
  assign n3723 = ~n367 & n2602 ;
  assign n3724 = n3723 ^ n2523 ^ n969 ;
  assign n3725 = n3724 ^ n3719 ^ 1'b0 ;
  assign n3726 = n2267 | n3725 ;
  assign n3727 = ~n306 & n2827 ;
  assign n3728 = n3727 ^ n2927 ^ 1'b0 ;
  assign n3729 = ( n347 & ~n2458 ) | ( n347 & n3728 ) | ( ~n2458 & n3728 ) ;
  assign n3730 = n494 | n1676 ;
  assign n3731 = n2768 & ~n3730 ;
  assign n3732 = n486 & n3731 ;
  assign n3733 = n2414 ^ n389 ^ 1'b0 ;
  assign n3734 = n3732 & ~n3733 ;
  assign n3735 = n932 & n3734 ;
  assign n3736 = n2400 & n3735 ;
  assign n3737 = n574 | n599 ;
  assign n3738 = n3737 ^ n1610 ^ 1'b0 ;
  assign n3739 = n3738 ^ x247 ^ 1'b0 ;
  assign n3740 = n1917 | n2841 ;
  assign n3741 = n3710 ^ n2218 ^ 1'b0 ;
  assign n3742 = n3308 & ~n3741 ;
  assign n3743 = x97 & n1371 ;
  assign n3744 = n3743 ^ n1473 ^ 1'b0 ;
  assign n3745 = n2464 | n3744 ;
  assign n3746 = n1989 ^ n334 ^ 1'b0 ;
  assign n3747 = n302 & ~n3746 ;
  assign n3748 = ~n3078 & n3747 ;
  assign n3749 = n3457 & n3748 ;
  assign n3750 = n1911 ^ n1765 ^ 1'b0 ;
  assign n3752 = n1149 ^ n400 ^ 1'b0 ;
  assign n3753 = n1590 | n3752 ;
  assign n3751 = n1535 & ~n2623 ;
  assign n3754 = n3753 ^ n3751 ^ n1001 ;
  assign n3755 = n1499 ^ n1125 ^ n366 ;
  assign n3756 = n2485 & n3755 ;
  assign n3757 = n3756 ^ n1603 ^ 1'b0 ;
  assign n3758 = ~n327 & n2745 ;
  assign n3759 = n3758 ^ n1099 ^ 1'b0 ;
  assign n3760 = n3287 & ~n3759 ;
  assign n3761 = x80 & ~n1716 ;
  assign n3762 = ~n2502 & n3761 ;
  assign n3763 = n2868 & ~n3762 ;
  assign n3769 = n510 ^ n300 ^ 1'b0 ;
  assign n3764 = n366 & ~n771 ;
  assign n3765 = n3764 ^ x26 ^ 1'b0 ;
  assign n3766 = ( n461 & n1097 ) | ( n461 & ~n3765 ) | ( n1097 & ~n3765 ) ;
  assign n3767 = n592 & ~n1695 ;
  assign n3768 = ~n3766 & n3767 ;
  assign n3770 = n3769 ^ n3768 ^ 1'b0 ;
  assign n3771 = n1884 | n3770 ;
  assign n3772 = n1123 & n3059 ;
  assign n3773 = n2846 ^ n1105 ^ 1'b0 ;
  assign n3774 = x134 & n262 ;
  assign n3775 = n3773 & n3774 ;
  assign n3776 = n3772 & n3775 ;
  assign n3777 = ~x25 & n3776 ;
  assign n3778 = n462 | n2710 ;
  assign n3779 = x132 & ~n1034 ;
  assign n3780 = n3778 & n3779 ;
  assign n3781 = n3780 ^ x163 ^ 1'b0 ;
  assign n3782 = ~n399 & n3781 ;
  assign n3783 = ~n3761 & n3782 ;
  assign n3784 = x252 & n1660 ;
  assign n3785 = ~x175 & n3784 ;
  assign n3786 = n260 & n3785 ;
  assign n3787 = n492 & n2998 ;
  assign n3788 = n1940 & n3787 ;
  assign n3789 = x146 & ~n2286 ;
  assign n3790 = n2595 & n3789 ;
  assign n3791 = ~n932 & n1185 ;
  assign n3792 = n3791 ^ n3040 ^ 1'b0 ;
  assign n3793 = n3790 | n3792 ;
  assign n3794 = n708 & ~n1152 ;
  assign n3795 = n3794 ^ n1643 ^ 1'b0 ;
  assign n3796 = ( ~n1465 & n2216 ) | ( ~n1465 & n3551 ) | ( n2216 & n3551 ) ;
  assign n3797 = n1032 | n2286 ;
  assign n3798 = n1091 ^ x236 ^ 1'b0 ;
  assign n3799 = ~x141 & n3798 ;
  assign n3800 = ~n606 & n2593 ;
  assign n3801 = n3800 ^ x46 ^ 1'b0 ;
  assign n3802 = n2900 | n3801 ;
  assign n3803 = n1393 & n2708 ;
  assign n3804 = n1772 & n3803 ;
  assign n3805 = n3804 ^ n3151 ^ 1'b0 ;
  assign n3808 = n477 & ~n3613 ;
  assign n3809 = n3293 & n3808 ;
  assign n3806 = n1148 ^ x216 ^ 1'b0 ;
  assign n3807 = n1721 & ~n3806 ;
  assign n3810 = n3809 ^ n3807 ^ 1'b0 ;
  assign n3811 = n2542 & n3543 ;
  assign n3812 = ~n3468 & n3811 ;
  assign n3813 = x174 & n732 ;
  assign n3814 = n585 & n3813 ;
  assign n3815 = n1342 ^ n272 ^ 1'b0 ;
  assign n3816 = n3815 ^ n3723 ^ 1'b0 ;
  assign n3817 = n1454 & ~n3816 ;
  assign n3818 = n3814 | n3817 ;
  assign n3819 = n2974 ^ n1554 ^ 1'b0 ;
  assign n3820 = n2823 | n3819 ;
  assign n3821 = n3818 & ~n3820 ;
  assign n3822 = ( x27 & n779 ) | ( x27 & ~n1169 ) | ( n779 & ~n1169 ) ;
  assign n3823 = x120 | n3822 ;
  assign n3824 = n1462 ^ n905 ^ 1'b0 ;
  assign n3825 = n3823 & n3824 ;
  assign n3828 = n728 ^ n283 ^ 1'b0 ;
  assign n3826 = x178 & ~n459 ;
  assign n3827 = n2746 & ~n3826 ;
  assign n3829 = n3828 ^ n3827 ^ 1'b0 ;
  assign n3834 = n1548 ^ n935 ^ 1'b0 ;
  assign n3830 = n1317 ^ n556 ^ 1'b0 ;
  assign n3831 = n909 & n1151 ;
  assign n3832 = n3831 ^ n1638 ^ 1'b0 ;
  assign n3833 = ~n3830 & n3832 ;
  assign n3835 = n3834 ^ n3833 ^ 1'b0 ;
  assign n3836 = x76 & ~n1071 ;
  assign n3837 = n2265 & n3836 ;
  assign n3838 = n3416 | n3837 ;
  assign n3839 = ~n2101 & n3838 ;
  assign n3840 = ( n564 & n2091 ) | ( n564 & n2526 ) | ( n2091 & n2526 ) ;
  assign n3841 = n466 & n3082 ;
  assign n3842 = ~n3671 & n3841 ;
  assign n3843 = n3842 ^ n1945 ^ 1'b0 ;
  assign n3844 = ~n1385 & n2196 ;
  assign n3845 = n790 & ~n1365 ;
  assign n3846 = ~n2231 & n2622 ;
  assign n3847 = n2176 | n3846 ;
  assign n3848 = x164 | n3847 ;
  assign n3849 = n3848 ^ n3372 ^ 1'b0 ;
  assign n3850 = ~n2569 & n3849 ;
  assign n3851 = ~n640 & n2927 ;
  assign n3852 = n1377 & ~n3851 ;
  assign n3853 = n3852 ^ n769 ^ 1'b0 ;
  assign n3854 = n1665 | n2701 ;
  assign n3855 = n3854 ^ x113 ^ 1'b0 ;
  assign n3856 = n2107 & ~n2837 ;
  assign n3857 = n3855 & n3856 ;
  assign n3858 = n3857 ^ n883 ^ 1'b0 ;
  assign n3859 = n3142 ^ n2804 ^ 1'b0 ;
  assign n3860 = x56 & ~n3859 ;
  assign n3861 = ( n1614 & n3858 ) | ( n1614 & ~n3860 ) | ( n3858 & ~n3860 ) ;
  assign n3862 = n2180 ^ n1174 ^ 1'b0 ;
  assign n3863 = n1234 & n3862 ;
  assign n3864 = n1791 | n3863 ;
  assign n3865 = ~n315 & n3864 ;
  assign n3866 = ~n1027 & n3865 ;
  assign n3867 = ( n2254 & n2798 ) | ( n2254 & ~n3866 ) | ( n2798 & ~n3866 ) ;
  assign n3868 = n2506 ^ x15 ^ 1'b0 ;
  assign n3869 = n542 & ~n2062 ;
  assign n3870 = n1536 & n1813 ;
  assign n3871 = n3870 ^ n801 ^ 1'b0 ;
  assign n3872 = ~n3869 & n3871 ;
  assign n3873 = n3872 ^ n2850 ^ 1'b0 ;
  assign n3874 = n3873 ^ n2434 ^ 1'b0 ;
  assign n3875 = n1656 | n2080 ;
  assign n3876 = n1854 & ~n2674 ;
  assign n3877 = ( ~n1333 & n3242 ) | ( ~n1333 & n3368 ) | ( n3242 & n3368 ) ;
  assign n3878 = n1242 | n2944 ;
  assign n3879 = ( ~x55 & n1070 ) | ( ~x55 & n1121 ) | ( n1070 & n1121 ) ;
  assign n3880 = n3879 ^ n1803 ^ 1'b0 ;
  assign n3881 = n3880 ^ n2325 ^ 1'b0 ;
  assign n3882 = ( n1286 & ~n1311 ) | ( n1286 & n1613 ) | ( ~n1311 & n1613 ) ;
  assign n3883 = n391 & ~n1185 ;
  assign n3884 = n2011 & n3883 ;
  assign n3885 = n451 & n3884 ;
  assign n3886 = n1599 & n2008 ;
  assign n3887 = n3886 ^ x19 ^ 1'b0 ;
  assign n3888 = n2348 ^ x150 ^ 1'b0 ;
  assign n3889 = n3888 ^ n3742 ^ n486 ;
  assign n3890 = n2047 ^ n876 ^ 1'b0 ;
  assign n3891 = x187 & ~n3890 ;
  assign n3892 = n886 & n3891 ;
  assign n3893 = n3892 ^ n3511 ^ n1933 ;
  assign n3894 = ~n1912 & n2039 ;
  assign n3895 = n3894 ^ n1084 ^ 1'b0 ;
  assign n3897 = n1730 & ~n2430 ;
  assign n3898 = n3897 ^ n1748 ^ 1'b0 ;
  assign n3896 = n1931 & n2258 ;
  assign n3899 = n3898 ^ n3896 ^ 1'b0 ;
  assign n3900 = ( ~n1114 & n1680 ) | ( ~n1114 & n1736 ) | ( n1680 & n1736 ) ;
  assign n3901 = n944 & ~n3900 ;
  assign n3902 = n3901 ^ n3035 ^ 1'b0 ;
  assign n3903 = n2256 & n3902 ;
  assign n3904 = ( n2569 & ~n3098 ) | ( n2569 & n3903 ) | ( ~n3098 & n3903 ) ;
  assign n3905 = ~n1317 & n2257 ;
  assign n3906 = n1550 & n3905 ;
  assign n3907 = n1788 & ~n3906 ;
  assign n3908 = n3907 ^ n3861 ^ 1'b0 ;
  assign n3909 = n807 | n1855 ;
  assign n3910 = n2027 & ~n3909 ;
  assign n3911 = n3910 ^ n1557 ^ 1'b0 ;
  assign n3912 = n3911 ^ n3119 ^ 1'b0 ;
  assign n3913 = n3225 ^ n1851 ^ 1'b0 ;
  assign n3914 = x61 & ~n2022 ;
  assign n3915 = n3914 ^ n262 ^ 1'b0 ;
  assign n3916 = n1366 & ~n1699 ;
  assign n3917 = n3916 ^ n880 ^ 1'b0 ;
  assign n3918 = x30 | n3917 ;
  assign n3919 = ~n2771 & n3747 ;
  assign n3920 = n281 & n3919 ;
  assign n3921 = n1539 | n3920 ;
  assign n3922 = n2150 | n3921 ;
  assign n3923 = n3922 ^ n1057 ^ 1'b0 ;
  assign n3924 = n449 & ~n3923 ;
  assign n3925 = n3918 & n3924 ;
  assign n3926 = ( x176 & ~n1734 ) | ( x176 & n1782 ) | ( ~n1734 & n1782 ) ;
  assign n3927 = n3926 ^ n2383 ^ 1'b0 ;
  assign n3928 = ~n3815 & n3927 ;
  assign n3929 = n3928 ^ n3922 ^ n2143 ;
  assign n3930 = n3925 | n3929 ;
  assign n3931 = n848 ^ x252 ^ 1'b0 ;
  assign n3932 = n3931 ^ n3011 ^ 1'b0 ;
  assign n3933 = n2287 ^ n2113 ^ n289 ;
  assign n3934 = n3932 & n3933 ;
  assign n3935 = n1048 & ~n2501 ;
  assign n3936 = n2190 ^ n1815 ^ n298 ;
  assign n3937 = n2354 ^ n1846 ^ 1'b0 ;
  assign n3938 = n2778 | n3937 ;
  assign n3939 = n3938 ^ n3245 ^ n2508 ;
  assign n3942 = ~n1397 & n1490 ;
  assign n3943 = n3942 ^ n3588 ^ 1'b0 ;
  assign n3944 = n1151 & ~n3943 ;
  assign n3940 = n1100 | n3250 ;
  assign n3941 = n3940 ^ n1680 ^ 1'b0 ;
  assign n3945 = n3944 ^ n3941 ^ 1'b0 ;
  assign n3946 = ~n1535 & n3886 ;
  assign n3947 = ( ~n774 & n2576 ) | ( ~n774 & n2889 ) | ( n2576 & n2889 ) ;
  assign n3948 = n3042 ^ n2827 ^ x139 ;
  assign n3949 = n3948 ^ n2887 ^ 1'b0 ;
  assign n3950 = n3947 & n3949 ;
  assign n3951 = n2950 ^ n1142 ^ 1'b0 ;
  assign n3952 = ( n1982 & n2958 ) | ( n1982 & n3951 ) | ( n2958 & n3951 ) ;
  assign n3953 = n1036 ^ x84 ^ 1'b0 ;
  assign n3954 = n786 & ~n3953 ;
  assign n3955 = x18 & n3954 ;
  assign n3956 = n1324 & n3955 ;
  assign n3957 = x212 | n3956 ;
  assign n3958 = ~n711 & n1796 ;
  assign n3959 = n894 | n1259 ;
  assign n3960 = n3223 ^ n2235 ^ 1'b0 ;
  assign n3961 = n3959 & ~n3960 ;
  assign n3962 = n1223 ^ n466 ^ 1'b0 ;
  assign n3963 = ( n3174 & ~n3961 ) | ( n3174 & n3962 ) | ( ~n3961 & n3962 ) ;
  assign n3964 = n1676 ^ n961 ^ n442 ;
  assign n3965 = n1901 & ~n3964 ;
  assign n3966 = n3965 ^ n1267 ^ 1'b0 ;
  assign n3967 = n1826 | n3357 ;
  assign n3968 = x79 & ~n2464 ;
  assign n3969 = n3968 ^ n2571 ^ 1'b0 ;
  assign n3970 = n2103 | n2714 ;
  assign n3971 = x238 & ~n3970 ;
  assign n3972 = n550 & n3971 ;
  assign n3973 = n3481 ^ n1731 ^ 1'b0 ;
  assign n3974 = n3973 ^ n3863 ^ n2827 ;
  assign n3975 = n3974 ^ n3410 ^ 1'b0 ;
  assign n3976 = n279 & n2433 ;
  assign n3977 = n3976 ^ n1060 ^ 1'b0 ;
  assign n3978 = n2725 ^ n2358 ^ x108 ;
  assign n3979 = n862 & ~n872 ;
  assign n3980 = ~x132 & n3979 ;
  assign n3981 = n3980 ^ n3116 ^ 1'b0 ;
  assign n3982 = ( n2739 & n3005 ) | ( n2739 & ~n3134 ) | ( n3005 & ~n3134 ) ;
  assign n3983 = n3974 ^ n1163 ^ 1'b0 ;
  assign n3984 = n828 | n3983 ;
  assign n3985 = n2526 ^ n2464 ^ n2248 ;
  assign n3992 = n3879 ^ n1276 ^ 1'b0 ;
  assign n3993 = n707 & ~n3992 ;
  assign n3986 = n1073 ^ x84 ^ 1'b0 ;
  assign n3987 = x40 & ~n264 ;
  assign n3988 = n3987 ^ x223 ^ 1'b0 ;
  assign n3989 = n1037 & ~n3988 ;
  assign n3990 = n1416 & n3989 ;
  assign n3991 = n3986 | n3990 ;
  assign n3994 = n3993 ^ n3991 ^ 1'b0 ;
  assign n3995 = ~n1994 & n3994 ;
  assign n3996 = n3995 ^ n2641 ^ 1'b0 ;
  assign n3997 = n2749 ^ n2319 ^ 1'b0 ;
  assign n3998 = n3997 ^ n2307 ^ 1'b0 ;
  assign n3999 = n1230 & ~n3998 ;
  assign n4000 = n2803 | n2967 ;
  assign n4001 = n4000 ^ x128 ^ 1'b0 ;
  assign n4002 = x14 & ~n475 ;
  assign n4003 = n2161 & n4002 ;
  assign n4004 = ~n776 & n4003 ;
  assign n4005 = n4004 ^ n2504 ^ 1'b0 ;
  assign n4007 = n2687 & n3607 ;
  assign n4008 = n4007 ^ n3532 ^ 1'b0 ;
  assign n4006 = n1922 & n2089 ;
  assign n4009 = n4008 ^ n4006 ^ 1'b0 ;
  assign n4012 = n391 & ~n1259 ;
  assign n4013 = n4012 ^ n813 ^ 1'b0 ;
  assign n4011 = ~n469 & n1651 ;
  assign n4010 = n1856 | n2502 ;
  assign n4014 = n4013 ^ n4011 ^ n4010 ;
  assign n4015 = ~n710 & n1606 ;
  assign n4016 = n2047 & n4015 ;
  assign n4017 = n933 & n1168 ;
  assign n4018 = n4016 & n4017 ;
  assign n4019 = n3431 ^ n1098 ^ 1'b0 ;
  assign n4020 = ( n2927 & ~n3296 ) | ( n2927 & n4019 ) | ( ~n3296 & n4019 ) ;
  assign n4021 = n446 ^ n436 ^ x239 ;
  assign n4022 = n4021 ^ n1278 ^ 1'b0 ;
  assign n4023 = x81 & ~n4022 ;
  assign n4024 = x201 & ~n399 ;
  assign n4025 = ~x104 & n4024 ;
  assign n4026 = x74 | n4025 ;
  assign n4027 = ( n691 & n1969 ) | ( n691 & n4026 ) | ( n1969 & n4026 ) ;
  assign n4028 = n4027 ^ x215 ^ 1'b0 ;
  assign n4029 = n1172 | n4028 ;
  assign n4030 = n4029 ^ x186 ^ 1'b0 ;
  assign n4031 = n1623 | n4030 ;
  assign n4032 = n4031 ^ n2990 ^ 1'b0 ;
  assign n4033 = ~x73 & x151 ;
  assign n4034 = n4033 ^ n1144 ^ 1'b0 ;
  assign n4035 = n1088 & n4034 ;
  assign n4036 = n4035 ^ n1820 ^ 1'b0 ;
  assign n4037 = ~n4003 & n4036 ;
  assign n4038 = n850 & ~n2963 ;
  assign n4039 = n1374 | n4038 ;
  assign n4040 = ~n2395 & n4039 ;
  assign n4041 = n842 & ~n3555 ;
  assign n4042 = n4041 ^ n1001 ^ 1'b0 ;
  assign n4043 = n553 & n916 ;
  assign n4044 = ~n1290 & n4043 ;
  assign n4045 = n1742 | n4044 ;
  assign n4046 = n260 & n291 ;
  assign n4047 = n2593 | n2975 ;
  assign n4051 = n1125 ^ x75 ^ 1'b0 ;
  assign n4052 = n3863 & n4051 ;
  assign n4053 = n4052 ^ n1070 ^ 1'b0 ;
  assign n4054 = n1809 | n4053 ;
  assign n4055 = n4054 ^ n618 ^ 1'b0 ;
  assign n4056 = n1073 ^ x22 ^ 1'b0 ;
  assign n4057 = n1969 ^ n1914 ^ 1'b0 ;
  assign n4058 = n1413 & ~n4057 ;
  assign n4059 = n395 & n4058 ;
  assign n4060 = n4056 & ~n4059 ;
  assign n4061 = ~n4055 & n4060 ;
  assign n4048 = x252 & n1312 ;
  assign n4049 = n4048 ^ n1001 ^ 1'b0 ;
  assign n4050 = ( n2211 & n3954 ) | ( n2211 & ~n4049 ) | ( n3954 & ~n4049 ) ;
  assign n4062 = n4061 ^ n4050 ^ 1'b0 ;
  assign n4064 = n1826 | n3114 ;
  assign n4065 = n1928 & ~n4064 ;
  assign n4063 = n2629 & n3887 ;
  assign n4066 = n4065 ^ n4063 ^ 1'b0 ;
  assign n4067 = ( n475 & n547 ) | ( n475 & n1894 ) | ( n547 & n1894 ) ;
  assign n4068 = n647 & n3453 ;
  assign n4069 = ~n1688 & n4068 ;
  assign n4070 = x40 & n4069 ;
  assign n4071 = n2507 ^ n1415 ^ 1'b0 ;
  assign n4072 = n2508 & ~n4071 ;
  assign n4073 = n1887 & n4072 ;
  assign n4074 = ~n4070 & n4073 ;
  assign n4075 = n1741 ^ n1028 ^ 1'b0 ;
  assign n4076 = n3795 | n4075 ;
  assign n4077 = n3313 & ~n4076 ;
  assign n4078 = n4077 ^ n2787 ^ 1'b0 ;
  assign n4079 = n4078 ^ n2269 ^ 1'b0 ;
  assign n4080 = ~n4074 & n4079 ;
  assign n4081 = n897 | n1382 ;
  assign n4082 = n3521 & ~n4081 ;
  assign n4083 = n3037 | n4082 ;
  assign n4087 = n4003 ^ x34 ^ 1'b0 ;
  assign n4088 = n1172 | n4087 ;
  assign n4084 = n657 | n817 ;
  assign n4085 = n3464 & n4084 ;
  assign n4086 = n4085 ^ n899 ^ 1'b0 ;
  assign n4089 = n4088 ^ n4086 ^ 1'b0 ;
  assign n4090 = ~n1073 & n4089 ;
  assign n4091 = ( n1926 & n2788 ) | ( n1926 & ~n4090 ) | ( n2788 & ~n4090 ) ;
  assign n4092 = n3801 ^ n2208 ^ n1039 ;
  assign n4093 = n2452 ^ n740 ^ 1'b0 ;
  assign n4094 = n2644 & n3203 ;
  assign n4095 = n4094 ^ x215 ^ 1'b0 ;
  assign n4096 = n2230 | n3333 ;
  assign n4097 = n291 & n2622 ;
  assign n4098 = n1980 & ~n2569 ;
  assign n4099 = ~n4097 & n4098 ;
  assign n4100 = n4099 ^ n1441 ^ 1'b0 ;
  assign n4101 = n4100 ^ n1647 ^ 1'b0 ;
  assign n4102 = ~n1720 & n4101 ;
  assign n4103 = n3191 ^ n2679 ^ 1'b0 ;
  assign n4104 = n1980 & n4103 ;
  assign n4105 = n4104 ^ n1362 ^ 1'b0 ;
  assign n4107 = n1851 ^ x231 ^ 1'b0 ;
  assign n4106 = n1665 | n3472 ;
  assign n4108 = n4107 ^ n4106 ^ 1'b0 ;
  assign n4109 = ( n944 & ~n3007 ) | ( n944 & n4108 ) | ( ~n3007 & n4108 ) ;
  assign n4112 = ~n498 & n3253 ;
  assign n4113 = n4112 ^ n953 ^ 1'b0 ;
  assign n4110 = n956 ^ n635 ^ 1'b0 ;
  assign n4111 = ~n1422 & n4110 ;
  assign n4114 = n4113 ^ n4111 ^ 1'b0 ;
  assign n4115 = n4114 ^ n1730 ^ x246 ;
  assign n4116 = n3372 & n4115 ;
  assign n4117 = ~n4109 & n4116 ;
  assign n4118 = n1802 & n3766 ;
  assign n4119 = n466 & n4118 ;
  assign n4120 = x92 & n1121 ;
  assign n4121 = n4120 ^ n1292 ^ 1'b0 ;
  assign n4122 = n3091 & n4121 ;
  assign n4123 = n3091 ^ n907 ^ 1'b0 ;
  assign n4124 = n992 ^ n625 ^ 1'b0 ;
  assign n4125 = n2576 & ~n4124 ;
  assign n4126 = ~n1340 & n1593 ;
  assign n4127 = n2331 & n4126 ;
  assign n4128 = n4127 ^ n3486 ^ 1'b0 ;
  assign n4129 = x124 & ~n369 ;
  assign n4130 = n4129 ^ n428 ^ 1'b0 ;
  assign n4131 = n4130 ^ n1080 ^ 1'b0 ;
  assign n4132 = n4131 ^ n3801 ^ n3367 ;
  assign n4133 = n1590 | n3400 ;
  assign n4134 = n4132 | n4133 ;
  assign n4135 = n3951 & ~n4134 ;
  assign n4136 = n2203 | n2890 ;
  assign n4137 = x237 & n1134 ;
  assign n4138 = n4137 ^ x138 ^ 1'b0 ;
  assign n4139 = ( n933 & ~n1585 ) | ( n933 & n2122 ) | ( ~n1585 & n2122 ) ;
  assign n4140 = n3248 ^ n2183 ^ 1'b0 ;
  assign n4141 = n1123 & n4140 ;
  assign n4142 = ~n3614 & n4141 ;
  assign n4143 = n1891 ^ n1321 ^ 1'b0 ;
  assign n4144 = ~n3990 & n4143 ;
  assign n4145 = ( ~n1600 & n3470 ) | ( ~n1600 & n3573 ) | ( n3470 & n3573 ) ;
  assign n4146 = ( ~n1398 & n1801 ) | ( ~n1398 & n3423 ) | ( n1801 & n3423 ) ;
  assign n4147 = n1238 & n1318 ;
  assign n4148 = n4147 ^ n3401 ^ 1'b0 ;
  assign n4149 = n2178 & ~n3771 ;
  assign n4150 = ( x68 & ~n634 ) | ( x68 & n2547 ) | ( ~n634 & n2547 ) ;
  assign n4151 = n2696 | n4150 ;
  assign n4152 = n1180 | n4151 ;
  assign n4153 = x114 | n2122 ;
  assign n4154 = ~n1249 & n4153 ;
  assign n4160 = x170 & n2465 ;
  assign n4161 = n1200 & n4160 ;
  assign n4155 = n2716 ^ n348 ^ 1'b0 ;
  assign n4156 = n486 & n675 ;
  assign n4157 = n4156 ^ n367 ^ 1'b0 ;
  assign n4158 = ~n3360 & n4157 ;
  assign n4159 = ~n4155 & n4158 ;
  assign n4162 = n4161 ^ n4159 ^ 1'b0 ;
  assign n4163 = ~n4154 & n4162 ;
  assign n4164 = ~n256 & n4163 ;
  assign n4165 = n1200 & n4164 ;
  assign n4166 = n537 & n3196 ;
  assign n4167 = ~n542 & n2655 ;
  assign n4168 = n1801 & n4167 ;
  assign n4169 = ~n673 & n4168 ;
  assign n4170 = n4169 ^ n3693 ^ n1422 ;
  assign n4171 = ~n3333 & n4170 ;
  assign n4172 = n4171 ^ n2184 ^ 1'b0 ;
  assign n4173 = n747 & ~n1993 ;
  assign n4174 = ( n1290 & ~n2224 ) | ( n1290 & n4173 ) | ( ~n2224 & n4173 ) ;
  assign n4175 = n3074 & n4174 ;
  assign n4176 = n2274 & ~n2730 ;
  assign n4177 = n4176 ^ n3098 ^ 1'b0 ;
  assign n4178 = n4177 ^ n3156 ^ n1261 ;
  assign n4179 = n1048 & n1230 ;
  assign n4180 = n4179 ^ n2382 ^ 1'b0 ;
  assign n4181 = n2392 ^ n2177 ^ n1457 ;
  assign n4182 = x36 | n4181 ;
  assign n4183 = n3831 & ~n4182 ;
  assign n4184 = n4183 ^ n3999 ^ 1'b0 ;
  assign n4185 = n3668 ^ n1491 ^ n963 ;
  assign n4186 = n2162 ^ n1027 ^ 1'b0 ;
  assign n4187 = x201 & n1062 ;
  assign n4188 = n1111 & ~n1809 ;
  assign n4189 = n2743 & n4188 ;
  assign n4190 = n1671 | n2785 ;
  assign n4191 = n1071 | n4190 ;
  assign n4192 = n4191 ^ n814 ^ 1'b0 ;
  assign n4193 = n3206 ^ n618 ^ 1'b0 ;
  assign n4194 = ~n905 & n2007 ;
  assign n4195 = ~n4010 & n4194 ;
  assign n4196 = n4195 ^ n1551 ^ n274 ;
  assign n4197 = n1500 & ~n3744 ;
  assign n4198 = x143 & ~n525 ;
  assign n4199 = n1653 ^ n1043 ^ 1'b0 ;
  assign n4200 = n4198 | n4199 ;
  assign n4201 = n1457 & ~n4200 ;
  assign n4202 = n4197 & n4201 ;
  assign n4203 = ~n1002 & n1098 ;
  assign n4204 = n2320 ^ n1632 ^ n1409 ;
  assign n4205 = n2788 & ~n4204 ;
  assign n4206 = n1495 & ~n4205 ;
  assign n4207 = n1333 ^ x155 ^ 1'b0 ;
  assign n4208 = n1142 | n1938 ;
  assign n4209 = ( ~n966 & n1776 ) | ( ~n966 & n2710 ) | ( n1776 & n2710 ) ;
  assign n4210 = n1752 | n2400 ;
  assign n4211 = n4210 ^ x107 ^ 1'b0 ;
  assign n4212 = n3886 & n4211 ;
  assign n4213 = n872 ^ n268 ^ x65 ;
  assign n4214 = n369 | n4213 ;
  assign n4215 = x67 & ~n923 ;
  assign n4216 = x38 ^ x8 ^ 1'b0 ;
  assign n4217 = n4216 ^ n991 ^ 1'b0 ;
  assign n4218 = n2164 & n4217 ;
  assign n4219 = n2974 & ~n4218 ;
  assign n4220 = ( n679 & n2190 ) | ( n679 & ~n4219 ) | ( n2190 & ~n4219 ) ;
  assign n4221 = n4215 & n4220 ;
  assign n4222 = n2234 & n4221 ;
  assign n4224 = n2699 & n3287 ;
  assign n4225 = n1671 & n4224 ;
  assign n4226 = n4225 ^ n2576 ^ n1877 ;
  assign n4223 = n863 | n1468 ;
  assign n4227 = n4226 ^ n4223 ^ 1'b0 ;
  assign n4228 = n3041 & ~n3888 ;
  assign n4229 = n4228 ^ n3908 ^ 1'b0 ;
  assign n4230 = n1060 ^ n277 ^ 1'b0 ;
  assign n4231 = n1085 & n2329 ;
  assign n4232 = ~n1496 & n4231 ;
  assign n4233 = n4232 ^ x231 ^ 1'b0 ;
  assign n4234 = n900 & ~n4233 ;
  assign n4235 = n3821 & n4234 ;
  assign n4236 = ~n4230 & n4235 ;
  assign n4237 = n4050 ^ n1255 ^ 1'b0 ;
  assign n4238 = ~n1519 & n4237 ;
  assign n4239 = x203 & n1877 ;
  assign n4240 = n4239 ^ n2320 ^ 1'b0 ;
  assign n4241 = n2530 ^ n1441 ^ 1'b0 ;
  assign n4242 = ~n1544 & n4241 ;
  assign n4243 = n4242 ^ n1867 ^ 1'b0 ;
  assign n4244 = n4240 & ~n4243 ;
  assign n4245 = x152 & ~n3954 ;
  assign n4246 = x143 & x150 ;
  assign n4247 = ~n4245 & n4246 ;
  assign n4248 = n2274 & n4247 ;
  assign n4249 = ( x48 & ~x132 ) | ( x48 & n2615 ) | ( ~x132 & n2615 ) ;
  assign n4250 = n3196 ^ n814 ^ 1'b0 ;
  assign n4251 = ~n1804 & n4250 ;
  assign n4252 = n4251 ^ n4240 ^ 1'b0 ;
  assign n4256 = n2560 ^ n1428 ^ 1'b0 ;
  assign n4253 = n1048 & n2133 ;
  assign n4254 = n4253 ^ n3147 ^ x60 ;
  assign n4255 = n4254 ^ n1682 ^ 1'b0 ;
  assign n4257 = n4256 ^ n4255 ^ n3814 ;
  assign n4258 = x178 ^ x2 ^ 1'b0 ;
  assign n4259 = ( n1639 & n1680 ) | ( n1639 & n4258 ) | ( n1680 & n4258 ) ;
  assign n4260 = n3754 ^ n2544 ^ n592 ;
  assign n4261 = n1192 ^ n481 ^ 1'b0 ;
  assign n4262 = n2868 ^ n2187 ^ 1'b0 ;
  assign n4263 = n776 | n4262 ;
  assign n4264 = n2250 ^ n634 ^ n440 ;
  assign n4265 = n4263 | n4264 ;
  assign n4266 = n4261 | n4265 ;
  assign n4267 = ( n2127 & n3978 ) | ( n2127 & n4266 ) | ( n3978 & n4266 ) ;
  assign n4268 = n4260 & n4267 ;
  assign n4269 = x125 & ~n2984 ;
  assign n4270 = ( n464 & n2883 ) | ( n464 & n4269 ) | ( n2883 & n4269 ) ;
  assign n4272 = n671 & n1174 ;
  assign n4273 = n4272 ^ n540 ^ 1'b0 ;
  assign n4274 = n3388 & ~n4273 ;
  assign n4275 = n709 & n4274 ;
  assign n4271 = ( n2472 & n3150 ) | ( n2472 & ~n3724 ) | ( n3150 & ~n3724 ) ;
  assign n4276 = n4275 ^ n4271 ^ 1'b0 ;
  assign n4277 = n1215 | n1219 ;
  assign n4278 = n3521 ^ n1192 ^ 1'b0 ;
  assign n4279 = ~n614 & n4278 ;
  assign n4280 = ( ~n3182 & n4277 ) | ( ~n3182 & n4279 ) | ( n4277 & n4279 ) ;
  assign n4281 = n342 | n2554 ;
  assign n4282 = n2001 & ~n4281 ;
  assign n4283 = n1032 & ~n4282 ;
  assign n4284 = n1069 & n4283 ;
  assign n4285 = n2823 & ~n3396 ;
  assign n4286 = n4166 & n4285 ;
  assign n4287 = n2785 ^ n638 ^ 1'b0 ;
  assign n4288 = n2620 ^ n628 ^ 1'b0 ;
  assign n4289 = n3070 ^ n1620 ^ 1'b0 ;
  assign n4290 = n1954 | n4289 ;
  assign n4291 = n357 & ~n4290 ;
  assign n4292 = ~x242 & n4291 ;
  assign n4293 = n1001 & n3203 ;
  assign n4294 = n4293 ^ n2408 ^ 1'b0 ;
  assign n4295 = n638 & n1175 ;
  assign n4296 = n3670 ^ n2403 ^ n258 ;
  assign n4297 = n871 | n2265 ;
  assign n4298 = n4297 ^ n3523 ^ 1'b0 ;
  assign n4299 = n983 | n3134 ;
  assign n4300 = n2035 & ~n4299 ;
  assign n4301 = ( ~n1462 & n2770 ) | ( ~n1462 & n2936 ) | ( n2770 & n2936 ) ;
  assign n4302 = n4301 ^ n3839 ^ 1'b0 ;
  assign n4303 = n3546 ^ n840 ^ 1'b0 ;
  assign n4304 = n2856 & ~n4117 ;
  assign n4305 = n4304 ^ x176 ^ 1'b0 ;
  assign n4306 = ( x181 & n789 ) | ( x181 & ~n4065 ) | ( n789 & ~n4065 ) ;
  assign n4307 = ( n374 & n1161 ) | ( n374 & n2194 ) | ( n1161 & n2194 ) ;
  assign n4308 = n4307 ^ n1848 ^ 1'b0 ;
  assign n4309 = ~n759 & n4308 ;
  assign n4313 = ( x115 & ~n1910 ) | ( x115 & n4232 ) | ( ~n1910 & n4232 ) ;
  assign n4314 = n4313 ^ n2926 ^ 1'b0 ;
  assign n4315 = ~n2993 & n4314 ;
  assign n4310 = n1692 | n1867 ;
  assign n4311 = n896 & ~n4310 ;
  assign n4312 = n523 & n4311 ;
  assign n4316 = n4315 ^ n4312 ^ 1'b0 ;
  assign n4317 = n2214 ^ x246 ^ 1'b0 ;
  assign n4318 = ~n2387 & n2801 ;
  assign n4319 = ~n917 & n4318 ;
  assign n4320 = n1259 | n4319 ;
  assign n4321 = n4320 ^ n2623 ^ 1'b0 ;
  assign n4322 = n3012 ^ x173 ^ 1'b0 ;
  assign n4323 = n409 & ~n4322 ;
  assign n4324 = n1039 ^ n571 ^ 1'b0 ;
  assign n4325 = n1588 & ~n4324 ;
  assign n4326 = n2719 | n4325 ;
  assign n4327 = ~n2585 & n3346 ;
  assign n4328 = n1653 & ~n4327 ;
  assign n4329 = x118 & ~n4328 ;
  assign n4330 = n957 | n4329 ;
  assign n4331 = n4330 ^ n2466 ^ 1'b0 ;
  assign n4332 = n3100 ^ n1985 ^ 1'b0 ;
  assign n4333 = n4331 | n4332 ;
  assign n4334 = x225 & n3951 ;
  assign n4335 = n4334 ^ n746 ^ 1'b0 ;
  assign n4336 = n2846 ^ n1756 ^ 1'b0 ;
  assign n4337 = n3491 & n4336 ;
  assign n4338 = n4337 ^ n4150 ^ n1151 ;
  assign n4340 = n503 & n1482 ;
  assign n4339 = n1489 | n2267 ;
  assign n4341 = n4340 ^ n4339 ^ 1'b0 ;
  assign n4342 = n2215 & n2819 ;
  assign n4343 = n3509 & ~n3828 ;
  assign n4344 = n2372 & ~n3047 ;
  assign n4345 = n4344 ^ n2469 ^ 1'b0 ;
  assign n4346 = n4345 ^ n3574 ^ 1'b0 ;
  assign n4347 = n2086 ^ n1828 ^ 1'b0 ;
  assign n4348 = n4347 ^ n3014 ^ n2378 ;
  assign n4349 = n2215 | n4348 ;
  assign n4350 = n4349 ^ n1167 ^ 1'b0 ;
  assign n4351 = ~n4316 & n4350 ;
  assign n4352 = n4351 ^ n3939 ^ 1'b0 ;
  assign n4353 = n2224 ^ x207 ^ 1'b0 ;
  assign n4354 = ~n3923 & n4353 ;
  assign n4355 = n4354 ^ n3317 ^ n2670 ;
  assign n4356 = ~n2679 & n3142 ;
  assign n4359 = ~n276 & n2047 ;
  assign n4357 = n801 & n2056 ;
  assign n4358 = n2317 & n4357 ;
  assign n4360 = n4359 ^ n4358 ^ 1'b0 ;
  assign n4361 = n2544 & n3260 ;
  assign n4362 = n4361 ^ n3663 ^ 1'b0 ;
  assign n4363 = n3829 & n4362 ;
  assign n4364 = ( ~n1303 & n4360 ) | ( ~n1303 & n4363 ) | ( n4360 & n4363 ) ;
  assign n4365 = n2106 | n4130 ;
  assign n4366 = n920 | n4365 ;
  assign n4367 = n4366 ^ n3001 ^ n2805 ;
  assign n4368 = ( n1148 & ~n3178 ) | ( n1148 & n4367 ) | ( ~n3178 & n4367 ) ;
  assign n4369 = n2631 ^ n1873 ^ x105 ;
  assign n4370 = n2858 ^ n1112 ^ 1'b0 ;
  assign n4371 = ~n842 & n1802 ;
  assign n4372 = n3319 & n4371 ;
  assign n4373 = n1121 & ~n2161 ;
  assign n4374 = n761 & n4373 ;
  assign n4375 = n4374 ^ n3890 ^ 1'b0 ;
  assign n4376 = n2844 ^ x157 ^ 1'b0 ;
  assign n4377 = n372 | n4376 ;
  assign n4378 = n2165 & ~n4377 ;
  assign n4379 = n4375 & n4378 ;
  assign n4380 = n3007 ^ n880 ^ 1'b0 ;
  assign n4381 = ~x107 & x252 ;
  assign n4382 = x193 & ~n603 ;
  assign n4383 = n4382 ^ n2485 ^ 1'b0 ;
  assign n4384 = n1763 & n2694 ;
  assign n4385 = n1244 ^ x32 ^ 1'b0 ;
  assign n4386 = x247 & ~n4385 ;
  assign n4387 = ( ~n445 & n3611 ) | ( ~n445 & n3877 ) | ( n3611 & n3877 ) ;
  assign n4388 = x198 & ~n718 ;
  assign n4389 = n1283 | n1975 ;
  assign n4390 = ~n4388 & n4389 ;
  assign n4391 = n4390 ^ n2904 ^ 1'b0 ;
  assign n4392 = n3640 | n4046 ;
  assign n4393 = n384 & ~n4392 ;
  assign n4394 = n1989 & ~n2712 ;
  assign n4395 = ~n294 & n4394 ;
  assign n4396 = n930 ^ x200 ^ 1'b0 ;
  assign n4397 = ~n3470 & n4396 ;
  assign n4398 = ~n574 & n1915 ;
  assign n4399 = n1547 & n4398 ;
  assign n4400 = n998 & ~n4399 ;
  assign n4401 = n4400 ^ n3027 ^ 1'b0 ;
  assign n4402 = n394 & n4401 ;
  assign n4403 = n4402 ^ x221 ^ 1'b0 ;
  assign n4404 = ~n4397 & n4403 ;
  assign n4405 = ~n1206 & n4150 ;
  assign n4406 = n845 & n4405 ;
  assign n4407 = n4406 ^ x187 ^ 1'b0 ;
  assign n4408 = n1168 & n1581 ;
  assign n4409 = ~n1133 & n4408 ;
  assign n4410 = n4409 ^ n2128 ^ n1710 ;
  assign n4411 = ~n2464 & n4410 ;
  assign n4412 = n2468 & n4397 ;
  assign n4413 = n4412 ^ n2001 ^ 1'b0 ;
  assign n4414 = n4394 ^ n3817 ^ 1'b0 ;
  assign n4415 = n4413 & n4414 ;
  assign n4416 = ~n1167 & n4415 ;
  assign n4417 = n710 & ~n1689 ;
  assign n4418 = ~n2264 & n3216 ;
  assign n4419 = n4418 ^ n357 ^ 1'b0 ;
  assign n4420 = ~n1940 & n4419 ;
  assign n4421 = n2040 | n2549 ;
  assign n4422 = n4421 ^ n486 ^ 1'b0 ;
  assign n4423 = x52 & n4422 ;
  assign n4424 = n4423 ^ n2654 ^ 1'b0 ;
  assign n4425 = n634 & ~n2389 ;
  assign n4426 = n1819 & n3359 ;
  assign n4427 = n4426 ^ n462 ^ 1'b0 ;
  assign n4428 = n2801 & n4427 ;
  assign n4429 = n3454 & ~n3938 ;
  assign n4430 = n376 & n4429 ;
  assign n4431 = n1135 | n4430 ;
  assign n4432 = n1513 & ~n4431 ;
  assign n4433 = n4432 ^ x212 ^ 1'b0 ;
  assign n4435 = ~n710 & n1433 ;
  assign n4436 = n4435 ^ n1151 ^ 1'b0 ;
  assign n4434 = n1119 | n1899 ;
  assign n4437 = n4436 ^ n4434 ^ n2812 ;
  assign n4438 = n2693 | n3005 ;
  assign n4439 = n3537 ^ n2706 ^ 1'b0 ;
  assign n4440 = n1756 & n3568 ;
  assign n4441 = n4440 ^ n1318 ^ 1'b0 ;
  assign n4442 = n1391 & ~n4441 ;
  assign n4443 = n2105 ^ x243 ^ 1'b0 ;
  assign n4444 = n2592 & n4443 ;
  assign n4445 = n4444 ^ n4150 ^ 1'b0 ;
  assign n4448 = n2010 ^ n328 ^ 1'b0 ;
  assign n4449 = n262 & ~n4448 ;
  assign n4450 = n4449 ^ n2410 ^ 1'b0 ;
  assign n4446 = n810 ^ x248 ^ 1'b0 ;
  assign n4447 = n4366 & ~n4446 ;
  assign n4451 = n4450 ^ n4447 ^ 1'b0 ;
  assign n4452 = ( n2264 & n4445 ) | ( n2264 & n4451 ) | ( n4445 & n4451 ) ;
  assign n4453 = n1606 ^ n1419 ^ n263 ;
  assign n4454 = x25 & n4453 ;
  assign n4455 = n1080 ^ n651 ^ 1'b0 ;
  assign n4456 = x72 & ~n4455 ;
  assign n4457 = x115 & ~n518 ;
  assign n4458 = n4457 ^ n2218 ^ 1'b0 ;
  assign n4459 = n2719 & n4458 ;
  assign n4460 = n3296 ^ n739 ^ 1'b0 ;
  assign n4461 = x13 & ~n2782 ;
  assign n4462 = n4461 ^ n1240 ^ 1'b0 ;
  assign n4463 = n1714 & ~n4462 ;
  assign n4464 = n642 | n2693 ;
  assign n4465 = n4464 ^ n2468 ^ 1'b0 ;
  assign n4466 = n2426 | n4019 ;
  assign n4467 = ~n3266 & n4466 ;
  assign n4468 = n4467 ^ n2443 ^ 1'b0 ;
  assign n4469 = n4468 ^ n2613 ^ 1'b0 ;
  assign n4470 = n4465 & n4469 ;
  assign n4471 = n984 & n1484 ;
  assign n4472 = n4471 ^ n485 ^ 1'b0 ;
  assign n4473 = n3461 ^ n550 ^ 1'b0 ;
  assign n4474 = n4472 | n4473 ;
  assign n4475 = n971 ^ n423 ^ 1'b0 ;
  assign n4476 = n1519 & ~n4475 ;
  assign n4477 = n2850 ^ n651 ^ 1'b0 ;
  assign n4478 = ~n2450 & n4477 ;
  assign n4479 = n1784 & ~n2218 ;
  assign n4480 = ~n1197 & n4479 ;
  assign n4481 = n4480 ^ n4225 ^ 1'b0 ;
  assign n4482 = n2093 ^ n877 ^ 1'b0 ;
  assign n4484 = n604 & ~n2718 ;
  assign n4483 = n485 | n2433 ;
  assign n4485 = n4484 ^ n4483 ^ 1'b0 ;
  assign n4486 = n4485 ^ n1968 ^ 1'b0 ;
  assign n4487 = n2109 | n4486 ;
  assign n4488 = n3140 ^ n1521 ^ 1'b0 ;
  assign n4496 = n3601 ^ n3152 ^ 1'b0 ;
  assign n4489 = n1471 ^ n1292 ^ 1'b0 ;
  assign n4490 = n1276 | n2763 ;
  assign n4491 = n4489 & ~n4490 ;
  assign n4492 = n1720 | n4491 ;
  assign n4493 = n2338 & ~n4492 ;
  assign n4494 = n2875 | n4493 ;
  assign n4495 = n4005 & n4494 ;
  assign n4497 = n4496 ^ n4495 ^ 1'b0 ;
  assign n4498 = n4121 ^ n1424 ^ 1'b0 ;
  assign n4499 = n973 & ~n1208 ;
  assign n4500 = n4499 ^ n1960 ^ 1'b0 ;
  assign n4501 = ~n2210 & n2830 ;
  assign n4502 = x171 & ~n1841 ;
  assign n4503 = n4107 & ~n4502 ;
  assign n4504 = n4503 ^ n2582 ^ 1'b0 ;
  assign n4505 = n3307 | n4504 ;
  assign n4506 = ~n3333 & n4505 ;
  assign n4507 = n510 & ~n889 ;
  assign n4508 = n4507 ^ x94 ^ 1'b0 ;
  assign n4509 = n672 & ~n4508 ;
  assign n4510 = n2946 ^ n2663 ^ n1039 ;
  assign n4511 = n2984 ^ n1854 ^ 1'b0 ;
  assign n4512 = n4511 ^ n608 ^ n424 ;
  assign n4513 = n3751 ^ n1775 ^ 1'b0 ;
  assign n4514 = ~n4512 & n4513 ;
  assign n4515 = n2383 & ~n2752 ;
  assign n4516 = n1952 | n4515 ;
  assign n4517 = n2140 ^ x185 ^ 1'b0 ;
  assign n4518 = n1351 | n4517 ;
  assign n4519 = x187 | n4518 ;
  assign n4520 = n830 & n1453 ;
  assign n4521 = n4520 ^ x239 ^ 1'b0 ;
  assign n4522 = n830 | n4521 ;
  assign n4523 = ~n1538 & n2592 ;
  assign n4524 = ~n3380 & n4523 ;
  assign n4525 = n364 | n946 ;
  assign n4526 = n4525 ^ n665 ^ 1'b0 ;
  assign n4527 = n1612 & ~n4526 ;
  assign n4528 = n1343 ^ x221 ^ 1'b0 ;
  assign n4529 = n424 & ~n4310 ;
  assign n4530 = ~n4528 & n4529 ;
  assign n4531 = n3326 | n4530 ;
  assign n4532 = n4531 ^ n3933 ^ 1'b0 ;
  assign n4533 = n4527 & n4532 ;
  assign n4534 = n312 & n4533 ;
  assign n4535 = n4132 ^ n1404 ^ 1'b0 ;
  assign n4536 = n4535 ^ n1581 ^ 1'b0 ;
  assign n4537 = x227 & n4536 ;
  assign n4538 = n3090 ^ n1125 ^ 1'b0 ;
  assign n4539 = n4537 & n4538 ;
  assign n4540 = n1803 ^ x182 ^ 1'b0 ;
  assign n4541 = n4540 ^ n2853 ^ 1'b0 ;
  assign n4543 = ~x27 & n353 ;
  assign n4544 = n1664 ^ x76 ^ 1'b0 ;
  assign n4545 = n4543 | n4544 ;
  assign n4542 = n2963 & ~n3357 ;
  assign n4546 = n4545 ^ n4542 ^ 1'b0 ;
  assign n4547 = n1466 & n4546 ;
  assign n4550 = n2376 ^ x133 ^ 1'b0 ;
  assign n4551 = n4550 ^ n3319 ^ 1'b0 ;
  assign n4548 = n971 | n2378 ;
  assign n4549 = x124 & ~n4548 ;
  assign n4552 = n4551 ^ n4549 ^ 1'b0 ;
  assign n4553 = n3345 ^ n676 ^ 1'b0 ;
  assign n4554 = n3963 | n4553 ;
  assign n4555 = n4554 ^ n2745 ^ 1'b0 ;
  assign n4556 = n4552 | n4555 ;
  assign n4557 = n1027 | n4556 ;
  assign n4558 = n759 & ~n4288 ;
  assign n4559 = ~n930 & n4558 ;
  assign n4560 = n459 & n984 ;
  assign n4561 = n4560 ^ x103 ^ 1'b0 ;
  assign n4562 = n4561 ^ n2790 ^ 1'b0 ;
  assign n4564 = n1398 | n4131 ;
  assign n4565 = n4564 ^ n1890 ^ 1'b0 ;
  assign n4563 = n2397 ^ n671 ^ 1'b0 ;
  assign n4566 = n4565 ^ n4563 ^ n3096 ;
  assign n4567 = x89 & ~x193 ;
  assign n4568 = x126 & ~n1623 ;
  assign n4569 = n4568 ^ n1092 ^ 1'b0 ;
  assign n4570 = x193 & x196 ;
  assign n4571 = n3262 & n4570 ;
  assign n4572 = n419 ^ x162 ^ 1'b0 ;
  assign n4573 = ~n338 & n786 ;
  assign n4574 = n4573 ^ n4502 ^ 1'b0 ;
  assign n4575 = n2953 ^ n1954 ^ n1837 ;
  assign n4576 = x115 | n4540 ;
  assign n4577 = ~n2188 & n3694 ;
  assign n4578 = n4577 ^ n1570 ^ 1'b0 ;
  assign n4582 = n3541 ^ n409 ^ 1'b0 ;
  assign n4583 = ~n744 & n4582 ;
  assign n4584 = n1156 & ~n4583 ;
  assign n4579 = n2625 ^ n1120 ^ 1'b0 ;
  assign n4580 = n4579 ^ n3659 ^ n2011 ;
  assign n4581 = ~n1362 & n4580 ;
  assign n4585 = n4584 ^ n4581 ^ 1'b0 ;
  assign n4591 = ( n419 & n445 ) | ( n419 & n1812 ) | ( n445 & n1812 ) ;
  assign n4592 = x241 | n3032 ;
  assign n4593 = n4591 & ~n4592 ;
  assign n4587 = x19 & ~n514 ;
  assign n4588 = ~n2004 & n4587 ;
  assign n4586 = x70 & ~n3111 ;
  assign n4589 = n4588 ^ n4586 ^ 1'b0 ;
  assign n4590 = ~n4409 & n4589 ;
  assign n4594 = n4593 ^ n4590 ^ 1'b0 ;
  assign n4595 = n4360 & n4594 ;
  assign n4596 = n2898 & ~n4595 ;
  assign n4597 = n3123 ^ n1896 ^ 1'b0 ;
  assign n4598 = n3272 & n4597 ;
  assign n4599 = n3108 ^ n1971 ^ 1'b0 ;
  assign n4600 = n2609 ^ n1465 ^ x224 ;
  assign n4601 = n2900 ^ n2161 ^ 1'b0 ;
  assign n4602 = ~n1368 & n4601 ;
  assign n4603 = n4602 ^ n3265 ^ 1'b0 ;
  assign n4604 = n4600 & n4603 ;
  assign n4605 = n539 & n4604 ;
  assign n4606 = x60 & ~n596 ;
  assign n4607 = n4606 ^ n638 ^ 1'b0 ;
  assign n4608 = n900 | n4607 ;
  assign n4609 = n3671 ^ n710 ^ 1'b0 ;
  assign n4610 = n4327 & n4609 ;
  assign n4611 = n4610 ^ n4409 ^ 1'b0 ;
  assign n4612 = ( n1140 & ~n2833 ) | ( n1140 & n3564 ) | ( ~n2833 & n3564 ) ;
  assign n4613 = ~n4611 & n4612 ;
  assign n4614 = n4613 ^ n3088 ^ 1'b0 ;
  assign n4615 = n4608 & ~n4614 ;
  assign n4616 = n4218 ^ n3124 ^ 1'b0 ;
  assign n4617 = n2159 & ~n4616 ;
  assign n4618 = n1101 ^ x89 ^ 1'b0 ;
  assign n4619 = n2353 & ~n4618 ;
  assign n4620 = n1144 ^ n1064 ^ 1'b0 ;
  assign n4621 = ~n4426 & n4620 ;
  assign n4622 = n4621 ^ n3679 ^ 1'b0 ;
  assign n4623 = ~n1704 & n4622 ;
  assign n4624 = ~n4619 & n4623 ;
  assign n4625 = n1433 ^ n804 ^ 1'b0 ;
  assign n4626 = n3790 | n4625 ;
  assign n4627 = ( n294 & n2572 ) | ( n294 & n4626 ) | ( n2572 & n4626 ) ;
  assign n4628 = n3168 | n4003 ;
  assign n4629 = n4627 | n4628 ;
  assign n4630 = n1922 & n4629 ;
  assign n4631 = n4630 ^ n1940 ^ 1'b0 ;
  assign n4632 = n4177 ^ n2926 ^ 1'b0 ;
  assign n4633 = x62 | n4632 ;
  assign n4634 = x1 & n450 ;
  assign n4635 = ~n262 & n1484 ;
  assign n4636 = n4635 ^ n985 ^ 1'b0 ;
  assign n4637 = n4634 & n4636 ;
  assign n4638 = ~n3001 & n4637 ;
  assign n4639 = n4409 ^ n2289 ^ 1'b0 ;
  assign n4640 = n1789 ^ n1638 ^ 1'b0 ;
  assign n4641 = x35 & n2443 ;
  assign n4642 = ~x91 & n4641 ;
  assign n4643 = n520 & n4642 ;
  assign n4644 = x204 ^ x103 ^ 1'b0 ;
  assign n4645 = n4643 | n4644 ;
  assign n4646 = n1619 ^ n653 ^ x223 ;
  assign n4647 = ~x57 & n4646 ;
  assign n4648 = n3757 & n4647 ;
  assign n4649 = n653 & n838 ;
  assign n4650 = n4649 ^ n716 ^ 1'b0 ;
  assign n4651 = n4650 ^ n3021 ^ 1'b0 ;
  assign n4652 = n1832 & ~n4651 ;
  assign n4653 = n1371 & n3551 ;
  assign n4654 = ~n4652 & n4653 ;
  assign n4655 = n689 & n3420 ;
  assign n4656 = n535 & n4655 ;
  assign n4657 = n4656 ^ n2177 ^ x120 ;
  assign n4658 = n1741 | n4657 ;
  assign n4659 = n4658 ^ n522 ^ 1'b0 ;
  assign n4660 = n615 | n4659 ;
  assign n4662 = n2763 | n3801 ;
  assign n4661 = n733 | n3039 ;
  assign n4663 = n4662 ^ n4661 ^ 1'b0 ;
  assign n4664 = n971 & ~n2841 ;
  assign n4665 = n4664 ^ n397 ^ 1'b0 ;
  assign n4666 = n4665 ^ n3348 ^ 1'b0 ;
  assign n4667 = n3405 & n4666 ;
  assign n4668 = n4667 ^ n891 ^ 1'b0 ;
  assign n4669 = ~n988 & n1993 ;
  assign n4670 = n628 ^ n433 ^ 1'b0 ;
  assign n4674 = n1605 ^ n475 ^ 1'b0 ;
  assign n4675 = ~n1197 & n4674 ;
  assign n4671 = n3332 ^ n1103 ^ 1'b0 ;
  assign n4672 = n3536 | n4671 ;
  assign n4673 = ( n985 & n2075 ) | ( n985 & n4672 ) | ( n2075 & n4672 ) ;
  assign n4676 = n4675 ^ n4673 ^ n1295 ;
  assign n4677 = ~n1545 & n4540 ;
  assign n4678 = n728 ^ x74 ^ 1'b0 ;
  assign n4679 = n1032 & n4678 ;
  assign n4680 = ~n595 & n724 ;
  assign n4681 = n4680 ^ n4611 ^ 1'b0 ;
  assign n4682 = n4679 & ~n4681 ;
  assign n4683 = n2051 ^ n1185 ^ 1'b0 ;
  assign n4684 = n794 & ~n4683 ;
  assign n4685 = n4267 & n4684 ;
  assign n4686 = n2317 ^ n1606 ^ n1405 ;
  assign n4687 = x242 & ~n346 ;
  assign n4688 = ~x40 & n4687 ;
  assign n4689 = n4688 ^ n2260 ^ 1'b0 ;
  assign n4690 = n3569 & n4689 ;
  assign n4691 = n4690 ^ n3349 ^ 1'b0 ;
  assign n4692 = n4136 ^ n2203 ^ 1'b0 ;
  assign n4693 = n694 & n4692 ;
  assign n4694 = n1307 & n1756 ;
  assign n4695 = n853 | n4694 ;
  assign n4696 = n3150 | n4695 ;
  assign n4703 = n4011 ^ n1059 ^ x88 ;
  assign n4697 = n863 ^ n416 ^ 1'b0 ;
  assign n4698 = n1812 | n4697 ;
  assign n4699 = ( ~x12 & n848 ) | ( ~x12 & n3042 ) | ( n848 & n3042 ) ;
  assign n4700 = n4699 ^ n1893 ^ 1'b0 ;
  assign n4701 = n4117 | n4700 ;
  assign n4702 = n4698 | n4701 ;
  assign n4704 = n4703 ^ n4702 ^ 1'b0 ;
  assign n4705 = n1154 | n2828 ;
  assign n4706 = n2442 & ~n4705 ;
  assign n4707 = n3382 ^ n904 ^ 1'b0 ;
  assign n4708 = ~n1648 & n4707 ;
  assign n4709 = n1543 ^ n318 ^ 1'b0 ;
  assign n4710 = n4708 & n4709 ;
  assign n4711 = n825 ^ n722 ^ 1'b0 ;
  assign n4712 = n3780 | n4711 ;
  assign n4713 = n941 ^ n556 ^ 1'b0 ;
  assign n4714 = n3034 | n4713 ;
  assign n4715 = n4714 ^ n357 ^ 1'b0 ;
  assign n4716 = n4482 | n4715 ;
  assign n4717 = ~n973 & n1635 ;
  assign n4718 = ~n4716 & n4717 ;
  assign n4719 = n3186 ^ n2692 ^ 1'b0 ;
  assign n4720 = n3546 | n4719 ;
  assign n4721 = ( x227 & n1730 ) | ( x227 & ~n2442 ) | ( n1730 & ~n2442 ) ;
  assign n4722 = ~x118 & n4721 ;
  assign n4723 = n4722 ^ n4494 ^ 1'b0 ;
  assign n4724 = ~n1999 & n2796 ;
  assign n4725 = n3025 & ~n4393 ;
  assign n4726 = ( x40 & n1071 ) | ( x40 & ~n4032 ) | ( n1071 & ~n4032 ) ;
  assign n4727 = n2093 ^ n1264 ^ 1'b0 ;
  assign n4728 = ~n3768 & n4727 ;
  assign n4729 = x84 & ~n571 ;
  assign n4730 = n4729 ^ n1592 ^ 1'b0 ;
  assign n4731 = n3864 & n4730 ;
  assign n4732 = n4731 ^ n2080 ^ 1'b0 ;
  assign n4735 = ~n306 & n2542 ;
  assign n4736 = n4735 ^ n2284 ^ 1'b0 ;
  assign n4737 = n4013 ^ n1558 ^ n1135 ;
  assign n4738 = n1727 ^ n906 ^ 1'b0 ;
  assign n4739 = n4737 | n4738 ;
  assign n4740 = n2622 & ~n4739 ;
  assign n4741 = n4736 | n4740 ;
  assign n4733 = n2203 ^ n932 ^ 1'b0 ;
  assign n4734 = ~n891 & n4733 ;
  assign n4742 = n4741 ^ n4734 ^ 1'b0 ;
  assign n4743 = n4724 ^ n778 ^ 1'b0 ;
  assign n4744 = n684 | n4743 ;
  assign n4745 = n3290 ^ n2542 ^ 1'b0 ;
  assign n4746 = n4300 ^ n613 ^ 1'b0 ;
  assign n4747 = n4745 & n4746 ;
  assign n4748 = ( ~x247 & n893 ) | ( ~x247 & n2900 ) | ( n893 & n2900 ) ;
  assign n4751 = n1093 ^ n957 ^ 1'b0 ;
  assign n4752 = ~n1545 & n4751 ;
  assign n4753 = n4752 ^ n2466 ^ n1861 ;
  assign n4754 = x99 & n4753 ;
  assign n4749 = n260 & n747 ;
  assign n4750 = n4749 ^ n2078 ^ 1'b0 ;
  assign n4755 = n4754 ^ n4750 ^ 1'b0 ;
  assign n4756 = n2896 & n4755 ;
  assign n4757 = n4748 & n4756 ;
  assign n4758 = x136 & n1440 ;
  assign n4761 = n844 & n1011 ;
  assign n4762 = n4761 ^ x207 ^ 1'b0 ;
  assign n4763 = n4543 | n4762 ;
  assign n4764 = n4763 ^ n1903 ^ 1'b0 ;
  assign n4759 = ( n1316 & ~n1332 ) | ( n1316 & n1590 ) | ( ~n1332 & n1590 ) ;
  assign n4760 = ~n2011 & n4759 ;
  assign n4765 = n4764 ^ n4760 ^ 1'b0 ;
  assign n4766 = n4758 | n4765 ;
  assign n4767 = n2582 ^ n2096 ^ 1'b0 ;
  assign n4768 = ( ~x111 & n1749 ) | ( ~x111 & n4767 ) | ( n1749 & n4767 ) ;
  assign n4769 = n4588 & ~n4768 ;
  assign n4770 = n4769 ^ n3881 ^ 1'b0 ;
  assign n4771 = n3790 ^ n784 ^ 1'b0 ;
  assign n4772 = n4771 ^ n752 ^ 1'b0 ;
  assign n4773 = x86 & ~n4772 ;
  assign n4777 = n754 | n3134 ;
  assign n4778 = n4777 ^ n1648 ^ 1'b0 ;
  assign n4774 = x224 & n402 ;
  assign n4775 = n312 & n4774 ;
  assign n4776 = n1671 | n4775 ;
  assign n4779 = n4778 ^ n4776 ^ 1'b0 ;
  assign n4780 = n4779 ^ n3425 ^ n1519 ;
  assign n4781 = n1914 & ~n2060 ;
  assign n4782 = ~n848 & n4781 ;
  assign n4783 = n4782 ^ n2045 ^ 1'b0 ;
  assign n4784 = n1750 ^ x229 ^ 1'b0 ;
  assign n4787 = x157 & ~n1424 ;
  assign n4785 = n575 & ~n792 ;
  assign n4786 = n4785 ^ n1342 ^ 1'b0 ;
  assign n4788 = n4787 ^ n4786 ^ n858 ;
  assign n4789 = n4788 ^ n1579 ^ 1'b0 ;
  assign n4790 = n4784 & ~n4789 ;
  assign n4791 = ~x202 & n477 ;
  assign n4792 = n3855 ^ n1899 ^ n428 ;
  assign n4793 = n784 & n4792 ;
  assign n4794 = n2276 ^ n759 ^ n637 ;
  assign n4795 = n3650 | n4794 ;
  assign n4796 = n928 & ~n3935 ;
  assign n4797 = ~n708 & n4796 ;
  assign n4798 = ~n1424 & n2294 ;
  assign n4799 = n4798 ^ n2618 ^ 1'b0 ;
  assign n4800 = n982 & n4799 ;
  assign n4801 = n4800 ^ n2618 ^ 1'b0 ;
  assign n4802 = n2995 | n4801 ;
  assign n4804 = n1523 ^ n971 ^ 1'b0 ;
  assign n4805 = n4804 ^ x198 ^ 1'b0 ;
  assign n4803 = n1232 | n2431 ;
  assign n4806 = n4805 ^ n4803 ^ n4219 ;
  assign n4807 = n1001 & n1735 ;
  assign n4808 = n4807 ^ n4165 ^ 1'b0 ;
  assign n4809 = ~n2397 & n4808 ;
  assign n4810 = n3257 & ~n3910 ;
  assign n4811 = ~x53 & n4810 ;
  assign n4812 = n3901 | n4811 ;
  assign n4813 = n1129 | n4812 ;
  assign n4814 = n4813 ^ n440 ^ 1'b0 ;
  assign n4815 = n2872 & ~n4814 ;
  assign n4816 = n1352 | n2763 ;
  assign n4817 = n2571 | n4816 ;
  assign n4818 = n4817 ^ n1349 ^ 1'b0 ;
  assign n4819 = n1590 | n3403 ;
  assign n4823 = n3121 ^ n1577 ^ 1'b0 ;
  assign n4824 = n367 & ~n4823 ;
  assign n4825 = n2750 & n4824 ;
  assign n4826 = n2916 & n4825 ;
  assign n4820 = n3238 & n3647 ;
  assign n4821 = n4820 ^ x48 ^ 1'b0 ;
  assign n4822 = n1318 & ~n4821 ;
  assign n4827 = n4826 ^ n4822 ^ 1'b0 ;
  assign n4828 = ( x192 & n3892 ) | ( x192 & n4827 ) | ( n3892 & n4827 ) ;
  assign n4829 = n710 | n4611 ;
  assign n4830 = n1636 | n4829 ;
  assign n4834 = ~n1036 & n1543 ;
  assign n4835 = n4834 ^ n2604 ^ 1'b0 ;
  assign n4831 = ~x88 & n3634 ;
  assign n4832 = ( n848 & ~n3506 ) | ( n848 & n4831 ) | ( ~n3506 & n4831 ) ;
  assign n4833 = ~n397 & n4832 ;
  assign n4836 = n4835 ^ n4833 ^ 1'b0 ;
  assign n4837 = n2424 ^ n1064 ^ x156 ;
  assign n4838 = n1958 & ~n4837 ;
  assign n4839 = n925 ^ x133 ^ 1'b0 ;
  assign n4840 = n4839 ^ n2310 ^ 1'b0 ;
  assign n4841 = n850 & ~n3835 ;
  assign n4842 = ~x84 & n4841 ;
  assign n4843 = n4580 ^ n2706 ^ 1'b0 ;
  assign n4844 = n3815 ^ n256 ^ 1'b0 ;
  assign n4845 = n3186 | n4107 ;
  assign n4846 = ( ~n4449 & n4844 ) | ( ~n4449 & n4845 ) | ( n4844 & n4845 ) ;
  assign n4847 = n1742 & ~n2900 ;
  assign n4848 = ~n4846 & n4847 ;
  assign n4849 = ~n885 & n4222 ;
  assign n4851 = n1221 & ~n1973 ;
  assign n4850 = n1227 | n3168 ;
  assign n4852 = n4851 ^ n4850 ^ 1'b0 ;
  assign n4853 = n3446 ^ x194 ^ 1'b0 ;
  assign n4854 = n653 | n1809 ;
  assign n4855 = n3603 & ~n4854 ;
  assign n4856 = n1440 | n4855 ;
  assign n4857 = n4856 ^ x75 ^ 1'b0 ;
  assign n4858 = n2032 ^ n779 ^ 1'b0 ;
  assign n4859 = ~n4292 & n4858 ;
  assign n4860 = n1968 ^ n466 ^ 1'b0 ;
  assign n4862 = n850 & ~n1311 ;
  assign n4863 = n1678 & ~n4862 ;
  assign n4864 = ~n1696 & n4863 ;
  assign n4861 = n3281 & ~n4775 ;
  assign n4865 = n4864 ^ n4861 ^ 1'b0 ;
  assign n4866 = n2208 & n4865 ;
  assign n4867 = n2456 & n4866 ;
  assign n4868 = ~n739 & n1610 ;
  assign n4869 = n1725 ^ x121 ^ 1'b0 ;
  assign n4870 = n3432 ^ n3027 ^ 1'b0 ;
  assign n4871 = ~n2715 & n4870 ;
  assign n4872 = ( n4868 & n4869 ) | ( n4868 & ~n4871 ) | ( n4869 & ~n4871 ) ;
  assign n4874 = n1200 | n1454 ;
  assign n4873 = n3340 | n3814 ;
  assign n4875 = n4874 ^ n4873 ^ 1'b0 ;
  assign n4876 = n655 | n2998 ;
  assign n4877 = n3895 ^ n3755 ^ 1'b0 ;
  assign n4878 = ~n1664 & n4877 ;
  assign n4879 = n2218 | n3091 ;
  assign n4880 = n4879 ^ n3977 ^ 1'b0 ;
  assign n4881 = x20 & ~n3845 ;
  assign n4882 = n2455 | n3415 ;
  assign n4883 = n4882 ^ n1676 ^ 1'b0 ;
  assign n4884 = n4883 ^ n2693 ^ 1'b0 ;
  assign n4885 = n1828 & n4884 ;
  assign n4886 = ~n1617 & n2146 ;
  assign n4887 = n4886 ^ n928 ^ 1'b0 ;
  assign n4888 = n3209 ^ n747 ^ n592 ;
  assign n4889 = n4888 ^ x60 ^ 1'b0 ;
  assign n4890 = n2633 & n4889 ;
  assign n4891 = n1238 & n1815 ;
  assign n4892 = ~n1156 & n4891 ;
  assign n4893 = n3326 ^ n494 ^ 1'b0 ;
  assign n4894 = x187 & n4893 ;
  assign n4895 = n4894 ^ n1318 ^ 1'b0 ;
  assign n4896 = n2326 ^ n336 ^ 1'b0 ;
  assign n4897 = n2972 | n4896 ;
  assign n4898 = n4897 ^ n3655 ^ 1'b0 ;
  assign n4899 = ~n2013 & n2446 ;
  assign n4900 = ( x219 & n4898 ) | ( x219 & ~n4899 ) | ( n4898 & ~n4899 ) ;
  assign n4901 = x197 & n547 ;
  assign n4902 = n4901 ^ n3087 ^ 1'b0 ;
  assign n4903 = n444 | n1198 ;
  assign n4904 = n1495 & n4903 ;
  assign n4905 = n1094 & n4904 ;
  assign n4906 = x130 | n1929 ;
  assign n4907 = n4905 | n4906 ;
  assign n4908 = n4907 ^ n853 ^ 1'b0 ;
  assign n4909 = n4902 & ~n4908 ;
  assign n4910 = n3150 & n3855 ;
  assign n4911 = n2262 ^ n1997 ^ x253 ;
  assign n4914 = x22 & n1182 ;
  assign n4912 = ~n2122 & n2538 ;
  assign n4913 = n4912 ^ n4386 ^ 1'b0 ;
  assign n4915 = n4914 ^ n4913 ^ 1'b0 ;
  assign n4916 = n4911 & ~n4915 ;
  assign n4917 = n1919 ^ n485 ^ 1'b0 ;
  assign n4918 = n1684 & ~n4917 ;
  assign n4919 = ~n643 & n4918 ;
  assign n4920 = n3967 | n4919 ;
  assign n4921 = n1290 | n4920 ;
  assign n4922 = n4360 ^ n3034 ^ 1'b0 ;
  assign n4924 = n430 & n1778 ;
  assign n4923 = n3546 ^ n1538 ^ 1'b0 ;
  assign n4925 = n4924 ^ n4923 ^ n2600 ;
  assign n4926 = n2807 & ~n4925 ;
  assign n4927 = ~n862 & n4926 ;
  assign n4928 = n1500 & ~n3670 ;
  assign n4929 = n4928 ^ n1467 ^ 1'b0 ;
  assign n4930 = n3296 ^ n2122 ^ 1'b0 ;
  assign n4931 = n4929 & ~n4930 ;
  assign n4932 = n3817 ^ n2006 ^ x241 ;
  assign n4933 = n4932 ^ n1286 ^ 1'b0 ;
  assign n4934 = n334 | n4933 ;
  assign n4935 = n4394 ^ n1772 ^ 1'b0 ;
  assign n4936 = ~n2431 & n4935 ;
  assign n4940 = x180 & n2378 ;
  assign n4937 = ~x78 & x83 ;
  assign n4938 = n1069 ^ n975 ^ x32 ;
  assign n4939 = n4937 & n4938 ;
  assign n4941 = n4940 ^ n4939 ^ 1'b0 ;
  assign n4942 = n4642 ^ n1494 ^ n746 ;
  assign n4943 = ~x204 & n4942 ;
  assign n4944 = ~n4842 & n4943 ;
  assign n4945 = x3 & ~n1539 ;
  assign n4946 = n4945 ^ n1097 ^ 1'b0 ;
  assign n4947 = n4946 ^ x129 ^ 1'b0 ;
  assign n4948 = n511 | n4947 ;
  assign n4949 = ( ~n444 & n4663 ) | ( ~n444 & n4948 ) | ( n4663 & n4948 ) ;
  assign n4950 = ~n276 & n1695 ;
  assign n4951 = ( n906 & n2183 ) | ( n906 & ~n4038 ) | ( n2183 & ~n4038 ) ;
  assign n4952 = n4950 & n4951 ;
  assign n4953 = n4952 ^ n1556 ^ 1'b0 ;
  assign n4954 = n3771 ^ n1219 ^ 1'b0 ;
  assign n4955 = ~n638 & n4824 ;
  assign n4956 = ~x157 & n4955 ;
  assign n4957 = n3121 | n3228 ;
  assign n4958 = n3861 & n4957 ;
  assign n4959 = ~n1420 & n3867 ;
  assign n4961 = n894 & n1091 ;
  assign n4962 = n2785 & n4961 ;
  assign n4963 = n2096 | n4962 ;
  assign n4964 = n4380 | n4963 ;
  assign n4960 = x6 & ~n1990 ;
  assign n4965 = n4964 ^ n4960 ^ 1'b0 ;
  assign n4966 = ~n2034 & n4871 ;
  assign n4967 = ~n1986 & n4580 ;
  assign n4968 = n4967 ^ x135 ^ 1'b0 ;
  assign n4969 = x137 & n579 ;
  assign n4970 = n2704 & n4969 ;
  assign n4971 = n1475 | n4970 ;
  assign n4972 = n4968 & ~n4971 ;
  assign n4973 = n4972 ^ x180 ^ 1'b0 ;
  assign n4974 = ~n1304 & n4973 ;
  assign n4975 = n336 & n3086 ;
  assign n4976 = n4975 ^ n1994 ^ 1'b0 ;
  assign n4977 = n2252 | n3342 ;
  assign n4978 = x50 & n4977 ;
  assign n4979 = n4978 ^ n3785 ^ 1'b0 ;
  assign n4980 = n4979 ^ n494 ^ 1'b0 ;
  assign n4981 = n4976 & ~n4980 ;
  assign n4982 = n1626 & n3568 ;
  assign n4983 = n4982 ^ x172 ^ 1'b0 ;
  assign n4984 = n4216 & n4983 ;
  assign n4985 = n4984 ^ n991 ^ 1'b0 ;
  assign n4986 = n4985 ^ n3352 ^ n1360 ;
  assign n4987 = n3340 | n3486 ;
  assign n4988 = n1775 & ~n4987 ;
  assign n4989 = n1707 ^ n710 ^ 1'b0 ;
  assign n4991 = n2780 & ~n3300 ;
  assign n4990 = x134 & n937 ;
  assign n4992 = n4991 ^ n4990 ^ 1'b0 ;
  assign n4993 = x142 & n3521 ;
  assign n4994 = n3549 & n4234 ;
  assign n4995 = n4993 & ~n4994 ;
  assign n4996 = n3496 & n4995 ;
  assign n4997 = n4996 ^ n2615 ^ 1'b0 ;
  assign n4998 = n4997 ^ n3537 ^ n3494 ;
  assign n4999 = n2935 ^ n865 ^ 1'b0 ;
  assign n5000 = n3300 | n4999 ;
  assign n5001 = n5000 ^ n937 ^ 1'b0 ;
  assign n5007 = n2013 ^ n260 ^ 1'b0 ;
  assign n5002 = n347 | n1386 ;
  assign n5003 = n2119 | n5002 ;
  assign n5004 = n3699 ^ n1763 ^ n1242 ;
  assign n5005 = n5004 ^ n2265 ^ 1'b0 ;
  assign n5006 = n5003 & n5005 ;
  assign n5008 = n5007 ^ n5006 ^ 1'b0 ;
  assign n5009 = n451 & ~n1237 ;
  assign n5010 = x17 | n1059 ;
  assign n5011 = n2803 | n2909 ;
  assign n5012 = n5010 & ~n5011 ;
  assign n5013 = n5009 & ~n5012 ;
  assign n5014 = n1760 & n5013 ;
  assign n5015 = n293 & n4622 ;
  assign n5016 = n5015 ^ n3607 ^ 1'b0 ;
  assign n5017 = n5016 ^ n4861 ^ 1'b0 ;
  assign n5018 = n2403 ^ n908 ^ x221 ;
  assign n5019 = n266 & ~n2970 ;
  assign n5020 = n2029 & n5019 ;
  assign n5021 = n4626 ^ n547 ^ 1'b0 ;
  assign n5022 = n2229 & n4631 ;
  assign n5023 = n2237 ^ n571 ^ x73 ;
  assign n5024 = x111 & n3504 ;
  assign n5025 = n1378 & n5024 ;
  assign n5026 = n991 & ~n1990 ;
  assign n5027 = ~n2542 & n5026 ;
  assign n5028 = n5027 ^ n3650 ^ n2893 ;
  assign n5029 = n4341 | n5028 ;
  assign n5030 = n5029 ^ n3588 ^ 1'b0 ;
  assign n5031 = n5025 | n5030 ;
  assign n5032 = n1335 & ~n3529 ;
  assign n5033 = ~n351 & n5032 ;
  assign n5034 = x138 & ~x226 ;
  assign n5035 = n4338 ^ n2852 ^ 1'b0 ;
  assign n5036 = ~n2018 & n5035 ;
  assign n5037 = x119 & ~n1725 ;
  assign n5038 = n3085 & n5037 ;
  assign n5039 = n4178 ^ x122 ^ x59 ;
  assign n5040 = n3202 & n5039 ;
  assign n5041 = n5038 & n5040 ;
  assign n5045 = n676 ^ n655 ^ 1'b0 ;
  assign n5046 = n1389 & ~n5045 ;
  assign n5044 = x107 & ~n1538 ;
  assign n5042 = n2268 ^ n488 ^ 1'b0 ;
  assign n5043 = n2615 & n5042 ;
  assign n5047 = n5046 ^ n5044 ^ n5043 ;
  assign n5048 = n951 & n2274 ;
  assign n5049 = n393 & n5048 ;
  assign n5050 = ( n1373 & n1649 ) | ( n1373 & n1707 ) | ( n1649 & n1707 ) ;
  assign n5051 = n395 & n1746 ;
  assign n5052 = n5050 | n5051 ;
  assign n5053 = n2187 & ~n2574 ;
  assign n5054 = n871 & n5053 ;
  assign n5055 = ( x83 & ~n1869 ) | ( x83 & n5054 ) | ( ~n1869 & n5054 ) ;
  assign n5056 = n5055 ^ n4708 ^ n853 ;
  assign n5057 = n5056 ^ n2030 ^ 1'b0 ;
  assign n5058 = n2779 & n5057 ;
  assign n5059 = ~n4306 & n5058 ;
  assign n5060 = n772 ^ n510 ^ 1'b0 ;
  assign n5061 = n5060 ^ n923 ^ 1'b0 ;
  assign n5062 = n5061 ^ n3875 ^ n3722 ;
  assign n5063 = n4935 ^ n4239 ^ 1'b0 ;
  assign n5064 = n1423 ^ x104 ^ 1'b0 ;
  assign n5065 = n4380 & n5064 ;
  assign n5066 = x13 | n2506 ;
  assign n5067 = n2868 & n4153 ;
  assign n5068 = x186 & ~n5067 ;
  assign n5069 = n5068 ^ n3425 ^ 1'b0 ;
  assign n5070 = ~n2452 & n5069 ;
  assign n5071 = ~n2948 & n5070 ;
  assign n5072 = ~n3235 & n5071 ;
  assign n5073 = n382 | n5072 ;
  assign n5074 = n2749 & ~n5073 ;
  assign n5075 = n4543 ^ n4268 ^ 1'b0 ;
  assign n5076 = n4525 & ~n4799 ;
  assign n5077 = n4368 ^ n3440 ^ 1'b0 ;
  assign n5078 = n3447 & n5077 ;
  assign n5079 = n2464 ^ n543 ^ 1'b0 ;
  assign n5080 = n2961 | n3370 ;
  assign n5081 = ( n1623 & ~n2746 ) | ( n1623 & n2903 ) | ( ~n2746 & n2903 ) ;
  assign n5082 = n5081 ^ n4572 ^ 1'b0 ;
  assign n5083 = n3577 & n4452 ;
  assign n5084 = n5083 ^ n260 ^ 1'b0 ;
  assign n5085 = n2076 & ~n3139 ;
  assign n5086 = n5085 ^ n2345 ^ 1'b0 ;
  assign n5087 = x150 & ~n708 ;
  assign n5088 = n2069 & n5087 ;
  assign n5089 = n5088 ^ n1830 ^ 1'b0 ;
  assign n5090 = n4389 ^ x174 ^ 1'b0 ;
  assign n5091 = n1947 & n5090 ;
  assign n5092 = n1095 | n1712 ;
  assign n5093 = n469 & ~n5092 ;
  assign n5094 = n5093 ^ n1894 ^ 1'b0 ;
  assign n5095 = n1398 & n4684 ;
  assign n5096 = n5094 | n5095 ;
  assign n5097 = n5096 ^ n2884 ^ 1'b0 ;
  assign n5098 = n3423 ^ n2567 ^ 1'b0 ;
  assign n5099 = n5097 | n5098 ;
  assign n5100 = x95 & n583 ;
  assign n5101 = n4804 ^ n336 ^ 1'b0 ;
  assign n5102 = ~n5100 & n5101 ;
  assign n5103 = n5102 ^ n4399 ^ 1'b0 ;
  assign n5104 = n637 | n4708 ;
  assign n5105 = n2905 & ~n4393 ;
  assign n5106 = n2040 ^ n679 ^ 1'b0 ;
  assign n5107 = n956 | n5106 ;
  assign n5108 = n5107 ^ x105 ^ 1'b0 ;
  assign n5109 = n3183 & n3235 ;
  assign n5110 = n2870 & n5109 ;
  assign n5111 = ~n3298 & n4354 ;
  assign n5112 = n772 ^ n754 ^ 1'b0 ;
  assign n5113 = n318 & n5112 ;
  assign n5114 = n4441 ^ n1245 ^ 1'b0 ;
  assign n5115 = n2725 ^ x252 ^ 1'b0 ;
  assign n5116 = ~n4450 & n5115 ;
  assign n5117 = n2817 & n4341 ;
  assign n5118 = n5117 ^ n2307 ^ 1'b0 ;
  assign n5122 = n3253 ^ n1737 ^ 1'b0 ;
  assign n5119 = n2968 ^ n2291 ^ 1'b0 ;
  assign n5120 = ( n1651 & n2341 ) | ( n1651 & ~n3903 ) | ( n2341 & ~n3903 ) ;
  assign n5121 = ( x190 & ~n5119 ) | ( x190 & n5120 ) | ( ~n5119 & n5120 ) ;
  assign n5123 = n5122 ^ n5121 ^ 1'b0 ;
  assign n5124 = n1495 & ~n3109 ;
  assign n5125 = n624 & n5124 ;
  assign n5131 = n3712 | n3801 ;
  assign n5132 = n2121 & ~n5131 ;
  assign n5126 = n869 ^ x249 ^ 1'b0 ;
  assign n5127 = ~n2403 & n5126 ;
  assign n5128 = n3302 ^ n1397 ^ 1'b0 ;
  assign n5129 = n5127 & n5128 ;
  assign n5130 = n294 & n5129 ;
  assign n5133 = n5132 ^ n5130 ^ 1'b0 ;
  assign n5134 = n3253 & ~n5133 ;
  assign n5135 = ~x91 & x188 ;
  assign n5138 = n4265 | n4622 ;
  assign n5136 = n900 & n1931 ;
  assign n5137 = n970 & ~n5136 ;
  assign n5139 = n5138 ^ n5137 ^ 1'b0 ;
  assign n5140 = ( x121 & ~n622 ) | ( x121 & n709 ) | ( ~n622 & n709 ) ;
  assign n5141 = ~x107 & n3150 ;
  assign n5142 = n1835 & n5141 ;
  assign n5143 = n274 & n831 ;
  assign n5144 = n5143 ^ n3290 ^ 1'b0 ;
  assign n5145 = n2148 & ~n5144 ;
  assign n5146 = n5145 ^ n2926 ^ 1'b0 ;
  assign n5147 = n5146 ^ n1381 ^ 1'b0 ;
  assign n5148 = n5142 | n5147 ;
  assign n5149 = n3887 ^ n1680 ^ 1'b0 ;
  assign n5150 = ~n4166 & n5149 ;
  assign n5151 = ~n1138 & n5150 ;
  assign n5152 = x140 & n2011 ;
  assign n5153 = n1737 & n3647 ;
  assign n5154 = ( n2170 & ~n3230 ) | ( n2170 & n5093 ) | ( ~n3230 & n5093 ) ;
  assign n5155 = n3206 & ~n5154 ;
  assign n5156 = n5155 ^ n4921 ^ 1'b0 ;
  assign n5159 = n1579 & ~n2321 ;
  assign n5160 = ~n1417 & n5159 ;
  assign n5161 = n5160 ^ n1183 ^ 1'b0 ;
  assign n5162 = n2087 & n5161 ;
  assign n5163 = n5162 ^ n3586 ^ 1'b0 ;
  assign n5157 = n2779 & n3233 ;
  assign n5158 = ~n2779 & n5157 ;
  assign n5164 = n5163 ^ n5158 ^ 1'b0 ;
  assign n5165 = n4305 ^ n479 ^ x244 ;
  assign n5166 = n5164 | n5165 ;
  assign n5167 = n5164 & ~n5166 ;
  assign n5168 = n2547 ^ x212 ^ 1'b0 ;
  assign n5169 = n4150 ^ n2330 ^ 1'b0 ;
  assign n5170 = n5169 ^ n4974 ^ n1877 ;
  assign n5171 = n2358 ^ n1571 ^ 1'b0 ;
  assign n5172 = ~n1473 & n5171 ;
  assign n5173 = n5172 ^ n3057 ^ 1'b0 ;
  assign n5174 = ~n2260 & n3704 ;
  assign n5175 = ~n5173 & n5174 ;
  assign n5177 = n766 & n4010 ;
  assign n5178 = n4093 ^ n3186 ^ 1'b0 ;
  assign n5179 = n5177 & ~n5178 ;
  assign n5176 = n2362 ^ n963 ^ 1'b0 ;
  assign n5180 = n5179 ^ n5176 ^ 1'b0 ;
  assign n5181 = n4018 & n4622 ;
  assign n5182 = n2657 ^ n2184 ^ 1'b0 ;
  assign n5183 = n2062 ^ x41 ^ 1'b0 ;
  assign n5184 = ( n1866 & ~n1913 ) | ( n1866 & n2655 ) | ( ~n1913 & n2655 ) ;
  assign n5185 = n5184 ^ n2200 ^ 1'b0 ;
  assign n5186 = ~n5183 & n5185 ;
  assign n5187 = x133 & ~n709 ;
  assign n5188 = n2355 ^ n569 ^ 1'b0 ;
  assign n5189 = n2196 & n5188 ;
  assign n5190 = ~n2474 & n4124 ;
  assign n5191 = ~n3627 & n5190 ;
  assign n5192 = n5189 & n5191 ;
  assign n5193 = n4696 ^ n4154 ^ n466 ;
  assign n5194 = n1822 & ~n3765 ;
  assign n5195 = n5194 ^ n385 ^ 1'b0 ;
  assign n5196 = n787 | n3335 ;
  assign n5197 = n5196 ^ n1373 ^ 1'b0 ;
  assign n5198 = n1371 & n5197 ;
  assign n5199 = n1656 & n5198 ;
  assign n5200 = n2532 & ~n4025 ;
  assign n5201 = n5200 ^ n2091 ^ 1'b0 ;
  assign n5202 = n1774 & ~n5201 ;
  assign n5203 = n5202 ^ n4676 ^ 1'b0 ;
  assign n5204 = n3678 ^ n1154 ^ 1'b0 ;
  assign n5205 = n1905 | n5204 ;
  assign n5206 = ( x245 & ~n432 ) | ( x245 & n2868 ) | ( ~n432 & n2868 ) ;
  assign n5207 = ~n5205 & n5206 ;
  assign n5209 = x143 | n1999 ;
  assign n5208 = n3038 ^ n2674 ^ 1'b0 ;
  assign n5210 = n5209 ^ n5208 ^ 1'b0 ;
  assign n5211 = n5210 ^ n3958 ^ 1'b0 ;
  assign n5212 = n4537 & ~n5211 ;
  assign n5213 = ~n2458 & n4929 ;
  assign n5214 = ( ~n1406 & n3137 ) | ( ~n1406 & n5213 ) | ( n3137 & n5213 ) ;
  assign n5215 = n2513 | n3777 ;
  assign n5216 = n5215 ^ n592 ^ 1'b0 ;
  assign n5217 = n527 ^ x187 ^ 1'b0 ;
  assign n5218 = n1417 & ~n5217 ;
  assign n5219 = ( n1762 & n1937 ) | ( n1762 & n5218 ) | ( n1937 & n5218 ) ;
  assign n5220 = n4327 ^ n446 ^ 1'b0 ;
  assign n5221 = n2848 | n5220 ;
  assign n5222 = n5219 | n5221 ;
  assign n5223 = n5222 ^ n1307 ^ 1'b0 ;
  assign n5224 = n2545 ^ n2301 ^ 1'b0 ;
  assign n5225 = n2853 | n5224 ;
  assign n5226 = n4379 ^ n4022 ^ 1'b0 ;
  assign n5227 = n4744 | n5226 ;
  assign n5228 = n707 & ~n889 ;
  assign n5229 = n5228 ^ x17 ^ 1'b0 ;
  assign n5230 = n4222 ^ n729 ^ 1'b0 ;
  assign n5231 = ~n5229 & n5230 ;
  assign n5232 = n4479 ^ n2141 ^ 1'b0 ;
  assign n5233 = n4659 ^ n3577 ^ 1'b0 ;
  assign n5234 = n5232 | n5233 ;
  assign n5235 = n1283 & n1615 ;
  assign n5236 = ( n4050 & n4867 ) | ( n4050 & ~n5235 ) | ( n4867 & ~n5235 ) ;
  assign n5237 = n2176 ^ n475 ^ 1'b0 ;
  assign n5238 = n5237 ^ n613 ^ 1'b0 ;
  assign n5239 = n4301 | n5238 ;
  assign n5240 = n5239 ^ n270 ^ 1'b0 ;
  assign n5241 = n4388 & ~n5231 ;
  assign n5242 = n3845 | n4122 ;
  assign n5243 = n389 | n4298 ;
  assign n5244 = n4380 & n5243 ;
  assign n5245 = n2387 & n5244 ;
  assign n5246 = ~n801 & n2840 ;
  assign n5247 = n5246 ^ x251 ^ 1'b0 ;
  assign n5248 = ~n2101 & n5247 ;
  assign n5249 = n5248 ^ n2314 ^ 1'b0 ;
  assign n5250 = n4708 & n5249 ;
  assign n5251 = ~n1036 & n5250 ;
  assign n5252 = n4238 & n5251 ;
  assign n5253 = n3411 ^ x198 ^ 1'b0 ;
  assign n5254 = n4489 ^ n2335 ^ 1'b0 ;
  assign n5255 = n3729 & n5254 ;
  assign n5256 = ~n801 & n5255 ;
  assign n5257 = ( x38 & n340 ) | ( x38 & n2582 ) | ( n340 & n2582 ) ;
  assign n5258 = n3977 ^ n3888 ^ 1'b0 ;
  assign n5259 = n5257 & n5258 ;
  assign n5261 = n943 & ~n1381 ;
  assign n5260 = n2328 & ~n5165 ;
  assign n5262 = n5261 ^ n5260 ^ 1'b0 ;
  assign n5265 = n842 ^ n719 ^ 1'b0 ;
  assign n5266 = n3590 & n5265 ;
  assign n5267 = n4779 | n5266 ;
  assign n5268 = n5267 ^ n850 ^ 1'b0 ;
  assign n5263 = n2438 ^ n1958 ^ n1335 ;
  assign n5264 = n2453 & ~n5263 ;
  assign n5269 = n5268 ^ n5264 ^ 1'b0 ;
  assign n5270 = n1360 ^ n961 ^ x14 ;
  assign n5271 = n4778 ^ x251 ^ 1'b0 ;
  assign n5272 = n5121 & ~n5271 ;
  assign n5273 = ~n2272 & n3593 ;
  assign n5274 = n3156 ^ n1562 ^ 1'b0 ;
  assign n5275 = n5095 ^ n1539 ^ 1'b0 ;
  assign n5276 = ~n5274 & n5275 ;
  assign n5277 = n1371 & n1538 ;
  assign n5278 = n2915 & n5277 ;
  assign n5283 = ~n1471 & n4033 ;
  assign n5284 = ~n2402 & n5283 ;
  assign n5279 = n3455 ^ n2570 ^ 1'b0 ;
  assign n5280 = x14 & ~n5279 ;
  assign n5281 = n4051 & n5280 ;
  assign n5282 = n5281 ^ n4360 ^ 1'b0 ;
  assign n5285 = n5284 ^ n5282 ^ 1'b0 ;
  assign n5286 = n5278 & ~n5285 ;
  assign n5287 = ~n1450 & n2362 ;
  assign n5288 = ( ~x53 & n2464 ) | ( ~x53 & n5287 ) | ( n2464 & n5287 ) ;
  assign n5290 = n3073 ^ n919 ^ n661 ;
  assign n5289 = n1151 & ~n1579 ;
  assign n5291 = n5290 ^ n5289 ^ 1'b0 ;
  assign n5292 = n5291 ^ n2367 ^ 1'b0 ;
  assign n5293 = n5003 ^ n1968 ^ 1'b0 ;
  assign n5294 = ( x13 & n1739 ) | ( x13 & n5293 ) | ( n1739 & n5293 ) ;
  assign n5295 = n5294 ^ n1813 ^ 1'b0 ;
  assign n5296 = n2776 | n4026 ;
  assign n5297 = n3321 & n4163 ;
  assign n5298 = ~n5296 & n5297 ;
  assign n5299 = n2455 | n3539 ;
  assign n5300 = n5299 ^ n2532 ^ 1'b0 ;
  assign n5301 = n5300 ^ n4521 ^ 1'b0 ;
  assign n5302 = n2337 | n2937 ;
  assign n5303 = n1786 | n4943 ;
  assign n5304 = ~n2867 & n3190 ;
  assign n5305 = n5304 ^ n3088 ^ 1'b0 ;
  assign n5306 = n4650 ^ n3947 ^ 1'b0 ;
  assign n5307 = n1565 & ~n5306 ;
  assign n5310 = x230 & ~n2473 ;
  assign n5308 = n483 | n4805 ;
  assign n5309 = n2369 & n5308 ;
  assign n5311 = n5310 ^ n5309 ^ n2853 ;
  assign n5312 = n5311 ^ n1736 ^ 1'b0 ;
  assign n5313 = n5307 & n5312 ;
  assign n5314 = n400 & ~n751 ;
  assign n5315 = n413 & n5314 ;
  assign n5316 = ~n2065 & n5315 ;
  assign n5317 = n3001 & n5316 ;
  assign n5318 = ~n262 & n2798 ;
  assign n5319 = n1295 & ~n1487 ;
  assign n5320 = n5318 & n5319 ;
  assign n5321 = n3890 ^ n2105 ^ 1'b0 ;
  assign n5322 = ~x204 & n5321 ;
  assign n5323 = n2048 & ~n3267 ;
  assign n5324 = ( x189 & ~n3680 ) | ( x189 & n5323 ) | ( ~n3680 & n5323 ) ;
  assign n5325 = ~n1018 & n5324 ;
  assign n5326 = n3425 ^ n2310 ^ 1'b0 ;
  assign n5327 = n1664 | n2763 ;
  assign n5328 = n679 & ~n5327 ;
  assign n5329 = x174 & n3467 ;
  assign n5330 = n5329 ^ n2694 ^ 1'b0 ;
  assign n5332 = x118 & ~n1707 ;
  assign n5333 = n2441 & n5332 ;
  assign n5331 = n2098 | n2617 ;
  assign n5334 = n5333 ^ n5331 ^ 1'b0 ;
  assign n5335 = n419 & ~n2743 ;
  assign n5336 = n3910 ^ n1470 ^ 1'b0 ;
  assign n5337 = x6 & n2691 ;
  assign n5338 = ~n2736 & n5337 ;
  assign n5339 = n5338 ^ n1758 ^ n780 ;
  assign n5340 = n3258 | n5339 ;
  assign n5341 = x60 & n2916 ;
  assign n5342 = n1220 ^ x164 ^ 1'b0 ;
  assign n5343 = x136 & ~n5342 ;
  assign n5344 = ~n737 & n5343 ;
  assign n5345 = n2232 ^ n1651 ^ 1'b0 ;
  assign n5346 = n4520 & ~n5345 ;
  assign n5347 = n5344 & n5346 ;
  assign n5348 = n5292 ^ n2949 ^ 1'b0 ;
  assign n5349 = ~n2399 & n5348 ;
  assign n5350 = x102 & n1010 ;
  assign n5351 = x54 & ~n1628 ;
  assign n5352 = n5351 ^ n1947 ^ 1'b0 ;
  assign n5353 = n3890 & ~n5352 ;
  assign n5354 = n5353 ^ n4275 ^ 1'b0 ;
  assign n5355 = ( n2794 & n5350 ) | ( n2794 & n5354 ) | ( n5350 & n5354 ) ;
  assign n5356 = n1534 & n4220 ;
  assign n5357 = n2708 ^ n1440 ^ n1367 ;
  assign n5358 = n2644 ^ n2403 ^ 1'b0 ;
  assign n5359 = n4911 & ~n5358 ;
  assign n5360 = n3610 & n5359 ;
  assign n5362 = n1366 & ~n4097 ;
  assign n5363 = n5054 | n5362 ;
  assign n5361 = ~n655 & n3335 ;
  assign n5364 = n5363 ^ n5361 ^ 1'b0 ;
  assign n5365 = n3572 ^ n3288 ^ 1'b0 ;
  assign n5366 = n5365 ^ n535 ^ 1'b0 ;
  assign n5367 = n2302 ^ n1512 ^ 1'b0 ;
  assign n5368 = ~n1768 & n3769 ;
  assign n5369 = n5367 & ~n5368 ;
  assign n5370 = ~n1556 & n3952 ;
  assign n5371 = n3256 & n5370 ;
  assign n5372 = n2542 & n2857 ;
  assign n5373 = ~x146 & n5372 ;
  assign n5374 = n5373 ^ n2792 ^ 1'b0 ;
  assign n5375 = n5374 ^ n3333 ^ 1'b0 ;
  assign n5376 = n5095 ^ n3116 ^ 1'b0 ;
  assign n5377 = n2370 | n5376 ;
  assign n5378 = n1561 & ~n1736 ;
  assign n5379 = n2267 & n5378 ;
  assign n5380 = n5377 & ~n5379 ;
  assign n5385 = x169 & ~n1374 ;
  assign n5381 = n1232 | n1443 ;
  assign n5382 = x179 | n5381 ;
  assign n5383 = ( n1828 & n2047 ) | ( n1828 & ~n5382 ) | ( n2047 & ~n5382 ) ;
  assign n5384 = ( x179 & ~n3272 ) | ( x179 & n5383 ) | ( ~n3272 & n5383 ) ;
  assign n5386 = n5385 ^ n5384 ^ 1'b0 ;
  assign n5387 = n3040 | n3258 ;
  assign n5388 = x135 | n5387 ;
  assign n5390 = n671 & ~n1092 ;
  assign n5391 = n5390 ^ n1499 ^ 1'b0 ;
  assign n5389 = n4359 & ~n4503 ;
  assign n5392 = n5391 ^ n5389 ^ 1'b0 ;
  assign n5393 = ~n2095 & n2571 ;
  assign n5394 = n3216 ^ n863 ^ 1'b0 ;
  assign n5395 = x184 & ~n5394 ;
  assign n5396 = n5395 ^ n4205 ^ n1674 ;
  assign n5397 = n5396 ^ n3488 ^ 1'b0 ;
  assign n5398 = n3925 ^ n1111 ^ 1'b0 ;
  assign n5399 = n5398 ^ n5356 ^ 1'b0 ;
  assign n5400 = n5397 & ~n5399 ;
  assign n5401 = n1822 & ~n2274 ;
  assign n5402 = ( n1406 & n1579 ) | ( n1406 & n4675 ) | ( n1579 & n4675 ) ;
  assign n5403 = n5302 & n5402 ;
  assign n5404 = n3074 & ~n5112 ;
  assign n5405 = n1032 & ~n5404 ;
  assign n5406 = n5405 ^ n2514 ^ 1'b0 ;
  assign n5407 = n3196 ^ n2286 ^ 1'b0 ;
  assign n5408 = n5407 ^ n3166 ^ n1001 ;
  assign n5409 = n3977 & ~n5408 ;
  assign n5410 = ( ~x86 & n3333 ) | ( ~x86 & n4979 ) | ( n3333 & n4979 ) ;
  assign n5411 = ~n4970 & n5410 ;
  assign n5412 = ~n4900 & n5411 ;
  assign n5413 = n1468 ^ n922 ^ 1'b0 ;
  assign n5414 = n3427 | n5413 ;
  assign n5415 = n1377 & n1810 ;
  assign n5416 = ~n2936 & n5415 ;
  assign n5417 = n2323 | n2951 ;
  assign n5418 = n5417 ^ n2641 ^ 1'b0 ;
  assign n5419 = n5418 ^ n4498 ^ 1'b0 ;
  assign n5420 = n5419 ^ n4571 ^ n4493 ;
  assign n5421 = n5420 ^ n2323 ^ 1'b0 ;
  assign n5422 = n4867 ^ n3622 ^ 1'b0 ;
  assign n5423 = ~n1598 & n2232 ;
  assign n5424 = n2415 & ~n3085 ;
  assign n5425 = n3457 & n5424 ;
  assign n5426 = n5407 & ~n5425 ;
  assign n5427 = ~n4652 & n5426 ;
  assign n5428 = n3823 ^ n941 ^ 1'b0 ;
  assign n5429 = n2540 ^ n2447 ^ 1'b0 ;
  assign n5430 = n4859 & ~n5429 ;
  assign n5431 = n5430 ^ n1509 ^ 1'b0 ;
  assign n5432 = ~n4126 & n4862 ;
  assign n5433 = x174 & ~n3319 ;
  assign n5434 = n3981 & n4554 ;
  assign n5435 = n2322 & n5434 ;
  assign n5436 = n3159 | n5435 ;
  assign n5437 = n5433 | n5436 ;
  assign n5438 = x232 & n1731 ;
  assign n5439 = n4652 ^ n3370 ^ 1'b0 ;
  assign n5440 = n260 & n5439 ;
  assign n5441 = n764 & ~n2464 ;
  assign n5442 = n1276 & n5441 ;
  assign n5444 = n529 & ~n5028 ;
  assign n5445 = n5444 ^ x26 ^ 1'b0 ;
  assign n5443 = x25 & n3413 ;
  assign n5446 = n5445 ^ n5443 ^ n2087 ;
  assign n5453 = x167 ^ x71 ^ 1'b0 ;
  assign n5452 = n2146 ^ n1055 ^ 1'b0 ;
  assign n5454 = n5453 ^ n5452 ^ 1'b0 ;
  assign n5447 = x145 & ~n874 ;
  assign n5448 = n5447 ^ n374 ^ 1'b0 ;
  assign n5449 = x117 & ~n2062 ;
  assign n5450 = ~n5448 & n5449 ;
  assign n5451 = n5169 & ~n5450 ;
  assign n5455 = n5454 ^ n5451 ^ 1'b0 ;
  assign n5456 = ( n1495 & n2538 ) | ( n1495 & ~n4216 ) | ( n2538 & ~n4216 ) ;
  assign n5457 = n5455 & n5456 ;
  assign n5458 = n5457 ^ n880 ^ 1'b0 ;
  assign n5468 = x200 & ~n3640 ;
  assign n5469 = n5468 ^ n1023 ^ 1'b0 ;
  assign n5467 = n4593 ^ n1254 ^ 1'b0 ;
  assign n5470 = n5469 ^ n5467 ^ 1'b0 ;
  assign n5459 = n1053 ^ x20 ^ 1'b0 ;
  assign n5460 = n5459 ^ n4076 ^ 1'b0 ;
  assign n5461 = n1774 & ~n5460 ;
  assign n5462 = ~n1653 & n5461 ;
  assign n5463 = ( n2077 & ~n5266 ) | ( n2077 & n5462 ) | ( ~n5266 & n5462 ) ;
  assign n5464 = ~n1391 & n5463 ;
  assign n5465 = ~n1125 & n5464 ;
  assign n5466 = n4838 & ~n5465 ;
  assign n5471 = n5470 ^ n5466 ^ 1'b0 ;
  assign n5472 = n3523 ^ n2337 ^ n900 ;
  assign n5473 = ~n2589 & n5472 ;
  assign n5474 = n1749 & n5300 ;
  assign n5475 = n2257 & n3502 ;
  assign n5476 = n5475 ^ n3595 ^ 1'b0 ;
  assign n5477 = n421 | n1632 ;
  assign n5478 = n5027 ^ n1383 ^ 1'b0 ;
  assign n5479 = ~n5477 & n5478 ;
  assign n5480 = n4449 & n4817 ;
  assign n5481 = n1981 & n5480 ;
  assign n5482 = ~n928 & n2571 ;
  assign n5483 = n2609 ^ n651 ^ 1'b0 ;
  assign n5484 = n279 & ~n5483 ;
  assign n5485 = n1379 & ~n5484 ;
  assign n5486 = x148 & x198 ;
  assign n5487 = n2754 & n5486 ;
  assign n5488 = n5487 ^ n5484 ^ 1'b0 ;
  assign n5489 = n3667 ^ n922 ^ 1'b0 ;
  assign n5490 = n2161 | n5489 ;
  assign n5491 = n1958 & n5490 ;
  assign n5492 = ~x222 & n5491 ;
  assign n5493 = ~n3007 & n5492 ;
  assign n5494 = ( n1219 & n5488 ) | ( n1219 & n5493 ) | ( n5488 & n5493 ) ;
  assign n5495 = x75 & n2542 ;
  assign n5496 = n842 & n5495 ;
  assign n5497 = n1250 & ~n5496 ;
  assign n5499 = ~n1869 & n4327 ;
  assign n5500 = n5499 ^ n4752 ^ 1'b0 ;
  assign n5501 = n5500 ^ n705 ^ 1'b0 ;
  assign n5502 = n5339 & ~n5501 ;
  assign n5498 = n4568 ^ n1123 ^ 1'b0 ;
  assign n5503 = n5502 ^ n5498 ^ 1'b0 ;
  assign n5504 = n2533 & n5503 ;
  assign n5505 = n3332 ^ n323 ^ 1'b0 ;
  assign n5506 = n5505 ^ n3329 ^ 1'b0 ;
  assign n5507 = n5504 & ~n5506 ;
  assign n5508 = ~n2585 & n5143 ;
  assign n5509 = n1639 | n5508 ;
  assign n5510 = n4286 ^ n928 ^ 1'b0 ;
  assign n5511 = n1376 | n3075 ;
  assign n5512 = n5511 ^ n2011 ^ 1'b0 ;
  assign n5513 = ( x116 & n2787 ) | ( x116 & ~n3114 ) | ( n2787 & ~n3114 ) ;
  assign n5514 = ~n3069 & n5513 ;
  assign n5515 = n5514 ^ n4316 ^ 1'b0 ;
  assign n5516 = n4035 ^ n908 ^ 1'b0 ;
  assign n5517 = n1389 & ~n5516 ;
  assign n5518 = x181 & n1522 ;
  assign n5519 = ~n271 & n5518 ;
  assign n5520 = x197 & n613 ;
  assign n5521 = n5519 & n5520 ;
  assign n5522 = n3860 & ~n5521 ;
  assign n5527 = n692 & n2087 ;
  assign n5528 = n5527 ^ n3140 ^ 1'b0 ;
  assign n5523 = ( ~n1172 & n1820 ) | ( ~n1172 & n3915 ) | ( n1820 & n3915 ) ;
  assign n5524 = n513 | n1487 ;
  assign n5525 = n5523 & ~n5524 ;
  assign n5526 = n1901 | n5525 ;
  assign n5529 = n5528 ^ n5526 ^ 1'b0 ;
  assign n5530 = n4744 ^ n3964 ^ 1'b0 ;
  assign n5531 = n2063 ^ x99 ^ 1'b0 ;
  assign n5532 = x38 & ~x217 ;
  assign n5533 = n2755 & n5532 ;
  assign n5534 = ~n5531 & n5533 ;
  assign n5535 = ( ~n3600 & n4400 ) | ( ~n3600 & n5534 ) | ( n4400 & n5534 ) ;
  assign n5536 = n1915 | n4766 ;
  assign n5537 = x48 & ~n3281 ;
  assign n5538 = n5537 ^ n1151 ^ 1'b0 ;
  assign n5539 = n3265 | n5538 ;
  assign n5540 = n1595 & ~n5414 ;
  assign n5541 = n417 & n5148 ;
  assign n5542 = n5541 ^ n1454 ^ n917 ;
  assign n5543 = n1336 ^ n308 ^ 1'b0 ;
  assign n5544 = n869 & n5543 ;
  assign n5545 = ~x180 & n5544 ;
  assign n5546 = x180 & n5545 ;
  assign n5547 = n2069 & n5546 ;
  assign n5548 = ~n2069 & n5547 ;
  assign n5549 = n5548 ^ n2304 ^ 1'b0 ;
  assign n5550 = n4918 ^ n1858 ^ 1'b0 ;
  assign n5551 = n4575 & ~n5550 ;
  assign n5552 = n5551 ^ n5528 ^ 1'b0 ;
  assign n5553 = n3647 & n5552 ;
  assign n5554 = ( n1393 & n1961 ) | ( n1393 & n3234 ) | ( n1961 & n3234 ) ;
  assign n5555 = n1404 | n2770 ;
  assign n5556 = n5555 ^ n2472 ^ 1'b0 ;
  assign n5557 = n534 ^ n325 ^ 1'b0 ;
  assign n5558 = ~n2248 & n5557 ;
  assign n5559 = n4210 & n5558 ;
  assign n5562 = n1272 ^ n1094 ^ 1'b0 ;
  assign n5563 = n3300 | n5562 ;
  assign n5564 = n2743 | n5563 ;
  assign n5565 = n869 | n5564 ;
  assign n5566 = n5565 ^ n2915 ^ 1'b0 ;
  assign n5560 = n2638 ^ x114 ^ 1'b0 ;
  assign n5561 = ~n810 & n5560 ;
  assign n5567 = n5566 ^ n5561 ^ 1'b0 ;
  assign n5568 = n904 & ~n5567 ;
  assign n5569 = ~n1206 & n4203 ;
  assign n5570 = n964 ^ x49 ^ 1'b0 ;
  assign n5571 = n3614 & ~n5570 ;
  assign n5572 = n5569 & ~n5571 ;
  assign n5573 = n1813 & n5572 ;
  assign n5574 = n2358 | n3494 ;
  assign n5575 = n1615 & ~n2135 ;
  assign n5576 = n5575 ^ n2870 ^ 1'b0 ;
  assign n5577 = n2528 ^ n1304 ^ 1'b0 ;
  assign n5578 = ~n2714 & n5577 ;
  assign n5579 = n2857 ^ n2326 ^ 1'b0 ;
  assign n5580 = n4197 ^ n2245 ^ n746 ;
  assign n5581 = n5579 & n5580 ;
  assign n5582 = n5581 ^ n3685 ^ x88 ;
  assign n5583 = ~n4264 & n5582 ;
  assign n5584 = n908 | n1203 ;
  assign n5585 = n5584 ^ n3806 ^ 1'b0 ;
  assign n5586 = n1861 & ~n2884 ;
  assign n5587 = n2306 ^ n2294 ^ 1'b0 ;
  assign n5588 = n5586 & n5587 ;
  assign n5589 = n4545 & n5588 ;
  assign n5590 = ~n1378 & n2365 ;
  assign n5591 = n1322 ^ x147 ^ 1'b0 ;
  assign n5592 = ~n5554 & n5591 ;
  assign n5593 = ~n5590 & n5592 ;
  assign n5594 = n5589 & n5593 ;
  assign n5595 = x44 & n3670 ;
  assign n5596 = ( x92 & ~x192 ) | ( x92 & n4415 ) | ( ~x192 & n4415 ) ;
  assign n5597 = n5596 ^ n4859 ^ 1'b0 ;
  assign n5598 = ~n755 & n5597 ;
  assign n5604 = n3866 ^ n300 ^ 1'b0 ;
  assign n5599 = ~n2112 & n2341 ;
  assign n5600 = n5599 ^ n3527 ^ 1'b0 ;
  assign n5601 = x6 & n5600 ;
  assign n5602 = n4025 & n5601 ;
  assign n5603 = n5367 | n5602 ;
  assign n5605 = n5604 ^ n5603 ^ 1'b0 ;
  assign n5606 = ( n1931 & n3579 ) | ( n1931 & n4686 ) | ( n3579 & n4686 ) ;
  assign n5607 = n986 ^ n680 ^ 1'b0 ;
  assign n5608 = n1471 | n4003 ;
  assign n5609 = n5608 ^ n3513 ^ 1'b0 ;
  assign n5610 = ~n3291 & n5609 ;
  assign n5611 = n1025 ^ n361 ^ 1'b0 ;
  assign n5612 = n1105 | n5611 ;
  assign n5613 = n5610 | n5612 ;
  assign n5614 = n5253 ^ n2309 ^ 1'b0 ;
  assign n5615 = n448 | n5165 ;
  assign n5616 = n3172 | n5615 ;
  assign n5617 = n838 & ~n5616 ;
  assign n5618 = ( n1725 & n2267 ) | ( n1725 & ~n2552 ) | ( n2267 & ~n2552 ) ;
  assign n5619 = n5618 ^ n1980 ^ 1'b0 ;
  assign n5620 = n4157 ^ n3966 ^ 1'b0 ;
  assign n5621 = ~n5619 & n5620 ;
  assign n5622 = n5621 ^ n453 ^ 1'b0 ;
  assign n5623 = n3744 ^ n2188 ^ 1'b0 ;
  assign n5624 = n5623 ^ x119 ^ 1'b0 ;
  assign n5625 = n3388 & ~n5624 ;
  assign n5626 = x204 | n4662 ;
  assign n5627 = n5626 ^ n844 ^ 1'b0 ;
  assign n5628 = n5627 ^ n2110 ^ 1'b0 ;
  assign n5629 = n1274 & ~n4678 ;
  assign n5630 = n4737 & n5629 ;
  assign n5631 = n4626 | n5630 ;
  assign n5632 = x61 | n5631 ;
  assign n5633 = n3593 ^ x234 ^ 1'b0 ;
  assign n5634 = ~n264 & n5633 ;
  assign n5635 = n2442 ^ x163 ^ 1'b0 ;
  assign n5636 = n5635 ^ n3258 ^ 1'b0 ;
  assign n5637 = n5206 | n5636 ;
  assign n5638 = n665 | n4150 ;
  assign n5639 = n2521 & ~n5638 ;
  assign n5640 = n496 & n5639 ;
  assign n5641 = n3251 | n5640 ;
  assign n5642 = n1439 & ~n5641 ;
  assign n5643 = ~n332 & n3161 ;
  assign n5644 = n2482 & ~n2873 ;
  assign n5645 = n5644 ^ n3986 ^ 1'b0 ;
  assign n5646 = n844 & ~n3108 ;
  assign n5647 = n914 & n5646 ;
  assign n5648 = ~n5645 & n5647 ;
  assign n5649 = ~n5643 & n5648 ;
  assign n5650 = n2442 & n5454 ;
  assign n5651 = n2883 ^ n1519 ^ 1'b0 ;
  assign n5652 = n1521 ^ n485 ^ 1'b0 ;
  assign n5653 = n4249 & n5652 ;
  assign n5654 = ~n5651 & n5653 ;
  assign n5655 = n1654 ^ n970 ^ 1'b0 ;
  assign n5656 = ~x163 & n739 ;
  assign n5657 = n5656 ^ n577 ^ 1'b0 ;
  assign n5658 = ~n4319 & n5657 ;
  assign n5659 = ~n5655 & n5658 ;
  assign n5660 = n2504 ^ n2130 ^ n711 ;
  assign n5661 = n1255 | n2403 ;
  assign n5662 = n348 & ~n5661 ;
  assign n5663 = n5662 ^ n5341 ^ 1'b0 ;
  assign n5664 = n5660 & ~n5663 ;
  assign n5665 = n3339 & ~n4786 ;
  assign n5666 = ~n320 & n3226 ;
  assign n5667 = n5666 ^ n1915 ^ 1'b0 ;
  assign n5668 = n5667 ^ n2829 ^ 1'b0 ;
  assign n5669 = x6 & n970 ;
  assign n5670 = n2081 | n2809 ;
  assign n5671 = n5670 ^ n931 ^ 1'b0 ;
  assign n5672 = n5669 & n5671 ;
  assign n5673 = n5672 ^ n1602 ^ 1'b0 ;
  assign n5674 = n5673 ^ n5320 ^ 1'b0 ;
  assign n5675 = n5240 | n5674 ;
  assign n5679 = n2143 ^ x61 ^ 1'b0 ;
  assign n5676 = n1981 & n3096 ;
  assign n5677 = n3961 ^ n1100 ^ 1'b0 ;
  assign n5678 = n5676 | n5677 ;
  assign n5680 = n5679 ^ n5678 ^ 1'b0 ;
  assign n5681 = n5680 ^ n2086 ^ 1'b0 ;
  assign n5682 = n1681 & n5681 ;
  assign n5683 = n5682 ^ n3534 ^ 1'b0 ;
  assign n5684 = n2740 & ~n5465 ;
  assign n5685 = n5229 & n5684 ;
  assign n5686 = n5540 ^ n1487 ^ n943 ;
  assign n5695 = x175 & n2974 ;
  assign n5694 = n2305 & n4470 ;
  assign n5696 = n5695 ^ n5694 ^ 1'b0 ;
  assign n5687 = n2037 ^ n1465 ^ 1'b0 ;
  assign n5688 = n2169 | n5687 ;
  assign n5689 = n5688 ^ n1633 ^ 1'b0 ;
  assign n5690 = ~n1952 & n5689 ;
  assign n5691 = n5690 ^ n718 ^ 1'b0 ;
  assign n5692 = n2722 & n5691 ;
  assign n5693 = n3454 & n5692 ;
  assign n5697 = n5696 ^ n5693 ^ 1'b0 ;
  assign n5698 = ~n2950 & n3087 ;
  assign n5699 = ~n302 & n5078 ;
  assign n5700 = n5699 ^ n4642 ^ 1'b0 ;
  assign n5701 = n1711 & ~n5307 ;
  assign n5702 = n5374 & ~n5701 ;
  assign n5703 = n5702 ^ n426 ^ 1'b0 ;
  assign n5705 = n2148 | n4399 ;
  assign n5706 = n909 & ~n5705 ;
  assign n5707 = n5706 ^ n3785 ^ 1'b0 ;
  assign n5704 = n4053 ^ n928 ^ 1'b0 ;
  assign n5708 = n5707 ^ n5704 ^ n3572 ;
  assign n5709 = n3786 & n5373 ;
  assign n5710 = n1001 ^ x219 ^ 1'b0 ;
  assign n5711 = ~n5709 & n5710 ;
  assign n5712 = n5711 ^ n1681 ^ 1'b0 ;
  assign n5713 = ~n3712 & n5712 ;
  assign n5714 = n327 | n3706 ;
  assign n5715 = n370 & ~n5714 ;
  assign n5716 = n5715 ^ n3298 ^ 1'b0 ;
  assign n5717 = n3942 & ~n5716 ;
  assign n5718 = n4460 & n4535 ;
  assign n5719 = n2837 & n5718 ;
  assign n5720 = n2807 ^ n977 ^ 1'b0 ;
  assign n5721 = n263 & ~n3237 ;
  assign n5722 = n5721 ^ n694 ^ 1'b0 ;
  assign n5723 = n5722 ^ n1720 ^ 1'b0 ;
  assign n5724 = n2735 & n5723 ;
  assign n5725 = n5724 ^ n5413 ^ 1'b0 ;
  assign n5726 = ~n5720 & n5725 ;
  assign n5727 = n5726 ^ n3213 ^ 1'b0 ;
  assign n5728 = n413 & n3776 ;
  assign n5729 = n4175 ^ n1371 ^ 1'b0 ;
  assign n5730 = n1528 ^ n514 ^ 1'b0 ;
  assign n5731 = n3765 | n5730 ;
  assign n5732 = n5731 ^ n1716 ^ 1'b0 ;
  assign n5733 = n4239 & ~n5732 ;
  assign n5734 = n4130 ^ n3042 ^ 1'b0 ;
  assign n5735 = n2064 & ~n5734 ;
  assign n5736 = n523 & n891 ;
  assign n5737 = n496 & n5736 ;
  assign n5738 = n2158 ^ x131 ^ 1'b0 ;
  assign n5739 = n5737 | n5738 ;
  assign n5741 = n423 | n3719 ;
  assign n5742 = n5741 ^ n3253 ^ 1'b0 ;
  assign n5740 = n621 & ~n3037 ;
  assign n5743 = n5742 ^ n5740 ^ 1'b0 ;
  assign n5744 = n5739 | n5743 ;
  assign n5745 = n3915 & ~n5744 ;
  assign n5746 = n1200 ^ n1168 ^ 1'b0 ;
  assign n5747 = n3734 ^ x252 ^ 1'b0 ;
  assign n5748 = ~n3702 & n5747 ;
  assign n5749 = n5473 ^ n1433 ^ 1'b0 ;
  assign n5750 = n4269 ^ n2376 ^ 1'b0 ;
  assign n5751 = n1547 & n5750 ;
  assign n5752 = n1010 & n5751 ;
  assign n5753 = n1780 ^ x145 ^ 1'b0 ;
  assign n5754 = n5560 & ~n5753 ;
  assign n5755 = ~n450 & n5754 ;
  assign n5756 = ~n5218 & n5755 ;
  assign n5757 = n3160 & ~n5756 ;
  assign n5758 = n5054 & n5757 ;
  assign n5759 = ( x187 & ~n5752 ) | ( x187 & n5758 ) | ( ~n5752 & n5758 ) ;
  assign n5760 = n2424 & ~n4473 ;
  assign n5761 = n5760 ^ n1379 ^ 1'b0 ;
  assign n5762 = n5759 & ~n5761 ;
  assign n5763 = ~n4937 & n5762 ;
  assign n5764 = n3885 ^ n3853 ^ 1'b0 ;
  assign n5765 = n1654 | n5764 ;
  assign n5766 = ~n863 & n4693 ;
  assign n5767 = n5766 ^ n4008 ^ 1'b0 ;
  assign n5768 = n5767 ^ n4553 ^ 1'b0 ;
  assign n5769 = x163 & n3116 ;
  assign n5770 = ( ~n1079 & n1371 ) | ( ~n1079 & n3196 ) | ( n1371 & n3196 ) ;
  assign n5771 = n5209 & n5770 ;
  assign n5772 = n2343 ^ n353 ^ 1'b0 ;
  assign n5773 = n1992 ^ x7 ^ 1'b0 ;
  assign n5774 = x8 & ~n3195 ;
  assign n5775 = n3451 ^ n613 ^ 1'b0 ;
  assign n5776 = x185 & n4047 ;
  assign n5777 = n4042 & n5776 ;
  assign n5778 = n5777 ^ n5442 ^ 1'b0 ;
  assign n5779 = ~n5775 & n5778 ;
  assign n5780 = ~n5066 & n5779 ;
  assign n5781 = n1965 ^ n1406 ^ 1'b0 ;
  assign n5782 = n3689 & n5781 ;
  assign n5783 = n5782 ^ n3668 ^ n890 ;
  assign n5784 = x252 & ~n4277 ;
  assign n5785 = ~n722 & n5784 ;
  assign n5786 = n5785 ^ n5350 ^ 1'b0 ;
  assign n5787 = n4209 ^ x78 ^ 1'b0 ;
  assign n5788 = n5786 & ~n5787 ;
  assign n5789 = n1459 ^ n1254 ^ 1'b0 ;
  assign n5790 = x108 & n5789 ;
  assign n5791 = n1798 & n5790 ;
  assign n5792 = n5791 ^ n5082 ^ 1'b0 ;
  assign n5793 = n2258 ^ n591 ^ 1'b0 ;
  assign n5794 = n5792 & n5793 ;
  assign n5795 = n2703 ^ n1654 ^ 1'b0 ;
  assign n5796 = n1441 ^ n961 ^ 1'b0 ;
  assign n5797 = ( ~n1067 & n5727 ) | ( ~n1067 & n5796 ) | ( n5727 & n5796 ) ;
  assign n5798 = n486 & n691 ;
  assign n5799 = ( n1389 & ~n2718 ) | ( n1389 & n3910 ) | ( ~n2718 & n3910 ) ;
  assign n5800 = ( n1213 & ~n5798 ) | ( n1213 & n5799 ) | ( ~n5798 & n5799 ) ;
  assign n5801 = n4572 & n5800 ;
  assign n5802 = n5801 ^ n714 ^ 1'b0 ;
  assign n5803 = n1615 & n5442 ;
  assign n5804 = n4296 ^ n3551 ^ n699 ;
  assign n5805 = n2767 & n5804 ;
  assign n5806 = ~n4788 & n5805 ;
  assign n5809 = n723 | n2878 ;
  assign n5810 = n5809 ^ n547 ^ 1'b0 ;
  assign n5808 = n491 | n4715 ;
  assign n5811 = n5810 ^ n5808 ^ 1'b0 ;
  assign n5807 = ~n2127 & n2414 ;
  assign n5812 = n5811 ^ n5807 ^ 1'b0 ;
  assign n5813 = n5812 ^ n3518 ^ 1'b0 ;
  assign n5814 = n387 & n1311 ;
  assign n5815 = n5814 ^ n1495 ^ 1'b0 ;
  assign n5816 = n3081 | n5815 ;
  assign n5817 = n1659 ^ x101 ^ 1'b0 ;
  assign n5818 = ~n2881 & n5817 ;
  assign n5819 = n2150 & n5818 ;
  assign n5820 = ~n732 & n5819 ;
  assign n5821 = n1086 & ~n5820 ;
  assign n5822 = n1135 & ~n5821 ;
  assign n5823 = ~n3614 & n5822 ;
  assign n5824 = n738 & n1909 ;
  assign n5825 = n5824 ^ n1864 ^ 1'b0 ;
  assign n5826 = n3085 ^ n3078 ^ 1'b0 ;
  assign n5827 = n5179 & n5826 ;
  assign n5828 = n1151 & ~n4553 ;
  assign n5829 = ~n5172 & n5828 ;
  assign n5830 = n369 & n575 ;
  assign n5831 = n5830 ^ n629 ^ 1'b0 ;
  assign n5832 = n992 ^ x153 ^ 1'b0 ;
  assign n5833 = n2615 & ~n5832 ;
  assign n5834 = n5831 & n5833 ;
  assign n5835 = ~n2633 & n5834 ;
  assign n5836 = n4977 | n5435 ;
  assign n5837 = n497 & n4914 ;
  assign n5838 = ~n899 & n1276 ;
  assign n5839 = n5069 ^ x86 ^ 1'b0 ;
  assign n5844 = n3377 ^ x187 ^ 1'b0 ;
  assign n5845 = ~n3300 & n5844 ;
  assign n5840 = ~n1593 & n2666 ;
  assign n5841 = n1219 & n5840 ;
  assign n5842 = ~n916 & n5841 ;
  assign n5843 = n4241 | n5842 ;
  assign n5846 = n5845 ^ n5843 ^ 1'b0 ;
  assign n5847 = n5846 ^ n2804 ^ n1206 ;
  assign n5848 = n3772 & n5847 ;
  assign n5849 = n5848 ^ n5425 ^ 1'b0 ;
  assign n5850 = n4125 & ~n5120 ;
  assign n5851 = ~n1803 & n5850 ;
  assign n5852 = n1558 & n3546 ;
  assign n5853 = ~n2466 & n5852 ;
  assign n5854 = ~n372 & n869 ;
  assign n5855 = n5854 ^ n391 ^ 1'b0 ;
  assign n5856 = x55 | n5855 ;
  assign n5857 = n1062 ^ n992 ^ 1'b0 ;
  assign n5858 = ~n3464 & n5857 ;
  assign n5859 = n3168 ^ n2026 ^ 1'b0 ;
  assign n5860 = n5858 & ~n5859 ;
  assign n5861 = n5856 & n5860 ;
  assign n5862 = n5853 | n5861 ;
  assign n5863 = n5284 ^ n3191 ^ 1'b0 ;
  assign n5864 = n2848 | n5863 ;
  assign n5865 = n1369 & ~n1413 ;
  assign n5866 = n2865 & ~n5135 ;
  assign n5867 = n1696 | n5156 ;
  assign n5868 = n5867 ^ n643 ^ 1'b0 ;
  assign n5869 = ~n1530 & n5868 ;
  assign n5870 = n1494 & n5365 ;
  assign n5871 = n431 & n1160 ;
  assign n5873 = n1905 ^ n357 ^ 1'b0 ;
  assign n5872 = n668 & ~n1254 ;
  assign n5874 = n5873 ^ n5872 ^ 1'b0 ;
  assign n5875 = ~n2310 & n5874 ;
  assign n5876 = n1071 & n5875 ;
  assign n5877 = n5871 & ~n5876 ;
  assign n5878 = n3470 & n5877 ;
  assign n5879 = n5878 ^ n3567 ^ n2462 ;
  assign n5880 = x189 & ~n3802 ;
  assign n5881 = n5880 ^ n1731 ^ 1'b0 ;
  assign n5882 = n5881 ^ n293 ^ 1'b0 ;
  assign n5883 = n4881 & n5882 ;
  assign n5884 = ( n425 & n1049 ) | ( n425 & n1422 ) | ( n1049 & n1422 ) ;
  assign n5885 = n3326 | n5884 ;
  assign n5886 = n5587 ^ n4911 ^ 1'b0 ;
  assign n5887 = ~n5885 & n5886 ;
  assign n5888 = ( n2143 & n2556 ) | ( n2143 & n5887 ) | ( n2556 & n5887 ) ;
  assign n5889 = n5888 ^ n3062 ^ 1'b0 ;
  assign n5890 = ~n3839 & n5889 ;
  assign n5891 = n5683 ^ n1698 ^ 1'b0 ;
  assign n5892 = n1623 | n2585 ;
  assign n5893 = n938 & ~n5892 ;
  assign n5894 = n5893 ^ n2110 ^ 1'b0 ;
  assign n5895 = n5457 ^ n4241 ^ 1'b0 ;
  assign n5896 = ( ~n1276 & n2095 ) | ( ~n1276 & n5659 ) | ( n2095 & n5659 ) ;
  assign n5897 = n287 | n370 ;
  assign n5898 = n2002 | n5897 ;
  assign n5899 = ~n2513 & n5898 ;
  assign n5900 = n899 & n5899 ;
  assign n5904 = n1575 ^ n915 ^ 1'b0 ;
  assign n5901 = x92 & n2353 ;
  assign n5902 = n5901 ^ n1960 ^ 1'b0 ;
  assign n5903 = n5902 ^ n5885 ^ 1'b0 ;
  assign n5905 = n5904 ^ n5903 ^ n3126 ;
  assign n5906 = ~n276 & n2367 ;
  assign n5907 = n2097 ^ x92 ^ 1'b0 ;
  assign n5908 = n5906 & ~n5907 ;
  assign n5909 = n2106 ^ n935 ^ x185 ;
  assign n5910 = ~n1867 & n5909 ;
  assign n5911 = n1727 & n5910 ;
  assign n5912 = n1561 ^ n1170 ^ 1'b0 ;
  assign n5913 = n2974 | n5912 ;
  assign n5914 = n3917 ^ n550 ^ 1'b0 ;
  assign n5915 = n649 & n5914 ;
  assign n5916 = n5915 ^ n1891 ^ 1'b0 ;
  assign n5917 = n2369 & ~n5916 ;
  assign n5918 = n2989 | n3328 ;
  assign n5919 = n5918 ^ n4236 ^ n413 ;
  assign n5920 = n2513 ^ x213 ^ 1'b0 ;
  assign n5921 = n812 | n5920 ;
  assign n5922 = x96 & n5921 ;
  assign n5923 = ~n5919 & n5922 ;
  assign n5924 = n5923 ^ n1081 ^ 1'b0 ;
  assign n5925 = n344 & n2625 ;
  assign n5926 = n5708 ^ n4742 ^ 1'b0 ;
  assign n5927 = n5925 | n5926 ;
  assign n5928 = n3010 & ~n4261 ;
  assign n5929 = n3754 ^ n2062 ^ 1'b0 ;
  assign n5930 = n2511 & n5929 ;
  assign n5931 = n1813 | n5798 ;
  assign n5932 = n2615 & n2657 ;
  assign n5933 = ~n5931 & n5932 ;
  assign n5934 = n5933 ^ n3265 ^ 1'b0 ;
  assign n5935 = x110 & n2779 ;
  assign n5936 = ~n5459 & n5935 ;
  assign n5937 = n2416 ^ n1381 ^ 1'b0 ;
  assign n5938 = n5937 ^ n2946 ^ 1'b0 ;
  assign n5939 = x13 & ~n5938 ;
  assign n5940 = ~n2843 & n4983 ;
  assign n5941 = n5940 ^ n4226 ^ 1'b0 ;
  assign n5942 = n1815 | n3419 ;
  assign n5943 = n5942 ^ n2604 ^ n891 ;
  assign n5944 = ~n604 & n2929 ;
  assign n5945 = n744 | n2337 ;
  assign n5946 = n3874 & ~n5945 ;
  assign n5947 = n1586 | n3900 ;
  assign n5948 = n3845 & ~n5947 ;
  assign n5949 = n5948 ^ n937 ^ 1'b0 ;
  assign n5950 = n5949 ^ n327 ^ 1'b0 ;
  assign n5951 = n5946 | n5950 ;
  assign n5952 = n2542 & n4708 ;
  assign n5953 = ~x75 & n5952 ;
  assign n5954 = n5953 ^ n2674 ^ 1'b0 ;
  assign n5955 = n5954 ^ x248 ^ 1'b0 ;
  assign n5956 = n5012 ^ n3339 ^ 1'b0 ;
  assign n5957 = n5955 | n5956 ;
  assign n5958 = n3210 ^ n2915 ^ 1'b0 ;
  assign n5959 = ( n1622 & ~n3352 ) | ( n1622 & n5958 ) | ( ~n3352 & n5958 ) ;
  assign n5960 = n3367 ^ n862 ^ 1'b0 ;
  assign n5961 = n3433 & ~n5960 ;
  assign n5962 = n707 & n3105 ;
  assign n5963 = ( ~x201 & n1553 ) | ( ~x201 & n4918 ) | ( n1553 & n4918 ) ;
  assign n5964 = n5963 ^ n4626 ^ 1'b0 ;
  assign n5965 = n3645 & n5964 ;
  assign n5966 = n5749 & ~n5965 ;
  assign n5967 = n3059 ^ n1312 ^ 1'b0 ;
  assign n5968 = n835 | n1575 ;
  assign n5969 = n5968 ^ n1086 ^ 1'b0 ;
  assign n5970 = n1333 & ~n5969 ;
  assign n5971 = n5970 ^ n3542 ^ 1'b0 ;
  assign n5972 = n2184 ^ n1219 ^ 1'b0 ;
  assign n5973 = n2775 & ~n5972 ;
  assign n5974 = n5973 ^ n4976 ^ 1'b0 ;
  assign n5975 = ~n5608 & n5974 ;
  assign n5976 = ( n488 & ~n1890 ) | ( n488 & n2655 ) | ( ~n1890 & n2655 ) ;
  assign n5977 = n2262 ^ n817 ^ 1'b0 ;
  assign n5978 = ~n1905 & n5977 ;
  assign n5979 = x248 & ~n4434 ;
  assign n5980 = n1147 & n5979 ;
  assign n5982 = n5569 ^ n4029 ^ 1'b0 ;
  assign n5983 = n5146 & ~n5982 ;
  assign n5981 = x116 & n2625 ;
  assign n5984 = n5983 ^ n5981 ^ 1'b0 ;
  assign n5985 = x118 & ~n5088 ;
  assign n5986 = n5985 ^ n4203 ^ 1'b0 ;
  assign n5987 = n1118 | n1306 ;
  assign n5988 = n5796 ^ n4615 ^ 1'b0 ;
  assign n5989 = ~n5987 & n5988 ;
  assign n5990 = ~n2633 & n5989 ;
  assign n5991 = n4372 | n5990 ;
  assign n5992 = n5991 ^ n1071 ^ 1'b0 ;
  assign n5993 = n1990 ^ n1925 ^ 1'b0 ;
  assign n5994 = ~n651 & n5993 ;
  assign n5995 = ( n4465 & ~n5742 ) | ( n4465 & n5994 ) | ( ~n5742 & n5994 ) ;
  assign n5996 = n1961 & n5273 ;
  assign n5998 = n2013 ^ n1230 ^ x69 ;
  assign n5997 = n2659 ^ n589 ^ 1'b0 ;
  assign n5999 = n5998 ^ n5997 ^ n1947 ;
  assign n6000 = n1776 & n5246 ;
  assign n6001 = ~n3647 & n6000 ;
  assign n6002 = n3407 & ~n6001 ;
  assign n6003 = ~n3362 & n6002 ;
  assign n6004 = n6003 ^ n724 ^ 1'b0 ;
  assign n6005 = n2424 & ~n6004 ;
  assign n6006 = n2161 ^ x115 ^ 1'b0 ;
  assign n6007 = n4347 ^ n2085 ^ 1'b0 ;
  assign n6008 = x243 | n6007 ;
  assign n6009 = n6008 ^ n5354 ^ 1'b0 ;
  assign n6010 = n5058 & n5234 ;
  assign n6011 = n1432 ^ n701 ^ 1'b0 ;
  assign n6012 = n5790 & ~n6011 ;
  assign n6013 = n975 & n6012 ;
  assign n6014 = n6013 ^ n4458 ^ 1'b0 ;
  assign n6015 = n5225 ^ n2816 ^ 1'b0 ;
  assign n6016 = ~n2109 & n2724 ;
  assign n6017 = n6016 ^ n4684 ^ 1'b0 ;
  assign n6018 = n6017 ^ n1980 ^ 1'b0 ;
  assign n6019 = n4718 ^ n3930 ^ x176 ;
  assign n6020 = ~n613 & n970 ;
  assign n6021 = n4925 ^ n2426 ^ 1'b0 ;
  assign n6022 = ~n6020 & n6021 ;
  assign n6023 = n2284 & n6022 ;
  assign n6024 = n3804 & n6023 ;
  assign n6025 = n2714 ^ n1478 ^ 1'b0 ;
  assign n6026 = x185 & n4213 ;
  assign n6027 = n1163 & n6026 ;
  assign n6029 = ~n638 & n1522 ;
  assign n6030 = n6029 ^ x201 ^ 1'b0 ;
  assign n6028 = n1983 & n4817 ;
  assign n6031 = n6030 ^ n6028 ^ 1'b0 ;
  assign n6032 = n1756 & ~n2410 ;
  assign n6033 = n5390 & n6032 ;
  assign n6034 = n6033 ^ n4975 ^ 1'b0 ;
  assign n6035 = n6031 & n6034 ;
  assign n6036 = ~n628 & n4944 ;
  assign n6037 = ~n1973 & n3486 ;
  assign n6038 = n2963 & ~n6037 ;
  assign n6039 = x85 & n6038 ;
  assign n6040 = n1958 & n6039 ;
  assign n6041 = ~n1579 & n4670 ;
  assign n6042 = n6041 ^ n847 ^ 1'b0 ;
  assign n6043 = n2989 ^ n1961 ^ 1'b0 ;
  assign n6044 = n5645 ^ n2602 ^ 1'b0 ;
  assign n6045 = n2157 & ~n6044 ;
  assign n6046 = n6045 ^ n3407 ^ 1'b0 ;
  assign n6047 = n2556 ^ n1521 ^ 1'b0 ;
  assign n6048 = n1947 & ~n6047 ;
  assign n6049 = n2458 ^ n2375 ^ n890 ;
  assign n6050 = n1190 & n6049 ;
  assign n6051 = ~n2767 & n6050 ;
  assign n6052 = n3755 & ~n6051 ;
  assign n6053 = ~n6048 & n6052 ;
  assign n6054 = n1671 & ~n6053 ;
  assign n6055 = n6054 ^ n5617 ^ 1'b0 ;
  assign n6056 = n1360 ^ n1034 ^ 1'b0 ;
  assign n6057 = n3110 & n6056 ;
  assign n6058 = n6057 ^ n3655 ^ n2010 ;
  assign n6059 = ( x84 & n1822 ) | ( x84 & ~n2807 ) | ( n1822 & ~n2807 ) ;
  assign n6060 = n1125 & n6059 ;
  assign n6061 = n3796 | n6060 ;
  assign n6062 = ~n1575 & n5333 ;
  assign n6063 = n5610 & ~n6062 ;
  assign n6064 = n6063 ^ n919 ^ 1'b0 ;
  assign n6065 = n6064 ^ n1039 ^ 1'b0 ;
  assign n6066 = ~n4138 & n6065 ;
  assign n6067 = n1219 ^ n466 ^ 1'b0 ;
  assign n6068 = n2086 | n3007 ;
  assign n6069 = n6067 & ~n6068 ;
  assign n6070 = n1105 ^ n547 ^ 1'b0 ;
  assign n6071 = n3348 | n6070 ;
  assign n6072 = n6069 & ~n6071 ;
  assign n6073 = n4227 ^ n2957 ^ n2172 ;
  assign n6074 = ~n2311 & n5729 ;
  assign n6075 = n6074 ^ n2182 ^ 1'b0 ;
  assign n6076 = n2262 & n5915 ;
  assign n6077 = ~x90 & n6076 ;
  assign n6078 = n3631 & ~n6077 ;
  assign n6079 = n6078 ^ n402 ^ 1'b0 ;
  assign n6080 = ( n970 & ~n5662 ) | ( n970 & n6079 ) | ( ~n5662 & n6079 ) ;
  assign n6081 = n6080 ^ n2183 ^ 1'b0 ;
  assign n6082 = x62 & ~n1931 ;
  assign n6083 = ~n1416 & n6082 ;
  assign n6084 = n2301 | n6083 ;
  assign n6085 = n6084 ^ n3419 ^ 1'b0 ;
  assign n6086 = n5922 ^ n2232 ^ 1'b0 ;
  assign n6088 = n2983 ^ x46 ^ 1'b0 ;
  assign n6089 = n4950 & ~n6088 ;
  assign n6090 = n3400 & n6089 ;
  assign n6087 = n2001 | n2975 ;
  assign n6091 = n6090 ^ n6087 ^ 1'b0 ;
  assign n6092 = n1696 & n2110 ;
  assign n6093 = n6092 ^ n2165 ^ 1'b0 ;
  assign n6094 = n455 ^ x43 ^ 1'b0 ;
  assign n6095 = n659 & ~n1272 ;
  assign n6096 = n6094 | n6095 ;
  assign n6097 = n6093 & ~n6096 ;
  assign n6098 = ( x138 & n2020 ) | ( x138 & ~n5848 ) | ( n2020 & ~n5848 ) ;
  assign n6099 = n1361 ^ n529 ^ 1'b0 ;
  assign n6100 = n854 & ~n6099 ;
  assign n6101 = n776 & n6100 ;
  assign n6102 = n6101 ^ n5160 ^ n1078 ;
  assign n6103 = n2840 | n2957 ;
  assign n6104 = n1937 & ~n6103 ;
  assign n6105 = n6104 ^ n1499 ^ 1'b0 ;
  assign n6106 = ~n1292 & n6105 ;
  assign n6107 = n930 & ~n2102 ;
  assign n6108 = n2747 & ~n6107 ;
  assign n6109 = ~n1466 & n6108 ;
  assign n6110 = n6109 ^ x19 ^ 1'b0 ;
  assign n6111 = n957 ^ x162 ^ 1'b0 ;
  assign n6112 = n6111 ^ n5124 ^ n2900 ;
  assign n6113 = n6110 & n6112 ;
  assign n6114 = n6106 & ~n6113 ;
  assign n6115 = ~n2348 & n3178 ;
  assign n6116 = n2406 ^ n2254 ^ 1'b0 ;
  assign n6117 = n6116 ^ n1244 ^ 1'b0 ;
  assign n6118 = ( n688 & ~n1733 ) | ( n688 & n2574 ) | ( ~n1733 & n2574 ) ;
  assign n6119 = n6118 ^ n1708 ^ 1'b0 ;
  assign n6120 = n6119 ^ n3606 ^ 1'b0 ;
  assign n6121 = x45 | n5963 ;
  assign n6122 = n2566 ^ n2262 ^ 1'b0 ;
  assign n6123 = n2385 | n5538 ;
  assign n6124 = n2738 & ~n6123 ;
  assign n6125 = ~n6122 & n6124 ;
  assign n6127 = n513 & n2137 ;
  assign n6126 = n2778 | n5398 ;
  assign n6128 = n6127 ^ n6126 ^ 1'b0 ;
  assign n6129 = n2845 ^ n1441 ^ 1'b0 ;
  assign n6130 = n6129 ^ n2580 ^ 1'b0 ;
  assign n6131 = ~n3822 & n6130 ;
  assign n6132 = n2122 ^ n491 ^ 1'b0 ;
  assign n6133 = ~n411 & n6132 ;
  assign n6134 = n6131 & n6133 ;
  assign n6135 = n560 & n1931 ;
  assign n6136 = n1125 & ~n6135 ;
  assign n6137 = ~n336 & n6136 ;
  assign n6138 = n4027 ^ n1812 ^ 1'b0 ;
  assign n6139 = ~n1684 & n6138 ;
  assign n6140 = ( x75 & n2070 ) | ( x75 & ~n2446 ) | ( n2070 & ~n2446 ) ;
  assign n6141 = n747 | n2103 ;
  assign n6142 = n6141 ^ n2622 ^ 1'b0 ;
  assign n6143 = n2614 | n6142 ;
  assign n6144 = ~n6140 & n6143 ;
  assign n6145 = n5138 ^ n3400 ^ n917 ;
  assign n6146 = n6049 & ~n6145 ;
  assign n6147 = n1585 | n2853 ;
  assign n6148 = n3007 & n6147 ;
  assign n6149 = n946 ^ n809 ^ 1'b0 ;
  assign n6150 = n2540 & n6149 ;
  assign n6151 = n6150 ^ n3126 ^ 1'b0 ;
  assign n6152 = n6151 ^ n2687 ^ 1'b0 ;
  assign n6153 = n854 | n871 ;
  assign n6154 = n6153 ^ n4238 ^ 1'b0 ;
  assign n6155 = n4502 ^ n1474 ^ 1'b0 ;
  assign n6156 = n1903 ^ n941 ^ 1'b0 ;
  assign n6157 = n6155 | n6156 ;
  assign n6158 = n6157 ^ n4826 ^ n2694 ;
  assign n6159 = n459 & ~n847 ;
  assign n6160 = n2044 & ~n6159 ;
  assign n6161 = n2714 ^ n1249 ^ 1'b0 ;
  assign n6162 = n3542 & ~n6161 ;
  assign n6163 = n6162 ^ n5175 ^ 1'b0 ;
  assign n6164 = n2064 & ~n3766 ;
  assign n6165 = n4843 ^ n1958 ^ 1'b0 ;
  assign n6166 = ~n3814 & n6165 ;
  assign n6167 = ~n473 & n3216 ;
  assign n6168 = n6167 ^ n3113 ^ 1'b0 ;
  assign n6169 = ( n1378 & n3126 ) | ( n1378 & ~n6168 ) | ( n3126 & ~n6168 ) ;
  assign n6170 = n6169 ^ n4178 ^ 1'b0 ;
  assign n6171 = n4827 & ~n6170 ;
  assign n6172 = ~n5094 & n6171 ;
  assign n6173 = n2967 & n6172 ;
  assign n6174 = n4673 ^ n2420 ^ 1'b0 ;
  assign n6175 = n4165 | n6174 ;
  assign n6176 = n5308 ^ n2240 ^ 1'b0 ;
  assign n6177 = n3493 & ~n6176 ;
  assign n6178 = n862 & ~n1566 ;
  assign n6179 = n3483 & n6178 ;
  assign n6180 = ( ~n579 & n2500 ) | ( ~n579 & n6179 ) | ( n2500 & n6179 ) ;
  assign n6181 = n1478 & ~n5010 ;
  assign n6182 = ~n6002 & n6181 ;
  assign n6183 = n4726 | n6182 ;
  assign n6184 = n4728 | n6183 ;
  assign n6188 = n621 & n3234 ;
  assign n6185 = n1606 & ~n5731 ;
  assign n6186 = n6185 ^ n1244 ^ 1'b0 ;
  assign n6187 = n560 & n6186 ;
  assign n6189 = n6188 ^ n6187 ^ 1'b0 ;
  assign n6190 = n4563 & n6189 ;
  assign n6191 = x143 | n6190 ;
  assign n6192 = n581 | n6191 ;
  assign n6193 = n1004 ^ x43 ^ 1'b0 ;
  assign n6194 = ~n471 & n6193 ;
  assign n6195 = n6194 ^ n2554 ^ 1'b0 ;
  assign n6196 = n3382 & n6195 ;
  assign n6197 = ~n6192 & n6196 ;
  assign n6198 = n4554 | n5461 ;
  assign n6199 = ( ~n1600 & n3160 ) | ( ~n1600 & n4698 ) | ( n3160 & n4698 ) ;
  assign n6200 = n3075 ^ n2070 ^ 1'b0 ;
  assign n6201 = n3293 ^ n1680 ^ 1'b0 ;
  assign n6202 = n776 & ~n3703 ;
  assign n6203 = ( n3149 & n6201 ) | ( n3149 & ~n6202 ) | ( n6201 & ~n6202 ) ;
  assign n6204 = n3460 & ~n3858 ;
  assign n6205 = ~n2203 & n3307 ;
  assign n6206 = n847 & n6205 ;
  assign n6207 = n3300 | n6206 ;
  assign n6208 = n2679 & n5357 ;
  assign n6209 = ~n2587 & n5356 ;
  assign n6210 = ~n809 & n6209 ;
  assign n6211 = n3696 ^ x32 ^ 1'b0 ;
  assign n6212 = n6211 ^ n1295 ^ x192 ;
  assign n6213 = n5611 ^ x87 ^ 1'b0 ;
  assign n6214 = n4496 & ~n6213 ;
  assign n6215 = n3745 & n6214 ;
  assign n6216 = n6215 ^ n4972 ^ 1'b0 ;
  assign n6217 = n6216 ^ n3395 ^ 1'b0 ;
  assign n6218 = n5925 | n6217 ;
  assign n6219 = n917 & ~n2622 ;
  assign n6220 = n5726 ^ n4141 ^ 1'b0 ;
  assign n6221 = n6220 ^ n4563 ^ 1'b0 ;
  assign n6222 = n4174 & n6221 ;
  assign n6223 = n850 ^ x157 ^ 1'b0 ;
  assign n6224 = x145 & n6223 ;
  assign n6225 = n6224 ^ n4080 ^ 1'b0 ;
  assign n6232 = n829 | n2710 ;
  assign n6233 = n6232 ^ x7 ^ 1'b0 ;
  assign n6234 = n6233 ^ n361 ^ 1'b0 ;
  assign n6235 = n2254 | n6234 ;
  assign n6236 = n1983 & n6235 ;
  assign n6229 = n5937 ^ n3728 ^ 1'b0 ;
  assign n6230 = x66 | n6229 ;
  assign n6226 = n5688 ^ n3845 ^ 1'b0 ;
  assign n6227 = n3213 ^ n1864 ^ n1799 ;
  assign n6228 = n6226 | n6227 ;
  assign n6231 = n6230 ^ n6228 ^ 1'b0 ;
  assign n6237 = n6236 ^ n6231 ^ 1'b0 ;
  assign n6238 = n1311 & ~n6237 ;
  assign n6239 = n2206 & ~n4166 ;
  assign n6240 = ~x183 & n6239 ;
  assign n6241 = n4595 & n6240 ;
  assign n6242 = n1879 & n5671 ;
  assign n6243 = ~n1065 & n6242 ;
  assign n6245 = n3086 | n3290 ;
  assign n6246 = n2710 & ~n6245 ;
  assign n6247 = n6246 ^ n3880 ^ 1'b0 ;
  assign n6248 = ~n928 & n6247 ;
  assign n6249 = ~n5842 & n6248 ;
  assign n6250 = n6249 ^ n5373 ^ 1'b0 ;
  assign n6244 = n1723 & ~n5769 ;
  assign n6251 = n6250 ^ n6244 ^ 1'b0 ;
  assign n6252 = n529 | n4657 ;
  assign n6253 = n3327 | n4572 ;
  assign n6254 = ( n445 & ~n6252 ) | ( n445 & n6253 ) | ( ~n6252 & n6253 ) ;
  assign n6255 = n3253 ^ n2296 ^ 1'b0 ;
  assign n6256 = ~x51 & n5646 ;
  assign n6259 = x159 & ~n3237 ;
  assign n6257 = n1720 ^ n1060 ^ x180 ;
  assign n6258 = ~n5390 & n6257 ;
  assign n6260 = n6259 ^ n6258 ^ 1'b0 ;
  assign n6261 = n6260 ^ n4222 ^ 1'b0 ;
  assign n6262 = ~n1583 & n6261 ;
  assign n6263 = n6256 & n6262 ;
  assign n6264 = n3651 & ~n4302 ;
  assign n6265 = n6264 ^ n3665 ^ 1'b0 ;
  assign n6266 = n5840 ^ n2157 ^ 1'b0 ;
  assign n6267 = n2678 & n6266 ;
  assign n6268 = n5887 & ~n6166 ;
  assign n6271 = n724 ^ x139 ^ 1'b0 ;
  assign n6272 = n450 | n6271 ;
  assign n6269 = n659 & ~n2484 ;
  assign n6270 = n6269 ^ n5153 ^ n2719 ;
  assign n6273 = n6272 ^ n6270 ^ 1'b0 ;
  assign n6274 = n854 | n1361 ;
  assign n6275 = n283 & ~n6274 ;
  assign n6276 = n6275 ^ n1710 ^ 1'b0 ;
  assign n6277 = n6273 & ~n6276 ;
  assign n6278 = ~x113 & n6277 ;
  assign n6279 = n606 | n1772 ;
  assign n6280 = n6279 ^ n2161 ^ 1'b0 ;
  assign n6281 = ~n4633 & n5827 ;
  assign n6282 = n3819 ^ n2589 ^ n1478 ;
  assign n6283 = ~n668 & n5350 ;
  assign n6284 = ~n6282 & n6283 ;
  assign n6285 = n1132 ^ n740 ^ 1'b0 ;
  assign n6286 = n2747 & n6285 ;
  assign n6287 = ~n5771 & n6286 ;
  assign n6288 = n6287 ^ n1880 ^ 1'b0 ;
  assign n6289 = n6284 & ~n6288 ;
  assign n6290 = x62 & ~n329 ;
  assign n6291 = n6290 ^ n5645 ^ 1'b0 ;
  assign n6292 = n6291 ^ n1101 ^ 1'b0 ;
  assign n6293 = ( ~n1720 & n2890 ) | ( ~n1720 & n6292 ) | ( n2890 & n6292 ) ;
  assign n6294 = ( x140 & n1001 ) | ( x140 & n1140 ) | ( n1001 & n1140 ) ;
  assign n6295 = ~n2577 & n6294 ;
  assign n6296 = n4942 & ~n6295 ;
  assign n6297 = n1206 & n6296 ;
  assign n6298 = n260 | n948 ;
  assign n6299 = ( n2360 & ~n4270 ) | ( n2360 & n6298 ) | ( ~n4270 & n6298 ) ;
  assign n6300 = ( ~n3796 & n4093 ) | ( ~n3796 & n5134 ) | ( n4093 & n5134 ) ;
  assign n6301 = ( x19 & ~n975 ) | ( x19 & n1837 ) | ( ~n975 & n1837 ) ;
  assign n6302 = n5544 ^ n444 ^ 1'b0 ;
  assign n6303 = n1344 & ~n6302 ;
  assign n6304 = n6301 & n6303 ;
  assign n6305 = ( ~n1032 & n2472 ) | ( ~n1032 & n6304 ) | ( n2472 & n6304 ) ;
  assign n6306 = n2045 ^ n1856 ^ n1426 ;
  assign n6307 = n1784 & ~n6306 ;
  assign n6308 = x85 & n2721 ;
  assign n6309 = n5242 & n6308 ;
  assign n6310 = n4218 ^ n2254 ^ 1'b0 ;
  assign n6311 = n3288 ^ n618 ^ 1'b0 ;
  assign n6312 = n2093 | n6311 ;
  assign n6313 = n4937 | n6312 ;
  assign n6314 = ~n3560 & n6313 ;
  assign n6315 = ~n6310 & n6314 ;
  assign n6316 = n411 | n638 ;
  assign n6317 = x143 | n6316 ;
  assign n6318 = ~n3673 & n6317 ;
  assign n6319 = n3317 ^ n2260 ^ 1'b0 ;
  assign n6320 = x80 & ~n2431 ;
  assign n6321 = ~n268 & n6320 ;
  assign n6322 = n2738 ^ n638 ^ 1'b0 ;
  assign n6323 = n6322 ^ n779 ^ 1'b0 ;
  assign n6324 = ~n3893 & n6323 ;
  assign n6325 = n2850 | n6324 ;
  assign n6326 = ( n953 & n4439 ) | ( n953 & ~n4892 ) | ( n4439 & ~n4892 ) ;
  assign n6327 = n4559 | n5363 ;
  assign n6328 = n5392 ^ n421 ^ 1'b0 ;
  assign n6329 = x111 & ~n6328 ;
  assign n6330 = ~n6175 & n6329 ;
  assign n6331 = n6330 ^ n2319 ^ 1'b0 ;
  assign n6332 = n752 & n4111 ;
  assign n6333 = n3929 ^ n1565 ^ 1'b0 ;
  assign n6334 = n5515 & n6333 ;
  assign n6335 = n6332 & n6334 ;
  assign n6336 = n903 | n3479 ;
  assign n6337 = n6336 ^ n3218 ^ 1'b0 ;
  assign n6338 = n3606 ^ n2013 ^ n694 ;
  assign n6339 = n4936 ^ n3415 ^ 1'b0 ;
  assign n6340 = n6339 ^ n1057 ^ 1'b0 ;
  assign n6341 = n417 & ~n4370 ;
  assign n6342 = n2614 ^ n510 ^ 1'b0 ;
  assign n6343 = n3044 ^ x157 ^ 1'b0 ;
  assign n6344 = n6342 & ~n6343 ;
  assign n6345 = n6252 & n6344 ;
  assign n6346 = n3420 ^ n1799 ^ n749 ;
  assign n6347 = n6346 ^ n1937 ^ 1'b0 ;
  assign n6348 = n2224 ^ n710 ^ 1'b0 ;
  assign n6349 = n3186 ^ n2029 ^ 1'b0 ;
  assign n6350 = ~n6348 & n6349 ;
  assign n6351 = n2534 ^ n2056 ^ 1'b0 ;
  assign n6352 = n1144 & n6351 ;
  assign n6353 = n4741 | n6352 ;
  assign n6354 = ( n2433 & n5237 ) | ( n2433 & ~n6042 ) | ( n5237 & ~n6042 ) ;
  assign n6355 = n466 | n5705 ;
  assign n6356 = ~n761 & n2534 ;
  assign n6357 = ~n1358 & n6356 ;
  assign n6358 = n1912 | n4109 ;
  assign n6359 = n2901 ^ n1733 ^ x158 ;
  assign n6360 = n6358 & n6359 ;
  assign n6361 = ~n6357 & n6360 ;
  assign n6362 = ~n2790 & n5996 ;
  assign n6363 = n6362 ^ x24 ^ 1'b0 ;
  assign n6364 = n2989 ^ n2514 ^ 1'b0 ;
  assign n6365 = n6364 ^ n3427 ^ 1'b0 ;
  assign n6366 = x195 & ~n6365 ;
  assign n6367 = n6366 ^ n3302 ^ 1'b0 ;
  assign n6368 = n5341 & n6367 ;
  assign n6369 = ~n6292 & n6368 ;
  assign n6370 = n5683 ^ n5422 ^ 1'b0 ;
  assign n6372 = n619 | n4543 ;
  assign n6373 = n6372 ^ n1766 ^ 1'b0 ;
  assign n6371 = n2798 & ~n2950 ;
  assign n6374 = n6373 ^ n6371 ^ 1'b0 ;
  assign n6375 = n6374 ^ n2883 ^ 1'b0 ;
  assign n6376 = n6370 & ~n6375 ;
  assign n6377 = ~n466 & n6376 ;
  assign n6378 = n6377 ^ n428 ^ 1'b0 ;
  assign n6380 = n1206 ^ x254 ^ 1'b0 ;
  assign n6381 = x101 & ~n6380 ;
  assign n6379 = n3620 & n4627 ;
  assign n6382 = n6381 ^ n6379 ^ 1'b0 ;
  assign n6383 = n1577 ^ n1030 ^ x34 ;
  assign n6384 = n3417 & n5265 ;
  assign n6385 = ~n6383 & n6384 ;
  assign n6386 = n6382 | n6385 ;
  assign n6388 = n5746 ^ n5463 ^ 1'b0 ;
  assign n6387 = ~n727 & n5082 ;
  assign n6389 = n6388 ^ n6387 ^ 1'b0 ;
  assign n6390 = n2335 ^ n1536 ^ 1'b0 ;
  assign n6391 = n3305 & n6390 ;
  assign n6392 = x192 & n6391 ;
  assign n6393 = ~n4347 & n6392 ;
  assign n6395 = n432 | n553 ;
  assign n6396 = ~n1936 & n6395 ;
  assign n6397 = n6396 ^ n1928 ^ 1'b0 ;
  assign n6394 = n4946 ^ n2966 ^ 1'b0 ;
  assign n6398 = n6397 ^ n6394 ^ n4256 ;
  assign n6399 = n6398 ^ n5980 ^ 1'b0 ;
  assign n6400 = ( x57 & n3114 ) | ( x57 & n4350 ) | ( n3114 & n4350 ) ;
  assign n6401 = n3499 & n6400 ;
  assign n6402 = ~n1997 & n6401 ;
  assign n6403 = n6216 ^ n6157 ^ 1'b0 ;
  assign n6404 = n6402 & ~n6403 ;
  assign n6405 = ( ~n3760 & n5883 ) | ( ~n3760 & n6404 ) | ( n5883 & n6404 ) ;
  assign n6406 = n1315 | n3379 ;
  assign n6407 = n2433 & ~n3674 ;
  assign n6408 = ~n3144 & n6407 ;
  assign n6409 = ( n1577 & n4754 ) | ( n1577 & n6408 ) | ( n4754 & n6408 ) ;
  assign n6410 = x193 | n3594 ;
  assign n6411 = n6410 ^ n4076 ^ 1'b0 ;
  assign n6412 = n5571 ^ n756 ^ 1'b0 ;
  assign n6414 = n1867 ^ n983 ^ 1'b0 ;
  assign n6413 = n2372 ^ x228 ^ 1'b0 ;
  assign n6415 = n6414 ^ n6413 ^ 1'b0 ;
  assign n6416 = n6415 ^ n3725 ^ 1'b0 ;
  assign n6417 = n5958 ^ x179 ^ 1'b0 ;
  assign n6418 = n5435 ^ n632 ^ 1'b0 ;
  assign n6419 = n2547 | n6418 ;
  assign n6420 = n2942 & n4898 ;
  assign n6421 = n4018 & n6420 ;
  assign n6422 = n1867 & ~n6421 ;
  assign n6423 = n6422 ^ n2294 ^ 1'b0 ;
  assign n6424 = x188 | n4200 ;
  assign n6425 = n6424 ^ n5094 ^ 1'b0 ;
  assign n6426 = n287 & ~n340 ;
  assign n6427 = n6426 ^ n3174 ^ 1'b0 ;
  assign n6428 = n6425 & ~n6427 ;
  assign n6429 = n6343 ^ n3659 ^ 1'b0 ;
  assign n6430 = n1016 | n1636 ;
  assign n6431 = x155 & n2529 ;
  assign n6432 = ( n3483 & ~n6304 ) | ( n3483 & n6431 ) | ( ~n6304 & n6431 ) ;
  assign n6433 = n6430 | n6432 ;
  assign n6434 = n6128 & ~n6327 ;
  assign n6435 = n1373 & ~n5848 ;
  assign n6436 = ~n2936 & n6435 ;
  assign n6437 = n4282 ^ n1630 ^ x188 ;
  assign n6438 = n3328 ^ n2708 ^ 1'b0 ;
  assign n6439 = n6437 | n6438 ;
  assign n6440 = n6439 ^ n4908 ^ 1'b0 ;
  assign n6441 = n5804 ^ n4109 ^ n3214 ;
  assign n6442 = n351 ^ n260 ^ 1'b0 ;
  assign n6443 = n6442 ^ n1929 ^ 1'b0 ;
  assign n6444 = n2308 ^ n409 ^ 1'b0 ;
  assign n6445 = n6443 & ~n6444 ;
  assign n6446 = ~n3958 & n6445 ;
  assign n6447 = n4918 ^ n1487 ^ n274 ;
  assign n6448 = n2198 ^ x63 ^ 1'b0 ;
  assign n6449 = n6448 ^ n4872 ^ 1'b0 ;
  assign n6450 = n6447 | n6449 ;
  assign n6451 = n2919 & ~n5284 ;
  assign n6452 = x96 & ~n1328 ;
  assign n6453 = n302 & n331 ;
  assign n6454 = ~n2144 & n6453 ;
  assign n6455 = n6452 & n6454 ;
  assign n6456 = n2801 | n5302 ;
  assign n6457 = n522 | n3230 ;
  assign n6458 = n6457 ^ n1471 ^ 1'b0 ;
  assign n6459 = n6458 ^ n5632 ^ 1'b0 ;
  assign n6460 = n6456 | n6459 ;
  assign n6461 = n6455 & ~n6460 ;
  assign n6462 = ~n6451 & n6461 ;
  assign n6463 = n1373 & ~n3795 ;
  assign n6464 = n6463 ^ n2666 ^ 1'b0 ;
  assign n6466 = n3023 ^ n2256 ^ 1'b0 ;
  assign n6465 = x22 & ~n2294 ;
  assign n6467 = n6466 ^ n6465 ^ 1'b0 ;
  assign n6468 = n4204 ^ n2082 ^ 1'b0 ;
  assign n6469 = x201 & ~n6468 ;
  assign n6470 = ~n3706 & n5309 ;
  assign n6471 = ~n6469 & n6470 ;
  assign n6472 = n1440 | n6188 ;
  assign n6473 = n6472 ^ n1190 ^ 1'b0 ;
  assign n6474 = n4069 ^ n1876 ^ n786 ;
  assign n6475 = n4271 & ~n6474 ;
  assign n6476 = n4489 ^ n2684 ^ 1'b0 ;
  assign n6477 = n3988 ^ n2948 ^ 1'b0 ;
  assign n6478 = n1120 & ~n6477 ;
  assign n6479 = ~n6476 & n6478 ;
  assign n6480 = n4786 ^ n455 ^ 1'b0 ;
  assign n6481 = n4737 | n6480 ;
  assign n6482 = n883 ^ x99 ^ 1'b0 ;
  assign n6483 = n1923 | n6482 ;
  assign n6484 = n2452 | n6483 ;
  assign n6485 = n6484 ^ n1506 ^ 1'b0 ;
  assign n6486 = ~n4767 & n6485 ;
  assign n6487 = n6486 ^ n2782 ^ 1'b0 ;
  assign n6488 = ~n1741 & n6487 ;
  assign n6489 = n6488 ^ n5683 ^ 1'b0 ;
  assign n6491 = x3 & ~n2321 ;
  assign n6492 = n6491 ^ n906 ^ 1'b0 ;
  assign n6490 = n2592 & n3221 ;
  assign n6493 = n6492 ^ n6490 ^ 1'b0 ;
  assign n6494 = n6493 ^ n3246 ^ 1'b0 ;
  assign n6495 = n1167 & n6494 ;
  assign n6496 = x243 ^ x6 ^ 1'b0 ;
  assign n6497 = n817 & n4473 ;
  assign n6498 = n3041 ^ n2122 ^ 1'b0 ;
  assign n6499 = ~n6497 & n6498 ;
  assign n6500 = n4561 | n5241 ;
  assign n6501 = x215 & ~n725 ;
  assign n6502 = n6501 ^ n6059 ^ 1'b0 ;
  assign n6503 = ( n1889 & n2670 ) | ( n1889 & ~n6502 ) | ( n2670 & ~n6502 ) ;
  assign n6504 = n6503 ^ x67 ^ 1'b0 ;
  assign n6505 = x140 & n4786 ;
  assign n6506 = n6505 ^ n4135 ^ 1'b0 ;
  assign n6507 = n2859 | n6506 ;
  assign n6508 = n6507 ^ n1450 ^ 1'b0 ;
  assign n6509 = n2590 & ~n6508 ;
  assign n6510 = ~n3750 & n6509 ;
  assign n6511 = n2426 ^ n274 ^ x48 ;
  assign n6512 = n6511 ^ n2106 ^ 1'b0 ;
  assign n6513 = n1654 | n5675 ;
  assign n6514 = n6513 ^ n2661 ^ 1'b0 ;
  assign n6515 = n2109 ^ n1495 ^ 1'b0 ;
  assign n6516 = n5274 | n6515 ;
  assign n6517 = n744 ^ n378 ^ 1'b0 ;
  assign n6518 = n2703 | n6517 ;
  assign n6519 = n3750 & ~n6518 ;
  assign n6520 = n6516 & n6519 ;
  assign n6521 = ( n266 & n4861 ) | ( n266 & n6520 ) | ( n4861 & n6520 ) ;
  assign n6522 = n3036 | n6521 ;
  assign n6523 = ~n819 & n4750 ;
  assign n6524 = n3969 & n6523 ;
  assign n6525 = n6359 & ~n6524 ;
  assign n6526 = ( ~n1210 & n3329 ) | ( ~n1210 & n5334 ) | ( n3329 & n5334 ) ;
  assign n6527 = n2304 ^ n2296 ^ 1'b0 ;
  assign n6534 = n2340 ^ n1089 ^ 1'b0 ;
  assign n6535 = n3425 | n6534 ;
  assign n6536 = n3491 | n6535 ;
  assign n6528 = ~n1791 & n2426 ;
  assign n6529 = ~n2918 & n6528 ;
  assign n6530 = n3911 | n6529 ;
  assign n6531 = n6530 ^ x115 ^ 1'b0 ;
  assign n6532 = ~n5033 & n6531 ;
  assign n6533 = n6532 ^ n2681 ^ 1'b0 ;
  assign n6537 = n6536 ^ n6533 ^ 1'b0 ;
  assign n6538 = ~n361 & n4236 ;
  assign n6539 = n6538 ^ n971 ^ 1'b0 ;
  assign n6540 = ~n2072 & n3383 ;
  assign n6541 = n6540 ^ n2951 ^ 1'b0 ;
  assign n6542 = x143 & ~n6541 ;
  assign n6544 = ~n4741 & n5931 ;
  assign n6545 = ~n2926 & n6544 ;
  assign n6543 = ~n1075 & n5800 ;
  assign n6546 = n6545 ^ n6543 ^ 1'b0 ;
  assign n6547 = n1600 & n6546 ;
  assign n6548 = x250 & n3139 ;
  assign n6549 = n1298 & n2125 ;
  assign n6550 = n2004 & ~n6549 ;
  assign n6551 = ( n705 & n2130 ) | ( n705 & ~n6550 ) | ( n2130 & ~n6550 ) ;
  assign n6552 = n6551 ^ n5771 ^ 1'b0 ;
  assign n6553 = ~n6548 & n6552 ;
  assign n6554 = n1432 | n2275 ;
  assign n6555 = ( x6 & ~x40 ) | ( x6 & n6554 ) | ( ~x40 & n6554 ) ;
  assign n6556 = n2516 & ~n5604 ;
  assign n6557 = n6556 ^ n3685 ^ 1'b0 ;
  assign n6558 = ~n4099 & n6557 ;
  assign n6559 = ~n2622 & n6558 ;
  assign n6560 = n5622 ^ n475 ^ 1'b0 ;
  assign n6561 = n1605 ^ n1070 ^ 1'b0 ;
  assign n6563 = ( n597 & n1069 ) | ( n597 & ~n1963 ) | ( n1069 & ~n1963 ) ;
  assign n6562 = n2367 | n2868 ;
  assign n6564 = n6563 ^ n6562 ^ 1'b0 ;
  assign n6565 = x120 | n6564 ;
  assign n6566 = ( n5848 & n6561 ) | ( n5848 & ~n6565 ) | ( n6561 & ~n6565 ) ;
  assign n6567 = n2165 ^ n2101 ^ n1575 ;
  assign n6568 = n2844 | n6567 ;
  assign n6569 = n1486 | n6568 ;
  assign n6570 = n1190 & n6569 ;
  assign n6571 = n6160 & n6570 ;
  assign n6572 = n365 | n3348 ;
  assign n6573 = x65 & ~n6572 ;
  assign n6574 = n3059 & n6573 ;
  assign n6575 = x206 & ~n3475 ;
  assign n6576 = n6575 ^ n2789 ^ 1'b0 ;
  assign n6577 = ~n3688 & n4787 ;
  assign n6578 = n5534 & n6577 ;
  assign n6579 = n6578 ^ n5201 ^ 1'b0 ;
  assign n6580 = n4356 & n6579 ;
  assign n6581 = n4584 ^ n4348 ^ 1'b0 ;
  assign n6582 = n2182 & ~n3225 ;
  assign n6583 = n5420 & n6582 ;
  assign n6584 = n4082 ^ n1662 ^ 1'b0 ;
  assign n6585 = n885 | n6584 ;
  assign n6586 = n634 ^ x246 ^ 1'b0 ;
  assign n6587 = ~n444 & n6586 ;
  assign n6588 = n2355 ^ x184 ^ 1'b0 ;
  assign n6589 = n6587 & n6588 ;
  assign n6590 = n6589 ^ n3000 ^ 1'b0 ;
  assign n6591 = n6585 & ~n6590 ;
  assign n6592 = n4038 ^ n686 ^ x164 ;
  assign n6593 = ~n3362 & n5465 ;
  assign n6594 = n2443 & ~n3749 ;
  assign n6595 = n6594 ^ n2881 ^ 1'b0 ;
  assign n6596 = n3099 & n6595 ;
  assign n6597 = ( ~n455 & n1295 ) | ( ~n455 & n6596 ) | ( n1295 & n6596 ) ;
  assign n6598 = n353 & ~n3393 ;
  assign n6599 = n6598 ^ x215 ^ 1'b0 ;
  assign n6600 = n2110 | n6182 ;
  assign n6601 = n5646 & n6600 ;
  assign n6602 = n6599 & n6601 ;
  assign n6603 = n5115 & ~n6602 ;
  assign n6604 = n1735 | n5093 ;
  assign n6605 = n4121 ^ n686 ^ 1'b0 ;
  assign n6606 = n3329 & ~n6193 ;
  assign n6607 = ~n1049 & n4725 ;
  assign n6608 = ( n1020 & n2002 ) | ( n1020 & ~n4672 ) | ( n2002 & ~n4672 ) ;
  assign n6609 = ~n384 & n739 ;
  assign n6610 = n2477 ^ n1215 ^ 1'b0 ;
  assign n6611 = ~n2249 & n6610 ;
  assign n6612 = ~n3183 & n6611 ;
  assign n6613 = n6609 | n6612 ;
  assign n6614 = n6608 & n6613 ;
  assign n6615 = n2492 & n6614 ;
  assign n6616 = n4480 | n4826 ;
  assign n6617 = n2428 & n6616 ;
  assign n6618 = ~n6580 & n6617 ;
  assign n6619 = ( ~n1393 & n4773 ) | ( ~n1393 & n6331 ) | ( n4773 & n6331 ) ;
  assign n6620 = n564 | n1505 ;
  assign n6621 = n6620 ^ n6159 ^ 1'b0 ;
  assign n6622 = n550 ^ n293 ^ 1'b0 ;
  assign n6623 = n3901 | n6622 ;
  assign n6624 = n420 & ~n6623 ;
  assign n6625 = n3427 ^ x17 ^ 1'b0 ;
  assign n6626 = n6624 & ~n6625 ;
  assign n6627 = n1672 & ~n2415 ;
  assign n6628 = n3877 & ~n6627 ;
  assign n6629 = n1728 | n6628 ;
  assign n6633 = n1844 | n3467 ;
  assign n6630 = n680 & ~n5390 ;
  assign n6631 = n6630 ^ n2466 ^ 1'b0 ;
  assign n6632 = n1190 & n6631 ;
  assign n6634 = n6633 ^ n6632 ^ 1'b0 ;
  assign n6635 = n6634 ^ n2188 ^ 1'b0 ;
  assign n6636 = ~n6629 & n6635 ;
  assign n6639 = ( n3319 & ~n3537 ) | ( n3319 & n5036 ) | ( ~n3537 & n5036 ) ;
  assign n6637 = n3425 & n4163 ;
  assign n6638 = n6637 ^ n5059 ^ 1'b0 ;
  assign n6640 = n6639 ^ n6638 ^ 1'b0 ;
  assign n6641 = n2523 | n4737 ;
  assign n6642 = n6641 ^ x72 ^ 1'b0 ;
  assign n6643 = x244 & n6642 ;
  assign n6644 = ~n991 & n6643 ;
  assign n6645 = n6644 ^ n2162 ^ 1'b0 ;
  assign n6646 = n501 & n6645 ;
  assign n6647 = n1252 & n6646 ;
  assign n6648 = n6647 ^ n3119 ^ 1'b0 ;
  assign n6649 = n1602 & n2514 ;
  assign n6650 = n3663 ^ n2039 ^ 1'b0 ;
  assign n6651 = ~n1192 & n6650 ;
  assign n6652 = ~n6649 & n6651 ;
  assign n6653 = n5961 ^ n3496 ^ 1'b0 ;
  assign n6654 = n1389 & ~n4598 ;
  assign n6655 = n5893 ^ n2297 ^ n970 ;
  assign n6656 = n547 | n6655 ;
  assign n6657 = n4357 | n6656 ;
  assign n6658 = n3802 ^ n574 ^ 1'b0 ;
  assign n6659 = n434 & n6658 ;
  assign n6660 = n3686 & n6659 ;
  assign n6661 = n2443 & n5714 ;
  assign n6662 = n5120 | n6661 ;
  assign n6663 = ~n1489 & n2466 ;
  assign n6664 = n4204 & n6663 ;
  assign n6665 = n1092 & ~n6664 ;
  assign n6666 = n5705 & n6665 ;
  assign n6667 = n406 & n4411 ;
  assign n6668 = ~n4801 & n6667 ;
  assign n6669 = n258 | n1499 ;
  assign n6670 = n1023 | n6669 ;
  assign n6671 = n4846 ^ n3929 ^ 1'b0 ;
  assign n6672 = ( x164 & ~n1195 ) | ( x164 & n6671 ) | ( ~n1195 & n6671 ) ;
  assign n6673 = ~x178 & n6204 ;
  assign n6674 = n6673 ^ n2082 ^ 1'b0 ;
  assign n6675 = ~n3517 & n5111 ;
  assign n6676 = n6675 ^ n1716 ^ 1'b0 ;
  assign n6677 = n2853 & n5715 ;
  assign n6678 = ( x225 & n867 ) | ( x225 & n5496 ) | ( n867 & n5496 ) ;
  assign n6679 = n6678 ^ n6339 ^ 1'b0 ;
  assign n6683 = n260 & n1964 ;
  assign n6684 = ~x123 & n6683 ;
  assign n6685 = n4666 ^ n1322 ^ 1'b0 ;
  assign n6686 = ~n780 & n6685 ;
  assign n6687 = n6684 & n6686 ;
  assign n6680 = n2294 ^ x230 ^ x16 ;
  assign n6681 = n6680 ^ n4943 ^ n2402 ;
  assign n6682 = ( n2272 & ~n3075 ) | ( n2272 & n6681 ) | ( ~n3075 & n6681 ) ;
  assign n6688 = n6687 ^ n6682 ^ 1'b0 ;
  assign n6689 = n4393 ^ n2210 ^ 1'b0 ;
  assign n6690 = n500 | n6689 ;
  assign n6691 = x87 & ~n2963 ;
  assign n6692 = n6691 ^ n1633 ^ 1'b0 ;
  assign n6693 = n6692 ^ n4784 ^ n260 ;
  assign n6694 = n2735 & n6693 ;
  assign n6695 = ( n1379 & n1513 ) | ( n1379 & n3676 ) | ( n1513 & n3676 ) ;
  assign n6696 = n1062 | n6695 ;
  assign n6697 = n3207 & n6696 ;
  assign n6698 = ~n883 & n6697 ;
  assign n6699 = ~n397 & n6698 ;
  assign n6700 = n2724 ^ n997 ^ 1'b0 ;
  assign n6701 = n6700 ^ n3684 ^ 1'b0 ;
  assign n6702 = n3179 ^ n2335 ^ 1'b0 ;
  assign n6703 = ~n5688 & n6702 ;
  assign n6704 = x243 & n2159 ;
  assign n6705 = ~n6703 & n6704 ;
  assign n6706 = n4874 | n5654 ;
  assign n6707 = n1006 | n6706 ;
  assign n6708 = n6473 ^ n2978 ^ 1'b0 ;
  assign n6709 = n6707 & n6708 ;
  assign n6710 = n617 & n2442 ;
  assign n6711 = n6710 ^ x243 ^ 1'b0 ;
  assign n6712 = ~n1636 & n6711 ;
  assign n6713 = n5763 & ~n6712 ;
  assign n6714 = n1025 & ~n6713 ;
  assign n6715 = n4543 ^ n3401 ^ 1'b0 ;
  assign n6716 = n1763 & n6715 ;
  assign n6717 = n4984 & n6716 ;
  assign n6718 = n6591 & n6717 ;
  assign n6719 = n2077 & ~n4255 ;
  assign n6721 = n2743 & ~n3119 ;
  assign n6720 = n946 & n2045 ;
  assign n6722 = n6721 ^ n6720 ^ 1'b0 ;
  assign n6723 = x115 & ~x119 ;
  assign n6724 = n3904 ^ n2065 ^ 1'b0 ;
  assign n6725 = ~n1593 & n6724 ;
  assign n6726 = n2371 ^ x101 ^ 1'b0 ;
  assign n6727 = n4508 & ~n6726 ;
  assign n6728 = n1272 | n2302 ;
  assign n6729 = n6727 | n6728 ;
  assign n6730 = n6725 | n6729 ;
  assign n6731 = n790 | n2239 ;
  assign n6733 = ( n1149 & n1335 ) | ( n1149 & n1958 ) | ( n1335 & n1958 ) ;
  assign n6734 = n5525 & n6733 ;
  assign n6732 = n2091 & ~n5756 ;
  assign n6735 = n6734 ^ n6732 ^ 1'b0 ;
  assign n6736 = n2984 ^ n2312 ^ 1'b0 ;
  assign n6737 = n2341 & n6736 ;
  assign n6738 = n399 | n1244 ;
  assign n6739 = n1278 | n6738 ;
  assign n6740 = ~n5028 & n6739 ;
  assign n6741 = ~n6737 & n6740 ;
  assign n6743 = ~n603 & n2534 ;
  assign n6744 = n1905 & n6743 ;
  assign n6745 = n2402 | n6744 ;
  assign n6742 = ~x166 & n860 ;
  assign n6746 = n6745 ^ n6742 ^ n2877 ;
  assign n6747 = n1928 | n5798 ;
  assign n6748 = n6746 & ~n6747 ;
  assign n6749 = n2609 & ~n2653 ;
  assign n6750 = n6748 & ~n6749 ;
  assign n6751 = n2702 ^ n1964 ^ 1'b0 ;
  assign n6752 = n4803 & n5462 ;
  assign n6753 = n3749 & n6752 ;
  assign n6754 = x69 & ~n3157 ;
  assign n6755 = ~n1295 & n6754 ;
  assign n6756 = ( x212 & ~n865 ) | ( x212 & n1132 ) | ( ~n865 & n1132 ) ;
  assign n6757 = ( ~n1826 & n2924 ) | ( ~n1826 & n3814 ) | ( n2924 & n3814 ) ;
  assign n6758 = n6757 ^ n4568 ^ 1'b0 ;
  assign n6759 = n6756 & ~n6758 ;
  assign n6760 = n5189 ^ n1157 ^ 1'b0 ;
  assign n6761 = n5221 | n6760 ;
  assign n6762 = ~n4372 & n5551 ;
  assign n6763 = n6761 & n6762 ;
  assign n6764 = n2852 ^ n328 ^ 1'b0 ;
  assign n6765 = n385 & n6764 ;
  assign n6766 = n3665 & ~n5821 ;
  assign n6767 = ~n6765 & n6766 ;
  assign n6768 = n5948 | n6767 ;
  assign n6769 = n6768 ^ x129 ^ 1'b0 ;
  assign n6770 = n2089 ^ n1900 ^ n1805 ;
  assign n6771 = n2756 & n6770 ;
  assign n6772 = n6771 ^ n5635 ^ 1'b0 ;
  assign n6773 = n1725 | n3226 ;
  assign n6774 = ( n1343 & ~n1590 ) | ( n1343 & n2202 ) | ( ~n1590 & n2202 ) ;
  assign n6775 = n6774 ^ n5775 ^ 1'b0 ;
  assign n6776 = n6773 & ~n6775 ;
  assign n6777 = ~n2265 & n6695 ;
  assign n6778 = n6471 & n6777 ;
  assign n6779 = n1570 | n4503 ;
  assign n6780 = n6779 ^ n281 ^ 1'b0 ;
  assign n6781 = n1294 | n6780 ;
  assign n6782 = ( x6 & ~n1830 ) | ( x6 & n5234 ) | ( ~n1830 & n5234 ) ;
  assign n6783 = n6782 ^ n4462 ^ 1'b0 ;
  assign n6784 = n1775 | n2995 ;
  assign n6785 = n6784 ^ n5679 ^ 1'b0 ;
  assign n6786 = n6785 ^ n4136 ^ 1'b0 ;
  assign n6787 = ~n1586 & n6701 ;
  assign n6788 = ~n6786 & n6787 ;
  assign n6789 = n4725 & ~n5856 ;
  assign n6790 = n2001 | n4333 ;
  assign n6791 = n6790 ^ x161 ^ 1'b0 ;
  assign n6792 = ~n1867 & n6791 ;
  assign n6793 = ~n2936 & n6792 ;
  assign n6794 = n6169 ^ n4656 ^ 1'b0 ;
  assign n6795 = n3046 ^ n473 ^ 1'b0 ;
  assign n6796 = n6794 & ~n6795 ;
  assign n6797 = n6796 ^ n634 ^ x227 ;
  assign n6798 = n871 ^ n571 ^ 1'b0 ;
  assign n6799 = n2264 | n6798 ;
  assign n6800 = n1762 & ~n6799 ;
  assign n6801 = n1774 & ~n3650 ;
  assign n6802 = n6801 ^ n2268 ^ 1'b0 ;
  assign n6803 = n6083 & ~n6802 ;
  assign n6804 = x166 & ~n6803 ;
  assign n6805 = n4266 & n6804 ;
  assign n6806 = n4249 & ~n6805 ;
  assign n6807 = n1376 & n6806 ;
  assign n6808 = ~x27 & n1154 ;
  assign n6809 = n6808 ^ n5700 ^ n4768 ;
  assign n6810 = n839 | n1620 ;
  assign n6811 = n6810 ^ n3378 ^ 1'b0 ;
  assign n6812 = n6811 ^ n3679 ^ 1'b0 ;
  assign n6813 = n285 ^ n264 ^ 1'b0 ;
  assign n6814 = x55 & n6813 ;
  assign n6815 = n6814 ^ n1780 ^ 1'b0 ;
  assign n6816 = n6815 ^ n4580 ^ 1'b0 ;
  assign n6817 = n6816 ^ n1014 ^ 1'b0 ;
  assign n6818 = ( ~n729 & n5277 ) | ( ~n729 & n6817 ) | ( n5277 & n6817 ) ;
  assign n6819 = ( ~x20 & n875 ) | ( ~x20 & n2925 ) | ( n875 & n2925 ) ;
  assign n6820 = ~n1906 & n6819 ;
  assign n6821 = ~n2458 & n3075 ;
  assign n6822 = n1514 ^ n378 ^ 1'b0 ;
  assign n6823 = n2511 & n6822 ;
  assign n6824 = n6823 ^ n4426 ^ 1'b0 ;
  assign n6825 = n3359 | n6824 ;
  assign n6826 = n6825 ^ n3633 ^ 1'b0 ;
  assign n6827 = n6826 ^ n4338 ^ 1'b0 ;
  assign n6828 = ( x160 & n333 ) | ( x160 & n1203 ) | ( n333 & n1203 ) ;
  assign n6829 = n830 | n6828 ;
  assign n6830 = n6827 & ~n6829 ;
  assign n6831 = ( ~n668 & n5992 ) | ( ~n668 & n6830 ) | ( n5992 & n6830 ) ;
  assign n6832 = n2133 & n4300 ;
  assign n6833 = n6832 ^ n1553 ^ 1'b0 ;
  assign n6837 = n1161 ^ n765 ^ 1'b0 ;
  assign n6838 = n1195 & ~n6837 ;
  assign n6835 = n1775 ^ n1458 ^ 1'b0 ;
  assign n6834 = ~n2785 & n3661 ;
  assign n6836 = n6835 ^ n6834 ^ n3982 ;
  assign n6839 = n6838 ^ n6836 ^ 1'b0 ;
  assign n6840 = n6347 | n6839 ;
  assign n6841 = ~n1489 & n2401 ;
  assign n6842 = n6841 ^ n5523 ^ 1'b0 ;
  assign n6843 = ~n1875 & n6842 ;
  assign n6844 = n6843 ^ n5772 ^ 1'b0 ;
  assign n6845 = n394 & ~n922 ;
  assign n6846 = n6845 ^ n3908 ^ 1'b0 ;
  assign n6847 = ~n761 & n6846 ;
  assign n6848 = n3725 ^ x148 ^ 1'b0 ;
  assign n6849 = n5294 & n6848 ;
  assign n6850 = n6847 & ~n6849 ;
  assign n6851 = n718 ^ x212 ^ 1'b0 ;
  assign n6852 = n5277 & ~n6851 ;
  assign n6853 = n3539 & n6852 ;
  assign n6854 = n4114 ^ n1762 ^ 1'b0 ;
  assign n6855 = n6744 ^ n2482 ^ 1'b0 ;
  assign n6856 = n4348 | n6855 ;
  assign n6857 = n6856 ^ n4968 ^ 1'b0 ;
  assign n6858 = n6857 ^ n2768 ^ 1'b0 ;
  assign n6859 = x89 | n6858 ;
  assign n6860 = ~n1215 & n6400 ;
  assign n6861 = ~n2420 & n6860 ;
  assign n6862 = n6220 ^ n2015 ^ 1'b0 ;
  assign n6863 = x120 & n990 ;
  assign n6864 = n6863 ^ n2276 ^ 1'b0 ;
  assign n6865 = n4894 & ~n6864 ;
  assign n6866 = n1204 ^ n351 ^ 1'b0 ;
  assign n6867 = n6866 ^ n1701 ^ 1'b0 ;
  assign n6868 = n2122 | n6867 ;
  assign n6871 = n994 | n1712 ;
  assign n6872 = n3279 & ~n6871 ;
  assign n6873 = ( n2670 & ~n4657 ) | ( n2670 & n6872 ) | ( ~n4657 & n6872 ) ;
  assign n6869 = n3837 ^ n1116 ^ 1'b0 ;
  assign n6870 = x108 & n6869 ;
  assign n6874 = n6873 ^ n6870 ^ 1'b0 ;
  assign n6875 = n2130 ^ n1552 ^ 1'b0 ;
  assign n6876 = x236 & n1659 ;
  assign n6877 = n6876 ^ n977 ^ 1'b0 ;
  assign n6878 = ~n3413 & n6877 ;
  assign n6879 = n6554 & n6878 ;
  assign n6880 = n3616 ^ x176 ^ 1'b0 ;
  assign n6881 = n6880 ^ x128 ^ 1'b0 ;
  assign n6885 = n668 | n1579 ;
  assign n6886 = n1238 | n6885 ;
  assign n6887 = ( ~n567 & n5618 ) | ( ~n567 & n6886 ) | ( n5618 & n6886 ) ;
  assign n6882 = n5127 ^ n1473 ^ 1'b0 ;
  assign n6883 = n671 & n6882 ;
  assign n6884 = ~n433 & n6883 ;
  assign n6888 = n6887 ^ n6884 ^ n6101 ;
  assign n6889 = n6888 ^ n1073 ^ 1'b0 ;
  assign n6890 = n5917 ^ n4149 ^ 1'b0 ;
  assign n6891 = ~n1368 & n6890 ;
  assign n6892 = n2105 | n4924 ;
  assign n6893 = n6892 ^ n2567 ^ 1'b0 ;
  assign n6894 = n4038 ^ n335 ^ 1'b0 ;
  assign n6895 = n2306 | n6894 ;
  assign n6896 = n415 & ~n6895 ;
  assign n6897 = ( n2101 & ~n2122 ) | ( n2101 & n4232 ) | ( ~n2122 & n4232 ) ;
  assign n6898 = x190 & n4359 ;
  assign n6899 = ~n3283 & n6898 ;
  assign n6900 = n6897 & n6899 ;
  assign n6901 = n5004 ^ n1238 ^ 1'b0 ;
  assign n6902 = n5771 | n6901 ;
  assign n6903 = n6781 ^ n1353 ^ 1'b0 ;
  assign n6906 = x250 & ~n1032 ;
  assign n6904 = n1261 | n2120 ;
  assign n6905 = n867 & ~n6904 ;
  assign n6907 = n6906 ^ n6905 ^ n5928 ;
  assign n6908 = n2782 ^ n809 ^ 1'b0 ;
  assign n6909 = n671 ^ x214 ^ 1'b0 ;
  assign n6910 = n1311 & n6909 ;
  assign n6911 = ~n2491 & n6910 ;
  assign n6912 = n6911 ^ n2433 ^ 1'b0 ;
  assign n6913 = n5726 ^ n5180 ^ 1'b0 ;
  assign n6914 = n6912 & ~n6913 ;
  assign n6915 = n3296 & ~n5492 ;
  assign n6916 = n6915 ^ n1763 ^ 1'b0 ;
  assign n6917 = n3676 ^ n3242 ^ 1'b0 ;
  assign n6918 = ~n2013 & n6917 ;
  assign n6919 = n5116 & n6918 ;
  assign n6920 = n2711 | n5973 ;
  assign n6921 = n5414 & n6920 ;
  assign n6922 = n723 | n6921 ;
  assign n6923 = n274 | n6922 ;
  assign n6924 = n6923 ^ n3287 ^ 1'b0 ;
  assign n6925 = n5898 & n6924 ;
  assign n6928 = n1570 ^ n679 ^ 1'b0 ;
  assign n6926 = n5410 & ~n5775 ;
  assign n6927 = n4988 & n6926 ;
  assign n6929 = n6928 ^ n6927 ^ 1'b0 ;
  assign n6930 = ~n1586 & n6929 ;
  assign n6931 = n6119 ^ n1195 ^ n684 ;
  assign n6932 = n6583 & ~n6931 ;
  assign n6933 = ~n2779 & n6932 ;
  assign n6934 = x159 & ~n302 ;
  assign n6935 = n3119 & ~n6934 ;
  assign n6936 = ~n1048 & n2514 ;
  assign n6937 = n6936 ^ n1795 ^ 1'b0 ;
  assign n6938 = n4357 ^ n2819 ^ 1'b0 ;
  assign n6939 = ~n6937 & n6938 ;
  assign n6940 = n4703 ^ n349 ^ 1'b0 ;
  assign n6941 = n6939 & n6940 ;
  assign n6942 = x226 & ~n473 ;
  assign n6943 = ~n5061 & n6942 ;
  assign n6944 = n490 | n6943 ;
  assign n6945 = n6944 ^ n1817 ^ 1'b0 ;
  assign n6946 = n1417 & ~n1447 ;
  assign n6947 = n2063 & n6946 ;
  assign n6948 = n1349 | n6947 ;
  assign n6949 = n6948 ^ n4543 ^ 1'b0 ;
  assign n6950 = n6949 ^ n839 ^ 1'b0 ;
  assign n6951 = n6945 & n6950 ;
  assign n6952 = x241 & n2002 ;
  assign n6953 = n6952 ^ n417 ^ 1'b0 ;
  assign n6954 = n911 & n6953 ;
  assign n6955 = n6954 ^ n2463 ^ 1'b0 ;
  assign n6956 = ~n1057 & n6955 ;
  assign n6957 = ( n697 & n5496 ) | ( n697 & ~n6077 ) | ( n5496 & ~n6077 ) ;
  assign n6958 = n5300 & ~n6957 ;
  assign n6959 = n6958 ^ n2096 ^ 1'b0 ;
  assign n6960 = n6959 ^ n3156 ^ 1'b0 ;
  assign n6961 = n4759 ^ n860 ^ 1'b0 ;
  assign n6962 = n5025 | n6961 ;
  assign n6963 = n6962 ^ n1558 ^ 1'b0 ;
  assign n6964 = n6963 ^ n471 ^ 1'b0 ;
  assign n6965 = x34 & ~n4146 ;
  assign n6966 = n2034 | n2341 ;
  assign n6967 = n6966 ^ n2710 ^ 1'b0 ;
  assign n6968 = ~n2711 & n6967 ;
  assign n6969 = n6968 ^ n3560 ^ 1'b0 ;
  assign n6970 = n4219 | n6969 ;
  assign n6971 = n968 & ~n6970 ;
  assign n6972 = x220 | n6741 ;
  assign n6973 = n2803 | n3038 ;
  assign n6974 = n6973 ^ n5878 ^ 1'b0 ;
  assign n6975 = ~n1933 & n3568 ;
  assign n6976 = x180 & n6975 ;
  assign n6977 = ~n3911 & n6454 ;
  assign n6978 = ~n6383 & n6977 ;
  assign n6981 = ~x72 & n781 ;
  assign n6979 = n1517 & n4994 ;
  assign n6980 = ~n479 & n6979 ;
  assign n6982 = n6981 ^ n6980 ^ 1'b0 ;
  assign n6983 = n2904 ^ n983 ^ 1'b0 ;
  assign n6984 = n3933 ^ n1807 ^ 1'b0 ;
  assign n6985 = n3670 | n6984 ;
  assign n6986 = ( n938 & ~n6840 ) | ( n938 & n6985 ) | ( ~n6840 & n6985 ) ;
  assign n6987 = n6703 ^ n1468 ^ n382 ;
  assign n6988 = n6987 ^ n5825 ^ 1'b0 ;
  assign n6989 = n5365 & ~n6988 ;
  assign n6990 = ~n2778 & n4543 ;
  assign n6991 = x201 | n2045 ;
  assign n6992 = n4491 & n6991 ;
  assign n6993 = n3235 ^ n325 ^ 1'b0 ;
  assign n6994 = n5459 & n6993 ;
  assign n6995 = n569 & n575 ;
  assign n6996 = n5084 & n6995 ;
  assign n6997 = n6996 ^ n5264 ^ 1'b0 ;
  assign n6998 = n6994 & ~n6997 ;
  assign n6999 = n3772 & ~n3844 ;
  assign n7000 = n5912 ^ n1020 ^ 1'b0 ;
  assign n7001 = ~n2008 & n4832 ;
  assign n7002 = n871 & n7001 ;
  assign n7003 = n810 ^ n289 ^ 1'b0 ;
  assign n7004 = n2312 & ~n7003 ;
  assign n7005 = ~n877 & n7004 ;
  assign n7006 = n5986 ^ n4520 ^ n3196 ;
  assign n7010 = n5915 ^ n3342 ^ 1'b0 ;
  assign n7011 = n954 & n7010 ;
  assign n7012 = n1481 & n7011 ;
  assign n7013 = n7012 ^ n1731 ^ 1'b0 ;
  assign n7014 = n4689 ^ x160 ^ 1'b0 ;
  assign n7015 = n7013 & n7014 ;
  assign n7016 = n1197 | n7015 ;
  assign n7007 = n5742 ^ n4027 ^ 1'b0 ;
  assign n7008 = n640 | n7007 ;
  assign n7009 = n5320 & ~n7008 ;
  assign n7017 = n7016 ^ n7009 ^ 1'b0 ;
  assign n7018 = n668 & n7017 ;
  assign n7019 = n3302 ^ n697 ^ 1'b0 ;
  assign n7020 = n267 | n2609 ;
  assign n7021 = x34 & ~n365 ;
  assign n7022 = ~n4787 & n7021 ;
  assign n7023 = n2922 | n7022 ;
  assign n7024 = n6225 & ~n7023 ;
  assign n7025 = n2011 & n7024 ;
  assign n7026 = n1215 & ~n3114 ;
  assign n7027 = n2174 & n7026 ;
  assign n7028 = ~x131 & n1573 ;
  assign n7029 = ~n2696 & n7028 ;
  assign n7030 = n5634 ^ n3682 ^ 1'b0 ;
  assign n7031 = n1965 & n7030 ;
  assign n7032 = ~n764 & n7031 ;
  assign n7034 = n436 & n2076 ;
  assign n7035 = ~n968 & n7034 ;
  assign n7033 = n4327 | n5342 ;
  assign n7036 = n7035 ^ n7033 ^ 1'b0 ;
  assign n7037 = n1525 | n7036 ;
  assign n7038 = n6442 | n7037 ;
  assign n7039 = n921 & n2677 ;
  assign n7040 = ~n826 & n7039 ;
  assign n7041 = n1404 & n7040 ;
  assign n7042 = n2771 ^ n483 ^ 1'b0 ;
  assign n7043 = n4543 ^ n4384 ^ 1'b0 ;
  assign n7044 = n7043 ^ n3106 ^ 1'b0 ;
  assign n7045 = ~n7042 & n7044 ;
  assign n7046 = n2684 ^ n1365 ^ 1'b0 ;
  assign n7047 = n1125 & ~n6639 ;
  assign n7048 = n7047 ^ n5707 ^ 1'b0 ;
  assign n7049 = n6672 ^ x141 ^ 1'b0 ;
  assign n7050 = n4528 & n7049 ;
  assign n7051 = n359 & ~n3440 ;
  assign n7052 = n1636 | n3739 ;
  assign n7053 = n4036 | n7052 ;
  assign n7054 = ~n1283 & n2649 ;
  assign n7055 = ~n462 & n7054 ;
  assign n7056 = n1630 & n7055 ;
  assign n7057 = ( ~n2615 & n7053 ) | ( ~n2615 & n7056 ) | ( n7053 & n7056 ) ;
  assign n7058 = n4919 ^ n1500 ^ 1'b0 ;
  assign n7059 = n7058 ^ n6695 ^ 1'b0 ;
  assign n7060 = n4708 ^ x248 ^ 1'b0 ;
  assign n7061 = n1219 & n7060 ;
  assign n7062 = x26 & n7061 ;
  assign n7063 = ~n7059 & n7062 ;
  assign n7064 = n4896 ^ n4745 ^ 1'b0 ;
  assign n7065 = n2112 | n7064 ;
  assign n7066 = n5500 & ~n7065 ;
  assign n7067 = n5273 ^ n2948 ^ n400 ;
  assign n7069 = ~n946 & n1254 ;
  assign n7070 = n2436 ^ x161 ^ 1'b0 ;
  assign n7071 = n7069 & n7070 ;
  assign n7068 = ~n2410 & n2903 ;
  assign n7072 = n7071 ^ n7068 ^ 1'b0 ;
  assign n7073 = n4593 & ~n7072 ;
  assign n7074 = n425 & ~n1846 ;
  assign n7075 = ~n2055 & n7074 ;
  assign n7076 = x208 & ~n1051 ;
  assign n7077 = ~n1931 & n7076 ;
  assign n7078 = n6798 & ~n7077 ;
  assign n7079 = n1716 ^ n838 ^ 1'b0 ;
  assign n7080 = n7079 ^ n5197 ^ 1'b0 ;
  assign n7081 = n2102 & ~n7080 ;
  assign n7082 = n7081 ^ n5402 ^ 1'b0 ;
  assign n7083 = n937 & n7082 ;
  assign n7084 = n7083 ^ n1120 ^ n625 ;
  assign n7085 = ~n863 & n903 ;
  assign n7086 = n7085 ^ n552 ^ 1'b0 ;
  assign n7087 = n567 & n935 ;
  assign n7088 = n4292 | n4856 ;
  assign n7089 = n7088 ^ n6410 ^ 1'b0 ;
  assign n7090 = n430 | n3440 ;
  assign n7091 = n1778 & ~n4008 ;
  assign n7092 = n7091 ^ n3521 ^ 1'b0 ;
  assign n7093 = n5756 & n7092 ;
  assign n7094 = n1193 | n5168 ;
  assign n7095 = x136 & x155 ;
  assign n7096 = n7095 ^ n4394 ^ 1'b0 ;
  assign n7097 = ~n3616 & n4708 ;
  assign n7098 = n2322 ^ n938 ^ 1'b0 ;
  assign n7099 = ~n3461 & n7098 ;
  assign n7100 = n7099 ^ n6222 ^ 1'b0 ;
  assign n7101 = n7097 & n7100 ;
  assign n7102 = ( n615 & ~n1739 ) | ( n615 & n6866 ) | ( ~n1739 & n6866 ) ;
  assign n7103 = n7102 ^ n2670 ^ x225 ;
  assign n7104 = ~n2975 & n7103 ;
  assign n7105 = n2774 ^ n1471 ^ 1'b0 ;
  assign n7106 = n7058 ^ n4260 ^ 1'b0 ;
  assign n7107 = ~n4288 & n7106 ;
  assign n7108 = n3961 ^ n3240 ^ 1'b0 ;
  assign n7109 = ~n2646 & n7108 ;
  assign n7110 = n7109 ^ n6211 ^ 1'b0 ;
  assign n7111 = ~n2550 & n5418 ;
  assign n7112 = ( ~n711 & n946 ) | ( ~n711 & n1770 ) | ( n946 & n1770 ) ;
  assign n7113 = n7111 | n7112 ;
  assign n7114 = x4 & n3645 ;
  assign n7115 = n7114 ^ n5752 ^ 1'b0 ;
  assign n7116 = n2870 & n7115 ;
  assign n7117 = n7116 ^ n1178 ^ 1'b0 ;
  assign n7118 = ( n638 & n708 ) | ( n638 & n4049 ) | ( n708 & n4049 ) ;
  assign n7119 = n7118 ^ n4792 ^ 1'b0 ;
  assign n7120 = ( n2030 & ~n4128 ) | ( n2030 & n7119 ) | ( ~n4128 & n7119 ) ;
  assign n7121 = n7120 ^ n2577 ^ 1'b0 ;
  assign n7122 = n4102 & n7121 ;
  assign n7123 = n2542 ^ n710 ^ 1'b0 ;
  assign n7124 = ~x0 & n4637 ;
  assign n7125 = n2176 | n7124 ;
  assign n7126 = n5122 & ~n7125 ;
  assign n7127 = n7126 ^ n5643 ^ 1'b0 ;
  assign n7128 = ~n7123 & n7127 ;
  assign n7129 = n618 | n1579 ;
  assign n7130 = n7129 ^ n1906 ^ 1'b0 ;
  assign n7131 = n5047 & ~n7130 ;
  assign n7132 = ~n7128 & n7131 ;
  assign n7133 = n4640 & ~n7132 ;
  assign n7134 = ~n6857 & n7133 ;
  assign n7135 = n3498 ^ n3052 ^ 1'b0 ;
  assign n7136 = n2472 | n5481 ;
  assign n7137 = n7135 | n7136 ;
  assign n7138 = ( n264 & ~n1017 ) | ( n264 & n2549 ) | ( ~n1017 & n2549 ) ;
  assign n7139 = n3973 ^ n1705 ^ 1'b0 ;
  assign n7140 = ~n7138 & n7139 ;
  assign n7141 = n911 & n1032 ;
  assign n7142 = n6780 ^ n1613 ^ 1'b0 ;
  assign n7143 = n7141 & n7142 ;
  assign n7147 = n2772 & n4640 ;
  assign n7144 = ~n1049 & n1316 ;
  assign n7145 = ~x160 & n7144 ;
  assign n7146 = n2866 & ~n7145 ;
  assign n7148 = n7147 ^ n7146 ^ 1'b0 ;
  assign n7149 = n2778 ^ n1763 ^ 1'b0 ;
  assign n7150 = n6725 & ~n7149 ;
  assign n7151 = n6621 & n6716 ;
  assign n7152 = n7151 ^ n733 ^ 1'b0 ;
  assign n7153 = n451 | n919 ;
  assign n7154 = n1213 | n7153 ;
  assign n7155 = n2663 | n4292 ;
  assign n7156 = n7155 ^ n2311 ^ 1'b0 ;
  assign n7157 = n1453 ^ n761 ^ 1'b0 ;
  assign n7158 = n1641 & ~n3894 ;
  assign n7159 = n1387 & n3291 ;
  assign n7160 = n680 & ~n7159 ;
  assign n7161 = ~n1219 & n2468 ;
  assign n7162 = n6442 ^ n5007 ^ n1632 ;
  assign n7163 = n2672 ^ n1397 ^ 1'b0 ;
  assign n7164 = ~n4491 & n7163 ;
  assign n7165 = ( n4185 & n7162 ) | ( n4185 & n7164 ) | ( n7162 & n7164 ) ;
  assign n7166 = n2105 ^ n449 ^ n256 ;
  assign n7167 = n3090 | n4027 ;
  assign n7168 = n7166 & ~n7167 ;
  assign n7169 = x92 & n1653 ;
  assign n7170 = n629 & n7169 ;
  assign n7171 = n4347 ^ n3367 ^ 1'b0 ;
  assign n7172 = n5604 | n7171 ;
  assign n7173 = ( ~n4409 & n7170 ) | ( ~n4409 & n7172 ) | ( n7170 & n7172 ) ;
  assign n7174 = n3860 & n4282 ;
  assign n7175 = n5241 | n7174 ;
  assign n7176 = n2299 & ~n5642 ;
  assign n7177 = ~n4128 & n7176 ;
  assign n7178 = n4279 ^ n3646 ^ n2559 ;
  assign n7179 = n4383 & ~n7178 ;
  assign n7180 = n6307 ^ n3778 ^ 1'b0 ;
  assign n7181 = n2035 ^ n1898 ^ 1'b0 ;
  assign n7182 = n3963 & n7181 ;
  assign n7183 = ~n3392 & n7182 ;
  assign n7184 = n2102 & ~n4593 ;
  assign n7185 = ( ~n836 & n1321 ) | ( ~n836 & n2030 ) | ( n1321 & n2030 ) ;
  assign n7186 = n7185 ^ n5893 ^ 1'b0 ;
  assign n7187 = n7184 & n7186 ;
  assign n7188 = x62 & ~x225 ;
  assign n7189 = n7188 ^ n4441 ^ 1'b0 ;
  assign n7190 = n7187 & n7189 ;
  assign n7191 = ~n4150 & n6402 ;
  assign n7192 = n5108 ^ n4016 ^ 1'b0 ;
  assign n7193 = n5208 & ~n7192 ;
  assign n7194 = x237 ^ x208 ^ 1'b0 ;
  assign n7195 = ~n3809 & n7194 ;
  assign n7196 = n2600 & n3840 ;
  assign n7197 = n1721 | n3085 ;
  assign n7198 = n2950 | n7197 ;
  assign n7199 = ( n1634 & ~n4832 ) | ( n1634 & n7198 ) | ( ~n4832 & n7198 ) ;
  assign n7200 = n4391 ^ n856 ^ 1'b0 ;
  assign n7201 = n6111 & ~n6118 ;
  assign n7202 = n7200 & n7201 ;
  assign n7203 = n6991 ^ n5569 ^ n2722 ;
  assign n7204 = n6168 & n6447 ;
  assign n7205 = n451 & ~n4512 ;
  assign n7206 = n5448 ^ n1728 ^ 1'b0 ;
  assign n7207 = x104 & ~n7206 ;
  assign n7208 = ~n1475 & n4271 ;
  assign n7209 = n7208 ^ n7124 ^ 1'b0 ;
  assign n7210 = n7209 ^ n5179 ^ 1'b0 ;
  assign n7211 = n7210 ^ n6061 ^ 1'b0 ;
  assign n7212 = n7207 & n7211 ;
  assign n7213 = n4327 & ~n4780 ;
  assign n7214 = n4902 & n7213 ;
  assign n7215 = n6447 ^ n1850 ^ 1'b0 ;
  assign n7216 = n3287 & ~n7215 ;
  assign n7217 = n7216 ^ n4403 ^ 1'b0 ;
  assign n7218 = ~n7214 & n7217 ;
  assign n7219 = n3785 ^ x123 ^ x41 ;
  assign n7220 = n6947 | n7219 ;
  assign n7221 = n431 ^ x244 ^ 1'b0 ;
  assign n7222 = n359 & n7221 ;
  assign n7223 = n2944 | n7222 ;
  assign n7224 = n7223 ^ n1462 ^ 1'b0 ;
  assign n7225 = n2883 | n5315 ;
  assign n7226 = n6134 | n7225 ;
  assign n7227 = ~n665 & n6442 ;
  assign n7228 = n7227 ^ n679 ^ 1'b0 ;
  assign n7229 = ( n2939 & ~n6187 ) | ( n2939 & n7228 ) | ( ~n6187 & n7228 ) ;
  assign n7230 = n5425 ^ n2681 ^ 1'b0 ;
  assign n7231 = n5720 | n7230 ;
  assign n7232 = n2646 & n4919 ;
  assign n7233 = x96 & n618 ;
  assign n7234 = ~n1591 & n7233 ;
  assign n7236 = n3269 ^ n1845 ^ 1'b0 ;
  assign n7237 = ~n5885 & n7236 ;
  assign n7238 = n1680 | n7237 ;
  assign n7235 = ~n3853 & n4276 ;
  assign n7239 = n7238 ^ n7235 ^ 1'b0 ;
  assign n7240 = ( ~n387 & n676 ) | ( ~n387 & n1664 ) | ( n676 & n1664 ) ;
  assign n7241 = n415 & n7240 ;
  assign n7242 = n7241 ^ n993 ^ 1'b0 ;
  assign n7243 = n7242 ^ n1230 ^ 1'b0 ;
  assign n7244 = n5116 ^ n3407 ^ 1'b0 ;
  assign n7245 = n5592 & n7244 ;
  assign n7246 = ~n2314 & n7245 ;
  assign n7247 = ( ~n4397 & n6905 ) | ( ~n4397 & n7011 ) | ( n6905 & n7011 ) ;
  assign n7248 = n1960 & ~n6094 ;
  assign n7249 = n7248 ^ n3296 ^ 1'b0 ;
  assign n7250 = ~n7247 & n7249 ;
  assign n7254 = n6332 ^ n4542 ^ 1'b0 ;
  assign n7255 = n3216 & n7254 ;
  assign n7256 = ~n860 & n7255 ;
  assign n7257 = n7256 ^ n4935 ^ 1'b0 ;
  assign n7258 = n4310 ^ n2143 ^ 1'b0 ;
  assign n7259 = n1630 | n7258 ;
  assign n7260 = n7259 ^ n2307 ^ 1'b0 ;
  assign n7261 = ~n4070 & n7260 ;
  assign n7262 = n7261 ^ n4248 ^ 1'b0 ;
  assign n7263 = n7257 | n7262 ;
  assign n7264 = n7263 ^ n4218 ^ n856 ;
  assign n7251 = ~n3307 & n4245 ;
  assign n7252 = n7251 ^ n1893 ^ 1'b0 ;
  assign n7253 = n1593 & ~n7252 ;
  assign n7265 = n7264 ^ n7253 ^ 1'b0 ;
  assign n7268 = n2081 | n2584 ;
  assign n7269 = n7268 ^ n589 ^ 1'b0 ;
  assign n7266 = n5590 & ~n7042 ;
  assign n7267 = n7252 & ~n7266 ;
  assign n7270 = n7269 ^ n7267 ^ 1'b0 ;
  assign n7271 = ( n481 & ~n1680 ) | ( n481 & n7028 ) | ( ~n1680 & n7028 ) ;
  assign n7272 = ( ~n274 & n416 ) | ( ~n274 & n6004 ) | ( n416 & n6004 ) ;
  assign n7273 = n1091 ^ n503 ^ 1'b0 ;
  assign n7274 = n7273 ^ n2418 ^ 1'b0 ;
  assign n7275 = ( n3421 & ~n5311 ) | ( n3421 & n7274 ) | ( ~n5311 & n7274 ) ;
  assign n7276 = n1660 & ~n6453 ;
  assign n7277 = n963 | n7276 ;
  assign n7278 = n7277 ^ n3532 ^ 1'b0 ;
  assign n7279 = n2172 | n3754 ;
  assign n7280 = ( n792 & n7278 ) | ( n792 & ~n7279 ) | ( n7278 & ~n7279 ) ;
  assign n7281 = ~n5654 & n5754 ;
  assign n7282 = n4198 & n7281 ;
  assign n7283 = n7280 | n7282 ;
  assign n7284 = ~n997 & n3588 ;
  assign n7285 = n7284 ^ n1603 ^ 1'b0 ;
  assign n7286 = n4470 ^ n3293 ^ n3235 ;
  assign n7289 = n716 | n1034 ;
  assign n7287 = n6059 ^ n2256 ^ 1'b0 ;
  assign n7288 = n4519 & n7287 ;
  assign n7290 = n7289 ^ n7288 ^ 1'b0 ;
  assign n7291 = n4056 ^ n3617 ^ 1'b0 ;
  assign n7292 = n7291 ^ n3272 ^ 1'b0 ;
  assign n7293 = n2047 | n2858 ;
  assign n7294 = n7293 ^ n4251 ^ 1'b0 ;
  assign n7295 = n5650 ^ n1292 ^ 1'b0 ;
  assign n7296 = ~n5959 & n7295 ;
  assign n7297 = n592 ^ n437 ^ 1'b0 ;
  assign n7298 = n875 & ~n7297 ;
  assign n7299 = n7298 ^ n3886 ^ 1'b0 ;
  assign n7300 = ~n2387 & n7299 ;
  assign n7301 = n258 & n7300 ;
  assign n7302 = n2722 & ~n3401 ;
  assign n7303 = n7302 ^ n1922 ^ 1'b0 ;
  assign n7304 = n7303 ^ n6112 ^ n4359 ;
  assign n7305 = n3157 & ~n3915 ;
  assign n7306 = n4659 & n7305 ;
  assign n7307 = ( n3255 & n5479 ) | ( n3255 & ~n6483 ) | ( n5479 & ~n6483 ) ;
  assign n7308 = n5840 ^ n399 ^ 1'b0 ;
  assign n7309 = ~n1336 & n2287 ;
  assign n7310 = ~x13 & n7309 ;
  assign n7311 = n917 & ~n7310 ;
  assign n7312 = n7311 ^ n2726 ^ 1'b0 ;
  assign n7313 = n617 & n7312 ;
  assign n7314 = n913 & n7313 ;
  assign n7315 = n2757 ^ n2402 ^ n1684 ;
  assign n7316 = n1894 & ~n2653 ;
  assign n7317 = n1619 & ~n7316 ;
  assign n7318 = n7317 ^ n890 ^ 1'b0 ;
  assign n7319 = ~n370 & n1385 ;
  assign n7320 = x53 & n7319 ;
  assign n7321 = ~n3642 & n7320 ;
  assign n7322 = n2771 ^ n1168 ^ 1'b0 ;
  assign n7323 = n729 & ~n7322 ;
  assign n7324 = n1298 & ~n4265 ;
  assign n7325 = n7324 ^ n3499 ^ 1'b0 ;
  assign n7326 = n1968 | n7325 ;
  assign n7327 = n4669 & ~n7326 ;
  assign n7328 = ~n7323 & n7327 ;
  assign n7329 = ~n7321 & n7328 ;
  assign n7330 = ~n1199 & n4583 ;
  assign n7331 = n7330 ^ n4386 ^ n2137 ;
  assign n7332 = ( n1450 & n1554 ) | ( n1450 & n2349 ) | ( n1554 & n2349 ) ;
  assign n7333 = n4994 ^ n453 ^ 1'b0 ;
  assign n7334 = n4935 & ~n7333 ;
  assign n7335 = ~n7332 & n7334 ;
  assign n7336 = n7335 ^ n7104 ^ 1'b0 ;
  assign n7337 = n7228 ^ n1838 ^ 1'b0 ;
  assign n7338 = ~n1163 & n7337 ;
  assign n7339 = n1417 & n2631 ;
  assign n7340 = n7339 ^ n3313 ^ 1'b0 ;
  assign n7341 = n4445 & ~n7340 ;
  assign n7342 = n7341 ^ x165 ^ 1'b0 ;
  assign n7343 = n7338 & ~n7342 ;
  assign n7344 = ~x74 & n7343 ;
  assign n7345 = n1411 | n7344 ;
  assign n7346 = n7330 ^ x229 ^ 1'b0 ;
  assign n7347 = n6695 & n7346 ;
  assign n7348 = ~n876 & n7347 ;
  assign n7349 = ~x95 & n7348 ;
  assign n7352 = n2710 ^ x240 ^ 1'b0 ;
  assign n7350 = ~x189 & n4093 ;
  assign n7351 = n7350 ^ n3703 ^ 1'b0 ;
  assign n7353 = n7352 ^ n7351 ^ 1'b0 ;
  assign n7354 = n6725 & n7353 ;
  assign n7355 = n7354 ^ n6534 ^ 1'b0 ;
  assign n7358 = n1871 ^ x206 ^ 1'b0 ;
  assign n7356 = n419 | n3577 ;
  assign n7357 = n1975 & ~n7356 ;
  assign n7359 = n7358 ^ n7357 ^ 1'b0 ;
  assign n7361 = ( x174 & n1623 ) | ( x174 & n3462 ) | ( n1623 & n3462 ) ;
  assign n7360 = x41 & n2392 ;
  assign n7362 = n7361 ^ n7360 ^ 1'b0 ;
  assign n7363 = ~n7359 & n7362 ;
  assign n7364 = n7067 ^ n3344 ^ 1'b0 ;
  assign n7365 = n6666 ^ n5022 ^ 1'b0 ;
  assign n7366 = n3450 & ~n4919 ;
  assign n7370 = n806 & n3427 ;
  assign n7367 = n2740 ^ x77 ^ 1'b0 ;
  assign n7368 = n1845 & n7367 ;
  assign n7369 = ~n4552 & n7368 ;
  assign n7371 = n7370 ^ n7369 ^ 1'b0 ;
  assign n7372 = n2430 & n4078 ;
  assign n7373 = n7372 ^ n779 ^ 1'b0 ;
  assign n7374 = ~x33 & x251 ;
  assign n7375 = n7374 ^ n6064 ^ 1'b0 ;
  assign n7381 = n1807 & n3980 ;
  assign n7382 = ( ~n2137 & n6567 ) | ( ~n2137 & n7381 ) | ( n6567 & n7381 ) ;
  assign n7376 = n1416 & ~n1997 ;
  assign n7377 = n7376 ^ n905 ^ 1'b0 ;
  assign n7378 = n707 & ~n7377 ;
  assign n7379 = ~n1053 & n7378 ;
  assign n7380 = ~n5903 & n7379 ;
  assign n7383 = n7382 ^ n7380 ^ 1'b0 ;
  assign n7384 = n1617 ^ n1133 ^ 1'b0 ;
  assign n7385 = n5114 & ~n5840 ;
  assign n7386 = n6008 ^ n1858 ^ 1'b0 ;
  assign n7388 = n5785 ^ n483 ^ 1'b0 ;
  assign n7387 = n5538 ^ n2884 ^ n2231 ;
  assign n7389 = n7388 ^ n7387 ^ n4719 ;
  assign n7390 = n1848 ^ n1765 ^ 1'b0 ;
  assign n7391 = n3400 & n7390 ;
  assign n7392 = n7391 ^ n2223 ^ 1'b0 ;
  assign n7393 = n5087 ^ n3884 ^ 1'b0 ;
  assign n7394 = n3214 & n7393 ;
  assign n7395 = n7394 ^ n485 ^ 1'b0 ;
  assign n7396 = n3440 ^ n3253 ^ 1'b0 ;
  assign n7397 = n6112 ^ n289 ^ 1'b0 ;
  assign n7398 = ~n535 & n1096 ;
  assign n7399 = n2970 ^ n1338 ^ 1'b0 ;
  assign n7400 = n6035 & n6670 ;
  assign n7401 = n7400 ^ n851 ^ 1'b0 ;
  assign n7402 = n7283 ^ n6014 ^ 1'b0 ;
  assign n7403 = n4872 ^ n3340 ^ 1'b0 ;
  assign n7404 = n2978 & n7403 ;
  assign n7405 = n7404 ^ n5536 ^ 1'b0 ;
  assign n7406 = n2308 ^ n1249 ^ 1'b0 ;
  assign n7407 = n1091 & n7406 ;
  assign n7408 = n2011 | n4736 ;
  assign n7409 = n7407 | n7408 ;
  assign n7410 = ~n2086 & n7409 ;
  assign n7411 = n6123 & n7410 ;
  assign n7412 = n7411 ^ n5504 ^ 1'b0 ;
  assign n7413 = n1383 & n1716 ;
  assign n7414 = ~n880 & n7413 ;
  assign n7415 = n7414 ^ n4232 ^ 1'b0 ;
  assign n7416 = x54 & n7415 ;
  assign n7417 = n4212 ^ n4009 ^ 1'b0 ;
  assign n7418 = ~n1632 & n7417 ;
  assign n7419 = n2595 & ~n6430 ;
  assign n7420 = n1230 | n3478 ;
  assign n7421 = ( x73 & ~n1521 ) | ( x73 & n2939 ) | ( ~n1521 & n2939 ) ;
  assign n7422 = n7421 ^ n4516 ^ 1'b0 ;
  assign n7423 = n3574 & n7422 ;
  assign n7424 = n619 & n847 ;
  assign n7425 = n5493 ^ n1718 ^ 1'b0 ;
  assign n7426 = ~n1352 & n7425 ;
  assign n7427 = n1665 & n2230 ;
  assign n7428 = n1053 ^ n593 ^ 1'b0 ;
  assign n7429 = n4794 & ~n7428 ;
  assign n7430 = n7429 ^ n4576 ^ 1'b0 ;
  assign n7431 = n4269 | n6104 ;
  assign n7432 = ~n672 & n977 ;
  assign n7433 = n7432 ^ n3981 ^ n492 ;
  assign n7434 = n6866 & ~n7433 ;
  assign n7435 = ~n4675 & n7434 ;
  assign n7436 = n3873 & n5556 ;
  assign n7437 = n7435 & n7436 ;
  assign n7438 = n382 | n3685 ;
  assign n7439 = n7438 ^ n4666 ^ 1'b0 ;
  assign n7440 = n5711 ^ x51 ^ 1'b0 ;
  assign n7441 = n7439 & n7440 ;
  assign n7442 = n4319 & n7441 ;
  assign n7443 = n467 | n1505 ;
  assign n7444 = n3319 & n5163 ;
  assign n7445 = n7444 ^ n647 ^ 1'b0 ;
  assign n7447 = ( n1985 & ~n4694 ) | ( n1985 & n5383 ) | ( ~n4694 & n5383 ) ;
  assign n7446 = n4227 | n6492 ;
  assign n7448 = n7447 ^ n7446 ^ 1'b0 ;
  assign n7449 = n7445 & ~n7448 ;
  assign n7450 = n597 | n7449 ;
  assign n7451 = x83 & n3399 ;
  assign n7452 = n7451 ^ x23 ^ 1'b0 ;
  assign n7453 = n1866 & n3939 ;
  assign n7454 = ~n3951 & n7453 ;
  assign n7455 = n7454 ^ n659 ^ 1'b0 ;
  assign n7456 = n3027 ^ n1894 ^ x154 ;
  assign n7457 = n7312 ^ n3417 ^ 1'b0 ;
  assign n7458 = ( n1371 & n2474 ) | ( n1371 & ~n3054 ) | ( n2474 & ~n3054 ) ;
  assign n7459 = n4374 ^ n3717 ^ 1'b0 ;
  assign n7460 = ~n6827 & n7459 ;
  assign n7461 = n7458 & n7460 ;
  assign n7462 = n7461 ^ n7448 ^ 1'b0 ;
  assign n7463 = ( n7456 & n7457 ) | ( n7456 & n7462 ) | ( n7457 & n7462 ) ;
  assign n7465 = n2641 & n4705 ;
  assign n7466 = n7465 ^ n5055 ^ 1'b0 ;
  assign n7467 = n7466 ^ n3134 ^ n2351 ;
  assign n7464 = ~n709 & n6631 ;
  assign n7468 = n7467 ^ n7464 ^ 1'b0 ;
  assign n7469 = n3421 & ~n7468 ;
  assign n7470 = n1328 ^ n419 ^ 1'b0 ;
  assign n7471 = n7470 ^ x40 ^ 1'b0 ;
  assign n7472 = ~n2194 & n7471 ;
  assign n7473 = n6563 ^ n353 ^ 1'b0 ;
  assign n7474 = ( n1347 & n4602 ) | ( n1347 & n7473 ) | ( n4602 & n7473 ) ;
  assign n7477 = n4993 ^ n532 ^ 1'b0 ;
  assign n7478 = n2879 & n7477 ;
  assign n7475 = x63 & ~n3140 ;
  assign n7476 = n7475 ^ n3588 ^ 1'b0 ;
  assign n7479 = n7478 ^ n7476 ^ 1'b0 ;
  assign n7480 = n3947 & n7479 ;
  assign n7481 = n3050 ^ n2076 ^ 1'b0 ;
  assign n7482 = n794 & ~n7481 ;
  assign n7483 = n3253 ^ n1492 ^ 1'b0 ;
  assign n7484 = x169 | n7483 ;
  assign n7485 = n4290 & ~n7484 ;
  assign n7486 = n7482 | n7485 ;
  assign n7487 = n7486 ^ n3458 ^ 1'b0 ;
  assign n7488 = n1494 & ~n2840 ;
  assign n7489 = n491 & n7488 ;
  assign n7490 = n7489 ^ n3045 ^ 1'b0 ;
  assign n7491 = ( n1923 & ~n3283 ) | ( n1923 & n3415 ) | ( ~n3283 & n3415 ) ;
  assign n7492 = n2091 & n7491 ;
  assign n7493 = n1395 | n3481 ;
  assign n7494 = n5743 & n7371 ;
  assign n7495 = n1365 ^ n335 ^ x107 ;
  assign n7496 = x181 & ~n7495 ;
  assign n7497 = n4400 ^ n3327 ^ 1'b0 ;
  assign n7498 = n2008 & ~n7497 ;
  assign n7499 = ~n7496 & n7498 ;
  assign n7500 = n6404 ^ n1956 ^ 1'b0 ;
  assign n7501 = n6796 & ~n7500 ;
  assign n7502 = n389 & n3169 ;
  assign n7503 = n3129 | n7502 ;
  assign n7504 = n7503 ^ n7423 ^ 1'b0 ;
  assign n7506 = n1954 & n2479 ;
  assign n7507 = n2631 & ~n7506 ;
  assign n7508 = x180 & n5560 ;
  assign n7509 = n7508 ^ n3657 ^ 1'b0 ;
  assign n7510 = n7507 | n7509 ;
  assign n7505 = x14 & n404 ;
  assign n7511 = n7510 ^ n7505 ^ 1'b0 ;
  assign n7512 = n6101 ^ n402 ^ 1'b0 ;
  assign n7513 = n6781 & ~n7512 ;
  assign n7514 = x6 | n1952 ;
  assign n7515 = x116 | n7514 ;
  assign n7516 = n3579 ^ n2164 ^ n2119 ;
  assign n7518 = n2208 & n2501 ;
  assign n7517 = n1032 & ~n2176 ;
  assign n7519 = n7518 ^ n7517 ^ 1'b0 ;
  assign n7520 = n1943 & ~n7519 ;
  assign n7521 = n5179 ^ n5034 ^ n1736 ;
  assign n7522 = n7520 & ~n7521 ;
  assign n7523 = n5560 ^ n1311 ^ 1'b0 ;
  assign n7524 = n4685 ^ n3666 ^ 1'b0 ;
  assign n7525 = n4591 | n4611 ;
  assign n7526 = n7525 ^ n4157 ^ 1'b0 ;
  assign n7527 = ~n3156 & n7526 ;
  assign n7528 = ~x1 & n7527 ;
  assign n7529 = n7059 ^ n2681 ^ 1'b0 ;
  assign n7530 = n5497 & n7529 ;
  assign n7531 = n1795 & n3879 ;
  assign n7532 = n7531 ^ n737 ^ 1'b0 ;
  assign n7533 = ~n2611 & n2935 ;
  assign n7534 = n7532 & n7533 ;
  assign n7535 = n2749 | n7534 ;
  assign n7536 = n2244 & ~n7535 ;
  assign n7537 = n7536 ^ x184 ^ 1'b0 ;
  assign n7538 = n2316 | n7537 ;
  assign n7539 = n5368 | n5465 ;
  assign n7540 = n518 & n4313 ;
  assign n7541 = n7282 & n7540 ;
  assign n7542 = n6010 ^ n2647 ^ 1'b0 ;
  assign n7546 = n3390 ^ n1016 ^ 1'b0 ;
  assign n7547 = ~n2975 & n7546 ;
  assign n7548 = n2767 & n7547 ;
  assign n7549 = n7548 ^ n1593 ^ 1'b0 ;
  assign n7544 = x26 & ~n5811 ;
  assign n7545 = n2769 & n7544 ;
  assign n7543 = n5913 ^ n2812 ^ 1'b0 ;
  assign n7550 = n7549 ^ n7545 ^ n7543 ;
  assign n7551 = n3367 ^ n3122 ^ 1'b0 ;
  assign n7552 = n893 | n7551 ;
  assign n7553 = n2404 & ~n7552 ;
  assign n7554 = x139 & n411 ;
  assign n7555 = n928 & n6342 ;
  assign n7556 = n274 & n7555 ;
  assign n7557 = n7170 & n7556 ;
  assign n7558 = n7190 ^ n5727 ^ 1'b0 ;
  assign n7559 = n5818 ^ n2582 ^ 1'b0 ;
  assign n7560 = ~n4206 & n7559 ;
  assign n7561 = n7560 ^ n4512 ^ 1'b0 ;
  assign n7562 = n5796 & ~n7178 ;
  assign n7563 = n375 & ~n7562 ;
  assign n7564 = n4710 ^ n4205 ^ 1'b0 ;
  assign n7565 = n6307 ^ x213 ^ 1'b0 ;
  assign n7566 = x144 & n754 ;
  assign n7567 = n7566 ^ n4948 ^ n2967 ;
  assign n7568 = n7567 ^ n5298 ^ n2453 ;
  assign n7569 = x169 | n5104 ;
  assign n7570 = n7419 ^ n1221 ^ 1'b0 ;
  assign n7571 = ( n461 & n1220 ) | ( n461 & ~n2144 ) | ( n1220 & ~n2144 ) ;
  assign n7572 = n453 & ~n7571 ;
  assign n7573 = n3878 & n7572 ;
  assign n7574 = n7573 ^ n4185 ^ 1'b0 ;
  assign n7575 = n4094 & n7574 ;
  assign n7576 = n3600 & ~n5559 ;
  assign n7577 = n1876 & n4754 ;
  assign n7578 = n7577 ^ n618 ^ 1'b0 ;
  assign n7579 = n7578 ^ n4780 ^ 1'b0 ;
  assign n7580 = n3627 ^ n2369 ^ 1'b0 ;
  assign n7581 = n7580 ^ n2247 ^ 1'b0 ;
  assign n7582 = n4845 & n6808 ;
  assign n7583 = n3313 & ~n5934 ;
  assign n7584 = ( n6666 & ~n7582 ) | ( n6666 & n7583 ) | ( ~n7582 & n7583 ) ;
  assign n7585 = n4076 ^ n1456 ^ 1'b0 ;
  assign n7586 = n4807 | n7585 ;
  assign n7587 = x116 | n7586 ;
  assign n7592 = ( ~n2634 & n4022 ) | ( ~n2634 & n6382 ) | ( n4022 & n6382 ) ;
  assign n7588 = n3147 ^ n2983 ^ 1'b0 ;
  assign n7589 = n2047 | n2663 ;
  assign n7590 = n1757 | n7589 ;
  assign n7591 = n7588 & n7590 ;
  assign n7593 = n7592 ^ n7591 ^ 1'b0 ;
  assign n7594 = n2672 ^ n2260 ^ n614 ;
  assign n7595 = n328 & ~n7594 ;
  assign n7596 = n7595 ^ n6115 ^ 1'b0 ;
  assign n7597 = ( n372 & ~n3890 ) | ( n372 & n5382 ) | ( ~n3890 & n5382 ) ;
  assign n7598 = n1802 & n7597 ;
  assign n7599 = n2631 & ~n3003 ;
  assign n7600 = ~x70 & n7599 ;
  assign n7601 = ~n3222 & n3349 ;
  assign n7602 = ( x149 & n680 ) | ( x149 & ~n7601 ) | ( n680 & ~n7601 ) ;
  assign n7603 = ( ~n1725 & n7600 ) | ( ~n1725 & n7602 ) | ( n7600 & n7602 ) ;
  assign n7604 = ~n2521 & n7603 ;
  assign n7605 = ~n7598 & n7604 ;
  assign n7606 = n6572 ^ n2122 ^ 1'b0 ;
  assign n7607 = ( n2098 & n5976 ) | ( n2098 & ~n7606 ) | ( n5976 & ~n7606 ) ;
  assign n7608 = n7607 ^ n2345 ^ 1'b0 ;
  assign n7609 = n2008 ^ n1353 ^ 1'b0 ;
  assign n7610 = n7609 ^ n896 ^ 1'b0 ;
  assign n7611 = n1548 & n7610 ;
  assign n7612 = n1387 & n5651 ;
  assign n7613 = n4588 & n7612 ;
  assign n7614 = n2227 ^ n970 ^ 1'b0 ;
  assign n7615 = ~n3419 & n7614 ;
  assign n7617 = n5127 ^ n1735 ^ 1'b0 ;
  assign n7618 = n7617 ^ n629 ^ 1'b0 ;
  assign n7619 = ~n2633 & n7618 ;
  assign n7620 = ~n4367 & n6350 ;
  assign n7621 = n7619 & n7620 ;
  assign n7622 = ~n4443 & n7621 ;
  assign n7616 = n2967 | n5452 ;
  assign n7623 = n7622 ^ n7616 ^ 1'b0 ;
  assign n7624 = ~x144 & n394 ;
  assign n7627 = n1373 | n2237 ;
  assign n7625 = x23 & x46 ;
  assign n7626 = n7625 ^ n2011 ^ 1'b0 ;
  assign n7628 = n7627 ^ n7626 ^ 1'b0 ;
  assign n7629 = ~n7624 & n7628 ;
  assign n7630 = x73 & n2306 ;
  assign n7631 = ( n1562 & n3649 ) | ( n1562 & n7630 ) | ( n3649 & n7630 ) ;
  assign n7632 = n692 & n7631 ;
  assign n7633 = n7632 ^ n752 ^ 1'b0 ;
  assign n7634 = n1605 | n7633 ;
  assign n7635 = n2905 ^ n2200 ^ 1'b0 ;
  assign n7636 = n7635 ^ n2798 ^ 1'b0 ;
  assign n7637 = n5374 & ~n7636 ;
  assign n7638 = n7637 ^ n5437 ^ n3504 ;
  assign n7639 = n3933 & ~n4663 ;
  assign n7640 = n7639 ^ n4515 ^ 1'b0 ;
  assign n7641 = ~n5170 & n7640 ;
  assign n7642 = n7141 ^ n4998 ^ 1'b0 ;
  assign n7643 = n357 & ~n7642 ;
  assign n7644 = n4434 & n7643 ;
  assign n7645 = n6816 ^ n4984 ^ 1'b0 ;
  assign n7646 = n7644 | n7645 ;
  assign n7647 = n7276 ^ n1326 ^ 1'b0 ;
  assign n7648 = n3454 ^ n2670 ^ 1'b0 ;
  assign n7649 = n4354 & n7648 ;
  assign n7650 = ~n7647 & n7649 ;
  assign n7651 = ( ~n713 & n5608 ) | ( ~n713 & n7650 ) | ( n5608 & n7650 ) ;
  assign n7652 = n5961 ^ n5525 ^ 1'b0 ;
  assign n7653 = n7652 ^ n2262 ^ n365 ;
  assign n7654 = n417 & ~n2736 ;
  assign n7656 = x115 & n1395 ;
  assign n7657 = n2901 & n7656 ;
  assign n7655 = n2063 ^ n968 ^ 1'b0 ;
  assign n7658 = n7657 ^ n7655 ^ 1'b0 ;
  assign n7659 = n2095 & ~n7658 ;
  assign n7660 = ( n1763 & n2403 ) | ( n1763 & n3944 ) | ( n2403 & n3944 ) ;
  assign n7661 = x41 & ~n4842 ;
  assign n7662 = ~n7660 & n7661 ;
  assign n7663 = n1008 & n7662 ;
  assign n7664 = n4638 ^ n274 ^ 1'b0 ;
  assign n7665 = n7664 ^ n6939 ^ n905 ;
  assign n7666 = ~n908 & n5925 ;
  assign n7667 = n6584 ^ n4736 ^ 1'b0 ;
  assign n7668 = n3614 | n7667 ;
  assign n7669 = n2574 ^ n1496 ^ 1'b0 ;
  assign n7670 = n1120 & ~n7669 ;
  assign n7671 = ( ~x140 & n1730 ) | ( ~x140 & n7670 ) | ( n1730 & n7670 ) ;
  assign n7672 = n4328 & ~n7671 ;
  assign n7673 = n7672 ^ n2732 ^ 1'b0 ;
  assign n7674 = n2125 | n7673 ;
  assign n7675 = x55 & ~x197 ;
  assign n7676 = n7675 ^ n359 ^ 1'b0 ;
  assign n7679 = n6700 ^ n2942 ^ 1'b0 ;
  assign n7677 = n1877 | n3817 ;
  assign n7678 = ~n532 & n7677 ;
  assign n7680 = n7679 ^ n7678 ^ 1'b0 ;
  assign n7681 = n3088 & ~n7680 ;
  assign n7682 = n4924 ^ n1430 ^ 1'b0 ;
  assign n7683 = n1219 & n7682 ;
  assign n7684 = n3040 ^ n514 ^ 1'b0 ;
  assign n7685 = n4235 & ~n7684 ;
  assign n7686 = ( n1114 & n7683 ) | ( n1114 & n7685 ) | ( n7683 & n7685 ) ;
  assign n7687 = n6723 | n7686 ;
  assign n7688 = n4166 ^ n2516 ^ 1'b0 ;
  assign n7689 = n2895 | n7688 ;
  assign n7690 = n2436 | n7689 ;
  assign n7691 = n7690 ^ n7029 ^ 1'b0 ;
  assign n7692 = n627 | n1711 ;
  assign n7693 = ( n1503 & n5431 ) | ( n1503 & ~n7692 ) | ( n5431 & ~n7692 ) ;
  assign n7694 = ~n466 & n1103 ;
  assign n7695 = n7694 ^ n4484 ^ 1'b0 ;
  assign n7696 = n1963 & n7361 ;
  assign n7697 = n7696 ^ n2085 ^ n2001 ;
  assign n7698 = n7695 & n7697 ;
  assign n7699 = n7698 ^ n6119 ^ 1'b0 ;
  assign n7700 = n2387 ^ n2097 ^ n274 ;
  assign n7701 = n7700 ^ n5803 ^ 1'b0 ;
  assign n7702 = n3931 ^ n2443 ^ x192 ;
  assign n7703 = n4929 & ~n5474 ;
  assign n7704 = ~n4094 & n5768 ;
  assign n7705 = n4832 ^ n409 ^ 1'b0 ;
  assign n7706 = x14 & n4139 ;
  assign n7707 = ( n6426 & ~n7705 ) | ( n6426 & n7706 ) | ( ~n7705 & n7706 ) ;
  assign n7708 = n1779 ^ n860 ^ 1'b0 ;
  assign n7709 = n2567 | n7708 ;
  assign n7710 = ~n716 & n7709 ;
  assign n7711 = ~n2306 & n7710 ;
  assign n7712 = n2975 & ~n6693 ;
  assign n7713 = ~n723 & n3223 ;
  assign n7714 = n7713 ^ n6402 ^ 1'b0 ;
  assign n7715 = n6322 | n7714 ;
  assign n7716 = n7715 ^ n5398 ^ 1'b0 ;
  assign n7717 = x18 & ~n6765 ;
  assign n7718 = n5076 | n7717 ;
  assign n7719 = n6343 & ~n7718 ;
  assign n7720 = n7719 ^ n4649 ^ 1'b0 ;
  assign n7721 = n1103 & n7720 ;
  assign n7722 = n7721 ^ x107 ^ 1'b0 ;
  assign n7723 = n2433 & n4515 ;
  assign n7724 = n2939 & n7723 ;
  assign n7725 = ~n4293 & n7724 ;
  assign n7726 = n7725 ^ n3868 ^ 1'b0 ;
  assign n7727 = n3704 ^ n2226 ^ 1'b0 ;
  assign n7728 = n5163 | n7727 ;
  assign n7729 = n7728 ^ n3287 ^ 1'b0 ;
  assign n7730 = n1303 ^ n409 ^ 1'b0 ;
  assign n7731 = n4208 & ~n7730 ;
  assign n7732 = ~n5060 & n7731 ;
  assign n7733 = n6972 ^ n2843 ^ 1'b0 ;
  assign n7734 = n7732 & ~n7733 ;
  assign n7735 = n2482 ^ n951 ^ 1'b0 ;
  assign n7736 = n3858 & n7735 ;
  assign n7737 = n1612 & ~n3462 ;
  assign n7738 = n7737 ^ n4688 ^ 1'b0 ;
  assign n7739 = ~n1848 & n3380 ;
  assign n7740 = n3532 ^ n560 ^ 1'b0 ;
  assign n7741 = n1657 | n7740 ;
  assign n7742 = ~n369 & n1198 ;
  assign n7743 = ( n3119 & n4432 ) | ( n3119 & n7742 ) | ( n4432 & n7742 ) ;
  assign n7744 = n1749 & ~n7743 ;
  assign n7745 = n6291 & n7744 ;
  assign n7746 = n3180 & ~n4169 ;
  assign n7747 = n1069 | n2011 ;
  assign n7748 = n7747 ^ n2462 ^ 1'b0 ;
  assign n7749 = ~n7606 & n7748 ;
  assign n7750 = ~n2039 & n7749 ;
  assign n7751 = n7750 ^ n2681 ^ 1'b0 ;
  assign n7752 = n1521 & ~n7751 ;
  assign n7753 = n4310 ^ n1958 ^ 1'b0 ;
  assign n7754 = n7015 & n7753 ;
  assign n7755 = n4811 ^ n3917 ^ 1'b0 ;
  assign n7756 = n809 & ~n1043 ;
  assign n7757 = n7756 ^ n2509 ^ 1'b0 ;
  assign n7758 = n1534 & n7757 ;
  assign n7759 = n7758 ^ n5579 ^ 1'b0 ;
  assign n7760 = n6559 | n7759 ;
  assign n7761 = n812 & ~n7760 ;
  assign n7762 = n7755 & ~n7761 ;
  assign n7763 = ~n4974 & n7762 ;
  assign n7764 = n765 | n7763 ;
  assign n7765 = n7764 ^ n3257 ^ 1'b0 ;
  assign n7766 = n7765 ^ n6834 ^ 1'b0 ;
  assign n7767 = n7473 ^ n3530 ^ 1'b0 ;
  assign n7768 = n6817 | n7767 ;
  assign n7769 = n6114 ^ n4248 ^ 1'b0 ;
  assign n7770 = ~n1225 & n7111 ;
  assign n7771 = n3508 & ~n4923 ;
  assign n7772 = n7771 ^ n7714 ^ 1'b0 ;
  assign n7775 = n3332 ^ n1413 ^ 1'b0 ;
  assign n7773 = n5062 ^ n3258 ^ 1'b0 ;
  assign n7774 = n1234 & n7773 ;
  assign n7776 = n7775 ^ n7774 ^ 1'b0 ;
  assign n7777 = n3116 ^ n1208 ^ 1'b0 ;
  assign n7778 = n1079 | n7777 ;
  assign n7779 = n433 | n1023 ;
  assign n7780 = n3942 & n7779 ;
  assign n7781 = n1116 & n7780 ;
  assign n7782 = n3942 ^ n2013 ^ 1'b0 ;
  assign n7783 = n400 & ~n7782 ;
  assign n7784 = n4453 & n7783 ;
  assign n7785 = n7784 ^ n1887 ^ 1'b0 ;
  assign n7786 = n7781 | n7785 ;
  assign n7787 = n7786 ^ n3990 ^ 1'b0 ;
  assign n7788 = ~n1279 & n7787 ;
  assign n7789 = x145 | n7265 ;
  assign n7790 = n611 | n2170 ;
  assign n7791 = n3446 | n7790 ;
  assign n7792 = n4031 ^ n3380 ^ 1'b0 ;
  assign n7793 = n5659 | n7792 ;
  assign n7794 = n7791 | n7793 ;
  assign n7795 = ~n3736 & n7794 ;
  assign n7796 = ~n3864 & n7795 ;
  assign n7797 = n7484 ^ x126 ^ 1'b0 ;
  assign n7798 = n3876 & ~n7797 ;
  assign n7799 = n7342 | n7798 ;
  assign n7800 = ~n716 & n4871 ;
  assign n7801 = n7800 ^ n2905 ^ 1'b0 ;
  assign n7802 = n5606 | n6357 ;
  assign n7803 = n7801 & ~n7802 ;
  assign n7804 = x193 & n3474 ;
  assign n7805 = n3404 & n7804 ;
  assign n7806 = ~n1921 & n6313 ;
  assign n7807 = ( n3534 & n6529 ) | ( n3534 & n6869 ) | ( n6529 & n6869 ) ;
  assign n7808 = ~n7806 & n7807 ;
  assign n7809 = n7808 ^ n4650 ^ 1'b0 ;
  assign n7810 = ( n2872 & n3145 ) | ( n2872 & n6381 ) | ( n3145 & n6381 ) ;
  assign n7811 = n7810 ^ n1848 ^ 1'b0 ;
  assign n7812 = n431 & n3710 ;
  assign n7813 = n3892 ^ n1653 ^ n733 ;
  assign n7814 = n4639 | n7813 ;
  assign n7815 = n2706 ^ n1763 ^ 1'b0 ;
  assign n7816 = n3362 & n5307 ;
  assign n7817 = n7816 ^ n4386 ^ 1'b0 ;
  assign n7818 = n7815 & n7817 ;
  assign n7819 = n293 & ~n4478 ;
  assign n7820 = n7819 ^ n3344 ^ 1'b0 ;
  assign n7821 = n3137 | n7820 ;
  assign n7822 = n1940 ^ n1443 ^ 1'b0 ;
  assign n7823 = n2206 & n7822 ;
  assign n7824 = n7823 ^ n1772 ^ 1'b0 ;
  assign n7825 = n1780 ^ n801 ^ 1'b0 ;
  assign n7826 = n7824 | n7825 ;
  assign n7827 = n5557 ^ n2653 ^ 1'b0 ;
  assign n7828 = n1681 ^ n1213 ^ 1'b0 ;
  assign n7829 = n3035 | n7828 ;
  assign n7830 = n7827 | n7829 ;
  assign n7831 = ~n4040 & n7830 ;
  assign n7832 = ~n1161 & n1322 ;
  assign n7833 = n604 & ~n7118 ;
  assign n7834 = ( n3596 & ~n4361 ) | ( n3596 & n7833 ) | ( ~n4361 & n7833 ) ;
  assign n7835 = n580 & n1195 ;
  assign n7836 = n7835 ^ n3332 ^ 1'b0 ;
  assign n7837 = n4033 ^ x145 ^ 1'b0 ;
  assign n7838 = n1833 & n7837 ;
  assign n7839 = ( x196 & n277 ) | ( x196 & n1513 ) | ( n277 & n1513 ) ;
  assign n7840 = n7839 ^ n6728 ^ n3648 ;
  assign n7841 = n7240 ^ n3892 ^ 1'b0 ;
  assign n7842 = n1610 & n7841 ;
  assign n7843 = n7842 ^ n4871 ^ 1'b0 ;
  assign n7844 = n7670 & n7843 ;
  assign n7845 = x150 & ~n2161 ;
  assign n7846 = n7845 ^ x184 ^ 1'b0 ;
  assign n7847 = n722 & n7846 ;
  assign n7848 = n7847 ^ n589 ^ 1'b0 ;
  assign n7849 = ( n998 & n1828 ) | ( n998 & n4698 ) | ( n1828 & n4698 ) ;
  assign n7850 = n4205 ^ n1494 ^ 1'b0 ;
  assign n7851 = n7849 & n7850 ;
  assign n7852 = n7851 ^ n2020 ^ 1'b0 ;
  assign n7853 = n1738 & ~n7852 ;
  assign n7854 = n1146 | n1876 ;
  assign n7855 = n973 & ~n7854 ;
  assign n7856 = ( n7848 & n7853 ) | ( n7848 & n7855 ) | ( n7853 & n7855 ) ;
  assign n7857 = ~n2897 & n7004 ;
  assign n7858 = ~n5393 & n7857 ;
  assign n7859 = n7858 ^ n2426 ^ 1'b0 ;
  assign n7860 = n4082 ^ n3172 ^ 1'b0 ;
  assign n7861 = n7177 & n7860 ;
  assign n7863 = ( n494 & n796 ) | ( n494 & ~n2077 ) | ( n796 & ~n2077 ) ;
  assign n7862 = n2968 | n4656 ;
  assign n7864 = n7863 ^ n7862 ^ 1'b0 ;
  assign n7865 = n7864 ^ n6583 ^ 1'b0 ;
  assign n7866 = n3929 & n7865 ;
  assign n7867 = n7210 ^ n2448 ^ 1'b0 ;
  assign n7868 = n4375 | n7648 ;
  assign n7869 = n587 & n7868 ;
  assign n7871 = ~n446 & n2595 ;
  assign n7872 = ( n4139 & ~n5416 ) | ( n4139 & n7871 ) | ( ~n5416 & n7871 ) ;
  assign n7870 = x25 & ~n7316 ;
  assign n7873 = n7872 ^ n7870 ^ 1'b0 ;
  assign n7874 = ~n1815 & n5176 ;
  assign n7875 = n7496 & ~n7874 ;
  assign n7876 = n4718 ^ n1276 ^ 1'b0 ;
  assign n7877 = n7876 ^ n4290 ^ 1'b0 ;
  assign n7878 = n7877 ^ n3218 ^ 1'b0 ;
  assign n7879 = n7875 & n7878 ;
  assign n7880 = n4209 ^ n2898 ^ 1'b0 ;
  assign n7881 = n2394 ^ n318 ^ 1'b0 ;
  assign n7882 = n5803 & ~n7881 ;
  assign n7883 = n511 ^ x10 ^ 1'b0 ;
  assign n7884 = n2782 | n7883 ;
  assign n7885 = n3942 & n6157 ;
  assign n7886 = n7884 & n7885 ;
  assign n7887 = n5713 ^ n5266 ^ 1'b0 ;
  assign n7888 = ( n851 & n916 ) | ( n851 & ~n1573 ) | ( n916 & ~n1573 ) ;
  assign n7889 = n7888 ^ n7404 ^ 1'b0 ;
  assign n7890 = n3683 | n7889 ;
  assign n7891 = ~n2620 & n7890 ;
  assign n7896 = ( n904 & ~n1496 ) | ( n904 & n2311 ) | ( ~n1496 & n2311 ) ;
  assign n7892 = n4170 & n6994 ;
  assign n7893 = n548 & n7892 ;
  assign n7894 = n6274 | n7759 ;
  assign n7895 = n7893 & ~n7894 ;
  assign n7897 = n7896 ^ n7895 ^ n3791 ;
  assign n7898 = n6015 ^ n3513 ^ 1'b0 ;
  assign n7899 = ~n589 & n7799 ;
  assign n7900 = n522 | n2067 ;
  assign n7901 = n3294 & n4918 ;
  assign n7902 = ~x146 & n7901 ;
  assign n7903 = n1039 | n7902 ;
  assign n7904 = ~n7657 & n7903 ;
  assign n7905 = n6582 ^ n4940 ^ 1'b0 ;
  assign n7906 = n7904 | n7905 ;
  assign n7907 = n5970 & n7906 ;
  assign n7908 = n7900 & n7907 ;
  assign n7909 = n400 & ~n3420 ;
  assign n7910 = n7909 ^ n7258 ^ x201 ;
  assign n7911 = ~n4616 & n7910 ;
  assign n7912 = n1789 & ~n7855 ;
  assign n7913 = n7912 ^ n2653 ^ 1'b0 ;
  assign n7914 = x91 & n7913 ;
  assign n7915 = n7914 ^ n7800 ^ 1'b0 ;
  assign n7916 = n7334 & ~n7915 ;
  assign n7917 = n4598 ^ n4132 ^ 1'b0 ;
  assign n7918 = n7294 ^ n2163 ^ 1'b0 ;
  assign n7919 = n1120 & ~n3721 ;
  assign n7920 = n7919 ^ n1001 ^ 1'b0 ;
  assign n7921 = ~n498 & n7920 ;
  assign n7922 = ~n4677 & n7921 ;
  assign n7923 = n3950 & n5497 ;
  assign n7924 = n7923 ^ n7664 ^ 1'b0 ;
  assign n7925 = ~n7372 & n7924 ;
  assign n7926 = n4432 ^ n3195 ^ 1'b0 ;
  assign n7927 = x115 & ~n7926 ;
  assign n7928 = n679 | n3472 ;
  assign n7929 = n4232 & ~n7928 ;
  assign n7930 = x183 & ~n7929 ;
  assign n7931 = n5316 ^ n5135 ^ 1'b0 ;
  assign n7932 = n7467 & ~n7931 ;
  assign n7933 = n1605 & n7932 ;
  assign n7934 = n4762 ^ n3600 ^ 1'b0 ;
  assign n7935 = ~n2291 & n6711 ;
  assign n7936 = n679 ^ x132 ^ 1'b0 ;
  assign n7937 = ~n7935 & n7936 ;
  assign n7938 = n3778 & n7937 ;
  assign n7939 = n5622 ^ n1956 ^ 1'b0 ;
  assign n7940 = n767 & n7939 ;
  assign n7941 = n3088 & ~n4506 ;
  assign n7942 = n3606 | n7166 ;
  assign n7943 = n3052 | n3102 ;
  assign n7944 = n7943 ^ n4093 ^ 1'b0 ;
  assign n7945 = n2919 ^ n1758 ^ 1'b0 ;
  assign n7946 = n537 & n7945 ;
  assign n7947 = ~n7944 & n7946 ;
  assign n7948 = ~n3014 & n7683 ;
  assign n7951 = ~n3345 & n6516 ;
  assign n7949 = ( n464 & ~n3156 ) | ( n464 & n4518 ) | ( ~n3156 & n4518 ) ;
  assign n7950 = n4402 & n7949 ;
  assign n7952 = n7951 ^ n7950 ^ 1'b0 ;
  assign n7953 = n7952 ^ n5450 ^ 1'b0 ;
  assign n7954 = n3728 & n7953 ;
  assign n7956 = ~n3427 & n7358 ;
  assign n7957 = ~n2823 & n7956 ;
  assign n7955 = ~n3685 & n5540 ;
  assign n7958 = n7957 ^ n7955 ^ 1'b0 ;
  assign n7959 = n7939 ^ n2058 ^ n733 ;
  assign n7960 = n3673 ^ n263 ^ 1'b0 ;
  assign n7961 = n1152 | n7960 ;
  assign n7962 = n7961 ^ n3751 ^ 1'b0 ;
  assign n7963 = ~n1148 & n1558 ;
  assign n7964 = n7963 ^ n5119 ^ n3417 ;
  assign n7968 = n2302 & n4936 ;
  assign n7965 = n3382 ^ x121 ^ 1'b0 ;
  assign n7966 = x184 & n7965 ;
  assign n7967 = n7966 ^ n2400 ^ x212 ;
  assign n7969 = n7968 ^ n7967 ^ 1'b0 ;
  assign n7970 = ( n725 & n5255 ) | ( n725 & n6006 ) | ( n5255 & n6006 ) ;
  assign n7971 = n7496 | n7970 ;
  assign n7972 = x87 & x153 ;
  assign n7973 = n7972 ^ n6009 ^ n1219 ;
  assign n7974 = n908 | n6276 ;
  assign n7975 = n7263 ^ n4935 ^ 1'b0 ;
  assign n7976 = n844 & n4992 ;
  assign n7977 = n7381 ^ n5532 ^ 1'b0 ;
  assign n7978 = n5767 & n7977 ;
  assign n7979 = n6873 & n7978 ;
  assign n7982 = n453 & ~n2772 ;
  assign n7983 = n2122 & n7982 ;
  assign n7980 = n5121 ^ n548 ^ 1'b0 ;
  assign n7981 = n4355 | n7980 ;
  assign n7984 = n7983 ^ n7981 ^ n920 ;
  assign n7985 = n7984 ^ n2086 ^ 1'b0 ;
  assign n7986 = ( x214 & n3055 ) | ( x214 & ~n6070 ) | ( n3055 & ~n6070 ) ;
  assign n7987 = n7985 & n7986 ;
  assign n7988 = n2424 ^ n1103 ^ 1'b0 ;
  assign n7989 = n1945 & ~n7988 ;
  assign n7990 = x9 & ~x211 ;
  assign n7991 = n665 | n1835 ;
  assign n7992 = n756 | n7991 ;
  assign n7993 = ~n1185 & n1393 ;
  assign n7994 = n3703 & n7993 ;
  assign n7995 = n4482 & ~n7994 ;
  assign n7996 = n7995 ^ n1257 ^ 1'b0 ;
  assign n7997 = n3458 & ~n6365 ;
  assign n7998 = n7997 ^ n990 ^ 1'b0 ;
  assign n7999 = ~n2311 & n5465 ;
  assign n8000 = n7999 ^ n7817 ^ 1'b0 ;
  assign n8001 = ~n2804 & n5632 ;
  assign n8002 = ~n1428 & n8001 ;
  assign n8003 = n5488 ^ n1606 ^ 1'b0 ;
  assign n8004 = n631 & n8003 ;
  assign n8005 = n2282 | n4438 ;
  assign n8006 = x169 | n496 ;
  assign n8007 = n8006 ^ x37 ^ 1'b0 ;
  assign n8008 = n5214 & n8007 ;
  assign n8009 = n2163 & ~n5438 ;
  assign n8014 = n1163 | n1167 ;
  assign n8015 = n2702 & ~n8014 ;
  assign n8013 = n2187 & n5385 ;
  assign n8016 = n8015 ^ n8013 ^ 1'b0 ;
  assign n8017 = n5218 ^ n3260 ^ 1'b0 ;
  assign n8018 = n8016 & ~n8017 ;
  assign n8010 = n3156 | n3171 ;
  assign n8011 = n3716 | n8010 ;
  assign n8012 = n8011 ^ n4968 ^ 1'b0 ;
  assign n8019 = n8018 ^ n8012 ^ 1'b0 ;
  assign n8020 = n5277 & ~n8019 ;
  assign n8021 = n1456 & ~n2711 ;
  assign n8022 = ~n4711 & n8021 ;
  assign n8023 = n2622 & ~n2895 ;
  assign n8024 = n8023 ^ n2146 ^ 1'b0 ;
  assign n8025 = n8024 ^ n7549 ^ 1'b0 ;
  assign n8026 = n7237 ^ n2668 ^ n1486 ;
  assign n8027 = n5833 & n7827 ;
  assign n8028 = ~n5339 & n8027 ;
  assign n8029 = n8026 | n8028 ;
  assign n8030 = n4264 ^ n1855 ^ 1'b0 ;
  assign n8031 = n1109 & ~n5020 ;
  assign n8032 = n923 & ~n993 ;
  assign n8033 = ~n2428 & n8032 ;
  assign n8034 = ~n2109 & n5885 ;
  assign n8035 = n8033 | n8034 ;
  assign n8036 = n7908 | n8035 ;
  assign n8037 = n3856 ^ n2710 ^ n1333 ;
  assign n8038 = n3050 & n8037 ;
  assign n8039 = n4323 & ~n8038 ;
  assign n8040 = n3046 ^ n1373 ^ 1'b0 ;
  assign n8041 = ~n1882 & n8040 ;
  assign n8042 = n4198 & n8041 ;
  assign n8043 = ~n3198 & n8042 ;
  assign n8044 = ( x128 & ~n7433 ) | ( x128 & n8043 ) | ( ~n7433 & n8043 ) ;
  assign n8045 = ~n810 & n7746 ;
  assign n8046 = n8045 ^ n3832 ^ 1'b0 ;
  assign n8047 = n6014 ^ n2525 ^ 1'b0 ;
  assign n8048 = ~n2878 & n8047 ;
  assign n8049 = n1163 & n7130 ;
  assign n8050 = n1593 ^ n742 ^ 1'b0 ;
  assign n8051 = n5054 | n5380 ;
  assign n8052 = n8050 | n8051 ;
  assign n8053 = n8052 ^ n7745 ^ 1'b0 ;
  assign n8054 = n5976 ^ n2062 ^ 1'b0 ;
  assign n8055 = n263 & n5626 ;
  assign n8056 = n8055 ^ n2390 ^ 1'b0 ;
  assign n8058 = n4935 & n6431 ;
  assign n8057 = n3975 & n8054 ;
  assign n8059 = n8058 ^ n8057 ^ 1'b0 ;
  assign n8060 = n2774 & n4270 ;
  assign n8061 = n8060 ^ n7172 ^ 1'b0 ;
  assign n8062 = n7426 & n8061 ;
  assign n8063 = n8062 ^ n3164 ^ 1'b0 ;
  assign n8067 = x244 ^ x9 ^ 1'b0 ;
  assign n8064 = ( n425 & ~n854 ) | ( n425 & n1993 ) | ( ~n854 & n1993 ) ;
  assign n8065 = n1933 ^ n1135 ^ 1'b0 ;
  assign n8066 = n8064 & ~n8065 ;
  assign n8068 = n8067 ^ n8066 ^ 1'b0 ;
  assign n8073 = ( x60 & ~x63 ) | ( x60 & n1937 ) | ( ~x63 & n1937 ) ;
  assign n8072 = n6765 ^ n5887 ^ 1'b0 ;
  assign n8070 = ( ~n496 & n1552 ) | ( ~n496 & n2604 ) | ( n1552 & n2604 ) ;
  assign n8069 = n986 | n6578 ;
  assign n8071 = n8070 ^ n8069 ^ 1'b0 ;
  assign n8074 = n8073 ^ n8072 ^ n8071 ;
  assign n8075 = n676 & n8074 ;
  assign n8076 = n1118 ^ n1114 ^ 1'b0 ;
  assign n8077 = n7264 & ~n8076 ;
  assign n8078 = ~n274 & n7378 ;
  assign n8079 = n8078 ^ n2735 ^ 1'b0 ;
  assign n8080 = n8079 ^ n6359 ^ 1'b0 ;
  assign n8081 = n6978 & ~n8080 ;
  assign n8082 = n1105 & n6745 ;
  assign n8083 = n8082 ^ n1519 ^ n826 ;
  assign n8084 = n7355 ^ n2355 ^ 1'b0 ;
  assign n8085 = n5457 ^ n1775 ^ 1'b0 ;
  assign n8086 = ~n2477 & n2609 ;
  assign n8087 = n8086 ^ n4394 ^ 1'b0 ;
  assign n8088 = n1099 ^ x228 ^ 1'b0 ;
  assign n8089 = n8088 ^ n1950 ^ 1'b0 ;
  assign n8090 = ~n2226 & n8089 ;
  assign n8091 = ~n2024 & n8090 ;
  assign n8092 = n8091 ^ n258 ^ 1'b0 ;
  assign n8093 = n8087 & n8092 ;
  assign n8094 = ~n1213 & n8093 ;
  assign n8095 = n8094 ^ n6278 ^ 1'b0 ;
  assign n8096 = ~n8085 & n8095 ;
  assign n8097 = n5028 ^ n3498 ^ 1'b0 ;
  assign n8098 = ~n1566 & n6112 ;
  assign n8099 = ~n932 & n4218 ;
  assign n8100 = ~n2674 & n8099 ;
  assign n8101 = n8100 ^ n2771 ^ 1'b0 ;
  assign n8103 = ( ~n2027 & n2718 ) | ( ~n2027 & n4656 ) | ( n2718 & n4656 ) ;
  assign n8102 = ~n3102 & n5177 ;
  assign n8104 = n8103 ^ n8102 ^ 1'b0 ;
  assign n8107 = n3012 ^ n425 ^ 1'b0 ;
  assign n8105 = n2732 & n6548 ;
  assign n8106 = ~n3793 & n8105 ;
  assign n8108 = n8107 ^ n8106 ^ 1'b0 ;
  assign n8109 = ~n8104 & n8108 ;
  assign n8110 = ~n2226 & n6574 ;
  assign n8111 = n2123 ^ n638 ^ 1'b0 ;
  assign n8112 = n6716 & n8111 ;
  assign n8113 = n8112 ^ n1726 ^ 1'b0 ;
  assign n8114 = n8113 ^ n6755 ^ n547 ;
  assign n8115 = n4083 ^ n1177 ^ 1'b0 ;
  assign n8116 = n6140 ^ n2839 ^ 1'b0 ;
  assign n8117 = n1699 ^ n1292 ^ 1'b0 ;
  assign n8119 = n4528 ^ n503 ^ 1'b0 ;
  assign n8120 = ~n3761 & n8119 ;
  assign n8121 = n4053 & n8120 ;
  assign n8122 = n4001 & ~n8121 ;
  assign n8123 = n8122 ^ n3064 ^ 1'b0 ;
  assign n8118 = n4248 ^ n3440 ^ x118 ;
  assign n8124 = n8123 ^ n8118 ^ 1'b0 ;
  assign n8125 = n8117 | n8124 ;
  assign n8126 = n3450 & ~n8125 ;
  assign n8127 = ~n4923 & n8126 ;
  assign n8128 = n8116 | n8127 ;
  assign n8129 = n8128 ^ n7009 ^ 1'b0 ;
  assign n8130 = n6856 ^ n3904 ^ 1'b0 ;
  assign n8131 = n5825 ^ n1788 ^ 1'b0 ;
  assign n8132 = ~n312 & n6138 ;
  assign n8133 = ~n2141 & n8132 ;
  assign n8134 = n4612 | n7170 ;
  assign n8135 = n4470 & ~n5089 ;
  assign n8136 = ~n5036 & n5062 ;
  assign n8137 = n2047 | n8136 ;
  assign n8138 = ( n2739 & n4267 ) | ( n2739 & n8022 ) | ( n4267 & n8022 ) ;
  assign n8139 = n395 & ~n3041 ;
  assign n8140 = ~n1344 & n8139 ;
  assign n8141 = n8140 ^ n4085 ^ n3721 ;
  assign n8142 = n8141 ^ n3721 ^ 1'b0 ;
  assign n8143 = n6069 | n8142 ;
  assign n8144 = n813 & ~n4975 ;
  assign n8145 = n8144 ^ n5420 ^ 1'b0 ;
  assign n8146 = ~n466 & n8145 ;
  assign n8147 = n8143 & n8146 ;
  assign n8148 = x173 & ~n3628 ;
  assign n8149 = n8148 ^ n5287 ^ 1'b0 ;
  assign n8150 = n4555 ^ n1346 ^ 1'b0 ;
  assign n8151 = n8150 ^ n2932 ^ 1'b0 ;
  assign n8152 = n449 & n6102 ;
  assign n8153 = n8152 ^ n4261 ^ 1'b0 ;
  assign n8154 = n871 | n7753 ;
  assign n8155 = n1053 | n8154 ;
  assign n8156 = n1261 | n2946 ;
  assign n8157 = n8156 ^ n3223 ^ 1'b0 ;
  assign n8158 = n924 ^ n809 ^ 1'b0 ;
  assign n8159 = ~n2901 & n8158 ;
  assign n8160 = n2218 | n8159 ;
  assign n8161 = n8160 ^ n5177 ^ 1'b0 ;
  assign n8162 = n4767 | n8161 ;
  assign n8163 = n1610 | n3853 ;
  assign n8164 = n8163 ^ n6238 ^ n1815 ;
  assign n8165 = n8041 ^ n4181 ^ 1'b0 ;
  assign n8166 = ( n1926 & n3142 ) | ( n1926 & ~n4460 ) | ( n3142 & ~n4460 ) ;
  assign n8167 = n8166 ^ n1124 ^ 1'b0 ;
  assign n8171 = ~n2501 & n2949 ;
  assign n8172 = n8171 ^ n6822 ^ 1'b0 ;
  assign n8173 = n7325 | n8172 ;
  assign n8174 = n5845 | n8173 ;
  assign n8168 = n1097 ^ n613 ^ 1'b0 ;
  assign n8169 = n1947 & n8168 ;
  assign n8170 = ~n1051 & n8169 ;
  assign n8175 = n8174 ^ n8170 ^ 1'b0 ;
  assign n8176 = n5268 ^ n3823 ^ 1'b0 ;
  assign n8177 = ~n853 & n8176 ;
  assign n8178 = n7110 & n8177 ;
  assign n8179 = n8178 ^ n8118 ^ 1'b0 ;
  assign n8180 = n8175 | n8179 ;
  assign n8184 = n787 | n2872 ;
  assign n8181 = n893 | n5175 ;
  assign n8182 = n2317 | n8181 ;
  assign n8183 = ~n5563 & n8182 ;
  assign n8185 = n8184 ^ n8183 ^ 1'b0 ;
  assign n8186 = n2538 ^ n1333 ^ 1'b0 ;
  assign n8187 = ~n6826 & n8186 ;
  assign n8188 = n4277 & n8187 ;
  assign n8189 = n6986 & n8188 ;
  assign n8190 = ~n4986 & n5046 ;
  assign n8191 = n8190 ^ n2047 ^ 1'b0 ;
  assign n8192 = n2569 & ~n3853 ;
  assign n8193 = n8192 ^ n7838 ^ 1'b0 ;
  assign n8194 = n5246 & n8193 ;
  assign n8195 = n1144 ^ x15 ^ 1'b0 ;
  assign n8196 = n8195 ^ n4611 ^ 1'b0 ;
  assign n8197 = n393 | n4706 ;
  assign n8198 = n5218 & ~n6310 ;
  assign n8199 = n1819 ^ n1365 ^ 1'b0 ;
  assign n8200 = n3879 & ~n8199 ;
  assign n8201 = n8200 ^ n4595 ^ 1'b0 ;
  assign n8202 = n1039 & ~n8201 ;
  assign n8203 = n4219 ^ n4139 ^ 1'b0 ;
  assign n8204 = ~n5911 & n8203 ;
  assign n8205 = n520 & n8204 ;
  assign n8206 = n5782 ^ n5511 ^ 1'b0 ;
  assign n8207 = n2946 | n8206 ;
  assign n8208 = n1919 & n4566 ;
  assign n8209 = n8208 ^ n5390 ^ 1'b0 ;
  assign n8210 = n8209 ^ n2530 ^ 1'b0 ;
  assign n8211 = ( n5815 & ~n6587 ) | ( n5815 & n7371 ) | ( ~n6587 & n7371 ) ;
  assign n8213 = n3359 | n6155 ;
  assign n8214 = n3598 & ~n8213 ;
  assign n8215 = n8214 ^ n3500 ^ n2663 ;
  assign n8216 = n8215 ^ n4708 ^ 1'b0 ;
  assign n8212 = x40 & ~n1492 ;
  assign n8217 = n8216 ^ n8212 ^ 1'b0 ;
  assign n8218 = ~n4493 & n5374 ;
  assign n8219 = n8218 ^ x121 ^ 1'b0 ;
  assign n8221 = x41 & n1989 ;
  assign n8222 = n2045 & n8221 ;
  assign n8220 = n3879 ^ n375 ^ 1'b0 ;
  assign n8223 = n8222 ^ n8220 ^ 1'b0 ;
  assign n8224 = ~n291 & n8223 ;
  assign n8225 = n5388 | n8224 ;
  assign n8226 = n1605 ^ n1219 ^ 1'b0 ;
  assign n8227 = n8226 ^ n7420 ^ 1'b0 ;
  assign n8228 = n8225 & n8227 ;
  assign n8229 = n3776 ^ n3233 ^ 1'b0 ;
  assign n8230 = n2257 & n8229 ;
  assign n8231 = n2830 ^ n1312 ^ 1'b0 ;
  assign n8232 = n729 & ~n8231 ;
  assign n8233 = n8232 ^ n591 ^ 1'b0 ;
  assign n8234 = n6336 ^ n5046 ^ n2798 ;
  assign n8235 = n6613 & n8234 ;
  assign n8236 = x233 | n461 ;
  assign n8237 = n8236 ^ x184 ^ 1'b0 ;
  assign n8238 = n6891 ^ n2845 ^ 1'b0 ;
  assign n8239 = n1474 | n8238 ;
  assign n8240 = ~n2501 & n4325 ;
  assign n8241 = n8240 ^ n3689 ^ 1'b0 ;
  assign n8242 = ~n7538 & n8241 ;
  assign n8243 = ( x20 & n992 ) | ( x20 & ~n3403 ) | ( n992 & ~n3403 ) ;
  assign n8244 = n8243 ^ n5093 ^ 1'b0 ;
  assign n8245 = n2817 & n5770 ;
  assign n8246 = ~n3738 & n8245 ;
  assign n8247 = n694 & ~n8246 ;
  assign n8248 = n8247 ^ n4936 ^ 1'b0 ;
  assign n8249 = ~n757 & n1965 ;
  assign n8250 = n3142 & ~n8249 ;
  assign n8251 = ~n2383 & n2909 ;
  assign n8252 = n6175 ^ n984 ^ 1'b0 ;
  assign n8253 = n8252 ^ n5330 ^ n2316 ;
  assign n8254 = ~n1720 & n4622 ;
  assign n8255 = n8254 ^ n807 ^ 1'b0 ;
  assign n8256 = n267 | n8255 ;
  assign n8257 = n2767 & ~n3205 ;
  assign n8258 = n8256 & n8257 ;
  assign n8259 = n5069 | n8258 ;
  assign n8260 = n8259 ^ n4090 ^ 1'b0 ;
  assign n8261 = ~n2990 & n4966 ;
  assign n8262 = n8261 ^ n3950 ^ 1'b0 ;
  assign n8263 = n3966 & n5152 ;
  assign n8264 = n8263 ^ n2665 ^ 1'b0 ;
  assign n8265 = n4379 ^ n2030 ^ n1528 ;
  assign n8266 = n3576 & ~n7161 ;
  assign n8267 = n8266 ^ n7579 ^ 1'b0 ;
  assign n8268 = n1684 ^ n1083 ^ 1'b0 ;
  assign n8269 = n1475 | n4313 ;
  assign n8270 = n8269 ^ n448 ^ 1'b0 ;
  assign n8271 = n8270 ^ n7779 ^ 1'b0 ;
  assign n8272 = n4109 & n8271 ;
  assign n8273 = n8268 | n8272 ;
  assign n8274 = n6609 ^ n752 ^ 1'b0 ;
  assign n8275 = n1259 | n8274 ;
  assign n8276 = ~n1125 & n8275 ;
  assign n8277 = n3134 ^ n2340 ^ 1'b0 ;
  assign n8278 = n3206 ^ x101 ^ 1'b0 ;
  assign n8279 = n6950 & ~n7753 ;
  assign n8280 = ( n2724 & n6325 ) | ( n2724 & n7825 ) | ( n6325 & n7825 ) ;
  assign n8281 = n8280 ^ n7427 ^ 1'b0 ;
  assign n8282 = n7001 ^ n723 ^ 1'b0 ;
  assign n8283 = n3853 & ~n8249 ;
  assign n8284 = n8282 & n8283 ;
  assign n8285 = n8284 ^ n629 ^ 1'b0 ;
  assign n8286 = n3614 & n8285 ;
  assign n8287 = n684 | n6713 ;
  assign n8288 = ~n2338 & n2514 ;
  assign n8289 = ~n4380 & n8288 ;
  assign n8290 = n6443 ^ n1442 ^ 1'b0 ;
  assign n8291 = n5626 & n8290 ;
  assign n8294 = n3840 ^ n2624 ^ 1'b0 ;
  assign n8295 = ~n3179 & n8294 ;
  assign n8296 = n8295 ^ n4266 ^ 1'b0 ;
  assign n8297 = n634 | n8296 ;
  assign n8292 = x154 & x237 ;
  assign n8293 = ~n3518 & n8292 ;
  assign n8298 = n8297 ^ n8293 ^ 1'b0 ;
  assign n8301 = n1230 & ~n1617 ;
  assign n8299 = n4542 | n5387 ;
  assign n8300 = n4733 | n8299 ;
  assign n8302 = n8301 ^ n8300 ^ 1'b0 ;
  assign n8303 = ~n917 & n1272 ;
  assign n8305 = n6581 ^ n3511 ^ 1'b0 ;
  assign n8306 = n8305 ^ n5295 ^ 1'b0 ;
  assign n8307 = n917 & n8306 ;
  assign n8304 = n1484 ^ n1293 ^ 1'b0 ;
  assign n8308 = n8307 ^ n8304 ^ x91 ;
  assign n8309 = ( n847 & n4368 ) | ( n847 & n8094 ) | ( n4368 & n8094 ) ;
  assign n8310 = n7392 & n8309 ;
  assign n8311 = n3589 & n8310 ;
  assign n8312 = n2644 & ~n6015 ;
  assign n8315 = n2651 | n3423 ;
  assign n8313 = n4693 ^ n3770 ^ 1'b0 ;
  assign n8314 = n8293 | n8313 ;
  assign n8316 = n8315 ^ n8314 ^ 1'b0 ;
  assign n8317 = n2868 | n8316 ;
  assign n8318 = n6233 ^ n446 ^ 1'b0 ;
  assign n8319 = n2569 | n8318 ;
  assign n8320 = x59 & ~n552 ;
  assign n8321 = ~x147 & n8320 ;
  assign n8322 = n4594 | n8321 ;
  assign n8323 = n8319 | n8322 ;
  assign n8324 = n6069 ^ n5208 ^ 1'b0 ;
  assign n8325 = n3956 | n8324 ;
  assign n8326 = x70 | n988 ;
  assign n8327 = ( ~x193 & n7089 ) | ( ~x193 & n8326 ) | ( n7089 & n8326 ) ;
  assign n8328 = n3272 ^ n3028 ^ 1'b0 ;
  assign n8329 = n6398 ^ n5864 ^ 1'b0 ;
  assign n8330 = ~n7650 & n8329 ;
  assign n8331 = n6094 ^ n2497 ^ n1148 ;
  assign n8332 = n8331 ^ n1749 ^ n581 ;
  assign n8333 = n8332 ^ n7496 ^ 1'b0 ;
  assign n8336 = ( n420 & n1841 ) | ( n420 & ~n7028 ) | ( n1841 & ~n7028 ) ;
  assign n8337 = n8336 ^ n3249 ^ 1'b0 ;
  assign n8338 = ~n4438 & n8337 ;
  assign n8339 = n8338 ^ n4741 ^ 1'b0 ;
  assign n8334 = n894 & n995 ;
  assign n8335 = n5829 | n8334 ;
  assign n8340 = n8339 ^ n8335 ^ 1'b0 ;
  assign n8341 = n1837 & ~n4439 ;
  assign n8342 = n8341 ^ n8141 ^ 1'b0 ;
  assign n8343 = n7359 ^ n925 ^ 1'b0 ;
  assign n8344 = n7766 & ~n8343 ;
  assign n8345 = n713 & n8344 ;
  assign n8346 = n8345 ^ n1432 ^ 1'b0 ;
  assign n8347 = n733 | n2615 ;
  assign n8348 = n5401 | n8347 ;
  assign n8349 = n8348 ^ n7851 ^ 1'b0 ;
  assign n8350 = ~n5492 & n8349 ;
  assign n8351 = n8350 ^ n7584 ^ 1'b0 ;
  assign n8352 = n4380 ^ n655 ^ 1'b0 ;
  assign n8353 = n6327 ^ n596 ^ 1'b0 ;
  assign n8354 = ~n8352 & n8353 ;
  assign n8357 = n2739 ^ x13 ^ 1'b0 ;
  assign n8358 = ~n5864 & n8357 ;
  assign n8355 = n3038 ^ n1147 ^ 1'b0 ;
  assign n8356 = n8355 ^ n5259 ^ 1'b0 ;
  assign n8359 = n8358 ^ n8356 ^ n308 ;
  assign n8360 = n3313 & ~n7674 ;
  assign n8361 = n8360 ^ n7929 ^ 1'b0 ;
  assign n8362 = n627 | n8361 ;
  assign n8365 = n6978 ^ n6451 ^ n4377 ;
  assign n8363 = n1360 | n7592 ;
  assign n8364 = n3332 | n8363 ;
  assign n8366 = n8365 ^ n8364 ^ 1'b0 ;
  assign n8367 = ~n8362 & n8366 ;
  assign n8368 = n8367 ^ n2587 ^ 1'b0 ;
  assign n8369 = x221 & n1154 ;
  assign n8370 = n5027 ^ n4790 ^ 1'b0 ;
  assign n8371 = n3554 | n8370 ;
  assign n8372 = n1437 | n8371 ;
  assign n8373 = n8372 ^ n2999 ^ 1'b0 ;
  assign n8374 = x133 & n556 ;
  assign n8375 = ~x62 & n8374 ;
  assign n8376 = n2726 | n8375 ;
  assign n8377 = n8376 ^ n4379 ^ 1'b0 ;
  assign n8378 = n5667 | n8377 ;
  assign n8379 = n8378 ^ x77 ^ 1'b0 ;
  assign n8380 = n7389 | n8379 ;
  assign n8381 = n8380 ^ n5896 ^ 1'b0 ;
  assign n8382 = n3474 & ~n7087 ;
  assign n8383 = n4972 | n8382 ;
  assign n8384 = n4593 & ~n8383 ;
  assign n8389 = n2164 ^ n1321 ^ 1'b0 ;
  assign n8390 = n272 & ~n8389 ;
  assign n8385 = n1814 & ~n3145 ;
  assign n8386 = ~n5544 & n8385 ;
  assign n8387 = n4675 ^ n2618 ^ 1'b0 ;
  assign n8388 = n8386 | n8387 ;
  assign n8391 = n8390 ^ n8388 ^ x96 ;
  assign n8392 = ~n6928 & n8391 ;
  assign n8393 = n2741 & n8392 ;
  assign n8394 = n713 & n5746 ;
  assign n8395 = ~x100 & n8394 ;
  assign n8396 = n7260 | n8395 ;
  assign n8397 = n8396 ^ n3313 ^ n903 ;
  assign n8398 = n6206 ^ n270 ^ 1'b0 ;
  assign n8399 = n344 | n8398 ;
  assign n8400 = n5750 ^ n529 ^ 1'b0 ;
  assign n8401 = n7670 & n8400 ;
  assign n8402 = n4867 & ~n5921 ;
  assign n8403 = ~n8401 & n8402 ;
  assign n8404 = n4920 | n6385 ;
  assign n8405 = n8404 ^ n1078 ^ 1'b0 ;
  assign n8406 = n453 & n8405 ;
  assign n8407 = ~n1525 & n8406 ;
  assign n8408 = n8407 ^ n2465 ^ 1'b0 ;
  assign n8409 = ~n1480 & n4095 ;
  assign n8410 = ~n5180 & n8409 ;
  assign n8411 = n8410 ^ n2633 ^ n1664 ;
  assign n8412 = ~n1467 & n3321 ;
  assign n8413 = n7185 & n8412 ;
  assign n8414 = n5606 ^ n3500 ^ n1903 ;
  assign n8415 = n3837 ^ n2745 ^ x157 ;
  assign n8416 = x119 & ~n1657 ;
  assign n8417 = ~n756 & n8416 ;
  assign n8418 = n879 & ~n8417 ;
  assign n8419 = n4875 | n8418 ;
  assign n8420 = n1220 & n6102 ;
  assign n8421 = n8420 ^ n3179 ^ 1'b0 ;
  assign n8422 = n4501 | n5403 ;
  assign n8423 = x216 ^ x59 ^ 1'b0 ;
  assign n8425 = n1284 | n3791 ;
  assign n8424 = n6062 ^ n357 ^ 1'b0 ;
  assign n8426 = n8425 ^ n8424 ^ n4003 ;
  assign n8427 = n5087 ^ n2988 ^ 1'b0 ;
  assign n8428 = n6739 & n8427 ;
  assign n8429 = ~n548 & n2984 ;
  assign n8430 = ~n7907 & n8429 ;
  assign n8431 = n2189 ^ n853 ^ 1'b0 ;
  assign n8432 = n778 & ~n3413 ;
  assign n8433 = n4264 & ~n8432 ;
  assign n8434 = n5079 & n8433 ;
  assign n8435 = n3248 & ~n8377 ;
  assign n8436 = n2401 & n2688 ;
  assign n8437 = n8436 ^ n7714 ^ 1'b0 ;
  assign n8438 = x153 & n8437 ;
  assign n8439 = n2027 | n2472 ;
  assign n8440 = n6413 & ~n8439 ;
  assign n8441 = n271 & n3620 ;
  assign n8442 = n8441 ^ n6020 ^ 1'b0 ;
  assign n8443 = n1230 & n8442 ;
  assign n8444 = n8440 & n8443 ;
  assign n8445 = x23 & ~n374 ;
  assign n8446 = n8445 ^ n2282 ^ 1'b0 ;
  assign n8447 = n618 ^ n300 ^ 1'b0 ;
  assign n8448 = n2127 ^ n1575 ^ 1'b0 ;
  assign n8449 = n8447 & n8448 ;
  assign n8450 = n8446 & n8449 ;
  assign n8451 = n1935 & n3665 ;
  assign n8452 = n8451 ^ n3576 ^ 1'b0 ;
  assign n8453 = n2183 & n2516 ;
  assign n8454 = n8453 ^ x20 ^ 1'b0 ;
  assign n8455 = n8454 ^ n6966 ^ x3 ;
  assign n8456 = ( n6561 & n8145 ) | ( n6561 & n8455 ) | ( n8145 & n8455 ) ;
  assign n8457 = n6122 ^ n2121 ^ n1727 ;
  assign n8458 = n1694 | n7029 ;
  assign n8459 = n8457 & ~n8458 ;
  assign n8460 = n7848 ^ n2538 ^ 1'b0 ;
  assign n8461 = n5642 ^ n3952 ^ 1'b0 ;
  assign n8462 = n4679 & ~n8461 ;
  assign n8463 = x64 | n6088 ;
  assign n8464 = n2073 & ~n8463 ;
  assign n8465 = n8464 ^ n1547 ^ 1'b0 ;
  assign n8466 = ~n5896 & n8117 ;
  assign n8467 = ~n8465 & n8466 ;
  assign n8468 = n6817 | n8467 ;
  assign n8470 = n3108 ^ n2144 ^ 1'b0 ;
  assign n8471 = ( n4851 & ~n8159 ) | ( n4851 & n8470 ) | ( ~n8159 & n8470 ) ;
  assign n8472 = n5909 & n8471 ;
  assign n8473 = n8472 ^ x153 ^ 1'b0 ;
  assign n8469 = n1714 | n4868 ;
  assign n8474 = n8473 ^ n8469 ^ 1'b0 ;
  assign n8475 = ( ~n1801 & n7524 ) | ( ~n1801 & n8474 ) | ( n7524 & n8474 ) ;
  assign n8476 = ( n1497 & n2027 ) | ( n1497 & ~n6609 ) | ( n2027 & ~n6609 ) ;
  assign n8477 = n6062 ^ n3451 ^ 1'b0 ;
  assign n8478 = n8476 | n8477 ;
  assign n8479 = n346 & ~n8478 ;
  assign n8480 = n5269 ^ n4645 ^ 1'b0 ;
  assign n8481 = n1091 & n8480 ;
  assign n8482 = n3041 & n5885 ;
  assign n8483 = ~n466 & n488 ;
  assign n8484 = x132 & ~n450 ;
  assign n8485 = n6728 & n8484 ;
  assign n8487 = n699 & ~n1147 ;
  assign n8486 = n2167 & ~n4381 ;
  assign n8488 = n8487 ^ n8486 ^ 1'b0 ;
  assign n8489 = ( n645 & n1480 ) | ( n645 & ~n3686 ) | ( n1480 & ~n3686 ) ;
  assign n8490 = ~n7157 & n8000 ;
  assign n8491 = n3644 | n8303 ;
  assign n8492 = n2715 | n2960 ;
  assign n8493 = n5667 | n8492 ;
  assign n8494 = n3614 & n3684 ;
  assign n8495 = n8494 ^ n2841 ^ 1'b0 ;
  assign n8496 = n5896 ^ n5016 ^ 1'b0 ;
  assign n8497 = n2694 & ~n8496 ;
  assign n8498 = ~n8495 & n8497 ;
  assign n8499 = n4380 ^ n3845 ^ 1'b0 ;
  assign n8500 = n8499 ^ n2613 ^ 1'b0 ;
  assign n8501 = n4701 | n8500 ;
  assign n8502 = n8501 ^ n6542 ^ n3209 ;
  assign n8503 = n4255 & n4474 ;
  assign n8504 = n4360 & ~n8284 ;
  assign n8505 = ( n2051 & n3160 ) | ( n2051 & ~n3674 ) | ( n3160 & ~n3674 ) ;
  assign n8506 = n8505 ^ n7264 ^ n2697 ;
  assign n8507 = n906 & n8201 ;
  assign n8508 = n8507 ^ n905 ^ 1'b0 ;
  assign n8509 = n2740 & ~n8508 ;
  assign n8510 = n5763 & n8509 ;
  assign n8511 = n4271 ^ n457 ^ 1'b0 ;
  assign n8512 = n1643 & ~n8511 ;
  assign n8513 = n6284 | n8512 ;
  assign n8514 = n8513 ^ x251 ^ 1'b0 ;
  assign n8515 = n3028 ^ n434 ^ 1'b0 ;
  assign n8516 = n6310 ^ n2263 ^ 1'b0 ;
  assign n8517 = n1345 | n8516 ;
  assign n8518 = n2023 | n4076 ;
  assign n8519 = n8518 ^ n6331 ^ 1'b0 ;
  assign n8520 = n6957 ^ n4861 ^ n819 ;
  assign n8521 = n2428 ^ n1393 ^ 1'b0 ;
  assign n8522 = ~n1894 & n8521 ;
  assign n8523 = n8522 ^ n4144 ^ 1'b0 ;
  assign n8524 = n7140 & ~n8523 ;
  assign n8525 = n6116 ^ n6033 ^ n1402 ;
  assign n8526 = n6868 | n8525 ;
  assign n8527 = n8526 ^ n6754 ^ 1'b0 ;
  assign n8528 = x50 & n2319 ;
  assign n8529 = n8528 ^ n6866 ^ 1'b0 ;
  assign n8530 = n1933 | n8529 ;
  assign n8531 = ( n433 & ~n6947 ) | ( n433 & n7600 ) | ( ~n6947 & n7600 ) ;
  assign n8532 = n6211 | n8531 ;
  assign n8533 = n618 & n1977 ;
  assign n8534 = n8533 ^ n619 ^ 1'b0 ;
  assign n8535 = n8534 ^ n2949 ^ 1'b0 ;
  assign n8536 = n3177 ^ n2450 ^ 1'b0 ;
  assign n8537 = n5531 & n6918 ;
  assign n8538 = ~n8536 & n8537 ;
  assign n8539 = n8538 ^ n2948 ^ 1'b0 ;
  assign n8540 = n921 & ~n8539 ;
  assign n8541 = n4341 ^ n2215 ^ n1160 ;
  assign n8542 = n3168 & n8541 ;
  assign n8543 = n8542 ^ n2715 ^ 1'b0 ;
  assign n8544 = n7112 ^ n2623 ^ 1'b0 ;
  assign n8545 = n3525 & n8544 ;
  assign n8546 = n1120 & n5408 ;
  assign n8547 = x42 & n1347 ;
  assign n8548 = ( x137 & n4038 ) | ( x137 & ~n4976 ) | ( n4038 & ~n4976 ) ;
  assign n8549 = n5803 & ~n8548 ;
  assign n8550 = n6782 & n8549 ;
  assign n8551 = n4977 ^ n1741 ^ n1575 ;
  assign n8552 = ~n5925 & n8551 ;
  assign n8553 = n8552 ^ n3806 ^ n1862 ;
  assign n8554 = n2798 & n3100 ;
  assign n8555 = n4252 & n8554 ;
  assign n8556 = ~n3686 & n8555 ;
  assign n8557 = ~n6157 & n7813 ;
  assign n8558 = n4964 & ~n7445 ;
  assign n8559 = n8258 ^ n1820 ^ 1'b0 ;
  assign n8560 = n505 | n5316 ;
  assign n8561 = n5195 & ~n8560 ;
  assign n8562 = n1340 | n4848 ;
  assign n8563 = n4848 & ~n8562 ;
  assign n8564 = ~n5505 & n7238 ;
  assign n8565 = ( n8058 & ~n8563 ) | ( n8058 & n8564 ) | ( ~n8563 & n8564 ) ;
  assign n8566 = n1973 ^ x186 ^ 1'b0 ;
  assign n8567 = n459 & n604 ;
  assign n8568 = ~n8566 & n8567 ;
  assign n8569 = n8568 ^ n4913 ^ 1'b0 ;
  assign n8570 = ~n6265 & n8569 ;
  assign n8571 = ~n1426 & n7742 ;
  assign n8572 = ( n4639 & n4839 ) | ( n4639 & n8571 ) | ( n4839 & n8571 ) ;
  assign n8573 = n8572 ^ n3588 ^ 1'b0 ;
  assign n8574 = n1281 ^ n997 ^ 1'b0 ;
  assign n8580 = n2286 & ~n8073 ;
  assign n8581 = ( x225 & ~n4447 ) | ( x225 & n8580 ) | ( ~n4447 & n8580 ) ;
  assign n8576 = n3180 | n8446 ;
  assign n8577 = n2369 | n8576 ;
  assign n8575 = n2396 & ~n7293 ;
  assign n8578 = n8577 ^ n8575 ^ 1'b0 ;
  assign n8579 = n2957 | n8578 ;
  assign n8582 = n8581 ^ n8579 ^ 1'b0 ;
  assign n8583 = n1554 & n2949 ;
  assign n8584 = n2781 | n8583 ;
  assign n8585 = n6206 ^ n4867 ^ 1'b0 ;
  assign n8586 = n572 & ~n1731 ;
  assign n8587 = n8586 ^ n1851 ^ 1'b0 ;
  assign n8588 = x68 & n6877 ;
  assign n8589 = ~n3440 & n8588 ;
  assign n8590 = ~n882 & n2360 ;
  assign n8591 = n8590 ^ n1810 ^ 1'b0 ;
  assign n8592 = x57 | n8591 ;
  assign n8593 = n8592 ^ n3345 ^ 1'b0 ;
  assign n8594 = n8589 | n8593 ;
  assign n8595 = ~n8587 & n8594 ;
  assign n8596 = x3 & n8595 ;
  assign n8597 = n2215 & n8596 ;
  assign n8598 = n3405 ^ x2 ^ 1'b0 ;
  assign n8599 = n3873 & ~n6632 ;
  assign n8600 = n5912 & n8599 ;
  assign n8601 = n8598 | n8600 ;
  assign n8602 = n8601 ^ n2467 ^ 1'b0 ;
  assign n8603 = n2509 & n3568 ;
  assign n8604 = n8603 ^ n7183 ^ 1'b0 ;
  assign n8605 = n8471 ^ x49 ^ 1'b0 ;
  assign n8606 = n4552 ^ n4380 ^ n3023 ;
  assign n8607 = n3637 ^ n2502 ^ 1'b0 ;
  assign n8608 = n732 & ~n8607 ;
  assign n8609 = ~n2482 & n8608 ;
  assign n8610 = n2110 & n5659 ;
  assign n8611 = n1471 ^ n1319 ^ 1'b0 ;
  assign n8612 = n2964 & ~n8611 ;
  assign n8613 = ~n2202 & n8612 ;
  assign n8614 = n7724 ^ n4509 ^ 1'b0 ;
  assign n8615 = ~n5856 & n7409 ;
  assign n8616 = ~n3001 & n8615 ;
  assign n8617 = n688 & n8341 ;
  assign n8618 = n8617 ^ n7749 ^ 1'b0 ;
  assign n8619 = n2135 ^ n455 ^ 1'b0 ;
  assign n8620 = n4600 | n8619 ;
  assign n8621 = n1969 | n8620 ;
  assign n8622 = n2978 | n8621 ;
  assign n8623 = ~n4045 & n5508 ;
  assign n8624 = ~n5325 & n8623 ;
  assign n8625 = n7077 ^ n2622 ^ 1'b0 ;
  assign n8626 = n2180 & n3397 ;
  assign n8627 = n2428 | n5775 ;
  assign n8628 = n8627 ^ n8591 ^ 1'b0 ;
  assign n8629 = n1379 & n8628 ;
  assign n8635 = ~n2321 & n6707 ;
  assign n8636 = n1651 & n8635 ;
  assign n8637 = n8636 ^ n2829 ^ 1'b0 ;
  assign n8638 = n4458 & n8637 ;
  assign n8631 = n796 & n1249 ;
  assign n8632 = n8100 & n8631 ;
  assign n8630 = n765 | n3938 ;
  assign n8633 = n8632 ^ n8630 ^ n6437 ;
  assign n8634 = ~n4568 & n8633 ;
  assign n8639 = n8638 ^ n8634 ^ 1'b0 ;
  assign n8640 = n1535 & ~n4409 ;
  assign n8641 = ~n2133 & n8640 ;
  assign n8644 = n587 | n804 ;
  assign n8645 = n3467 | n8644 ;
  assign n8642 = n708 & ~n7209 ;
  assign n8643 = n8552 & ~n8642 ;
  assign n8646 = n8645 ^ n8643 ^ 1'b0 ;
  assign n8647 = n4273 ^ n4165 ^ 1'b0 ;
  assign n8648 = ~n1244 & n2868 ;
  assign n8649 = n8648 ^ n3729 ^ 1'b0 ;
  assign n8650 = n8649 ^ n5479 ^ 1'b0 ;
  assign n8651 = n682 | n8650 ;
  assign n8652 = n6824 ^ n3670 ^ 1'b0 ;
  assign n8653 = n3558 | n8652 ;
  assign n8654 = x7 & ~n3539 ;
  assign n8655 = n8654 ^ n2276 ^ 1'b0 ;
  assign n8656 = ~n716 & n8655 ;
  assign n8657 = n4352 | n8656 ;
  assign n8658 = n8529 ^ n5900 ^ 1'b0 ;
  assign n8659 = n8015 ^ n7105 ^ 1'b0 ;
  assign n8661 = ~x13 & n318 ;
  assign n8662 = n1775 & n8661 ;
  assign n8660 = n631 ^ x213 ^ 1'b0 ;
  assign n8663 = n8662 ^ n8660 ^ 1'b0 ;
  assign n8664 = ~n963 & n3293 ;
  assign n8665 = n548 | n2098 ;
  assign n8666 = n6116 ^ n3180 ^ n3023 ;
  assign n8667 = n4516 | n8666 ;
  assign n8668 = n8667 ^ n5089 ^ n1626 ;
  assign n8669 = ~n8665 & n8668 ;
  assign n8670 = n8669 ^ n8627 ^ 1'b0 ;
  assign n8671 = n4285 | n5839 ;
  assign n8672 = n8671 ^ n1980 ^ 1'b0 ;
  assign n8673 = n2306 | n8672 ;
  assign n8675 = n3493 ^ x50 ^ 1'b0 ;
  assign n8676 = ~n1321 & n8675 ;
  assign n8674 = n5848 ^ n2584 ^ 1'b0 ;
  assign n8677 = n8676 ^ n8674 ^ 1'b0 ;
  assign n8678 = n1197 | n6203 ;
  assign n8679 = ~n7530 & n7815 ;
  assign n8680 = n7657 ^ n2787 ^ 1'b0 ;
  assign n8681 = n2959 & n8680 ;
  assign n8682 = n8660 ^ n917 ^ 1'b0 ;
  assign n8683 = n7058 & n8682 ;
  assign n8684 = n5187 ^ n2998 ^ 1'b0 ;
  assign n8685 = n274 ^ x70 ^ 1'b0 ;
  assign n8686 = n8685 ^ n6340 ^ 1'b0 ;
  assign n8687 = n8684 & n8686 ;
  assign n8689 = x160 & x211 ;
  assign n8690 = n2638 & n8689 ;
  assign n8688 = n2101 | n4425 ;
  assign n8691 = n8690 ^ n8688 ^ 1'b0 ;
  assign n8692 = n6854 ^ n6470 ^ 1'b0 ;
  assign n8693 = n1690 | n8692 ;
  assign n8694 = ~n733 & n8378 ;
  assign n8695 = n2011 & ~n2944 ;
  assign n8696 = n1801 | n4333 ;
  assign n8697 = n8696 ^ n2289 ^ 1'b0 ;
  assign n8698 = n8697 ^ n346 ^ 1'b0 ;
  assign n8699 = n4367 ^ n1884 ^ n421 ;
  assign n8700 = n8699 ^ n3631 ^ n1521 ;
  assign n8701 = n7224 ^ n527 ^ 1'b0 ;
  assign n8702 = n6496 & ~n8701 ;
  assign n8709 = n4906 ^ n4747 ^ n3915 ;
  assign n8703 = n7549 ^ n3288 ^ 1'b0 ;
  assign n8704 = n1395 & n8703 ;
  assign n8705 = n3317 & n8704 ;
  assign n8706 = n5703 ^ n722 ^ 1'b0 ;
  assign n8707 = ~n2730 & n8706 ;
  assign n8708 = ~n8705 & n8707 ;
  assign n8710 = n8709 ^ n8708 ^ 1'b0 ;
  assign n8716 = x125 & x226 ;
  assign n8717 = n8716 ^ n1047 ^ 1'b0 ;
  assign n8718 = n2054 | n8717 ;
  assign n8713 = n3648 ^ n954 ^ 1'b0 ;
  assign n8711 = n5928 & ~n6684 ;
  assign n8712 = n8711 ^ n4474 ^ 1'b0 ;
  assign n8714 = n8713 ^ n8712 ^ n973 ;
  assign n8715 = n8714 ^ n8209 ^ n6043 ;
  assign n8719 = n8718 ^ n8715 ^ 1'b0 ;
  assign n8720 = n1548 & ~n8719 ;
  assign n8721 = n6842 ^ n3757 ^ 1'b0 ;
  assign n8722 = n1283 | n8721 ;
  assign n8723 = n1854 ^ x238 ^ 1'b0 ;
  assign n8724 = n1165 & ~n4045 ;
  assign n8725 = n2718 ^ x92 ^ 1'b0 ;
  assign n8726 = ( x37 & ~n7273 ) | ( x37 & n8725 ) | ( ~n7273 & n8725 ) ;
  assign n8727 = n1312 & ~n3074 ;
  assign n8728 = ~n5616 & n8727 ;
  assign n8729 = n8186 | n8728 ;
  assign n8730 = n481 | n4369 ;
  assign n8731 = n8730 ^ n7952 ^ n3230 ;
  assign n8732 = n3233 & ~n5088 ;
  assign n8733 = n8732 ^ x226 ^ 1'b0 ;
  assign n8734 = n1583 & n8733 ;
  assign n8735 = n714 & n8734 ;
  assign n8736 = ~n1841 & n2239 ;
  assign n8737 = n2895 | n8736 ;
  assign n8738 = n8737 ^ n2015 ^ 1'b0 ;
  assign n8739 = n2924 | n8738 ;
  assign n8740 = n5734 ^ n3297 ^ 1'b0 ;
  assign n8741 = n1550 | n7536 ;
  assign n8742 = n3666 | n8741 ;
  assign n8743 = n1611 ^ n904 ^ 1'b0 ;
  assign n8744 = n1903 & n8743 ;
  assign n8745 = n5587 & n8744 ;
  assign n8746 = n2819 & n7846 ;
  assign n8747 = ( n865 & ~n4896 ) | ( n865 & n8011 ) | ( ~n4896 & n8011 ) ;
  assign n8748 = ~n8746 & n8747 ;
  assign n8749 = n8748 ^ n8735 ^ 1'b0 ;
  assign n8750 = n756 ^ x63 ^ 1'b0 ;
  assign n8751 = ~n2560 & n8750 ;
  assign n8752 = ( n1404 & n1824 ) | ( n1404 & n8751 ) | ( n1824 & n8751 ) ;
  assign n8753 = n8752 ^ n1950 ^ 1'b0 ;
  assign n8754 = ~n2831 & n8753 ;
  assign n8755 = n4844 ^ n2706 ^ 1'b0 ;
  assign n8756 = n4220 & n4258 ;
  assign n8759 = n4750 ^ x152 ^ 1'b0 ;
  assign n8760 = n3206 ^ n935 ^ 1'b0 ;
  assign n8761 = n2140 ^ n752 ^ 1'b0 ;
  assign n8762 = n8760 & n8761 ;
  assign n8763 = ( n5286 & ~n8759 ) | ( n5286 & n8762 ) | ( ~n8759 & n8762 ) ;
  assign n8757 = n5025 ^ n4622 ^ 1'b0 ;
  assign n8758 = n6991 | n8757 ;
  assign n8764 = n8763 ^ n8758 ^ n2249 ;
  assign n8765 = n5154 ^ n4871 ^ n4540 ;
  assign n8766 = n8765 ^ n2310 ^ 1'b0 ;
  assign n8767 = n3626 ^ n2954 ^ 1'b0 ;
  assign n8768 = ~n1075 & n8767 ;
  assign n8769 = x249 & n8768 ;
  assign n8770 = n8769 ^ n1387 ^ 1'b0 ;
  assign n8771 = ~n1728 & n7617 ;
  assign n8772 = n4890 & ~n8771 ;
  assign n8773 = n5831 ^ n5325 ^ 1'b0 ;
  assign n8774 = n5973 & n8773 ;
  assign n8775 = n1356 & n1926 ;
  assign n8776 = ~n1541 & n8775 ;
  assign n8777 = n1509 & n8776 ;
  assign n8778 = ( n2356 & n3537 ) | ( n2356 & n7979 ) | ( n3537 & n7979 ) ;
  assign n8779 = n6140 ^ n917 ^ 1'b0 ;
  assign n8780 = n2856 & ~n8779 ;
  assign n8781 = ~n5884 & n7588 ;
  assign n8782 = n5746 ^ n1749 ^ 1'b0 ;
  assign n8783 = ~n5630 & n8782 ;
  assign n8784 = ( ~n8315 & n8781 ) | ( ~n8315 & n8783 ) | ( n8781 & n8783 ) ;
  assign n8785 = n1180 & n2131 ;
  assign n8786 = ( n4172 & n8352 ) | ( n4172 & n8785 ) | ( n8352 & n8785 ) ;
  assign n8787 = n8786 ^ x247 ^ 1'b0 ;
  assign n8788 = n8784 & n8787 ;
  assign n8789 = ( n1432 & ~n6017 ) | ( n1432 & n7538 ) | ( ~n6017 & n7538 ) ;
  assign n8792 = n897 ^ x77 ^ 1'b0 ;
  assign n8793 = n8792 ^ n5536 ^ n3035 ;
  assign n8790 = x176 & n4313 ;
  assign n8791 = n8790 ^ n5551 ^ 1'b0 ;
  assign n8794 = n8793 ^ n8791 ^ n6900 ;
  assign n8795 = n3551 ^ n1180 ^ 1'b0 ;
  assign n8796 = ~n393 & n8795 ;
  assign n8797 = n4279 & ~n5735 ;
  assign n8798 = ~n8351 & n8797 ;
  assign n8799 = n1788 ^ n1698 ^ n1611 ;
  assign n8800 = ~n498 & n2609 ;
  assign n8801 = n8800 ^ n5047 ^ 1'b0 ;
  assign n8802 = n4117 & ~n8801 ;
  assign n8804 = ( n387 & n2788 ) | ( n387 & ~n5054 ) | ( n2788 & ~n5054 ) ;
  assign n8803 = n3044 & ~n7626 ;
  assign n8805 = n8804 ^ n8803 ^ 1'b0 ;
  assign n8806 = n2919 | n8805 ;
  assign n8807 = n1596 | n7592 ;
  assign n8808 = x116 & n4014 ;
  assign n8809 = n8808 ^ n1799 ^ 1'b0 ;
  assign n8810 = n1989 & n8809 ;
  assign n8811 = n8810 ^ n5913 ^ 1'b0 ;
  assign n8812 = n5238 ^ n3145 ^ 1'b0 ;
  assign n8813 = ~n2755 & n8812 ;
  assign n8814 = n8813 ^ n4876 ^ 1'b0 ;
  assign n8815 = x89 & ~n3228 ;
  assign n8816 = n8815 ^ n7462 ^ 1'b0 ;
  assign n8817 = ~n1198 & n8418 ;
  assign n8818 = n3670 & n8817 ;
  assign n8819 = n3288 | n7214 ;
  assign n8820 = n8818 & ~n8819 ;
  assign n8821 = ~n1261 & n6604 ;
  assign n8822 = n389 | n2281 ;
  assign n8823 = n1306 | n8822 ;
  assign n8824 = n7409 & ~n8823 ;
  assign n8825 = ( x14 & n8821 ) | ( x14 & n8824 ) | ( n8821 & n8824 ) ;
  assign n8826 = n3462 ^ n2056 ^ 1'b0 ;
  assign n8827 = n583 | n8826 ;
  assign n8828 = n4423 & ~n4793 ;
  assign n8829 = n8827 & n8828 ;
  assign n8830 = n3912 ^ n587 ^ 1'b0 ;
  assign n8831 = n2448 ^ n1680 ^ 1'b0 ;
  assign n8832 = n8831 ^ n3012 ^ 1'b0 ;
  assign n8833 = n8735 & ~n8832 ;
  assign n8834 = n6155 & n8833 ;
  assign n8835 = n2450 ^ n2187 ^ 1'b0 ;
  assign n8836 = n2582 ^ n2170 ^ 1'b0 ;
  assign n8837 = n8835 & ~n8836 ;
  assign n8838 = n992 & ~n3901 ;
  assign n8839 = ~n6748 & n8838 ;
  assign n8840 = n5535 ^ n498 ^ 1'b0 ;
  assign n8841 = n4571 | n8840 ;
  assign n8842 = n2929 & n4342 ;
  assign n8843 = x176 ^ x154 ^ 1'b0 ;
  assign n8844 = ~n550 & n8843 ;
  assign n8845 = n4347 | n6095 ;
  assign n8846 = n8845 ^ n1137 ^ 1'b0 ;
  assign n8847 = n1264 | n8846 ;
  assign n8848 = n8844 | n8847 ;
  assign n8849 = n8842 | n8848 ;
  assign n8850 = n5616 ^ n699 ^ 1'b0 ;
  assign n8851 = n1147 & ~n8850 ;
  assign n8852 = n2452 ^ x81 ^ 1'b0 ;
  assign n8853 = n7018 & ~n8852 ;
  assign n8854 = ~n1374 & n5646 ;
  assign n8855 = n8854 ^ n3367 ^ 1'b0 ;
  assign n8856 = n8855 ^ n6949 ^ n5494 ;
  assign n8857 = ( n3293 & n8853 ) | ( n3293 & n8856 ) | ( n8853 & n8856 ) ;
  assign n8858 = n5775 ^ n617 ^ 1'b0 ;
  assign n8859 = n8858 ^ n3959 ^ 1'b0 ;
  assign n8860 = n8859 ^ n6803 ^ n3174 ;
  assign n8861 = ( n2589 & n4552 ) | ( n2589 & ~n6095 ) | ( n4552 & ~n6095 ) ;
  assign n8862 = n8861 ^ n5473 ^ 1'b0 ;
  assign n8863 = n1725 | n3309 ;
  assign n8864 = n8141 & ~n8863 ;
  assign n8865 = n6933 ^ n1995 ^ 1'b0 ;
  assign n8866 = n6668 ^ n4913 ^ 1'b0 ;
  assign n8867 = n1611 & n3296 ;
  assign n8868 = ~n2531 & n8867 ;
  assign n8876 = n4416 ^ n2666 ^ 1'b0 ;
  assign n8877 = n7247 | n8876 ;
  assign n8869 = ( n2567 & n2682 ) | ( n2567 & n7368 ) | ( n2682 & n7368 ) ;
  assign n8870 = ( n490 & ~n1739 ) | ( n490 & n6529 ) | ( ~n1739 & n6529 ) ;
  assign n8871 = n8870 ^ n4067 ^ 1'b0 ;
  assign n8872 = ~n1402 & n8871 ;
  assign n8873 = n4242 & n8872 ;
  assign n8874 = n7130 & ~n8873 ;
  assign n8875 = n8869 & ~n8874 ;
  assign n8878 = n8877 ^ n8875 ^ 1'b0 ;
  assign n8880 = ~n1125 & n4180 ;
  assign n8881 = n8880 ^ n5845 ^ n2975 ;
  assign n8882 = n814 & ~n8881 ;
  assign n8879 = n708 & ~n5662 ;
  assign n8883 = n8882 ^ n8879 ^ 1'b0 ;
  assign n8884 = n7952 ^ n5836 ^ 1'b0 ;
  assign n8885 = n8884 ^ n4862 ^ n325 ;
  assign n8887 = n264 | n1261 ;
  assign n8888 = n8887 ^ n3197 ^ 1'b0 ;
  assign n8886 = n4299 ^ n3622 ^ 1'b0 ;
  assign n8889 = n8888 ^ n8886 ^ 1'b0 ;
  assign n8890 = x159 & ~n4008 ;
  assign n8891 = n8890 ^ n6934 ^ 1'b0 ;
  assign n8892 = n8754 ^ n2721 ^ 1'b0 ;
  assign n8893 = n1442 & ~n3762 ;
  assign n8894 = n8893 ^ n1206 ^ 1'b0 ;
  assign n8895 = n1132 & ~n8894 ;
  assign n8896 = n1276 ^ x189 ^ 1'b0 ;
  assign n8897 = n5984 | n8896 ;
  assign n8898 = n611 | n8897 ;
  assign n8899 = n4042 & ~n8898 ;
  assign n8900 = n1353 | n3846 ;
  assign n8901 = n2915 & n8900 ;
  assign n8902 = ~n6119 & n8901 ;
  assign n8903 = n6242 ^ n5264 ^ 1'b0 ;
  assign n8904 = ~n8902 & n8903 ;
  assign n8905 = n2618 ^ n1921 ^ 1'b0 ;
  assign n8906 = ~n1777 & n7564 ;
  assign n8907 = ~n4070 & n8906 ;
  assign n8908 = ~n1527 & n4325 ;
  assign n8909 = n7575 & n8908 ;
  assign n8910 = n1001 & ~n5884 ;
  assign n8911 = n4497 & n8910 ;
  assign n8912 = ( ~x145 & n2108 ) | ( ~x145 & n8911 ) | ( n2108 & n8911 ) ;
  assign n8913 = n5508 ^ n3044 ^ 1'b0 ;
  assign n8914 = n8912 | n8913 ;
  assign n8915 = n2949 & ~n7187 ;
  assign n8916 = ( n1077 & n5626 ) | ( n1077 & ~n8915 ) | ( n5626 & ~n8915 ) ;
  assign n8917 = n4786 & ~n6763 ;
  assign n8918 = n8917 ^ n2930 ^ 1'b0 ;
  assign n8919 = x136 & ~n8918 ;
  assign n8920 = n7759 ^ n2755 ^ 1'b0 ;
  assign n8921 = x6 & n8920 ;
  assign n8922 = n6383 & n8921 ;
  assign n8923 = n8922 ^ n7275 ^ 1'b0 ;
  assign n8924 = n4104 & n6129 ;
  assign n8925 = n8845 ^ n3104 ^ 1'b0 ;
  assign n8926 = ( n7190 & n8924 ) | ( n7190 & n8925 ) | ( n8924 & n8925 ) ;
  assign n8927 = n8105 ^ n5765 ^ 1'b0 ;
  assign n8928 = n6976 & ~n8927 ;
  assign n8937 = n7042 ^ n2506 ^ 1'b0 ;
  assign n8938 = n8937 ^ n1069 ^ 1'b0 ;
  assign n8929 = n1368 ^ x247 ^ 1'b0 ;
  assign n8930 = n1898 | n8929 ;
  assign n8931 = n8930 ^ n1432 ^ n1036 ;
  assign n8932 = x152 & n8931 ;
  assign n8933 = ~n1879 & n8932 ;
  assign n8934 = n8933 ^ n4908 ^ 1'b0 ;
  assign n8935 = n2154 & n8934 ;
  assign n8936 = n8935 ^ n1020 ^ 1'b0 ;
  assign n8939 = n8938 ^ n8936 ^ n8194 ;
  assign n8940 = ( n2366 & ~n6778 ) | ( n2366 & n8939 ) | ( ~n6778 & n8939 ) ;
  assign n8941 = n908 | n4082 ;
  assign n8942 = ~n514 & n1500 ;
  assign n8943 = n8942 ^ n3385 ^ 1'b0 ;
  assign n8944 = ~n3615 & n8041 ;
  assign n8945 = n8944 ^ n5463 ^ 1'b0 ;
  assign n8947 = n6358 ^ n501 ^ 1'b0 ;
  assign n8946 = n2705 & n3267 ;
  assign n8948 = n8947 ^ n8946 ^ 1'b0 ;
  assign n8949 = n1845 & n8270 ;
  assign n8950 = n8949 ^ n6872 ^ 1'b0 ;
  assign n8951 = n3444 & n3819 ;
  assign n8952 = ~x112 & n3631 ;
  assign n8953 = n6920 & n8952 ;
  assign n8954 = n8953 ^ n5715 ^ 1'b0 ;
  assign n8955 = n3421 ^ n875 ^ 1'b0 ;
  assign n8956 = x53 | n2464 ;
  assign n8957 = n3772 & ~n8956 ;
  assign n8958 = n2809 & ~n8957 ;
  assign n8959 = ( n739 & n8955 ) | ( n739 & ~n8958 ) | ( n8955 & ~n8958 ) ;
  assign n8961 = ~n4316 & n7954 ;
  assign n8962 = n372 & n8961 ;
  assign n8960 = n440 | n1051 ;
  assign n8963 = n8962 ^ n8960 ^ 1'b0 ;
  assign n8964 = n2190 & ~n3944 ;
  assign n8965 = n4627 & n7350 ;
  assign n8966 = ~n8964 & n8965 ;
  assign n8967 = n2224 | n6116 ;
  assign n8968 = ~n471 & n1449 ;
  assign n8969 = n8967 & n8968 ;
  assign n8970 = n863 & ~n1351 ;
  assign n8971 = n5680 & n8970 ;
  assign n8972 = ( n2228 & n4433 ) | ( n2228 & ~n8028 ) | ( n4433 & ~n8028 ) ;
  assign n8973 = n8972 ^ n1830 ^ 1'b0 ;
  assign n8974 = n5560 & ~n7016 ;
  assign n8975 = n3541 & ~n5511 ;
  assign n8976 = n8975 ^ n501 ^ 1'b0 ;
  assign n8977 = ~n3778 & n6051 ;
  assign n8978 = ( n5613 & n8976 ) | ( n5613 & ~n8977 ) | ( n8976 & ~n8977 ) ;
  assign n8979 = n3637 | n4011 ;
  assign n8980 = n8979 ^ n8506 ^ 1'b0 ;
  assign n8981 = ( n8974 & n8978 ) | ( n8974 & n8980 ) | ( n8978 & n8980 ) ;
  assign n8983 = ( n666 & n3325 ) | ( n666 & ~n3948 ) | ( n3325 & ~n3948 ) ;
  assign n8982 = n4562 & ~n7447 ;
  assign n8984 = n8983 ^ n8982 ^ n1749 ;
  assign n8986 = n1001 | n4811 ;
  assign n8987 = n787 & ~n8986 ;
  assign n8985 = n1958 & n3267 ;
  assign n8988 = n8987 ^ n8985 ^ 1'b0 ;
  assign n8989 = n7015 & ~n8988 ;
  assign n8990 = n3416 & ~n8989 ;
  assign n8991 = ( n469 & ~n1238 ) | ( n469 & n3465 ) | ( ~n1238 & n3465 ) ;
  assign n8992 = n1220 & ~n3060 ;
  assign n8993 = n8992 ^ n4616 ^ 1'b0 ;
  assign n8994 = n4876 | n8993 ;
  assign n8995 = n4780 | n8994 ;
  assign n8996 = n8995 ^ n3962 ^ 1'b0 ;
  assign n8997 = ( n6412 & n8991 ) | ( n6412 & n8996 ) | ( n8991 & n8996 ) ;
  assign n8998 = n4282 | n8997 ;
  assign n8999 = n3812 & ~n8583 ;
  assign n9000 = n556 & n8999 ;
  assign n9001 = n9000 ^ x217 ^ 1'b0 ;
  assign n9002 = n5350 & n5420 ;
  assign n9003 = n1595 | n2670 ;
  assign n9004 = n4292 & ~n9003 ;
  assign n9005 = n9004 ^ n3345 ^ 1'b0 ;
  assign n9006 = n9002 & n9005 ;
  assign n9007 = n9001 | n9006 ;
  assign n9008 = ~n2975 & n7580 ;
  assign n9009 = n9008 ^ n2850 ^ 1'b0 ;
  assign n9010 = ( n3272 & n3498 ) | ( n3272 & ~n4811 ) | ( n3498 & ~n4811 ) ;
  assign n9011 = x218 & ~n4377 ;
  assign n9012 = ~n9010 & n9011 ;
  assign n9013 = n3477 ^ x90 ^ 1'b0 ;
  assign n9014 = ( n3543 & ~n6490 ) | ( n3543 & n9013 ) | ( ~n6490 & n9013 ) ;
  assign n9015 = n9014 ^ n3970 ^ 1'b0 ;
  assign n9016 = ( n865 & ~n9012 ) | ( n865 & n9015 ) | ( ~n9012 & n9015 ) ;
  assign n9017 = n9016 ^ n7853 ^ n1395 ;
  assign n9018 = n5481 ^ n5425 ^ 1'b0 ;
  assign n9019 = ~n4091 & n9018 ;
  assign n9020 = n7261 & n7423 ;
  assign n9021 = n9020 ^ n5136 ^ 1'b0 ;
  assign n9022 = n1995 | n2900 ;
  assign n9023 = n3262 | n4301 ;
  assign n9024 = n9022 | n9023 ;
  assign n9025 = ~n834 & n4420 ;
  assign n9026 = n9025 ^ n6458 ^ 1'b0 ;
  assign n9027 = n9026 ^ n8630 ^ 1'b0 ;
  assign n9028 = n6414 ^ n6179 ^ n2919 ;
  assign n9029 = n2075 | n9028 ;
  assign n9030 = n4384 | n9029 ;
  assign n9031 = n7902 | n9030 ;
  assign n9037 = n2566 ^ n1134 ^ 1'b0 ;
  assign n9032 = n4988 ^ n4187 ^ 1'b0 ;
  assign n9033 = n4657 ^ x77 ^ 1'b0 ;
  assign n9034 = ~n6017 & n9033 ;
  assign n9035 = n9034 ^ n8064 ^ 1'b0 ;
  assign n9036 = n9032 & n9035 ;
  assign n9038 = n9037 ^ n9036 ^ 1'b0 ;
  assign n9039 = ~n4764 & n6745 ;
  assign n9040 = n3237 | n5458 ;
  assign n9041 = n2309 | n9040 ;
  assign n9042 = ~n4757 & n9041 ;
  assign n9043 = n9042 ^ n1613 ^ 1'b0 ;
  assign n9044 = ~n9039 & n9043 ;
  assign n9045 = n7110 & n9044 ;
  assign n9046 = n5837 ^ n4617 ^ 1'b0 ;
  assign n9047 = n4566 & n8976 ;
  assign n9048 = n2291 & n9047 ;
  assign n9049 = ( x238 & n4360 ) | ( x238 & n9048 ) | ( n4360 & n9048 ) ;
  assign n9050 = n1298 & n8947 ;
  assign n9051 = n9050 ^ n1147 ^ 1'b0 ;
  assign n9052 = n5086 & n9051 ;
  assign n9053 = n9049 & n9052 ;
  assign n9056 = n315 | n867 ;
  assign n9054 = ( ~x107 & n4115 ) | ( ~x107 & n9012 ) | ( n4115 & n9012 ) ;
  assign n9055 = ~n8820 & n9054 ;
  assign n9057 = n9056 ^ n9055 ^ 1'b0 ;
  assign n9058 = n8408 ^ n2936 ^ 1'b0 ;
  assign n9059 = n1333 & ~n9058 ;
  assign n9060 = n3926 ^ n3260 ^ 1'b0 ;
  assign n9061 = n1276 ^ x14 ^ 1'b0 ;
  assign n9062 = n9061 ^ n2986 ^ 1'b0 ;
  assign n9063 = n3077 | n3977 ;
  assign n9064 = n8996 & ~n9063 ;
  assign n9065 = n8996 ^ n4767 ^ 1'b0 ;
  assign n9066 = n7478 ^ n569 ^ 1'b0 ;
  assign n9067 = n1001 | n9066 ;
  assign n9068 = x64 & ~n9067 ;
  assign n9069 = n4642 & n7099 ;
  assign n9070 = n9069 ^ n4650 ^ 1'b0 ;
  assign n9071 = ~n9068 & n9070 ;
  assign n9072 = n9071 ^ n5252 ^ 1'b0 ;
  assign n9073 = n276 | n411 ;
  assign n9074 = n9073 ^ n2828 ^ 1'b0 ;
  assign n9075 = n9072 | n9074 ;
  assign n9077 = n4230 ^ n2309 ^ 1'b0 ;
  assign n9078 = n7407 & n9077 ;
  assign n9079 = n722 & ~n4328 ;
  assign n9080 = ( n997 & n9078 ) | ( n997 & n9079 ) | ( n9078 & n9079 ) ;
  assign n9076 = ~n1817 & n2092 ;
  assign n9081 = n9080 ^ n9076 ^ 1'b0 ;
  assign n9082 = n5667 ^ n3925 ^ 1'b0 ;
  assign n9083 = n9081 & n9082 ;
  assign n9084 = ~n8529 & n9083 ;
  assign n9085 = ~n5570 & n9084 ;
  assign n9086 = n466 & ~n5649 ;
  assign n9087 = ~n9085 & n9086 ;
  assign n9088 = n9087 ^ n957 ^ 1'b0 ;
  assign n9089 = n5586 ^ x91 ^ 1'b0 ;
  assign n9090 = ~n291 & n9089 ;
  assign n9093 = n1739 & n5179 ;
  assign n9092 = n1552 & ~n5768 ;
  assign n9094 = n9093 ^ n9092 ^ 1'b0 ;
  assign n9091 = n569 & ~n921 ;
  assign n9095 = n9094 ^ n9091 ^ n2462 ;
  assign n9096 = ~n9090 & n9095 ;
  assign n9097 = x185 & n3016 ;
  assign n9098 = n6278 & n9097 ;
  assign n9099 = n1264 & n1671 ;
  assign n9100 = n1206 ^ n682 ^ 1'b0 ;
  assign n9101 = n9099 & n9100 ;
  assign n9102 = n9101 ^ n3888 ^ 1'b0 ;
  assign n9103 = ~n4543 & n9102 ;
  assign n9104 = ~n6031 & n9103 ;
  assign n9105 = n6018 ^ n1186 ^ 1'b0 ;
  assign n9106 = n5881 & n9105 ;
  assign n9107 = n9106 ^ n7407 ^ 1'b0 ;
  assign n9108 = ~n3109 & n6467 ;
  assign n9109 = n7266 & n9108 ;
  assign n9113 = n1318 & n4666 ;
  assign n9112 = ~n507 & n5476 ;
  assign n9114 = n9113 ^ n9112 ^ 1'b0 ;
  assign n9110 = n1301 & ~n4780 ;
  assign n9111 = n9110 ^ n585 ^ 1'b0 ;
  assign n9115 = n9114 ^ n9111 ^ 1'b0 ;
  assign n9117 = n8877 ^ n5728 ^ 1'b0 ;
  assign n9116 = ( n615 & n1028 ) | ( n615 & n5412 ) | ( n1028 & n5412 ) ;
  assign n9118 = n9117 ^ n9116 ^ 1'b0 ;
  assign n9119 = ~n5452 & n9118 ;
  assign n9120 = ~n1071 & n2533 ;
  assign n9121 = n9120 ^ n2382 ^ 1'b0 ;
  assign n9122 = x106 & ~n3215 ;
  assign n9123 = ~n9121 & n9122 ;
  assign n9124 = n3500 & ~n9123 ;
  assign n9125 = n9124 ^ n1653 ^ 1'b0 ;
  assign n9126 = n4016 | n9125 ;
  assign n9127 = n7994 ^ n3003 ^ 1'b0 ;
  assign n9128 = ~n2029 & n9127 ;
  assign n9129 = n9128 ^ n3786 ^ 1'b0 ;
  assign n9130 = ~n9126 & n9129 ;
  assign n9136 = ~x180 & n4357 ;
  assign n9137 = n4042 & n9136 ;
  assign n9131 = n3304 | n4004 ;
  assign n9132 = n4310 & ~n9131 ;
  assign n9133 = n2966 | n9132 ;
  assign n9134 = n2881 & ~n9133 ;
  assign n9135 = n4892 | n9134 ;
  assign n9138 = n9137 ^ n9135 ^ 1'b0 ;
  assign n9139 = n2456 | n3344 ;
  assign n9140 = n3888 & ~n9139 ;
  assign n9141 = n8997 & ~n9140 ;
  assign n9142 = n9141 ^ n7306 ^ 1'b0 ;
  assign n9143 = ~n1910 & n2091 ;
  assign n9144 = ~n2520 & n9143 ;
  assign n9145 = n1048 ^ x97 ^ 1'b0 ;
  assign n9146 = n2622 & n9145 ;
  assign n9147 = n3643 & n9146 ;
  assign n9148 = ~n9144 & n9147 ;
  assign n9149 = n5450 & n9148 ;
  assign n9150 = n6902 | n7558 ;
  assign n9151 = n9150 ^ n4844 ^ 1'b0 ;
  assign n9152 = x181 & n3607 ;
  assign n9153 = ~n2110 & n9152 ;
  assign n9154 = n9153 ^ n4153 ^ 1'b0 ;
  assign n9155 = ( n2972 & n7361 ) | ( n2972 & n9154 ) | ( n7361 & n9154 ) ;
  assign n9156 = n2925 | n4515 ;
  assign n9157 = n9156 ^ n4861 ^ 1'b0 ;
  assign n9158 = ~n9155 & n9157 ;
  assign n9159 = ~n2110 & n9158 ;
  assign n9160 = n3926 ^ x218 ^ 1'b0 ;
  assign n9161 = n3118 | n9160 ;
  assign n9162 = n9161 ^ n4861 ^ x142 ;
  assign n9169 = n1442 & n5902 ;
  assign n9170 = n9169 ^ n4607 ^ 1'b0 ;
  assign n9167 = n7923 ^ n6805 ^ n2178 ;
  assign n9166 = n4325 & n4443 ;
  assign n9168 = n9167 ^ n9166 ^ 1'b0 ;
  assign n9163 = ~n498 & n5413 ;
  assign n9164 = n1215 & n9163 ;
  assign n9165 = n3429 & n9164 ;
  assign n9171 = n9170 ^ n9168 ^ n9165 ;
  assign n9172 = n7484 ^ n4267 ^ 1'b0 ;
  assign n9173 = n1932 ^ x223 ^ 1'b0 ;
  assign n9174 = n3226 & n9173 ;
  assign n9175 = n9174 ^ n3703 ^ 1'b0 ;
  assign n9176 = n9175 ^ x127 ^ 1'b0 ;
  assign n9177 = n2182 & n9176 ;
  assign n9178 = n9177 ^ n2401 ^ 1'b0 ;
  assign n9179 = n9172 & n9178 ;
  assign n9180 = n5685 | n7515 ;
  assign n9181 = n1633 & n3772 ;
  assign n9182 = n4542 ^ n1909 ^ 1'b0 ;
  assign n9183 = n6385 | n9182 ;
  assign n9184 = n3059 ^ n1943 ^ 1'b0 ;
  assign n9185 = n3416 & ~n9184 ;
  assign n9186 = n9185 ^ n8052 ^ n7355 ;
  assign n9188 = n5970 ^ n2105 ^ 1'b0 ;
  assign n9189 = x175 & ~n9188 ;
  assign n9187 = n5996 ^ n2320 ^ 1'b0 ;
  assign n9190 = n9189 ^ n9187 ^ n8166 ;
  assign n9191 = n2450 ^ n973 ^ 1'b0 ;
  assign n9192 = ~n713 & n9191 ;
  assign n9193 = n6311 ^ n3650 ^ 1'b0 ;
  assign n9194 = ( n720 & n2040 ) | ( n720 & ~n2319 ) | ( n2040 & ~n2319 ) ;
  assign n9195 = n9194 ^ n4400 ^ 1'b0 ;
  assign n9196 = x162 & ~n1020 ;
  assign n9197 = n9196 ^ n336 ^ 1'b0 ;
  assign n9198 = n9195 & ~n9197 ;
  assign n9199 = n4553 ^ n3258 ^ 1'b0 ;
  assign n9200 = ~n6411 & n9199 ;
  assign n9201 = x212 & n9200 ;
  assign n9202 = n9201 ^ n4571 ^ 1'b0 ;
  assign n9203 = n1608 ^ n1028 ^ 1'b0 ;
  assign n9204 = n4696 & n9203 ;
  assign n9205 = n9204 ^ n8270 ^ n4524 ;
  assign n9206 = n9205 ^ n5065 ^ n4011 ;
  assign n9207 = n2735 & n3830 ;
  assign n9208 = x49 & n1133 ;
  assign n9209 = n9208 ^ n1445 ^ 1'b0 ;
  assign n9210 = n9207 & n9209 ;
  assign n9211 = n6177 ^ n5786 ^ 1'b0 ;
  assign n9212 = ~n486 & n3850 ;
  assign n9213 = n2859 ^ n1042 ^ 1'b0 ;
  assign n9214 = n9212 | n9213 ;
  assign n9215 = n9214 ^ n5163 ^ 1'b0 ;
  assign n9218 = n5269 ^ n1471 ^ 1'b0 ;
  assign n9216 = n2701 ^ n2221 ^ 1'b0 ;
  assign n9217 = ~n2097 & n9216 ;
  assign n9219 = n9218 ^ n9217 ^ 1'b0 ;
  assign n9220 = n5229 | n6313 ;
  assign n9221 = ~n7448 & n9220 ;
  assign n9222 = n6927 ^ n882 ^ 1'b0 ;
  assign n9223 = n9221 & n9222 ;
  assign n9224 = ~n1089 & n5017 ;
  assign n9225 = n826 & n9224 ;
  assign n9226 = ~n1353 & n1579 ;
  assign n9227 = ~n1119 & n7742 ;
  assign n9228 = ( n4788 & n8219 ) | ( n4788 & n9227 ) | ( n8219 & n9227 ) ;
  assign n9229 = n8253 ^ n4768 ^ 1'b0 ;
  assign n9230 = ~n3164 & n9229 ;
  assign n9231 = ~n3481 & n7031 ;
  assign n9232 = n9231 ^ n3003 ^ 1'b0 ;
  assign n9234 = ~n1936 & n2055 ;
  assign n9235 = n2754 & n9234 ;
  assign n9233 = n842 & ~n4159 ;
  assign n9236 = n9235 ^ n9233 ^ 1'b0 ;
  assign n9237 = n4807 ^ n940 ^ 1'b0 ;
  assign n9238 = n2622 & ~n3251 ;
  assign n9239 = n7433 & n9238 ;
  assign n9240 = n6291 | n7240 ;
  assign n9241 = n9240 ^ n4276 ^ 1'b0 ;
  assign n9242 = n2011 | n6037 ;
  assign n9243 = n2705 | n9242 ;
  assign n9244 = n6367 & n9243 ;
  assign n9245 = n9244 ^ n4033 ^ 1'b0 ;
  assign n9246 = n9245 ^ n4638 ^ 1'b0 ;
  assign n9247 = n7779 & ~n8624 ;
  assign n9248 = ~n4835 & n9247 ;
  assign n9249 = n8647 ^ n1874 ^ 1'b0 ;
  assign n9250 = x96 & n9249 ;
  assign n9251 = n7761 ^ n5749 ^ 1'b0 ;
  assign n9252 = n9251 ^ n3903 ^ 1'b0 ;
  assign n9253 = n6246 ^ n4649 ^ 1'b0 ;
  assign n9254 = n1913 & n9253 ;
  assign n9255 = ~n1219 & n9254 ;
  assign n9256 = n7700 ^ n2884 ^ 1'b0 ;
  assign n9257 = n8933 ^ n7819 ^ 1'b0 ;
  assign n9258 = n4329 | n9257 ;
  assign n9259 = n8544 ^ n1710 ^ 1'b0 ;
  assign n9260 = n5261 ^ n2529 ^ 1'b0 ;
  assign n9261 = n9260 ^ n8577 ^ 1'b0 ;
  assign n9262 = n4056 & n9261 ;
  assign n9263 = n3819 | n9262 ;
  assign n9271 = n3595 & n4222 ;
  assign n9272 = n9271 ^ n8822 ^ 1'b0 ;
  assign n9273 = ~n4094 & n9272 ;
  assign n9265 = n1118 & ~n2770 ;
  assign n9266 = ~x104 & n9265 ;
  assign n9267 = n9212 & ~n9266 ;
  assign n9268 = n9267 ^ n2867 ^ n839 ;
  assign n9264 = n5324 & ~n5705 ;
  assign n9269 = n9268 ^ n9264 ^ 1'b0 ;
  assign n9270 = n8030 & ~n9269 ;
  assign n9274 = n9273 ^ n9270 ^ 1'b0 ;
  assign n9275 = ~n3554 & n9274 ;
  assign n9276 = ~n2516 & n9275 ;
  assign n9279 = n1536 & ~n1851 ;
  assign n9280 = ~n4039 & n9279 ;
  assign n9277 = n2247 & ~n4161 ;
  assign n9278 = n9277 ^ n925 ^ 1'b0 ;
  assign n9281 = n9280 ^ n9278 ^ 1'b0 ;
  assign n9282 = n3936 & ~n9281 ;
  assign n9283 = n9282 ^ n1017 ^ 1'b0 ;
  assign n9284 = n611 & ~n973 ;
  assign n9285 = n2462 & n9284 ;
  assign n9286 = n1975 & n9285 ;
  assign n9287 = ~n5355 & n9286 ;
  assign n9288 = n3619 & ~n6638 ;
  assign n9289 = n6192 ^ n1030 ^ 1'b0 ;
  assign n9290 = ( n1048 & n1437 ) | ( n1048 & n6815 ) | ( n1437 & n6815 ) ;
  assign n9291 = n2274 & ~n9290 ;
  assign n9292 = ( ~n378 & n4434 ) | ( ~n378 & n9291 ) | ( n4434 & n9291 ) ;
  assign n9293 = n2746 | n9292 ;
  assign n9294 = n2741 | n5469 ;
  assign n9295 = ~n6678 & n6981 ;
  assign n9298 = ~n1126 & n4669 ;
  assign n9296 = ( n749 & ~n4599 ) | ( n749 & n5587 ) | ( ~n4599 & n5587 ) ;
  assign n9297 = ~n893 & n9296 ;
  assign n9299 = n9298 ^ n9297 ^ 1'b0 ;
  assign n9301 = n606 & ~n5737 ;
  assign n9300 = ~x6 & n1111 ;
  assign n9302 = n9301 ^ n9300 ^ 1'b0 ;
  assign n9303 = ( n761 & ~n3039 ) | ( n761 & n6947 ) | ( ~n3039 & n6947 ) ;
  assign n9304 = n9303 ^ n6974 ^ 1'b0 ;
  assign n9305 = ~n5617 & n8112 ;
  assign n9306 = n9305 ^ n9078 ^ 1'b0 ;
  assign n9307 = n9260 & ~n9306 ;
  assign n9313 = ~n725 & n2508 ;
  assign n9309 = n2394 ^ n2331 ^ 1'b0 ;
  assign n9310 = x83 & ~n9309 ;
  assign n9308 = n509 | n4704 ;
  assign n9311 = n9310 ^ n9308 ^ 1'b0 ;
  assign n9312 = ~n4342 & n9311 ;
  assign n9314 = n9313 ^ n9312 ^ 1'b0 ;
  assign n9315 = n1441 & ~n1505 ;
  assign n9316 = n9315 ^ x68 ^ 1'b0 ;
  assign n9317 = n4693 ^ n1799 ^ 1'b0 ;
  assign n9318 = n9317 ^ n2976 ^ 1'b0 ;
  assign n9319 = n9316 | n9318 ;
  assign n9320 = n8346 ^ n5018 ^ 1'b0 ;
  assign n9321 = n2939 | n9320 ;
  assign n9323 = n4259 & ~n5475 ;
  assign n9324 = ~n4888 & n9323 ;
  assign n9322 = ( n518 & n2587 ) | ( n518 & ~n8738 ) | ( n2587 & ~n8738 ) ;
  assign n9325 = n9324 ^ n9322 ^ 1'b0 ;
  assign n9326 = n6319 ^ n2935 ^ 1'b0 ;
  assign n9327 = n9232 & n9326 ;
  assign n9333 = ~n2095 & n2853 ;
  assign n9331 = x100 | n1805 ;
  assign n9332 = n7361 & ~n9331 ;
  assign n9334 = n9333 ^ n9332 ^ 1'b0 ;
  assign n9328 = ~n1369 & n3059 ;
  assign n9329 = n9328 ^ x113 ^ 1'b0 ;
  assign n9330 = ~n5951 & n9329 ;
  assign n9335 = n9334 ^ n9330 ^ n4485 ;
  assign n9337 = n3165 | n5241 ;
  assign n9338 = n1415 | n1905 ;
  assign n9339 = n9338 ^ n8401 ^ n4942 ;
  assign n9340 = ~n9337 & n9339 ;
  assign n9336 = n3892 | n4296 ;
  assign n9341 = n9340 ^ n9336 ^ 1'b0 ;
  assign n9342 = ~n514 & n9341 ;
  assign n9343 = x46 & ~n9342 ;
  assign n9344 = n5293 ^ n3319 ^ 1'b0 ;
  assign n9345 = n8718 | n9344 ;
  assign n9348 = ( ~n1667 & n3631 ) | ( ~n1667 & n4739 ) | ( n3631 & n4739 ) ;
  assign n9349 = n9348 ^ x6 ^ 1'b0 ;
  assign n9350 = ~n5608 & n9349 ;
  assign n9351 = ( n614 & n2641 ) | ( n614 & ~n9350 ) | ( n2641 & ~n9350 ) ;
  assign n9352 = n9351 ^ n6192 ^ 1'b0 ;
  assign n9346 = n7496 ^ n5967 ^ 1'b0 ;
  assign n9347 = n1975 & ~n9346 ;
  assign n9353 = n9352 ^ n9347 ^ n2267 ;
  assign n9354 = n9126 ^ n4216 ^ 1'b0 ;
  assign n9355 = n5055 ^ n3890 ^ 1'b0 ;
  assign n9356 = n4855 ^ n2993 ^ 1'b0 ;
  assign n9357 = n2434 & n9356 ;
  assign n9358 = n3287 | n3851 ;
  assign n9359 = ( ~x157 & n1901 ) | ( ~x157 & n9358 ) | ( n1901 & n9358 ) ;
  assign n9360 = ( n4612 & n9357 ) | ( n4612 & n9359 ) | ( n9357 & n9359 ) ;
  assign n9365 = ( n799 & n2572 ) | ( n799 & ~n2705 ) | ( n2572 & ~n2705 ) ;
  assign n9366 = n9365 ^ n9066 ^ 1'b0 ;
  assign n9361 = n2026 | n5038 ;
  assign n9362 = n9361 ^ n1680 ^ 1'b0 ;
  assign n9363 = ~n1258 & n9362 ;
  assign n9364 = n2500 & n9363 ;
  assign n9367 = n9366 ^ n9364 ^ 1'b0 ;
  assign n9368 = n1914 & ~n6148 ;
  assign n9369 = ~n529 & n9368 ;
  assign n9370 = ~n9368 & n9369 ;
  assign n9371 = n5119 ^ n1257 ^ 1'b0 ;
  assign n9372 = n2209 | n3513 ;
  assign n9373 = n9371 & ~n9372 ;
  assign n9374 = ~n2354 & n6595 ;
  assign n9375 = n618 & n9374 ;
  assign n9376 = n2796 | n6639 ;
  assign n9377 = n9375 & ~n9376 ;
  assign n9378 = n9373 & ~n9377 ;
  assign n9379 = n988 | n2867 ;
  assign n9380 = n4431 & ~n9379 ;
  assign n9381 = n7096 & ~n9380 ;
  assign n9382 = n9381 ^ n1200 ^ 1'b0 ;
  assign n9384 = n1008 & n5998 ;
  assign n9385 = n5623 & n9384 ;
  assign n9383 = n1352 ^ n710 ^ 1'b0 ;
  assign n9386 = n9385 ^ n9383 ^ 1'b0 ;
  assign n9387 = n4366 ^ n3052 ^ 1'b0 ;
  assign n9388 = n6671 & ~n9387 ;
  assign n9389 = n4880 ^ x47 ^ 1'b0 ;
  assign n9390 = n9389 ^ n6155 ^ n2345 ;
  assign n9391 = n9390 ^ n3070 ^ 1'b0 ;
  assign n9392 = x175 & n3018 ;
  assign n9393 = ~n2208 & n9392 ;
  assign n9394 = n4540 | n9393 ;
  assign n9395 = n2225 & ~n9394 ;
  assign n9396 = n2064 & ~n9395 ;
  assign n9397 = ~n6810 & n9396 ;
  assign n9398 = n9397 ^ n6168 ^ n1851 ;
  assign n9399 = ~n992 & n6231 ;
  assign n9400 = n9399 ^ n7087 ^ 1'b0 ;
  assign n9401 = ( x182 & n274 ) | ( x182 & n3368 ) | ( n274 & n3368 ) ;
  assign n9402 = n2861 & n7904 ;
  assign n9403 = n6222 ^ n1869 ^ 1'b0 ;
  assign n9404 = n9402 | n9403 ;
  assign n9405 = n8573 & ~n9404 ;
  assign n9406 = n4892 & n9405 ;
  assign n9407 = n8819 ^ n3704 ^ 1'b0 ;
  assign n9408 = n385 & n9407 ;
  assign n9410 = n6991 ^ n4288 ^ 1'b0 ;
  assign n9411 = ~n8073 & n9410 ;
  assign n9409 = n951 & n3372 ;
  assign n9412 = n9411 ^ n9409 ^ 1'b0 ;
  assign n9413 = ~n5236 & n9412 ;
  assign n9414 = n3222 & ~n3514 ;
  assign n9415 = n9414 ^ n4580 ^ 1'b0 ;
  assign n9416 = ( n4481 & n6055 ) | ( n4481 & ~n9415 ) | ( n6055 & ~n9415 ) ;
  assign n9417 = n8276 ^ n5063 ^ 1'b0 ;
  assign n9418 = n562 & n9417 ;
  assign n9419 = n6294 ^ n4503 ^ n2509 ;
  assign n9420 = n3818 & n8063 ;
  assign n9421 = n3319 ^ n1657 ^ 1'b0 ;
  assign n9422 = ~n7428 & n9421 ;
  assign n9423 = n4591 & n8594 ;
  assign n9430 = n4047 ^ n3956 ^ 1'b0 ;
  assign n9431 = n4498 | n9430 ;
  assign n9429 = n483 & n4716 ;
  assign n9424 = n1344 ^ n1030 ^ 1'b0 ;
  assign n9425 = n2484 & n9424 ;
  assign n9426 = n9425 ^ n2711 ^ 1'b0 ;
  assign n9427 = n8957 | n9426 ;
  assign n9428 = ( n3475 & ~n6415 ) | ( n3475 & n9427 ) | ( ~n6415 & n9427 ) ;
  assign n9432 = n9431 ^ n9429 ^ n9428 ;
  assign n9433 = n3703 & ~n5563 ;
  assign n9434 = ( ~n294 & n2768 ) | ( ~n294 & n3255 ) | ( n2768 & n3255 ) ;
  assign n9440 = n4335 ^ n2468 ^ n642 ;
  assign n9441 = ~n6780 & n9440 ;
  assign n9442 = n4617 & n9441 ;
  assign n9435 = ~n2061 & n2721 ;
  assign n9436 = ~x106 & n9435 ;
  assign n9437 = n1568 & n9436 ;
  assign n9438 = n9437 ^ n3087 ^ 1'b0 ;
  assign n9439 = n9438 ^ n2215 ^ 1'b0 ;
  assign n9443 = n9442 ^ n9439 ^ x1 ;
  assign n9444 = n7345 & ~n9443 ;
  assign n9445 = n3156 ^ x30 ^ 1'b0 ;
  assign n9446 = n689 & ~n9445 ;
  assign n9447 = n7910 ^ n5001 ^ x16 ;
  assign n9448 = n8723 ^ n7099 ^ n5773 ;
  assign n9449 = x128 & ~n1219 ;
  assign n9450 = n7022 & n9449 ;
  assign n9451 = n9450 ^ n2752 ^ 1'b0 ;
  assign n9452 = ~n1276 & n9451 ;
  assign n9453 = n380 & ~n1557 ;
  assign n9454 = n9453 ^ x241 ^ 1'b0 ;
  assign n9455 = n4025 ^ n2871 ^ 1'b0 ;
  assign n9456 = n9015 & ~n9455 ;
  assign n9457 = n4547 ^ n338 ^ 1'b0 ;
  assign n9458 = n9457 ^ n3961 ^ 1'b0 ;
  assign n9459 = n9456 | n9458 ;
  assign n9460 = n1851 ^ n680 ^ 1'b0 ;
  assign n9461 = ~n2704 & n9460 ;
  assign n9462 = n323 & n9461 ;
  assign n9463 = n3258 & n9462 ;
  assign n9464 = n1151 & ~n2081 ;
  assign n9465 = ~x70 & n9464 ;
  assign n9466 = n7569 ^ n1313 ^ 1'b0 ;
  assign n9467 = ~n3592 & n3595 ;
  assign n9468 = ~n900 & n9467 ;
  assign n9469 = ~n787 & n2167 ;
  assign n9470 = n9469 ^ n9093 ^ 1'b0 ;
  assign n9471 = n4130 ^ n3034 ^ 1'b0 ;
  assign n9472 = n9471 ^ n3498 ^ 1'b0 ;
  assign n9473 = n9470 & ~n9472 ;
  assign n9474 = n523 & n2210 ;
  assign n9475 = n1165 & n9474 ;
  assign n9476 = n9475 ^ n1264 ^ n363 ;
  assign n9477 = n9476 ^ n5969 ^ n4165 ;
  assign n9478 = n4418 & n5377 ;
  assign n9479 = n4494 ^ x88 ^ 1'b0 ;
  assign n9480 = ~n9478 & n9479 ;
  assign n9481 = n5136 & n9480 ;
  assign n9482 = n2011 & ~n2039 ;
  assign n9483 = n9482 ^ n1590 ^ 1'b0 ;
  assign n9484 = n8815 ^ n1186 ^ x208 ;
  assign n9485 = n4933 & n9484 ;
  assign n9486 = n9485 ^ n5286 ^ 1'b0 ;
  assign n9487 = ~n2027 & n8366 ;
  assign n9488 = n9487 ^ n5374 ^ 1'b0 ;
  assign n9489 = n1662 & n9488 ;
  assign n9490 = ( x22 & n262 ) | ( x22 & ~n449 ) | ( n262 & ~n449 ) ;
  assign n9491 = ~n8276 & n9490 ;
  assign n9492 = n9491 ^ n1019 ^ 1'b0 ;
  assign n9493 = n3325 | n9492 ;
  assign n9494 = ( n766 & n1267 ) | ( n766 & ~n3258 ) | ( n1267 & ~n3258 ) ;
  assign n9495 = ( n2602 & n8869 ) | ( n2602 & ~n9494 ) | ( n8869 & ~n9494 ) ;
  assign n9496 = ~n3271 & n3823 ;
  assign n9498 = n8666 ^ n2455 ^ 1'b0 ;
  assign n9497 = n1290 & ~n2937 ;
  assign n9499 = n9498 ^ n9497 ^ 1'b0 ;
  assign n9500 = n9499 ^ n7799 ^ 1'b0 ;
  assign n9501 = x143 & ~n9500 ;
  assign n9502 = ( n1519 & ~n4599 ) | ( n1519 & n9501 ) | ( ~n4599 & n9501 ) ;
  assign n9503 = n442 | n1577 ;
  assign n9504 = n9503 ^ n2574 ^ 1'b0 ;
  assign n9505 = n5933 & ~n9504 ;
  assign n9506 = n3600 | n3975 ;
  assign n9507 = n9506 ^ n527 ^ 1'b0 ;
  assign n9508 = n4474 ^ n3399 ^ 1'b0 ;
  assign n9509 = n7838 & n9508 ;
  assign n9510 = n9507 & n9509 ;
  assign n9511 = n663 ^ n553 ^ 1'b0 ;
  assign n9512 = n2213 | n9511 ;
  assign n9513 = n4251 & n8945 ;
  assign n9514 = n5937 ^ n5063 ^ 1'b0 ;
  assign n9515 = n4070 & ~n4491 ;
  assign n9516 = ~n3622 & n4742 ;
  assign n9517 = n9516 ^ n8337 ^ 1'b0 ;
  assign n9518 = n9515 & n9517 ;
  assign n9520 = n407 & n2141 ;
  assign n9519 = n5431 & n7347 ;
  assign n9521 = n9520 ^ n9519 ^ 1'b0 ;
  assign n9522 = n9359 ^ n8660 ^ 1'b0 ;
  assign n9523 = x122 & ~n2883 ;
  assign n9524 = n4861 ^ n2622 ^ 1'b0 ;
  assign n9525 = n2570 & n9524 ;
  assign n9526 = n5229 ^ n3085 ^ 1'b0 ;
  assign n9527 = ~n2552 & n9526 ;
  assign n9528 = ~n1185 & n1822 ;
  assign n9529 = n9528 ^ n1763 ^ 1'b0 ;
  assign n9530 = x217 & ~n9529 ;
  assign n9531 = n9530 ^ n951 ^ 1'b0 ;
  assign n9532 = ~n444 & n6561 ;
  assign n9533 = n3149 ^ n2081 ^ 1'b0 ;
  assign n9534 = n5241 | n9533 ;
  assign n9535 = n1481 ^ n1124 ^ 1'b0 ;
  assign n9536 = n933 & n9535 ;
  assign n9537 = ~n3814 & n9536 ;
  assign n9538 = n9537 ^ n6910 ^ 1'b0 ;
  assign n9539 = ( n516 & n4605 ) | ( n516 & ~n6982 ) | ( n4605 & ~n6982 ) ;
  assign n9540 = n9461 ^ n5898 ^ n5342 ;
  assign n9541 = n4487 ^ n2400 ^ 1'b0 ;
  assign n9542 = x78 & n9541 ;
  assign n9543 = ~n7655 & n9542 ;
  assign n9544 = n5488 & n9543 ;
  assign n9545 = n8988 ^ n1001 ^ n529 ;
  assign n9546 = n963 & ~n9545 ;
  assign n9547 = ~n3328 & n3823 ;
  assign n9548 = n2809 & n9547 ;
  assign n9549 = ( n399 & n5061 ) | ( n399 & n7407 ) | ( n5061 & n7407 ) ;
  assign n9550 = n1660 & n9549 ;
  assign n9551 = n9548 & n9550 ;
  assign n9552 = n3263 & n5379 ;
  assign n9553 = ~n3012 & n9552 ;
  assign n9554 = n9551 & n9553 ;
  assign n9555 = n1858 | n3486 ;
  assign n9556 = n9555 ^ n1185 ^ 1'b0 ;
  assign n9557 = n3274 & n7219 ;
  assign n9558 = ( ~n1624 & n2180 ) | ( ~n1624 & n9557 ) | ( n2180 & n9557 ) ;
  assign n9559 = n9558 ^ n5648 ^ 1'b0 ;
  assign n9560 = ~n2081 & n9559 ;
  assign n9561 = n5080 ^ n2375 ^ 1'b0 ;
  assign n9562 = n9560 & n9561 ;
  assign n9563 = n3498 & ~n3768 ;
  assign n9564 = n8144 & n9563 ;
  assign n9565 = n9562 & ~n9564 ;
  assign n9566 = ~n4049 & n9565 ;
  assign n9568 = n6925 ^ n4920 ^ 1'b0 ;
  assign n9567 = n1610 & ~n4185 ;
  assign n9569 = n9568 ^ n9567 ^ 1'b0 ;
  assign n9570 = n1346 ^ x162 ^ 1'b0 ;
  assign n9571 = n9569 & n9570 ;
  assign n9572 = n5920 ^ n4768 ^ 1'b0 ;
  assign n9573 = ~n1415 & n3377 ;
  assign n9574 = n9573 ^ n2701 ^ 1'b0 ;
  assign n9575 = n587 | n9574 ;
  assign n9576 = n9575 ^ n817 ^ 1'b0 ;
  assign n9577 = ( ~n6578 & n7319 ) | ( ~n6578 & n7638 ) | ( n7319 & n7638 ) ;
  assign n9578 = n7222 ^ n4290 ^ 1'b0 ;
  assign n9579 = n9578 ^ n8673 ^ 1'b0 ;
  assign n9580 = ~n7290 & n9579 ;
  assign n9581 = ~n5608 & n6865 ;
  assign n9582 = n9581 ^ n2237 ^ 1'b0 ;
  assign n9583 = n9582 ^ x164 ^ 1'b0 ;
  assign n9584 = n1324 & n9583 ;
  assign n9585 = x189 & ~n1911 ;
  assign n9586 = n9585 ^ n2172 ^ 1'b0 ;
  assign n9587 = ( ~n606 & n8366 ) | ( ~n606 & n9586 ) | ( n8366 & n9586 ) ;
  assign n9588 = ~n320 & n2545 ;
  assign n9589 = n9588 ^ x89 ^ 1'b0 ;
  assign n9590 = n9589 ^ x6 ^ 1'b0 ;
  assign n9594 = n8305 ^ n1065 ^ n851 ;
  assign n9591 = x70 & ~n2883 ;
  assign n9592 = n9591 ^ n5112 ^ 1'b0 ;
  assign n9593 = ~n4892 & n9592 ;
  assign n9595 = n9594 ^ n9593 ^ 1'b0 ;
  assign n9596 = x7 & ~n3035 ;
  assign n9597 = ~x37 & n9596 ;
  assign n9598 = n1600 & ~n9597 ;
  assign n9599 = ~n8011 & n9598 ;
  assign n9600 = ( n2592 & n5210 ) | ( n2592 & ~n7775 ) | ( n5210 & ~n7775 ) ;
  assign n9601 = n4029 ^ n1065 ^ 1'b0 ;
  assign n9602 = n3817 ^ n1257 ^ 1'b0 ;
  assign n9603 = n369 | n9602 ;
  assign n9604 = n627 & ~n9603 ;
  assign n9605 = ~n9601 & n9604 ;
  assign n9606 = x112 & ~n9605 ;
  assign n9607 = n9606 ^ n6295 ^ 1'b0 ;
  assign n9608 = ~x113 & n510 ;
  assign n9617 = n7635 ^ n4938 ^ 1'b0 ;
  assign n9609 = ~n806 & n951 ;
  assign n9610 = n9609 ^ n1086 ^ n333 ;
  assign n9611 = n9610 ^ n3110 ^ 1'b0 ;
  assign n9612 = x244 & n4138 ;
  assign n9613 = n2424 & ~n9612 ;
  assign n9614 = n5777 & n9613 ;
  assign n9615 = n6506 & ~n9614 ;
  assign n9616 = ~n9611 & n9615 ;
  assign n9618 = n9617 ^ n9616 ^ 1'b0 ;
  assign n9619 = x236 & n1667 ;
  assign n9620 = n2735 & ~n9619 ;
  assign n9621 = x41 & ~x42 ;
  assign n9622 = n9621 ^ n9461 ^ 1'b0 ;
  assign n9623 = n659 & ~n9622 ;
  assign n9624 = n7752 ^ n5831 ^ 1'b0 ;
  assign n9625 = n6391 | n8622 ;
  assign n9626 = ~n1204 & n2219 ;
  assign n9627 = n1492 & n9626 ;
  assign n9628 = n1121 & ~n9627 ;
  assign n9629 = ~n1925 & n9173 ;
  assign n9630 = ~n2073 & n9629 ;
  assign n9631 = n1307 | n4588 ;
  assign n9632 = n2372 | n9631 ;
  assign n9633 = ~n9630 & n9632 ;
  assign n9634 = n5050 & n9633 ;
  assign n9635 = n1371 & n8360 ;
  assign n9636 = ( x239 & n4438 ) | ( x239 & n9635 ) | ( n4438 & n9635 ) ;
  assign n9637 = n7454 ^ n1254 ^ 1'b0 ;
  assign n9638 = ~n1931 & n9637 ;
  assign n9639 = n727 | n3179 ;
  assign n9640 = n9638 | n9639 ;
  assign n9641 = n444 | n7338 ;
  assign n9642 = n1820 | n4764 ;
  assign n9643 = n8311 & n9642 ;
  assign n9644 = x248 & n3908 ;
  assign n9645 = n3429 & ~n9644 ;
  assign n9646 = n9645 ^ n5465 ^ 1'b0 ;
  assign n9647 = n4424 & ~n5797 ;
  assign n9648 = n9647 ^ n1802 ^ 1'b0 ;
  assign n9649 = n8682 & n9648 ;
  assign n9650 = n4519 & ~n9649 ;
  assign n9651 = n9650 ^ n2785 ^ 1'b0 ;
  assign n9652 = n1435 & ~n5274 ;
  assign n9653 = n1820 & n3339 ;
  assign n9654 = ~n9652 & n9653 ;
  assign n9655 = n5782 ^ n3589 ^ 1'b0 ;
  assign n9656 = n1393 & n2064 ;
  assign n9657 = ~n9655 & n9656 ;
  assign n9658 = n946 & ~n8487 ;
  assign n9659 = n9658 ^ n3228 ^ 1'b0 ;
  assign n9660 = x16 & ~n2898 ;
  assign n9661 = n9659 & ~n9660 ;
  assign n9662 = n5440 ^ n3424 ^ 1'b0 ;
  assign n9663 = ~n920 & n6722 ;
  assign n9664 = n7289 & ~n9663 ;
  assign n9665 = n6138 & ~n6695 ;
  assign n9666 = ~n1185 & n1861 ;
  assign n9667 = n9666 ^ x231 ^ 1'b0 ;
  assign n9668 = n6400 & ~n9667 ;
  assign n9669 = n9668 ^ n6405 ^ 1'b0 ;
  assign n9670 = ( n385 & n2500 ) | ( n385 & n9669 ) | ( n2500 & n9669 ) ;
  assign n9671 = ~n426 & n2577 ;
  assign n9672 = n9671 ^ n2936 ^ 1'b0 ;
  assign n9673 = n9672 ^ n1004 ^ 1'b0 ;
  assign n9674 = n4865 & ~n9673 ;
  assign n9676 = n3989 & ~n8007 ;
  assign n9677 = n2582 & ~n9676 ;
  assign n9678 = n529 & n9677 ;
  assign n9675 = n769 & n3810 ;
  assign n9679 = n9678 ^ n9675 ^ 1'b0 ;
  assign n9680 = n6566 | n7025 ;
  assign n9683 = n4566 ^ n680 ^ 1'b0 ;
  assign n9682 = ~n1680 & n4635 ;
  assign n9684 = n9683 ^ n9682 ^ 1'b0 ;
  assign n9681 = n5461 & n5763 ;
  assign n9685 = n9684 ^ n9681 ^ 1'b0 ;
  assign n9686 = ~n9680 & n9685 ;
  assign n9687 = n7304 & ~n9686 ;
  assign n9688 = ( ~n8307 & n9679 ) | ( ~n8307 & n9687 ) | ( n9679 & n9687 ) ;
  assign n9689 = n1568 & ~n1741 ;
  assign n9690 = n9689 ^ n4107 ^ 1'b0 ;
  assign n9691 = ~n420 & n9690 ;
  assign n9692 = ~n263 & n3099 ;
  assign n9693 = n2714 ^ n593 ^ 1'b0 ;
  assign n9694 = n4574 | n6902 ;
  assign n9695 = n668 & n2443 ;
  assign n9696 = n9695 ^ n5119 ^ n3201 ;
  assign n9697 = n9696 ^ n9513 ^ 1'b0 ;
  assign n9698 = n8578 | n9697 ;
  assign n9699 = n6110 | n7947 ;
  assign n9700 = n3845 & n6813 ;
  assign n9701 = n7658 ^ n387 ^ 1'b0 ;
  assign n9702 = n6822 & n9701 ;
  assign n9703 = n8114 ^ n7379 ^ n6471 ;
  assign n9704 = n7967 ^ n3930 ^ 1'b0 ;
  assign n9705 = n7923 ^ n4887 ^ 1'b0 ;
  assign n9708 = n8580 ^ x13 ^ 1'b0 ;
  assign n9706 = ~x213 & n3728 ;
  assign n9707 = n2167 & ~n9706 ;
  assign n9709 = n9708 ^ n9707 ^ 1'b0 ;
  assign n9710 = ~n2255 & n4178 ;
  assign n9711 = n9710 ^ n9492 ^ 1'b0 ;
  assign n9714 = n1223 ^ n992 ^ 1'b0 ;
  assign n9715 = n657 | n9714 ;
  assign n9712 = n7456 ^ n5551 ^ 1'b0 ;
  assign n9713 = n4142 & ~n9712 ;
  assign n9716 = n9715 ^ n9713 ^ 1'b0 ;
  assign n9717 = n946 & ~n9716 ;
  assign n9721 = n2785 ^ n426 ^ 1'b0 ;
  assign n9718 = n1593 & ~n4568 ;
  assign n9719 = n761 & n9718 ;
  assign n9720 = n2763 & ~n9719 ;
  assign n9722 = n9721 ^ n9720 ^ n6311 ;
  assign n9723 = n389 | n1125 ;
  assign n9724 = n9722 | n9723 ;
  assign n9725 = n2949 ^ x205 ^ x159 ;
  assign n9726 = n4411 ^ n1175 ^ 1'b0 ;
  assign n9727 = n9725 | n9726 ;
  assign n9728 = n9727 ^ n6676 ^ n973 ;
  assign n9729 = ~n4883 & n7773 ;
  assign n9730 = ~n3635 & n8305 ;
  assign n9731 = ~n2827 & n5965 ;
  assign n9732 = ~n615 & n6745 ;
  assign n9733 = n1562 & n9732 ;
  assign n9734 = n3696 & ~n6827 ;
  assign n9735 = n9733 & ~n9734 ;
  assign n9736 = n9731 | n9735 ;
  assign n9737 = n8822 ^ n5475 ^ 1'b0 ;
  assign n9738 = n6361 & ~n9737 ;
  assign n9739 = ~n518 & n1912 ;
  assign n9740 = n3795 & ~n8276 ;
  assign n9742 = n3411 ^ n1786 ^ 1'b0 ;
  assign n9741 = n3226 & n5709 ;
  assign n9743 = n9742 ^ n9741 ^ 1'b0 ;
  assign n9744 = n9740 & n9743 ;
  assign n9745 = n5255 & ~n5640 ;
  assign n9746 = x212 & ~n1369 ;
  assign n9747 = n3576 & ~n5237 ;
  assign n9748 = n6120 & n9747 ;
  assign n9749 = ~n9746 & n9748 ;
  assign n9757 = n7115 ^ n3770 ^ 1'b0 ;
  assign n9758 = n1817 | n9757 ;
  assign n9754 = n2770 ^ x156 ^ 1'b0 ;
  assign n9750 = n665 ^ x187 ^ 1'b0 ;
  assign n9751 = x198 & ~n9750 ;
  assign n9752 = n638 & ~n5151 ;
  assign n9753 = ~n9751 & n9752 ;
  assign n9755 = n9754 ^ n9753 ^ 1'b0 ;
  assign n9756 = ~n3722 & n9755 ;
  assign n9759 = n9758 ^ n9756 ^ 1'b0 ;
  assign n9760 = ~n1043 & n7655 ;
  assign n9761 = n9760 ^ n9014 ^ 1'b0 ;
  assign n9762 = n1714 & n4787 ;
  assign n9763 = n7232 | n9762 ;
  assign n9764 = n8351 | n9763 ;
  assign n9765 = ~n5903 & n7291 ;
  assign n9766 = ~n7846 & n9765 ;
  assign n9767 = n2176 & ~n9766 ;
  assign n9768 = n7450 & n9767 ;
  assign n9769 = n9768 ^ n8471 ^ 1'b0 ;
  assign n9770 = n4484 | n6604 ;
  assign n9771 = n4665 | n5229 ;
  assign n9772 = n7286 & ~n9727 ;
  assign n9773 = ~n9771 & n9772 ;
  assign n9774 = ~n1400 & n9773 ;
  assign n9776 = n3744 & ~n4238 ;
  assign n9777 = n9776 ^ n6952 ^ 1'b0 ;
  assign n9775 = n966 ^ n597 ^ 1'b0 ;
  assign n9778 = n9777 ^ n9775 ^ 1'b0 ;
  assign n9779 = n7558 ^ n3586 ^ 1'b0 ;
  assign n9780 = n9779 ^ n7799 ^ 1'b0 ;
  assign n9781 = n8025 ^ n5418 ^ 1'b0 ;
  assign n9782 = n9144 ^ x63 ^ 1'b0 ;
  assign n9786 = n3593 & n4417 ;
  assign n9787 = ~n6186 & n9786 ;
  assign n9788 = n9787 ^ n5921 ^ 1'b0 ;
  assign n9789 = n9788 ^ n2119 ^ 1'b0 ;
  assign n9790 = n366 & ~n9789 ;
  assign n9783 = n436 | n1309 ;
  assign n9784 = ~n919 & n4114 ;
  assign n9785 = n9783 | n9784 ;
  assign n9791 = n9790 ^ n9785 ^ 1'b0 ;
  assign n9792 = n2538 & n5277 ;
  assign n9793 = n9792 ^ n6821 ^ n2545 ;
  assign n9794 = n2252 & n4837 ;
  assign n9796 = n8657 ^ n5183 ^ 1'b0 ;
  assign n9797 = n3195 & n9796 ;
  assign n9798 = ~n1776 & n9797 ;
  assign n9795 = ~n1709 & n7910 ;
  assign n9799 = n9798 ^ n9795 ^ 1'b0 ;
  assign n9800 = n4117 & ~n5604 ;
  assign n9801 = n3036 & n9800 ;
  assign n9802 = n8200 ^ n860 ^ 1'b0 ;
  assign n9805 = n5385 ^ n4521 ^ 1'b0 ;
  assign n9806 = n2992 & ~n9805 ;
  assign n9803 = ~n4316 & n8956 ;
  assign n9804 = ~n4108 & n9803 ;
  assign n9807 = n9806 ^ n9804 ^ 1'b0 ;
  assign n9808 = n2271 | n9807 ;
  assign n9809 = n9771 ^ n1633 ^ 1'b0 ;
  assign n9812 = x96 & n920 ;
  assign n9813 = n733 & n9812 ;
  assign n9810 = n1681 ^ n523 ^ 1'b0 ;
  assign n9811 = n933 & n9810 ;
  assign n9814 = n9813 ^ n9811 ^ n1338 ;
  assign n9815 = n9809 & n9814 ;
  assign n9816 = n3586 ^ n367 ^ 1'b0 ;
  assign n9817 = n9816 ^ n7864 ^ 1'b0 ;
  assign n9818 = n4805 ^ n2234 ^ 1'b0 ;
  assign n9819 = ~n9817 & n9818 ;
  assign n9820 = x100 & ~n5667 ;
  assign n9821 = n8026 & n9820 ;
  assign n9822 = x27 & n880 ;
  assign n9823 = n8067 & n9822 ;
  assign n9824 = ~n1654 & n9823 ;
  assign n9825 = n3642 & ~n4169 ;
  assign n9826 = ~n9824 & n9825 ;
  assign n9827 = n4555 ^ n1633 ^ 1'b0 ;
  assign n9828 = n2986 & ~n3695 ;
  assign n9829 = n6687 ^ n2265 ^ 1'b0 ;
  assign n9830 = ~n423 & n7384 ;
  assign n9831 = n6432 ^ n4503 ^ 1'b0 ;
  assign n9832 = ~n3571 & n9831 ;
  assign n9833 = ~n589 & n3123 ;
  assign n9834 = x0 & n9833 ;
  assign n9835 = ~n9771 & n9834 ;
  assign n9836 = ~n3701 & n4679 ;
  assign n9837 = ( n296 & n4310 ) | ( n296 & n9836 ) | ( n4310 & n9836 ) ;
  assign n9838 = ~x195 & n3493 ;
  assign n9839 = ~n6367 & n9838 ;
  assign n9840 = n3822 & ~n9839 ;
  assign n9841 = n1312 & ~n2139 ;
  assign n9843 = n4105 ^ n908 ^ 1'b0 ;
  assign n9844 = n432 | n9843 ;
  assign n9845 = n4937 ^ n4498 ^ 1'b0 ;
  assign n9846 = n9844 | n9845 ;
  assign n9842 = n2804 ^ x128 ^ 1'b0 ;
  assign n9847 = n9846 ^ n9842 ^ 1'b0 ;
  assign n9848 = n8346 ^ n7826 ^ n3685 ;
  assign n9849 = n2153 & n4421 ;
  assign n9850 = ~n6228 & n9849 ;
  assign n9851 = n2595 | n4004 ;
  assign n9852 = n9851 ^ n3557 ^ 1'b0 ;
  assign n9853 = ( n2644 & n5342 ) | ( n2644 & n7502 ) | ( n5342 & n7502 ) ;
  assign n9854 = n5336 & ~n9853 ;
  assign n9855 = ~n6972 & n9854 ;
  assign n9856 = n6466 ^ n2174 ^ n1134 ;
  assign n9857 = n1180 & ~n9856 ;
  assign n9858 = n4321 & n9857 ;
  assign n9859 = ~n7307 & n9858 ;
  assign n9860 = n2477 & n6874 ;
  assign n9861 = n9860 ^ n2043 ^ 1'b0 ;
  assign n9862 = n6793 | n9861 ;
  assign n9863 = n2835 & n4849 ;
  assign n9864 = n1919 & n9863 ;
  assign n9865 = n1730 & ~n8455 ;
  assign n9866 = n917 ^ n467 ^ 1'b0 ;
  assign n9867 = n9866 ^ n6574 ^ 1'b0 ;
  assign n9868 = n1301 & n5544 ;
  assign n9869 = n9868 ^ n2509 ^ 1'b0 ;
  assign n9870 = ~n1255 & n9869 ;
  assign n9871 = n9870 ^ n9048 ^ 1'b0 ;
  assign n9872 = n2148 & ~n9871 ;
  assign n9873 = n3853 & n4122 ;
  assign n9874 = n5720 ^ n4163 ^ 1'b0 ;
  assign n9878 = ~n333 & n5448 ;
  assign n9875 = n2577 & n9792 ;
  assign n9876 = n9875 ^ n984 ^ 1'b0 ;
  assign n9877 = n6761 | n9876 ;
  assign n9879 = n9878 ^ n9877 ^ 1'b0 ;
  assign n9880 = n5961 & ~n8930 ;
  assign n9881 = n9880 ^ n5395 ^ 1'b0 ;
  assign n9882 = n3046 & ~n9881 ;
  assign n9883 = n2995 & n9882 ;
  assign n9884 = n5061 ^ n3837 ^ 1'b0 ;
  assign n9885 = n9883 | n9884 ;
  assign n9886 = n3508 & ~n4662 ;
  assign n9887 = n6300 & n9886 ;
  assign n9888 = n8436 ^ n6991 ^ 1'b0 ;
  assign n9889 = n4197 | n9888 ;
  assign n9890 = n7407 & n7700 ;
  assign n9891 = ~n2271 & n4528 ;
  assign n9892 = n9891 ^ n5452 ^ 1'b0 ;
  assign n9893 = n6770 ^ n2747 ^ 1'b0 ;
  assign n9894 = ~n3086 & n9893 ;
  assign n9895 = ( n688 & n1326 ) | ( n688 & ~n2646 ) | ( n1326 & ~n2646 ) ;
  assign n9896 = n9895 ^ n3102 ^ 1'b0 ;
  assign n9897 = n9644 | n9896 ;
  assign n9898 = n4069 | n9897 ;
  assign n9899 = n7979 | n9898 ;
  assign n9900 = n7745 & ~n9899 ;
  assign n9902 = n3000 & ~n7700 ;
  assign n9903 = n9902 ^ n7838 ^ 1'b0 ;
  assign n9901 = n7366 ^ n5452 ^ 1'b0 ;
  assign n9904 = n9903 ^ n9901 ^ x110 ;
  assign n9905 = n2552 ^ n1558 ^ 1'b0 ;
  assign n9906 = n9905 ^ n3551 ^ 1'b0 ;
  assign n9907 = n6291 | n9260 ;
  assign n9908 = n8237 ^ n7109 ^ 1'b0 ;
  assign n9909 = n9907 & ~n9908 ;
  assign n9910 = n5067 ^ x128 ^ 1'b0 ;
  assign n9911 = n3114 | n9910 ;
  assign n9912 = ~n9130 & n9250 ;
  assign n9913 = ~n2178 & n8337 ;
  assign n9914 = n9913 ^ x25 ^ 1'b0 ;
  assign n9915 = ~n1780 & n7141 ;
  assign n9916 = n9914 & n9915 ;
  assign n9917 = n9916 ^ n9281 ^ 1'b0 ;
  assign n9918 = ~n571 & n3588 ;
  assign n9919 = n9918 ^ n7557 ^ 1'b0 ;
  assign n9920 = n7830 & ~n9919 ;
  assign n9921 = n4450 ^ n1172 ^ 1'b0 ;
  assign n9922 = n9797 ^ n6786 ^ n4451 ;
  assign n9923 = n1335 & ~n2473 ;
  assign n9924 = ~n6121 & n9923 ;
  assign n9925 = n4132 & n9419 ;
  assign n9926 = n9925 ^ n3190 ^ 1'b0 ;
  assign n9927 = n3642 | n7077 ;
  assign n9928 = n8512 ^ n6746 ^ 1'b0 ;
  assign n9929 = n7737 & ~n9928 ;
  assign n9930 = ( ~n1211 & n3499 ) | ( ~n1211 & n3915 ) | ( n3499 & n3915 ) ;
  assign n9931 = n3855 & ~n9930 ;
  assign n9932 = n7219 ^ n2122 ^ 1'b0 ;
  assign n9933 = n9931 | n9932 ;
  assign n9934 = n4025 & ~n8620 ;
  assign n9935 = ~n9933 & n9934 ;
  assign n9936 = n4673 ^ n1835 ^ n1130 ;
  assign n9937 = ~n1119 & n1829 ;
  assign n9938 = ~n547 & n9937 ;
  assign n9939 = n457 | n6826 ;
  assign n9940 = n9938 & ~n9939 ;
  assign n9941 = n6854 | n9940 ;
  assign n9942 = n9941 ^ n8277 ^ 1'b0 ;
  assign n9943 = n2366 & ~n3258 ;
  assign n9944 = n9943 ^ n2614 ^ 1'b0 ;
  assign n9945 = n3884 ^ n2163 ^ 1'b0 ;
  assign n9946 = n2473 | n9945 ;
  assign n9947 = n2065 | n9946 ;
  assign n9948 = n9947 ^ n6910 ^ 1'b0 ;
  assign n9949 = n4827 & n8784 ;
  assign n9950 = n4851 ^ n3932 ^ x27 ;
  assign n9951 = ( n613 & n2504 ) | ( n613 & n3039 ) | ( n2504 & n3039 ) ;
  assign n9952 = n4062 & n5600 ;
  assign n9953 = ~n9951 & n9952 ;
  assign n9954 = n2684 ^ n516 ^ 1'b0 ;
  assign n9955 = n3348 | n9954 ;
  assign n9956 = n9955 ^ n4150 ^ 1'b0 ;
  assign n9957 = n3012 & ~n9956 ;
  assign n9958 = n996 ^ n806 ^ n699 ;
  assign n9959 = n2830 & ~n9958 ;
  assign n9960 = n821 & n9959 ;
  assign n9961 = n9960 ^ n1326 ^ 1'b0 ;
  assign n9962 = n262 & ~n9739 ;
  assign n9963 = ~n9961 & n9962 ;
  assign n9964 = n7976 ^ n7449 ^ n4878 ;
  assign n9965 = n9964 ^ n3848 ^ 1'b0 ;
  assign n9966 = n4346 | n5758 ;
  assign n9967 = n7024 | n9966 ;
  assign n9968 = n6292 ^ n5874 ^ n4846 ;
  assign n9969 = n1919 & ~n5589 ;
  assign n9970 = n9969 ^ n8291 ^ 1'b0 ;
  assign n9971 = ( n9967 & n9968 ) | ( n9967 & n9970 ) | ( n9968 & n9970 ) ;
  assign n9982 = n5310 ^ n3610 ^ 1'b0 ;
  assign n9972 = x142 & ~n2748 ;
  assign n9973 = ~n268 & n9972 ;
  assign n9974 = n9973 ^ n2139 ^ 1'b0 ;
  assign n9975 = n9974 ^ n6454 ^ 1'b0 ;
  assign n9976 = ~n2724 & n9975 ;
  assign n9977 = n9976 ^ n5888 ^ n5742 ;
  assign n9978 = n961 & n9175 ;
  assign n9979 = ~n7508 & n9978 ;
  assign n9980 = n9977 | n9979 ;
  assign n9981 = n6887 | n9980 ;
  assign n9983 = n9982 ^ n9981 ^ 1'b0 ;
  assign n9984 = n2360 & n9983 ;
  assign n9985 = n3298 & n9759 ;
  assign n9986 = n5469 | n7430 ;
  assign n9987 = n5391 ^ x229 ^ 1'b0 ;
  assign n9988 = n9987 ^ n8730 ^ n5505 ;
  assign n9989 = n9492 & ~n9988 ;
  assign n9990 = n6186 ^ n5497 ^ n1846 ;
  assign n9994 = n7423 ^ n5067 ^ 1'b0 ;
  assign n9991 = n589 | n2890 ;
  assign n9992 = n9991 ^ n3884 ^ 1'b0 ;
  assign n9993 = n9992 ^ n7632 ^ 1'b0 ;
  assign n9995 = n9994 ^ n9993 ^ 1'b0 ;
  assign n9996 = ~n720 & n1619 ;
  assign n9997 = ~n7521 & n9996 ;
  assign n9998 = n2741 & n9997 ;
  assign n9999 = ~n2287 & n6963 ;
  assign n10000 = n3856 & ~n6313 ;
  assign n10001 = n10000 ^ n4187 ^ n2224 ;
  assign n10002 = ~n2502 & n6576 ;
  assign n10003 = n10002 ^ n9012 ^ 1'b0 ;
  assign n10004 = n5616 ^ n1053 ^ 1'b0 ;
  assign n10005 = x196 & ~n2602 ;
  assign n10006 = ~n5407 & n10005 ;
  assign n10007 = ( n1611 & n4793 ) | ( n1611 & n6930 ) | ( n4793 & n6930 ) ;
  assign n10008 = ( n4215 & n10006 ) | ( n4215 & ~n10007 ) | ( n10006 & ~n10007 ) ;
  assign n10009 = n10008 ^ n7361 ^ n686 ;
  assign n10010 = n4565 ^ n2267 ^ n481 ;
  assign n10011 = n6318 & ~n10010 ;
  assign n10012 = n5648 & n10011 ;
  assign n10013 = n10012 ^ n1142 ^ 1'b0 ;
  assign n10014 = n2369 & ~n10013 ;
  assign n10015 = n7464 & n10014 ;
  assign n10016 = n2018 | n3215 ;
  assign n10017 = ~n2813 & n10016 ;
  assign n10018 = n10017 ^ n769 ^ 1'b0 ;
  assign n10019 = n4139 | n10018 ;
  assign n10024 = n597 & ~n4566 ;
  assign n10021 = n3420 ^ n1645 ^ 1'b0 ;
  assign n10022 = ~n1544 & n10021 ;
  assign n10020 = n1377 & n7597 ;
  assign n10023 = n10022 ^ n10020 ^ 1'b0 ;
  assign n10025 = n10024 ^ n10023 ^ 1'b0 ;
  assign n10026 = n1739 | n10025 ;
  assign n10027 = n7989 ^ n1315 ^ 1'b0 ;
  assign n10028 = n5237 & ~n10027 ;
  assign n10029 = n2735 & n6930 ;
  assign n10030 = n10029 ^ n375 ^ 1'b0 ;
  assign n10031 = n575 & ~n1245 ;
  assign n10032 = n10031 ^ n9848 ^ 1'b0 ;
  assign n10033 = n10030 | n10032 ;
  assign n10034 = n5287 & ~n6386 ;
  assign n10037 = ~n270 & n3087 ;
  assign n10038 = n10037 ^ n7185 ^ 1'b0 ;
  assign n10039 = n2443 & ~n10038 ;
  assign n10035 = ~n8275 & n9191 ;
  assign n10036 = n9823 & n10035 ;
  assign n10040 = n10039 ^ n10036 ^ n6018 ;
  assign n10041 = x169 & n3723 ;
  assign n10042 = n5898 ^ n2646 ^ 1'b0 ;
  assign n10043 = n10042 ^ n7148 ^ 1'b0 ;
  assign n10044 = n10041 & n10043 ;
  assign n10045 = x13 & x247 ;
  assign n10046 = n10045 ^ n529 ^ 1'b0 ;
  assign n10047 = n3362 & ~n10046 ;
  assign n10048 = n927 | n1126 ;
  assign n10049 = n10048 ^ n7301 ^ n4703 ;
  assign n10061 = n809 & n4999 ;
  assign n10062 = n10061 ^ n1909 ^ 1'b0 ;
  assign n10050 = n5571 ^ n1416 ^ 1'b0 ;
  assign n10051 = ~n3081 & n10050 ;
  assign n10054 = n449 ^ n328 ^ 1'b0 ;
  assign n10055 = x26 & n10054 ;
  assign n10056 = n486 & n5005 ;
  assign n10057 = n10055 & n10056 ;
  assign n10052 = x40 & n1726 ;
  assign n10053 = n4654 & n10052 ;
  assign n10058 = n10057 ^ n10053 ^ 1'b0 ;
  assign n10059 = n10051 & ~n10058 ;
  assign n10060 = n4296 & n10059 ;
  assign n10063 = n10062 ^ n10060 ^ 1'b0 ;
  assign n10064 = n3627 ^ x114 ^ 1'b0 ;
  assign n10065 = n899 | n7094 ;
  assign n10066 = n882 & ~n2848 ;
  assign n10067 = n1989 & n4058 ;
  assign n10068 = n10067 ^ x180 ^ 1'b0 ;
  assign n10069 = ( n4704 & n6352 ) | ( n4704 & ~n10068 ) | ( n6352 & ~n10068 ) ;
  assign n10070 = n882 & ~n10069 ;
  assign n10071 = n5007 ^ n2287 ^ 1'b0 ;
  assign n10072 = x73 & n673 ;
  assign n10073 = n2092 | n3765 ;
  assign n10074 = n10072 | n10073 ;
  assign n10075 = n10071 & n10074 ;
  assign n10076 = n2387 | n6655 ;
  assign n10077 = n10076 ^ n8783 ^ 1'b0 ;
  assign n10078 = n7958 & n10077 ;
  assign n10079 = n810 & n10078 ;
  assign n10080 = n3362 & ~n10079 ;
  assign n10081 = n10080 ^ n1541 ^ 1'b0 ;
  assign n10082 = n3038 ^ n1979 ^ 1'b0 ;
  assign n10083 = ~n3486 & n10082 ;
  assign n10084 = n3078 & n10083 ;
  assign n10085 = n3257 & n4890 ;
  assign n10086 = n5580 | n10085 ;
  assign n10087 = n915 & n1111 ;
  assign n10088 = n10087 ^ n5270 ^ 1'b0 ;
  assign n10089 = ( n908 & ~n1023 ) | ( n908 & n4502 ) | ( ~n1023 & n4502 ) ;
  assign n10090 = n10089 ^ n3978 ^ n2937 ;
  assign n10091 = n10090 ^ n2508 ^ 1'b0 ;
  assign n10092 = n5290 | n10091 ;
  assign n10093 = n8945 & ~n10092 ;
  assign n10094 = n3059 & n10093 ;
  assign n10095 = n3326 & n9951 ;
  assign n10096 = n1185 | n7932 ;
  assign n10097 = n425 & n3613 ;
  assign n10098 = x123 & n2801 ;
  assign n10099 = ~n10097 & n10098 ;
  assign n10100 = n4232 & ~n5969 ;
  assign n10101 = n8860 ^ n7019 ^ 1'b0 ;
  assign n10102 = n585 | n6674 ;
  assign n10103 = n5532 & n5554 ;
  assign n10104 = n7103 & ~n10103 ;
  assign n10105 = n5896 & n10104 ;
  assign n10106 = n9024 ^ n6553 ^ 1'b0 ;
  assign n10107 = n3416 & ~n4029 ;
  assign n10108 = n10107 ^ n1161 ^ 1'b0 ;
  assign n10109 = n3574 & ~n10108 ;
  assign n10110 = ~n1300 & n10109 ;
  assign n10111 = n10110 ^ n3195 ^ 1'b0 ;
  assign n10112 = n2712 ^ n1699 ^ 1'b0 ;
  assign n10113 = n3321 & ~n10112 ;
  assign n10114 = n2367 ^ n666 ^ 1'b0 ;
  assign n10115 = n776 | n3941 ;
  assign n10116 = n3571 & ~n10115 ;
  assign n10117 = n1512 & ~n9355 ;
  assign n10118 = ~n3999 & n10117 ;
  assign n10119 = n10118 ^ n5097 ^ 1'b0 ;
  assign n10120 = ~n10116 & n10119 ;
  assign n10121 = ~n8738 & n10120 ;
  assign n10122 = n10121 ^ n6307 ^ 1'b0 ;
  assign n10123 = n1614 & n6633 ;
  assign n10124 = ~n9686 & n10123 ;
  assign n10125 = n9100 ^ n8053 ^ 1'b0 ;
  assign n10126 = n6339 & n10125 ;
  assign n10127 = ~n6508 & n10126 ;
  assign n10128 = n1620 & n2964 ;
  assign n10129 = n10128 ^ n3886 ^ 1'b0 ;
  assign n10130 = n9961 ^ n9864 ^ 1'b0 ;
  assign n10131 = n9083 & n10130 ;
  assign n10132 = n10131 ^ n2961 ^ 1'b0 ;
  assign n10133 = n4676 & ~n10132 ;
  assign n10134 = n618 & ~n908 ;
  assign n10135 = n10134 ^ n4976 ^ 1'b0 ;
  assign n10136 = n5250 & ~n9468 ;
  assign n10137 = n10136 ^ n1756 ^ 1'b0 ;
  assign n10138 = n2944 | n5004 ;
  assign n10139 = n10138 ^ x48 ^ 1'b0 ;
  assign n10140 = n10139 ^ n8026 ^ 1'b0 ;
  assign n10141 = n10140 ^ n4011 ^ 1'b0 ;
  assign n10142 = n3337 | n10141 ;
  assign n10143 = n2668 & n10142 ;
  assign n10145 = ( n518 & n4400 ) | ( n518 & n7358 ) | ( n4400 & n7358 ) ;
  assign n10144 = n4468 ^ n2287 ^ 1'b0 ;
  assign n10146 = n10145 ^ n10144 ^ n2108 ;
  assign n10147 = n1921 & ~n10146 ;
  assign n10163 = ~n1198 & n3569 ;
  assign n10164 = n10163 ^ x211 ^ 1'b0 ;
  assign n10165 = ( n5362 & n6739 ) | ( n5362 & ~n10164 ) | ( n6739 & ~n10164 ) ;
  assign n10160 = ~n1193 & n1867 ;
  assign n10161 = n746 & n10160 ;
  assign n10154 = n4325 & ~n5602 ;
  assign n10155 = n10154 ^ n6483 ^ 1'b0 ;
  assign n10156 = n3981 & n10155 ;
  assign n10157 = n10156 ^ n1716 ^ 1'b0 ;
  assign n10149 = n1628 ^ n274 ^ 1'b0 ;
  assign n10148 = n4126 & n6067 ;
  assign n10150 = n10149 ^ n10148 ^ n1952 ;
  assign n10151 = ~n3555 & n5393 ;
  assign n10152 = n3552 & n10151 ;
  assign n10153 = n10150 & ~n10152 ;
  assign n10158 = n10157 ^ n10153 ^ 1'b0 ;
  assign n10159 = ~n6937 & n10158 ;
  assign n10162 = n10161 ^ n10159 ^ 1'b0 ;
  assign n10166 = n10165 ^ n10162 ^ 1'b0 ;
  assign n10167 = ~n1956 & n10166 ;
  assign n10168 = n8952 ^ n3110 ^ 1'b0 ;
  assign n10169 = n8990 | n10168 ;
  assign n10171 = n1708 ^ n780 ^ 1'b0 ;
  assign n10172 = n277 | n10171 ;
  assign n10170 = n492 ^ n274 ^ 1'b0 ;
  assign n10173 = n10172 ^ n10170 ^ 1'b0 ;
  assign n10174 = ~n6873 & n10173 ;
  assign n10175 = n10174 ^ n8912 ^ 1'b0 ;
  assign n10176 = ( ~x243 & n1671 ) | ( ~x243 & n5563 ) | ( n1671 & n5563 ) ;
  assign n10177 = ( x158 & ~x237 ) | ( x158 & n10176 ) | ( ~x237 & n10176 ) ;
  assign n10178 = n815 & n6844 ;
  assign n10179 = n8756 ^ n7298 ^ 1'b0 ;
  assign n10180 = n3875 & ~n5365 ;
  assign n10186 = ~n1705 & n2007 ;
  assign n10187 = n10186 ^ x132 ^ 1'b0 ;
  assign n10188 = n7111 | n10187 ;
  assign n10189 = n10188 ^ n5921 ^ 1'b0 ;
  assign n10181 = n1900 & ~n6991 ;
  assign n10182 = n10181 ^ n6745 ^ 1'b0 ;
  assign n10183 = n5581 ^ n3288 ^ 1'b0 ;
  assign n10184 = ~n10182 & n10183 ;
  assign n10185 = n1077 & n10184 ;
  assign n10190 = n10189 ^ n10185 ^ 1'b0 ;
  assign n10191 = ( n432 & ~n1999 ) | ( n432 & n2083 ) | ( ~n1999 & n2083 ) ;
  assign n10192 = n5815 ^ n2592 ^ 1'b0 ;
  assign n10193 = n9186 | n10192 ;
  assign n10194 = n10191 & n10193 ;
  assign n10195 = n1373 & ~n4238 ;
  assign n10196 = ~n5187 & n10195 ;
  assign n10197 = ~n615 & n2328 ;
  assign n10198 = ~x210 & n10197 ;
  assign n10199 = n7936 ^ n4021 ^ 1'b0 ;
  assign n10200 = ~n10198 & n10199 ;
  assign n10201 = ( x127 & n8249 ) | ( x127 & ~n10200 ) | ( n8249 & ~n10200 ) ;
  assign n10202 = n5976 & ~n10201 ;
  assign n10203 = n3830 & n10202 ;
  assign n10204 = n7243 | n10203 ;
  assign n10205 = n10196 & ~n10204 ;
  assign n10206 = n1083 & ~n5130 ;
  assign n10207 = n10206 ^ n3608 ^ 1'b0 ;
  assign n10208 = n8728 ^ n2798 ^ n904 ;
  assign n10209 = ~n406 & n10208 ;
  assign n10214 = n9806 ^ n7387 ^ 1'b0 ;
  assign n10215 = n5069 | n10214 ;
  assign n10216 = ( n535 & n3174 ) | ( n535 & n10215 ) | ( n3174 & n10215 ) ;
  assign n10217 = n10216 ^ n6023 ^ 1'b0 ;
  assign n10210 = ~n797 & n3073 ;
  assign n10211 = n10210 ^ n361 ^ 1'b0 ;
  assign n10212 = n10211 ^ n1019 ^ 1'b0 ;
  assign n10213 = n8225 | n10212 ;
  assign n10218 = n10217 ^ n10213 ^ 1'b0 ;
  assign n10219 = n3331 | n4699 ;
  assign n10220 = n2925 & ~n9255 ;
  assign n10221 = ~n10219 & n10220 ;
  assign n10222 = n3677 ^ n991 ^ n961 ;
  assign n10223 = ( n1193 & n3119 ) | ( n1193 & ~n10222 ) | ( n3119 & ~n10222 ) ;
  assign n10228 = n2523 ^ n1114 ^ 1'b0 ;
  assign n10229 = n4894 & n10228 ;
  assign n10230 = n359 & ~n4663 ;
  assign n10231 = ~n10229 & n10230 ;
  assign n10224 = n2332 ^ n274 ^ 1'b0 ;
  assign n10225 = ~n5435 & n10224 ;
  assign n10226 = ~n4553 & n10225 ;
  assign n10227 = ~n6416 & n10226 ;
  assign n10232 = n10231 ^ n10227 ^ 1'b0 ;
  assign n10233 = n3070 & ~n8268 ;
  assign n10234 = n10233 ^ n6042 ^ 1'b0 ;
  assign n10235 = n2334 & n10234 ;
  assign n10236 = n1791 & n10235 ;
  assign n10237 = n4058 | n10236 ;
  assign n10238 = n7532 ^ n2013 ^ 1'b0 ;
  assign n10239 = ~n6563 & n10238 ;
  assign n10240 = ~n1599 & n10239 ;
  assign n10241 = ~n4023 & n6116 ;
  assign n10242 = n5742 ^ n4949 ^ 1'b0 ;
  assign n10243 = n10241 & ~n10242 ;
  assign n10244 = ~n3948 & n7069 ;
  assign n10245 = n8395 ^ n1855 ^ 1'b0 ;
  assign n10246 = n6838 & n10245 ;
  assign n10247 = n10244 & ~n10246 ;
  assign n10248 = n1393 & ~n10247 ;
  assign n10249 = n1735 ^ n266 ^ 1'b0 ;
  assign n10250 = n10249 ^ n1676 ^ 1'b0 ;
  assign n10251 = n10250 ^ n3966 ^ 1'b0 ;
  assign n10252 = n3651 & ~n10251 ;
  assign n10253 = n10252 ^ n7557 ^ 1'b0 ;
  assign n10254 = n5210 ^ n2171 ^ 1'b0 ;
  assign n10255 = x73 & x147 ;
  assign n10256 = ~n5163 & n10255 ;
  assign n10257 = n3957 & ~n9574 ;
  assign n10258 = n10257 ^ n10036 ^ 1'b0 ;
  assign n10259 = ~x48 & n1634 ;
  assign n10260 = n2587 | n6363 ;
  assign n10261 = n3651 | n10260 ;
  assign n10262 = n3772 & n10261 ;
  assign n10263 = n4021 & n8512 ;
  assign n10264 = n10263 ^ n4487 ^ 1'b0 ;
  assign n10265 = n9074 ^ n5849 ^ 1'b0 ;
  assign n10266 = n10264 & ~n10265 ;
  assign n10267 = n3957 & ~n10266 ;
  assign n10268 = n627 | n2006 ;
  assign n10269 = x81 & ~n10268 ;
  assign n10270 = ~n4049 & n10269 ;
  assign n10271 = n10270 ^ n2473 ^ 1'b0 ;
  assign n10272 = n10271 ^ n7071 ^ 1'b0 ;
  assign n10273 = ( n1332 & n3933 ) | ( n1332 & n7163 ) | ( n3933 & n7163 ) ;
  assign n10274 = n10273 ^ n9623 ^ 1'b0 ;
  assign n10275 = n4213 & ~n10274 ;
  assign n10276 = ~n1283 & n4308 ;
  assign n10277 = n6458 | n10276 ;
  assign n10278 = n8618 ^ n4425 ^ 1'b0 ;
  assign n10279 = n6364 & ~n10278 ;
  assign n10290 = n7243 ^ n6742 ^ n6059 ;
  assign n10287 = n1945 & n5302 ;
  assign n10288 = n1667 & ~n10287 ;
  assign n10289 = n10148 & ~n10288 ;
  assign n10280 = n1553 & n7908 ;
  assign n10283 = n1796 ^ n1620 ^ 1'b0 ;
  assign n10281 = n3822 ^ n2572 ^ n1385 ;
  assign n10282 = n10281 ^ x174 ^ 1'b0 ;
  assign n10284 = n10283 ^ n10282 ^ 1'b0 ;
  assign n10285 = ~n4663 & n10284 ;
  assign n10286 = n10280 | n10285 ;
  assign n10291 = n10290 ^ n10289 ^ n10286 ;
  assign n10292 = n10291 ^ n5420 ^ 1'b0 ;
  assign n10293 = ( ~n784 & n1374 ) | ( ~n784 & n2641 ) | ( n1374 & n2641 ) ;
  assign n10294 = x143 & ~n10293 ;
  assign n10295 = x31 & ~n5366 ;
  assign n10296 = n4845 ^ n3795 ^ 1'b0 ;
  assign n10297 = ( n640 & n3157 ) | ( n640 & ~n10189 ) | ( n3157 & ~n10189 ) ;
  assign n10298 = n657 & ~n4198 ;
  assign n10299 = ~n2677 & n9532 ;
  assign n10302 = n4225 ^ n4046 ^ 1'b0 ;
  assign n10303 = n613 & n10302 ;
  assign n10300 = n765 | n1928 ;
  assign n10301 = n9870 | n10300 ;
  assign n10304 = n10303 ^ n10301 ^ 1'b0 ;
  assign n10305 = ~n4909 & n10304 ;
  assign n10306 = ~n1193 & n7414 ;
  assign n10307 = n3815 & ~n10306 ;
  assign n10308 = n5811 | n8935 ;
  assign n10309 = n9543 ^ n2759 ^ 1'b0 ;
  assign n10310 = ( n724 & ~n2283 ) | ( n724 & n5745 ) | ( ~n2283 & n5745 ) ;
  assign n10311 = ( n1676 & ~n4399 ) | ( n1676 & n10310 ) | ( ~n4399 & n10310 ) ;
  assign n10312 = n6650 & ~n10311 ;
  assign n10313 = n7264 & ~n9053 ;
  assign n10314 = n8258 | n9273 ;
  assign n10315 = n3508 & ~n10314 ;
  assign n10316 = n3209 | n3684 ;
  assign n10317 = n9228 & n10316 ;
  assign n10318 = n2276 & ~n7015 ;
  assign n10319 = n6231 & ~n9957 ;
  assign n10320 = n6698 & n10319 ;
  assign n10321 = n4957 ^ n2688 ^ 1'b0 ;
  assign n10322 = n10321 ^ n8784 ^ 1'b0 ;
  assign n10323 = n4680 & n10322 ;
  assign n10324 = ~n3263 & n10323 ;
  assign n10326 = n2349 & ~n4122 ;
  assign n10327 = n4284 & n10326 ;
  assign n10325 = n5009 & n8673 ;
  assign n10328 = n10327 ^ n10325 ^ 1'b0 ;
  assign n10329 = n8998 & n10328 ;
  assign n10330 = n3190 & ~n3771 ;
  assign n10331 = ~n4995 & n10330 ;
  assign n10332 = ~n5627 & n7608 ;
  assign n10333 = n10332 ^ n2513 ^ 1'b0 ;
  assign n10334 = n4910 & n10333 ;
  assign n10335 = n2901 & n10334 ;
  assign n10336 = n3738 & ~n5835 ;
  assign n10337 = x217 & n759 ;
  assign n10338 = n5003 ^ n1626 ^ 1'b0 ;
  assign n10339 = ~n986 & n10338 ;
  assign n10340 = n10339 ^ n9931 ^ 1'b0 ;
  assign n10341 = n10211 ^ n5207 ^ x66 ;
  assign n10342 = n3211 | n10341 ;
  assign n10343 = n6846 ^ n5333 ^ 1'b0 ;
  assign n10344 = n5328 ^ n2622 ^ 1'b0 ;
  assign n10345 = n8851 & ~n10344 ;
  assign n10346 = ~n1772 & n2736 ;
  assign n10347 = n3357 & n10346 ;
  assign n10348 = n10347 ^ n1981 ^ 1'b0 ;
  assign n10349 = ~n1073 & n10348 ;
  assign n10350 = n6043 | n10349 ;
  assign n10351 = n475 | n10350 ;
  assign n10352 = n9284 ^ n8386 ^ n1295 ;
  assign n10353 = n937 & n9154 ;
  assign n10355 = n442 ^ x159 ^ 1'b0 ;
  assign n10356 = n957 | n10355 ;
  assign n10354 = n1490 & n1617 ;
  assign n10357 = n10356 ^ n10354 ^ n318 ;
  assign n10358 = n10339 ^ n1324 ^ 1'b0 ;
  assign n10359 = n448 & ~n10358 ;
  assign n10360 = n10357 & n10359 ;
  assign n10361 = n5087 ^ n1736 ^ 1'b0 ;
  assign n10362 = n9378 ^ n3525 ^ 1'b0 ;
  assign n10363 = n10361 & ~n10362 ;
  assign n10364 = ~n4502 & n7903 ;
  assign n10365 = n10364 ^ n8499 ^ 1'b0 ;
  assign n10366 = n4665 ^ n4061 ^ 1'b0 ;
  assign n10367 = n4610 & n10366 ;
  assign n10368 = n3468 & ~n7432 ;
  assign n10369 = n10368 ^ n10066 ^ n1210 ;
  assign n10370 = n8039 ^ n2948 ^ 1'b0 ;
  assign n10371 = n8138 | n10370 ;
  assign n10372 = x73 & n2788 ;
  assign n10373 = n10372 ^ n2216 ^ 1'b0 ;
  assign n10374 = n759 & ~n1523 ;
  assign n10375 = ~n8802 & n10374 ;
  assign n10376 = n10375 ^ x46 ^ 1'b0 ;
  assign n10377 = ~n2054 & n4099 ;
  assign n10378 = n2148 | n10377 ;
  assign n10379 = n9221 ^ n8326 ^ 1'b0 ;
  assign n10380 = ~n1680 & n10379 ;
  assign n10381 = n10380 ^ n3379 ^ 1'b0 ;
  assign n10382 = n4242 ^ n2487 ^ 1'b0 ;
  assign n10383 = ~n425 & n10382 ;
  assign n10384 = n3023 | n4515 ;
  assign n10385 = n10384 ^ n1032 ^ 1'b0 ;
  assign n10386 = ~n4767 & n10385 ;
  assign n10387 = n10386 ^ n9302 ^ 1'b0 ;
  assign n10388 = n3577 ^ x113 ^ 1'b0 ;
  assign n10389 = ~n697 & n10388 ;
  assign n10390 = ( ~n6424 & n9665 ) | ( ~n6424 & n10389 ) | ( n9665 & n10389 ) ;
  assign n10393 = n692 | n8746 ;
  assign n10394 = n10393 ^ x3 ^ 1'b0 ;
  assign n10395 = n10394 ^ n4082 ^ 1'b0 ;
  assign n10391 = n7251 ^ n2289 ^ 1'b0 ;
  assign n10392 = n1400 | n10391 ;
  assign n10396 = n10395 ^ n10392 ^ 1'b0 ;
  assign n10397 = ~n6833 & n10396 ;
  assign n10398 = ( x18 & n1796 ) | ( x18 & n4069 ) | ( n1796 & n4069 ) ;
  assign n10399 = n10398 ^ n8877 ^ n589 ;
  assign n10400 = n5029 & ~n10399 ;
  assign n10401 = n2464 & n10400 ;
  assign n10402 = ~n4959 & n5478 ;
  assign n10403 = n5001 & n10402 ;
  assign n10404 = ( n2904 & n2951 ) | ( n2904 & ~n3926 ) | ( n2951 & ~n3926 ) ;
  assign n10405 = n10403 & ~n10404 ;
  assign n10406 = ~n1261 & n10405 ;
  assign n10407 = n10406 ^ n1775 ^ 1'b0 ;
  assign n10408 = n1694 & n9536 ;
  assign n10409 = n10407 & ~n10408 ;
  assign n10410 = ~n9684 & n10409 ;
  assign n10411 = n4417 ^ n2404 ^ 1'b0 ;
  assign n10412 = n9709 & n10411 ;
  assign n10413 = n5123 & ~n7428 ;
  assign n10414 = ~n3362 & n10413 ;
  assign n10415 = n1577 | n5302 ;
  assign n10416 = n2719 & ~n10415 ;
  assign n10417 = x98 & ~n5132 ;
  assign n10418 = n10416 & n10417 ;
  assign n10419 = ~n828 & n8386 ;
  assign n10424 = ( n2701 & n7853 ) | ( n2701 & ~n8219 ) | ( n7853 & ~n8219 ) ;
  assign n10420 = x229 & ~n498 ;
  assign n10421 = n1393 & n1833 ;
  assign n10422 = n10421 ^ n10085 ^ 1'b0 ;
  assign n10423 = n10420 & ~n10422 ;
  assign n10425 = n10424 ^ n10423 ^ 1'b0 ;
  assign n10426 = n9617 ^ n3942 ^ n1579 ;
  assign n10427 = n2687 & ~n8870 ;
  assign n10428 = n1699 & n10427 ;
  assign n10429 = n10428 ^ n6959 ^ 1'b0 ;
  assign n10430 = ~n888 & n1936 ;
  assign n10431 = n814 & ~n10430 ;
  assign n10432 = n9739 ^ n628 ^ 1'b0 ;
  assign n10433 = ( ~n424 & n1242 ) | ( ~n424 & n10432 ) | ( n1242 & n10432 ) ;
  assign n10434 = ~n5705 & n7930 ;
  assign n10435 = n10434 ^ n4566 ^ 1'b0 ;
  assign n10436 = n10435 ^ n448 ^ 1'b0 ;
  assign n10437 = n10436 ^ n9714 ^ 1'b0 ;
  assign n10438 = n318 & ~n1049 ;
  assign n10439 = n10438 ^ n888 ^ 1'b0 ;
  assign n10440 = n1983 & n10439 ;
  assign n10441 = n10440 ^ n2502 ^ 1'b0 ;
  assign n10447 = n1943 ^ n1698 ^ 1'b0 ;
  assign n10448 = n9316 | n10447 ;
  assign n10442 = n1986 ^ x20 ^ 1'b0 ;
  assign n10443 = n1585 & n2489 ;
  assign n10444 = n6155 ^ n1437 ^ 1'b0 ;
  assign n10445 = n10443 & n10444 ;
  assign n10446 = n10442 & n10445 ;
  assign n10449 = n10448 ^ n10446 ^ 1'b0 ;
  assign n10450 = n2944 | n3057 ;
  assign n10451 = n10450 ^ n1140 ^ 1'b0 ;
  assign n10456 = n3855 & n7130 ;
  assign n10457 = ~n3855 & n10456 ;
  assign n10458 = n2609 & n6700 ;
  assign n10459 = n10457 & n10458 ;
  assign n10452 = n1413 ^ n503 ^ 1'b0 ;
  assign n10453 = n8688 ^ n6569 ^ 1'b0 ;
  assign n10454 = n10055 & ~n10453 ;
  assign n10455 = ~n10452 & n10454 ;
  assign n10460 = n10459 ^ n10455 ^ 1'b0 ;
  assign n10461 = n848 & n3275 ;
  assign n10462 = ~n3275 & n10461 ;
  assign n10463 = n1630 | n5392 ;
  assign n10464 = n5392 & ~n10463 ;
  assign n10465 = n10464 ^ n2697 ^ 1'b0 ;
  assign n10466 = n10462 | n10465 ;
  assign n10467 = n4554 & n4951 ;
  assign n10468 = n10466 | n10467 ;
  assign n10469 = n10460 | n10468 ;
  assign n10470 = n5203 ^ n4740 ^ 1'b0 ;
  assign n10471 = ~n5559 & n10470 ;
  assign n10472 = n9302 ^ n7473 ^ 1'b0 ;
  assign n10473 = n4480 ^ n1440 ^ 1'b0 ;
  assign n10474 = n1570 | n10473 ;
  assign n10475 = n3542 & n10474 ;
  assign n10476 = n10475 ^ n4337 ^ 1'b0 ;
  assign n10477 = n3499 ^ n1874 ^ 1'b0 ;
  assign n10478 = n3115 & ~n5608 ;
  assign n10479 = ~n5928 & n10478 ;
  assign n10480 = n10479 ^ n10225 ^ 1'b0 ;
  assign n10481 = x119 & ~n10480 ;
  assign n10482 = n10477 & ~n10481 ;
  assign n10483 = ~n2797 & n10482 ;
  assign n10484 = ~n3964 & n7168 ;
  assign n10485 = n5537 ^ n2069 ^ 1'b0 ;
  assign n10486 = n5421 ^ x36 ^ 1'b0 ;
  assign n10487 = n4025 & n10486 ;
  assign n10488 = n4839 & n10487 ;
  assign n10489 = n10488 ^ n692 ^ 1'b0 ;
  assign n10490 = ( n3887 & n8485 ) | ( n3887 & ~n9336 ) | ( n8485 & ~n9336 ) ;
  assign n10491 = n8867 ^ n4505 ^ 1'b0 ;
  assign n10492 = n2370 & ~n4522 ;
  assign n10493 = ( n964 & n3370 ) | ( n964 & n9592 ) | ( n3370 & n9592 ) ;
  assign n10494 = ~n2958 & n7630 ;
  assign n10495 = ~n5382 & n10494 ;
  assign n10496 = n1371 & ~n10495 ;
  assign n10497 = n10496 ^ n3400 ^ 1'b0 ;
  assign n10498 = ~n5726 & n7282 ;
  assign n10499 = ~n6551 & n9078 ;
  assign n10500 = n10499 ^ n6780 ^ 1'b0 ;
  assign n10501 = ~n799 & n10500 ;
  assign n10502 = n4309 & ~n4449 ;
  assign n10503 = n7545 ^ n1645 ^ 1'b0 ;
  assign n10504 = ~n10502 & n10503 ;
  assign n10505 = ~n8052 & n10504 ;
  assign n10506 = n2481 & ~n10505 ;
  assign n10507 = n7373 & ~n10506 ;
  assign n10508 = n5420 & ~n6307 ;
  assign n10509 = n4327 & n5645 ;
  assign n10510 = ( n845 & ~n5962 ) | ( n845 & n9860 ) | ( ~n5962 & n9860 ) ;
  assign n10511 = n3639 | n4094 ;
  assign n10512 = n10511 ^ n10369 ^ 1'b0 ;
  assign n10513 = n10356 ^ n4226 ^ 1'b0 ;
  assign n10514 = n1552 & n10513 ;
  assign n10515 = n10514 ^ n6533 ^ 1'b0 ;
  assign n10516 = n10515 ^ n8614 ^ n4061 ;
  assign n10517 = ~n2785 & n8192 ;
  assign n10518 = n9501 ^ n4360 ^ 1'b0 ;
  assign n10521 = n5307 ^ n4295 ^ 1'b0 ;
  assign n10522 = n3461 | n10521 ;
  assign n10523 = n2047 & ~n10522 ;
  assign n10524 = ( ~n4104 & n5865 ) | ( ~n4104 & n10523 ) | ( n5865 & n10523 ) ;
  assign n10519 = n5831 ^ n3342 ^ 1'b0 ;
  assign n10520 = ~n4094 & n10519 ;
  assign n10525 = n10524 ^ n10520 ^ 1'b0 ;
  assign n10526 = n1018 & ~n10525 ;
  assign n10531 = n3225 ^ n2073 ^ 1'b0 ;
  assign n10532 = n7310 | n10531 ;
  assign n10527 = n4950 ^ n1956 ^ 1'b0 ;
  assign n10528 = ~n2098 & n10527 ;
  assign n10529 = n10528 ^ n7672 ^ 1'b0 ;
  assign n10530 = n7627 & n10529 ;
  assign n10533 = n10532 ^ n10530 ^ 1'b0 ;
  assign n10534 = ~n1147 & n10533 ;
  assign n10535 = n6241 | n10534 ;
  assign n10536 = x42 & ~n9211 ;
  assign n10537 = n10522 ^ n6425 ^ 1'b0 ;
  assign n10538 = n713 & ~n10418 ;
  assign n10540 = ( n375 & n6057 ) | ( n375 & ~n6470 ) | ( n6057 & ~n6470 ) ;
  assign n10541 = ~n2724 & n10540 ;
  assign n10539 = n2730 | n4871 ;
  assign n10542 = n10541 ^ n10539 ^ 1'b0 ;
  assign n10545 = n3539 & ~n4222 ;
  assign n10543 = n2654 ^ n395 ^ 1'b0 ;
  assign n10544 = n3994 & n10543 ;
  assign n10546 = n10545 ^ n10544 ^ 1'b0 ;
  assign n10547 = n4426 | n10402 ;
  assign n10548 = n6533 | n10547 ;
  assign n10549 = n10548 ^ n331 ^ 1'b0 ;
  assign n10550 = n749 & ~n2078 ;
  assign n10551 = n10550 ^ n6681 ^ 1'b0 ;
  assign n10552 = ( n547 & n7838 ) | ( n547 & n10551 ) | ( n7838 & n10551 ) ;
  assign n10553 = n645 | n1775 ;
  assign n10554 = n9543 & ~n10553 ;
  assign n10555 = n6632 ^ n5613 ^ 1'b0 ;
  assign n10556 = n2649 & n10555 ;
  assign n10557 = n1138 ^ n1112 ^ n867 ;
  assign n10558 = ~n1405 & n10557 ;
  assign n10559 = n10558 ^ n8252 ^ 1'b0 ;
  assign n10560 = ~n274 & n4696 ;
  assign n10561 = n2471 | n10560 ;
  assign n10562 = ( ~n1338 & n2482 ) | ( ~n1338 & n3882 ) | ( n2482 & n3882 ) ;
  assign n10563 = n1083 & n9538 ;
  assign n10564 = n10562 & n10563 ;
  assign n10565 = n1796 & ~n4150 ;
  assign n10566 = n10565 ^ n4202 ^ 1'b0 ;
  assign n10567 = n10566 ^ n5821 ^ 1'b0 ;
  assign n10568 = n7430 | n9383 ;
  assign n10569 = n10568 ^ n5722 ^ 1'b0 ;
  assign n10570 = ~n6731 & n6920 ;
  assign n10571 = ~n9873 & n10570 ;
  assign n10572 = n3047 ^ n2668 ^ 1'b0 ;
  assign n10573 = n6140 ^ n4522 ^ 1'b0 ;
  assign n10574 = n1610 & n10573 ;
  assign n10575 = n5116 | n10001 ;
  assign n10576 = n3903 ^ n689 ^ 1'b0 ;
  assign n10577 = ~n3027 & n10576 ;
  assign n10578 = n7755 ^ n2204 ^ 1'b0 ;
  assign n10579 = ~n1948 & n6293 ;
  assign n10580 = ~n10578 & n10579 ;
  assign n10581 = x180 & ~n1432 ;
  assign n10582 = n10580 & n10581 ;
  assign n10583 = n10577 & ~n10582 ;
  assign n10584 = n6974 & n10583 ;
  assign n10585 = n6187 ^ n4311 ^ 1'b0 ;
  assign n10586 = n10584 | n10585 ;
  assign n10587 = ~n2165 & n3723 ;
  assign n10588 = n10587 ^ n1002 ^ 1'b0 ;
  assign n10589 = n8880 ^ n359 ^ 1'b0 ;
  assign n10590 = n10589 ^ n8011 ^ 1'b0 ;
  assign n10591 = n10588 & ~n10590 ;
  assign n10594 = n794 & ~n8331 ;
  assign n10595 = n1960 | n4485 ;
  assign n10596 = n10594 | n10595 ;
  assign n10592 = n361 | n1505 ;
  assign n10593 = n10592 ^ n9727 ^ 1'b0 ;
  assign n10597 = n10596 ^ n10593 ^ 1'b0 ;
  assign n10598 = n2348 | n10597 ;
  assign n10599 = n7013 ^ n6243 ^ n3151 ;
  assign n10600 = ~n2618 & n3257 ;
  assign n10601 = n3258 & n10600 ;
  assign n10602 = ~n333 & n5049 ;
  assign n10603 = ~n3974 & n10602 ;
  assign n10604 = n3271 ^ x247 ^ 1'b0 ;
  assign n10605 = n5134 & n10604 ;
  assign n10606 = n10605 ^ n1255 ^ 1'b0 ;
  assign n10609 = ~n2047 & n4920 ;
  assign n10607 = n3844 ^ n2665 ^ 1'b0 ;
  assign n10608 = n4354 & ~n10607 ;
  assign n10610 = n10609 ^ n10608 ^ n4602 ;
  assign n10611 = n8747 & n10610 ;
  assign n10612 = n9494 | n10611 ;
  assign n10613 = n10612 ^ n3693 ^ 1'b0 ;
  assign n10614 = n10606 & n10613 ;
  assign n10615 = n6627 ^ n3975 ^ 1'b0 ;
  assign n10616 = n10615 ^ n1114 ^ 1'b0 ;
  assign n10617 = n10313 & n10616 ;
  assign n10618 = n10617 ^ n5919 ^ 1'b0 ;
  assign n10621 = x6 & n9974 ;
  assign n10622 = n1664 & n10621 ;
  assign n10623 = ( ~n2562 & n7323 ) | ( ~n2562 & n10622 ) | ( n7323 & n10622 ) ;
  assign n10624 = n5069 ^ n682 ^ 1'b0 ;
  assign n10625 = n10623 & n10624 ;
  assign n10619 = n9080 ^ n7846 ^ 1'b0 ;
  assign n10620 = n8000 & n10619 ;
  assign n10626 = n10625 ^ n10620 ^ 1'b0 ;
  assign n10627 = n5325 & ~n7301 ;
  assign n10628 = n10627 ^ n296 ^ 1'b0 ;
  assign n10629 = n6425 ^ n5216 ^ 1'b0 ;
  assign n10630 = n10629 ^ n1250 ^ 1'b0 ;
  assign n10631 = n5528 & n9886 ;
  assign n10632 = ~n10630 & n10631 ;
  assign n10633 = n2276 & ~n10632 ;
  assign n10634 = n1630 & n10633 ;
  assign n10635 = n10634 ^ n8823 ^ 1'b0 ;
  assign n10636 = n10628 & n10635 ;
  assign n10637 = ~n1078 & n4694 ;
  assign n10638 = n973 | n9674 ;
  assign n10639 = n2937 & ~n10638 ;
  assign n10640 = n2378 | n5454 ;
  assign n10641 = n10640 ^ n8030 ^ 1'b0 ;
  assign n10642 = ~n10639 & n10641 ;
  assign n10643 = n10642 ^ n1558 ^ 1'b0 ;
  assign n10644 = n3791 | n8056 ;
  assign n10645 = n5750 ^ n1688 ^ 1'b0 ;
  assign n10646 = n353 & n10645 ;
  assign n10650 = n4567 ^ n1244 ^ 1'b0 ;
  assign n10647 = x3 & n2868 ;
  assign n10648 = n10647 ^ n4232 ^ 1'b0 ;
  assign n10649 = ~n4503 & n10648 ;
  assign n10651 = n10650 ^ n10649 ^ 1'b0 ;
  assign n10652 = n2653 & n9350 ;
  assign n10653 = ( n500 & n2953 ) | ( n500 & ~n5373 ) | ( n2953 & ~n5373 ) ;
  assign n10654 = n10652 & ~n10653 ;
  assign n10655 = n7301 ^ n374 ^ 1'b0 ;
  assign n10656 = n6424 | n7199 ;
  assign n10657 = n9294 | n10656 ;
  assign n10658 = ~n1901 & n8524 ;
  assign n10659 = n10658 ^ x146 ^ 1'b0 ;
  assign n10660 = n4325 & ~n9973 ;
  assign n10661 = n10660 ^ n5396 ^ 1'b0 ;
  assign n10662 = n5183 & n10661 ;
  assign n10663 = n4747 & ~n7959 ;
  assign n10664 = n1802 & ~n6235 ;
  assign n10665 = x180 & n10664 ;
  assign n10666 = n9829 & n10665 ;
  assign n10667 = n4494 & ~n6873 ;
  assign n10668 = n10667 ^ n3757 ^ 1'b0 ;
  assign n10669 = n7874 ^ n2116 ^ 1'b0 ;
  assign n10670 = n4090 & ~n10669 ;
  assign n10671 = n5870 & ~n9586 ;
  assign n10672 = ~n2959 & n10671 ;
  assign n10673 = ( n2192 & n5775 ) | ( n2192 & ~n9212 ) | ( n5775 & ~n9212 ) ;
  assign n10674 = n10673 ^ n2291 ^ n580 ;
  assign n10675 = n2472 | n3331 ;
  assign n10676 = n8759 & ~n10675 ;
  assign n10677 = n6506 & ~n7963 ;
  assign n10678 = n1948 & n10677 ;
  assign n10679 = n5523 ^ n709 ^ 1'b0 ;
  assign n10680 = n1528 ^ n724 ^ 1'b0 ;
  assign n10681 = x128 & x236 ;
  assign n10682 = ~n8471 & n10681 ;
  assign n10683 = x13 | n2870 ;
  assign n10684 = n5046 | n10683 ;
  assign n10685 = n619 | n3331 ;
  assign n10686 = n7318 ^ n1456 ^ 1'b0 ;
  assign n10687 = ~n10685 & n10686 ;
  assign n10688 = n3542 & ~n7522 ;
  assign n10689 = n10688 ^ n4402 ^ 1'b0 ;
  assign n10690 = n10689 ^ n9648 ^ n3080 ;
  assign n10691 = n10051 & ~n10690 ;
  assign n10692 = n9739 ^ n5515 ^ n2054 ;
  assign n10693 = n1575 | n1725 ;
  assign n10694 = n1636 & ~n10693 ;
  assign n10695 = n10694 ^ n4797 ^ 1'b0 ;
  assign n10698 = n1632 & ~n7203 ;
  assign n10696 = n520 & n2286 ;
  assign n10697 = n539 | n10696 ;
  assign n10699 = n10698 ^ n10697 ^ 1'b0 ;
  assign n10700 = ~n2078 & n3830 ;
  assign n10701 = n3183 & n10700 ;
  assign n10702 = n10701 ^ n7813 ^ 1'b0 ;
  assign n10703 = n3653 ^ n3453 ^ 1'b0 ;
  assign n10704 = n5519 | n10703 ;
  assign n10705 = n10704 ^ n3494 ^ 1'b0 ;
  assign n10706 = ~n666 & n6819 ;
  assign n10707 = n2964 & ~n3935 ;
  assign n10708 = n10707 ^ n3686 ^ 1'b0 ;
  assign n10709 = n6022 & n10708 ;
  assign n10710 = ( ~n2008 & n10242 ) | ( ~n2008 & n10709 ) | ( n10242 & n10709 ) ;
  assign n10711 = n8276 ^ n7930 ^ 1'b0 ;
  assign n10712 = n10711 ^ n4313 ^ 1'b0 ;
  assign n10713 = n7650 | n10712 ;
  assign n10714 = n8829 ^ n7270 ^ 1'b0 ;
  assign n10715 = n993 | n10074 ;
  assign n10716 = ~n8189 & n8351 ;
  assign n10717 = n10716 ^ n4732 ^ 1'b0 ;
  assign n10718 = n9806 & n10717 ;
  assign n10719 = n8881 & n10718 ;
  assign n10720 = n8309 ^ n4509 ^ 1'b0 ;
  assign n10721 = ~n993 & n10720 ;
  assign n10722 = n7515 & ~n10721 ;
  assign n10723 = n9990 ^ n6077 ^ 1'b0 ;
  assign n10724 = n1657 | n10723 ;
  assign n10725 = n6112 & ~n6805 ;
  assign n10726 = ~n1624 & n10725 ;
  assign n10727 = n7183 ^ n3589 ^ 1'b0 ;
  assign n10728 = ~n10726 & n10727 ;
  assign n10729 = ~n530 & n4752 ;
  assign n10730 = n1165 & n4335 ;
  assign n10731 = ~n10729 & n10730 ;
  assign n10732 = n10731 ^ n9412 ^ 1'b0 ;
  assign n10733 = n8853 ^ n835 ^ 1'b0 ;
  assign n10734 = x139 & n1124 ;
  assign n10735 = n10734 ^ n4851 ^ 1'b0 ;
  assign n10736 = n6688 | n10735 ;
  assign n10737 = n8607 & ~n10736 ;
  assign n10738 = n3684 & ~n3931 ;
  assign n10739 = x113 & ~n10738 ;
  assign n10740 = ~x113 & n10739 ;
  assign n10741 = n7350 ^ n6359 ^ 1'b0 ;
  assign n10743 = ~n1023 & n3499 ;
  assign n10742 = n3413 | n5333 ;
  assign n10744 = n10743 ^ n10742 ^ n4563 ;
  assign n10745 = n5243 & ~n9393 ;
  assign n10746 = n10745 ^ n5231 ^ 1'b0 ;
  assign n10747 = n2091 & n8861 ;
  assign n10748 = n10747 ^ n1178 ^ 1'b0 ;
  assign n10749 = n7513 & ~n10748 ;
  assign n10750 = n3904 & n10749 ;
  assign n10751 = n4434 | n9334 ;
  assign n10752 = n4754 | n10751 ;
  assign n10753 = n2340 & n10752 ;
  assign n10754 = n10753 ^ n6490 ^ 1'b0 ;
  assign n10755 = ~n2433 & n9872 ;
  assign n10756 = x136 & n7801 ;
  assign n10757 = ~n270 & n9209 ;
  assign n10758 = ~n5782 & n10757 ;
  assign n10759 = n2338 ^ n1319 ^ 1'b0 ;
  assign n10760 = n2950 & ~n3628 ;
  assign n10761 = n10760 ^ n2868 ^ 1'b0 ;
  assign n10762 = n10761 ^ n10345 ^ 1'b0 ;
  assign n10763 = n3848 ^ n3604 ^ 1'b0 ;
  assign n10764 = n2141 & ~n2770 ;
  assign n10765 = n10764 ^ n10448 ^ 1'b0 ;
  assign n10766 = ~n6682 & n10765 ;
  assign n10767 = n1137 & n4280 ;
  assign n10768 = ~n3988 & n10767 ;
  assign n10769 = n7627 ^ n3328 ^ 1'b0 ;
  assign n10770 = n7914 & n10769 ;
  assign n10771 = ~n10768 & n10770 ;
  assign n10775 = ~n1406 & n3886 ;
  assign n10772 = n1653 ^ n708 ^ 1'b0 ;
  assign n10773 = n4258 & n10772 ;
  assign n10774 = ~n2387 & n10773 ;
  assign n10776 = n10775 ^ n10774 ^ 1'b0 ;
  assign n10777 = ~n4970 & n10776 ;
  assign n10778 = n3810 & ~n10010 ;
  assign n10779 = n391 & ~n3290 ;
  assign n10780 = n10779 ^ n10619 ^ 1'b0 ;
  assign n10781 = n5034 & ~n8616 ;
  assign n10782 = n10780 | n10781 ;
  assign n10783 = n8033 & ~n10782 ;
  assign n10784 = n10778 & ~n10783 ;
  assign n10785 = n2117 & ~n8216 ;
  assign n10786 = ~n4404 & n4919 ;
  assign n10787 = ~n7791 & n10786 ;
  assign n10788 = n4739 | n10787 ;
  assign n10789 = n10788 ^ n4099 ^ 1'b0 ;
  assign n10790 = n5278 ^ n3238 ^ 1'b0 ;
  assign n10791 = ~n2203 & n8755 ;
  assign n10792 = n5422 & n10791 ;
  assign n10793 = n4876 ^ n2322 ^ 1'b0 ;
  assign n10794 = ~n5756 & n10793 ;
  assign n10795 = n10391 & n10794 ;
  assign n10796 = n421 & n2443 ;
  assign n10797 = n10796 ^ n4115 ^ 1'b0 ;
  assign n10798 = n7473 ^ n2693 ^ 1'b0 ;
  assign n10799 = n2165 & n8525 ;
  assign n10800 = ~n7839 & n10799 ;
  assign n10801 = n10800 ^ n4754 ^ 1'b0 ;
  assign n10802 = ~n7606 & n10801 ;
  assign n10803 = n8248 & n10802 ;
  assign n10804 = n5649 ^ n2982 ^ n1648 ;
  assign n10805 = ~n1851 & n8088 ;
  assign n10806 = n348 | n10805 ;
  assign n10807 = n10806 ^ n6785 ^ 1'b0 ;
  assign n10808 = n10807 ^ n1328 ^ 1'b0 ;
  assign n10809 = ~n3719 & n4855 ;
  assign n10810 = ~n10164 & n10809 ;
  assign n10811 = n10055 ^ n7330 ^ 1'b0 ;
  assign n10812 = n4511 | n10811 ;
  assign n10813 = n10812 ^ n7197 ^ 1'b0 ;
  assign n10814 = n3549 | n8742 ;
  assign n10815 = n366 & n1947 ;
  assign n10816 = n10815 ^ n4003 ^ 1'b0 ;
  assign n10817 = n10816 ^ n2993 ^ 1'b0 ;
  assign n10818 = n6624 ^ n1696 ^ 1'b0 ;
  assign n10819 = n5318 | n10818 ;
  assign n10820 = n10817 | n10819 ;
  assign n10821 = n6551 | n8041 ;
  assign n10822 = x73 & n5136 ;
  assign n10823 = n7401 ^ n2397 ^ 1'b0 ;
  assign n10824 = n4659 | n5851 ;
  assign n10825 = n10824 ^ n5954 ^ 1'b0 ;
  assign n10826 = n10825 ^ n1605 ^ 1'b0 ;
  assign n10827 = n5046 ^ n3564 ^ 1'b0 ;
  assign n10828 = n747 & n10827 ;
  assign n10829 = ~n3576 & n10828 ;
  assign n10830 = n5705 ^ n4222 ^ 1'b0 ;
  assign n10831 = n5310 & n10830 ;
  assign n10832 = n10831 ^ n7678 ^ n3098 ;
  assign n10833 = n1788 ^ n1306 ^ 1'b0 ;
  assign n10834 = n5602 | n10833 ;
  assign n10835 = x81 & n1826 ;
  assign n10836 = n3814 | n10835 ;
  assign n10837 = n6548 & ~n10836 ;
  assign n10838 = ~n4226 & n10403 ;
  assign n10839 = n8022 & n10838 ;
  assign n10840 = n10837 & ~n10839 ;
  assign n10841 = n8651 ^ n6327 ^ 1'b0 ;
  assign n10842 = n5556 & ~n7896 ;
  assign n10843 = n10842 ^ n8088 ^ 1'b0 ;
  assign n10844 = n10721 ^ n3352 ^ 1'b0 ;
  assign n10845 = n10843 & n10844 ;
  assign n10846 = n4209 ^ n3150 ^ 1'b0 ;
  assign n10847 = n4044 & ~n10846 ;
  assign n10848 = n7705 ^ n2322 ^ 1'b0 ;
  assign n10849 = n10848 ^ n10675 ^ n3091 ;
  assign n10850 = n4175 | n10849 ;
  assign n10851 = n10850 ^ n9667 ^ 1'b0 ;
  assign n10852 = n3209 ^ n2302 ^ n325 ;
  assign n10853 = n7753 ^ n496 ^ 1'b0 ;
  assign n10854 = n9708 & n10853 ;
  assign n10855 = ~n3724 & n10089 ;
  assign n10861 = n7356 ^ n7276 ^ 1'b0 ;
  assign n10856 = n2112 ^ n1757 ^ 1'b0 ;
  assign n10857 = n7393 & ~n10856 ;
  assign n10858 = ~n2692 & n3834 ;
  assign n10859 = n10857 & ~n10858 ;
  assign n10860 = ~n3951 & n10859 ;
  assign n10862 = n10861 ^ n10860 ^ 1'b0 ;
  assign n10863 = n749 & ~n3137 ;
  assign n10864 = ~n3021 & n10863 ;
  assign n10865 = n10864 ^ n10042 ^ n5954 ;
  assign n10866 = n466 | n2085 ;
  assign n10867 = n10866 ^ n703 ^ 1'b0 ;
  assign n10868 = n10867 ^ n7709 ^ 1'b0 ;
  assign n10869 = n4168 | n10868 ;
  assign n10870 = n10865 & ~n10869 ;
  assign n10871 = n8243 & n10870 ;
  assign n10872 = n1379 & ~n3057 ;
  assign n10873 = n3417 ^ n409 ^ 1'b0 ;
  assign n10874 = ~n9720 & n10873 ;
  assign n10875 = ~n1797 & n2691 ;
  assign n10876 = n10875 ^ n1585 ^ 1'b0 ;
  assign n10877 = ( ~n10872 & n10874 ) | ( ~n10872 & n10876 ) | ( n10874 & n10876 ) ;
  assign n10878 = n8994 & n9958 ;
  assign n10880 = n4121 ^ n1947 ^ n970 ;
  assign n10881 = n6923 ^ n4659 ^ 1'b0 ;
  assign n10882 = n10880 & ~n10881 ;
  assign n10883 = n3802 | n9365 ;
  assign n10884 = n9128 | n10883 ;
  assign n10885 = n10882 & ~n10884 ;
  assign n10879 = n991 & ~n5618 ;
  assign n10886 = n10885 ^ n10879 ^ 1'b0 ;
  assign n10887 = n1094 | n5165 ;
  assign n10888 = n1032 | n10887 ;
  assign n10889 = n5004 & n6453 ;
  assign n10890 = n10888 & ~n10889 ;
  assign n10891 = n10890 ^ n2915 ^ 1'b0 ;
  assign n10892 = n10891 ^ n1627 ^ 1'b0 ;
  assign n10893 = n5511 | n10892 ;
  assign n10894 = n5067 ^ n3751 ^ 1'b0 ;
  assign n10895 = n6437 ^ n1080 ^ 1'b0 ;
  assign n10896 = n8424 | n10895 ;
  assign n10897 = n7355 & ~n10896 ;
  assign n10898 = n3903 & ~n6695 ;
  assign n10899 = n10898 ^ n1932 ^ 1'b0 ;
  assign n10900 = ~x216 & n10899 ;
  assign n10901 = n9186 & ~n9914 ;
  assign n10902 = ~n994 & n10901 ;
  assign n10903 = n10902 ^ n6633 ^ 1'b0 ;
  assign n10904 = n4608 ^ n3771 ^ 1'b0 ;
  assign n10905 = n2102 & ~n10904 ;
  assign n10906 = ~n5227 & n10905 ;
  assign n10907 = n347 & n10906 ;
  assign n10908 = n7271 ^ n7179 ^ n5206 ;
  assign n10909 = n5909 & ~n10648 ;
  assign n10910 = n10909 ^ n7038 ^ 1'b0 ;
  assign n10911 = n3648 & ~n10910 ;
  assign n10912 = ~n277 & n10911 ;
  assign n10913 = ~n4035 & n10912 ;
  assign n10914 = n4044 ^ n937 ^ 1'b0 ;
  assign n10915 = n10914 ^ n8286 ^ 1'b0 ;
  assign n10916 = n6471 | n10915 ;
  assign n10917 = n10916 ^ n7427 ^ 1'b0 ;
  assign n10918 = n9271 & n10917 ;
  assign n10919 = ~n1871 & n6485 ;
  assign n10920 = ~x111 & n10919 ;
  assign n10921 = n4791 | n10920 ;
  assign n10922 = n8999 | n10921 ;
  assign n10923 = n1966 | n8844 ;
  assign n10924 = n4584 ^ n858 ^ 1'b0 ;
  assign n10925 = ~n3653 & n10924 ;
  assign n10926 = n5504 & ~n10925 ;
  assign n10927 = n8092 ^ n6842 ^ 1'b0 ;
  assign n10928 = n537 & n10927 ;
  assign n10929 = ~n6340 & n8988 ;
  assign n10930 = n10928 & n10929 ;
  assign n10931 = n6655 ^ n5404 ^ 1'b0 ;
  assign n10932 = n4634 & ~n10931 ;
  assign n10933 = n7569 & n10932 ;
  assign n10934 = n10933 ^ n10653 ^ 1'b0 ;
  assign n10935 = n6781 & n7439 ;
  assign n10936 = n5944 ^ n5771 ^ 1'b0 ;
  assign n10937 = n7977 & ~n10936 ;
  assign n10938 = n3603 ^ n2967 ^ 1'b0 ;
  assign n10939 = ~n7231 & n10938 ;
  assign n10940 = ~n10937 & n10939 ;
  assign n10946 = n4368 ^ n2281 ^ 1'b0 ;
  assign n10941 = n3703 | n5626 ;
  assign n10942 = n6813 & ~n10941 ;
  assign n10943 = ( n256 & n4849 ) | ( n256 & ~n6045 ) | ( n4849 & ~n6045 ) ;
  assign n10944 = ~n2242 & n10943 ;
  assign n10945 = n10942 | n10944 ;
  assign n10947 = n10946 ^ n10945 ^ 1'b0 ;
  assign n10948 = n988 | n1036 ;
  assign n10949 = n10948 ^ x66 ^ 1'b0 ;
  assign n10950 = n3568 & ~n10949 ;
  assign n10951 = n1478 ^ x213 ^ 1'b0 ;
  assign n10952 = ~n1516 & n10951 ;
  assign n10953 = n10952 ^ n897 ^ 1'b0 ;
  assign n10954 = n3970 | n10953 ;
  assign n10955 = n10196 & ~n10954 ;
  assign n10956 = n2148 & ~n4383 ;
  assign n10957 = n10956 ^ n4059 ^ 1'b0 ;
  assign n10958 = n10957 ^ n2178 ^ 1'b0 ;
  assign n10959 = n9473 & n10958 ;
  assign n10960 = n9911 ^ n4111 ^ 1'b0 ;
  assign n10961 = n4099 ^ n1388 ^ 1'b0 ;
  assign n10962 = n677 & ~n10961 ;
  assign n10963 = n8574 & n10962 ;
  assign n10964 = n3483 | n4086 ;
  assign n10965 = n4423 | n10964 ;
  assign n10966 = ( n3251 & ~n5948 ) | ( n3251 & n10965 ) | ( ~n5948 & n10965 ) ;
  assign n10967 = n2932 ^ n2034 ^ 1'b0 ;
  assign n10968 = n2741 | n10967 ;
  assign n10969 = n2528 & ~n10968 ;
  assign n10970 = n6778 ^ n458 ^ 1'b0 ;
  assign n10971 = n4394 & ~n10970 ;
  assign n10981 = ~n3801 & n5840 ;
  assign n10972 = n938 | n5274 ;
  assign n10973 = n10972 ^ n2655 ^ 1'b0 ;
  assign n10974 = n10973 ^ n2953 ^ n2310 ;
  assign n10975 = n3518 & n3895 ;
  assign n10976 = n10975 ^ n3529 ^ 1'b0 ;
  assign n10977 = n5488 & n10976 ;
  assign n10978 = n270 & n10977 ;
  assign n10979 = n10974 | n10978 ;
  assign n10980 = n891 & ~n10979 ;
  assign n10982 = n10981 ^ n10980 ^ 1'b0 ;
  assign n10983 = n8919 ^ n6272 ^ 1'b0 ;
  assign n10984 = n4400 | n10983 ;
  assign n10985 = n9526 ^ n5476 ^ 1'b0 ;
  assign n10986 = n10985 ^ n10756 ^ 1'b0 ;
  assign n10987 = n1481 & ~n5450 ;
  assign n10988 = n4391 & n10987 ;
  assign n10989 = n10062 ^ n1333 ^ 1'b0 ;
  assign n10990 = ~n10988 & n10989 ;
  assign n10992 = n1725 | n8704 ;
  assign n10991 = n5087 | n6338 ;
  assign n10993 = n10992 ^ n10991 ^ 1'b0 ;
  assign n10994 = n2724 & n10993 ;
  assign n10995 = n5261 ^ n5097 ^ n2213 ;
  assign n10996 = n10995 ^ n876 ^ 1'b0 ;
  assign n10997 = x1 & n2184 ;
  assign n10998 = n10997 ^ x113 ^ 1'b0 ;
  assign n10999 = n6080 & n10998 ;
  assign n11005 = n2170 | n6346 ;
  assign n11006 = n2441 & ~n11005 ;
  assign n11007 = n732 & n11006 ;
  assign n11000 = n5322 ^ n4852 ^ n4070 ;
  assign n11001 = n3300 ^ n1931 ^ x168 ;
  assign n11002 = n11001 ^ n3768 ^ 1'b0 ;
  assign n11003 = n11000 | n11002 ;
  assign n11004 = n11003 ^ n4726 ^ 1'b0 ;
  assign n11008 = n11007 ^ n11004 ^ 1'b0 ;
  assign n11009 = n4146 ^ n2615 ^ 1'b0 ;
  assign n11010 = ~n4649 & n11009 ;
  assign n11014 = n1376 | n7307 ;
  assign n11013 = n6753 ^ n5561 ^ n1324 ;
  assign n11015 = n11014 ^ n11013 ^ 1'b0 ;
  assign n11011 = ~n3386 & n6387 ;
  assign n11012 = n6343 & n11011 ;
  assign n11016 = n11015 ^ n11012 ^ n9911 ;
  assign n11017 = n9350 & n11016 ;
  assign n11018 = n11017 ^ n1352 ^ 1'b0 ;
  assign n11019 = n9737 & ~n11018 ;
  assign n11020 = n3994 ^ n2120 ^ 1'b0 ;
  assign n11021 = ~n3765 & n9199 ;
  assign n11022 = n11021 ^ n2286 ^ 1'b0 ;
  assign n11026 = n498 & ~n511 ;
  assign n11023 = n1911 | n2390 ;
  assign n11024 = n6090 & ~n11023 ;
  assign n11025 = n11024 ^ n1534 ^ 1'b0 ;
  assign n11027 = n11026 ^ n11025 ^ 1'b0 ;
  assign n11028 = n11022 & n11027 ;
  assign n11029 = n2529 & ~n10471 ;
  assign n11030 = x88 & ~x97 ;
  assign n11031 = ~n2110 & n8557 ;
  assign n11032 = n11031 ^ n8700 ^ 1'b0 ;
  assign n11033 = ~n3327 & n11032 ;
  assign n11034 = n11033 ^ n5221 ^ 1'b0 ;
  assign n11035 = n2844 & ~n8712 ;
  assign n11036 = n4752 ^ n2192 ^ 1'b0 ;
  assign n11037 = n1807 & ~n11036 ;
  assign n11038 = n998 ^ x163 ^ 1'b0 ;
  assign n11039 = n1389 ^ n850 ^ 1'b0 ;
  assign n11040 = n3867 & n11039 ;
  assign n11041 = n11040 ^ x46 ^ 1'b0 ;
  assign n11042 = n11041 ^ n10046 ^ n6387 ;
  assign n11043 = ( ~n11037 & n11038 ) | ( ~n11037 & n11042 ) | ( n11038 & n11042 ) ;
  assign n11044 = ~n4639 & n11043 ;
  assign n11045 = n3393 ^ n3326 ^ 1'b0 ;
  assign n11046 = x245 & n11045 ;
  assign n11047 = n6802 & ~n8642 ;
  assign n11048 = ~n860 & n7972 ;
  assign n11049 = n11048 ^ n4905 ^ 1'b0 ;
  assign n11050 = n10880 ^ n6282 ^ 1'b0 ;
  assign n11051 = n11049 & n11050 ;
  assign n11052 = n11051 ^ n2018 ^ 1'b0 ;
  assign n11053 = n2193 ^ n548 ^ 1'b0 ;
  assign n11054 = x100 | n6001 ;
  assign n11055 = n11054 ^ x41 ^ 1'b0 ;
  assign n11056 = n10593 | n11055 ;
  assign n11057 = n4330 | n11056 ;
  assign n11058 = n4676 & n10690 ;
  assign n11059 = ~n11057 & n11058 ;
  assign n11060 = n1328 & n2334 ;
  assign n11061 = n11060 ^ n668 ^ 1'b0 ;
  assign n11062 = n2858 & n11061 ;
  assign n11063 = n11062 ^ n4374 ^ 1'b0 ;
  assign n11064 = ~n1725 & n11063 ;
  assign n11065 = n11064 ^ n1450 ^ 1'b0 ;
  assign n11067 = n8594 ^ n1298 ^ 1'b0 ;
  assign n11068 = n11067 ^ n5701 ^ 1'b0 ;
  assign n11069 = n11068 ^ n8340 ^ n3379 ;
  assign n11066 = n3389 & ~n6088 ;
  assign n11070 = n11069 ^ n11066 ^ 1'b0 ;
  assign n11071 = ~n11065 & n11070 ;
  assign n11072 = n8224 ^ n4276 ^ n458 ;
  assign n11073 = n9017 ^ n5009 ^ 1'b0 ;
  assign n11074 = n2764 & ~n11073 ;
  assign n11075 = n3096 & n9100 ;
  assign n11076 = n11075 ^ n7541 ^ 1'b0 ;
  assign n11077 = ~n3211 & n11076 ;
  assign n11078 = n8084 ^ n3564 ^ 1'b0 ;
  assign n11079 = n4537 ^ n1729 ^ 1'b0 ;
  assign n11080 = n3603 | n11079 ;
  assign n11081 = ~n2711 & n2958 ;
  assign n11082 = n4216 & ~n9774 ;
  assign n11083 = n11082 ^ n3910 ^ 1'b0 ;
  assign n11084 = n274 & ~n2304 ;
  assign n11085 = ~n2013 & n4229 ;
  assign n11086 = n11085 ^ n2180 ^ 1'b0 ;
  assign n11087 = n7588 ^ n2265 ^ 1'b0 ;
  assign n11088 = n5410 ^ n2445 ^ 1'b0 ;
  assign n11089 = ~n7484 & n11088 ;
  assign n11090 = n2203 ^ n1189 ^ 1'b0 ;
  assign n11091 = n11089 & n11090 ;
  assign n11092 = n11087 & n11091 ;
  assign n11093 = n11086 & n11092 ;
  assign n11094 = n3121 ^ n511 ^ 1'b0 ;
  assign n11095 = n6476 & n10679 ;
  assign n11096 = n11095 ^ n9618 ^ 1'b0 ;
  assign n11101 = n459 & ~n3003 ;
  assign n11102 = ~n5459 & n11101 ;
  assign n11097 = n6886 ^ n2706 ^ x101 ;
  assign n11098 = n5921 | n11097 ;
  assign n11099 = n11098 ^ n2584 ^ 1'b0 ;
  assign n11100 = ~n9634 & n11099 ;
  assign n11103 = n11102 ^ n11100 ^ 1'b0 ;
  assign n11107 = n853 | n1369 ;
  assign n11108 = n11107 ^ n4306 ^ 1'b0 ;
  assign n11106 = ~n899 & n1889 ;
  assign n11104 = n799 | n4768 ;
  assign n11105 = n6448 | n11104 ;
  assign n11109 = n11108 ^ n11106 ^ n11105 ;
  assign n11110 = n9721 ^ n2614 ^ n1032 ;
  assign n11111 = n5685 & ~n6618 ;
  assign n11112 = n11111 ^ n2472 ^ 1'b0 ;
  assign n11113 = n3951 & ~n6151 ;
  assign n11114 = n11113 ^ n1822 ^ 1'b0 ;
  assign n11115 = n2240 ^ n1964 ^ 1'b0 ;
  assign n11116 = n2442 & n11115 ;
  assign n11117 = n8380 ^ n2234 ^ 1'b0 ;
  assign n11118 = n11116 & n11117 ;
  assign n11119 = n6045 ^ n5714 ^ 1'b0 ;
  assign n11120 = n312 | n4310 ;
  assign n11121 = n11120 ^ n5261 ^ 1'b0 ;
  assign n11122 = n4292 & ~n11121 ;
  assign n11123 = n7156 ^ n2062 ^ 1'b0 ;
  assign n11124 = ~n627 & n11123 ;
  assign n11125 = n2015 & ~n11124 ;
  assign n11126 = ~n4867 & n7160 ;
  assign n11127 = n11126 ^ n3795 ^ 1'b0 ;
  assign n11128 = n3001 & n11127 ;
  assign n11129 = n1116 | n2736 ;
  assign n11130 = n276 | n11129 ;
  assign n11131 = n9478 ^ n4906 ^ 1'b0 ;
  assign n11132 = ~n5369 & n11131 ;
  assign n11133 = n11132 ^ n3624 ^ 1'b0 ;
  assign n11134 = n8592 & n11133 ;
  assign n11135 = n6585 ^ n3508 ^ n579 ;
  assign n11136 = ~n9487 & n10529 ;
  assign n11137 = ~n3321 & n11136 ;
  assign n11138 = n11137 ^ n7433 ^ 1'b0 ;
  assign n11140 = x168 & n4876 ;
  assign n11139 = n7107 | n8955 ;
  assign n11141 = n11140 ^ n11139 ^ 1'b0 ;
  assign n11142 = n4388 | n5958 ;
  assign n11143 = n5448 | n7484 ;
  assign n11144 = n2951 | n11143 ;
  assign n11145 = n6547 & n7467 ;
  assign n11146 = n11145 ^ n10968 ^ 1'b0 ;
  assign n11147 = ( n5667 & n9351 ) | ( n5667 & n11146 ) | ( n9351 & n11146 ) ;
  assign n11148 = n1826 | n6964 ;
  assign n11151 = n423 | n1160 ;
  assign n11149 = n4070 | n9407 ;
  assign n11150 = n5457 & n11149 ;
  assign n11152 = n11151 ^ n11150 ^ 1'b0 ;
  assign n11153 = n11152 ^ n7002 ^ 1'b0 ;
  assign n11154 = n1466 | n6001 ;
  assign n11155 = ( n904 & n1870 ) | ( n904 & ~n5540 ) | ( n1870 & ~n5540 ) ;
  assign n11156 = ~n5227 & n11155 ;
  assign n11157 = n11154 & n11156 ;
  assign n11158 = n11157 ^ n5016 ^ n4509 ;
  assign n11159 = n6049 ^ n4993 ^ 1'b0 ;
  assign n11160 = x148 & n10442 ;
  assign n11161 = n11159 & n11160 ;
  assign n11162 = n11161 ^ n1258 ^ 1'b0 ;
  assign n11163 = n11162 ^ n5908 ^ 1'b0 ;
  assign n11164 = n8645 & n11163 ;
  assign n11166 = n2670 ^ n2282 ^ 1'b0 ;
  assign n11165 = n1219 & n4303 ;
  assign n11167 = n11166 ^ n11165 ^ 1'b0 ;
  assign n11168 = ~n1639 & n6338 ;
  assign n11169 = x156 & ~n1227 ;
  assign n11170 = ~x73 & n11169 ;
  assign n11171 = n1085 & ~n1728 ;
  assign n11172 = n11170 & n11171 ;
  assign n11173 = n8498 ^ n5303 ^ 1'b0 ;
  assign n11174 = n4509 & n11173 ;
  assign n11176 = ~n2229 & n7602 ;
  assign n11177 = n11176 ^ n1926 ^ 1'b0 ;
  assign n11178 = n4197 & ~n11177 ;
  assign n11175 = n8850 ^ n5165 ^ n534 ;
  assign n11179 = n11178 ^ n11175 ^ 1'b0 ;
  assign n11180 = n1721 & ~n5156 ;
  assign n11181 = n11180 ^ n4612 ^ 1'b0 ;
  assign n11182 = n11181 ^ n3502 ^ 1'b0 ;
  assign n11183 = n2796 ^ n913 ^ 1'b0 ;
  assign n11184 = n890 & n11183 ;
  assign n11185 = n3288 ^ n2096 ^ 1'b0 ;
  assign n11186 = n1710 & ~n11185 ;
  assign n11190 = n6033 ^ n3910 ^ 1'b0 ;
  assign n11191 = ~n5234 & n11190 ;
  assign n11187 = n9268 ^ n6495 ^ 1'b0 ;
  assign n11188 = n2371 | n11187 ;
  assign n11189 = n11188 ^ n8952 ^ 1'b0 ;
  assign n11192 = n11191 ^ n11189 ^ 1'b0 ;
  assign n11193 = n2331 & n11192 ;
  assign n11194 = ~n1281 & n11193 ;
  assign n11195 = ~n10378 & n11194 ;
  assign n11196 = ~n4232 & n9013 ;
  assign n11197 = ( n1678 & n8978 ) | ( n1678 & ~n11196 ) | ( n8978 & ~n11196 ) ;
  assign n11198 = n6582 & ~n8832 ;
  assign n11199 = n11198 ^ n1911 ^ 1'b0 ;
  assign n11200 = n6292 & n11199 ;
  assign n11201 = n11200 ^ n334 ^ 1'b0 ;
  assign n11202 = n11201 ^ n1342 ^ 1'b0 ;
  assign n11203 = n11197 & ~n11202 ;
  assign n11204 = n5655 | n10733 ;
  assign n11205 = n328 & n3372 ;
  assign n11206 = n5665 & n11205 ;
  assign n11207 = n1599 & ~n11206 ;
  assign n11208 = n11207 ^ n2964 ^ 1'b0 ;
  assign n11215 = n1756 & ~n4518 ;
  assign n11216 = n4518 & n11215 ;
  assign n11217 = n428 & ~n11216 ;
  assign n11218 = n11216 & n11217 ;
  assign n11219 = n446 | n7466 ;
  assign n11220 = n7466 & ~n11219 ;
  assign n11221 = n11220 ^ n5933 ^ 1'b0 ;
  assign n11222 = ~n11218 & n11221 ;
  assign n11211 = n380 | n1649 ;
  assign n11212 = ~n9132 & n11211 ;
  assign n11213 = ~n11211 & n11212 ;
  assign n11209 = n471 | n956 ;
  assign n11210 = n471 & ~n11209 ;
  assign n11214 = n11213 ^ n11210 ^ 1'b0 ;
  assign n11223 = n11222 ^ n11214 ^ 1'b0 ;
  assign n11224 = ~n10724 & n11223 ;
  assign n11225 = n503 & n4416 ;
  assign n11226 = n11225 ^ n4948 ^ 1'b0 ;
  assign n11227 = ( n1714 & ~n5746 ) | ( n1714 & n11226 ) | ( ~n5746 & n11226 ) ;
  assign n11228 = n7130 ^ n404 ^ 1'b0 ;
  assign n11229 = ~n6678 & n11228 ;
  assign n11230 = n2428 ^ n2122 ^ x172 ;
  assign n11231 = n11230 ^ n4959 ^ 1'b0 ;
  assign n11232 = n11229 | n11231 ;
  assign n11233 = n4603 & ~n11232 ;
  assign n11234 = n11227 & n11233 ;
  assign n11235 = n1867 & n4895 ;
  assign n11236 = x8 & n8900 ;
  assign n11237 = n6228 & n11236 ;
  assign n11238 = n7116 & n8768 ;
  assign n11239 = n5446 & n11238 ;
  assign n11240 = ~n4766 & n11013 ;
  assign n11241 = n8072 & n11240 ;
  assign n11242 = x25 & ~n7351 ;
  assign n11243 = ~n7179 & n11242 ;
  assign n11244 = n11243 ^ n11030 ^ n4563 ;
  assign n11245 = n8784 ^ n7342 ^ 1'b0 ;
  assign n11246 = n9736 ^ n5369 ^ 1'b0 ;
  assign n11247 = n1004 | n11246 ;
  assign n11248 = n8355 ^ n1621 ^ 1'b0 ;
  assign n11249 = n6726 | n11248 ;
  assign n11250 = ~n665 & n3240 ;
  assign n11251 = n11250 ^ n5634 ^ 1'b0 ;
  assign n11252 = n11251 ^ n6133 ^ 1'b0 ;
  assign n11253 = n287 | n11252 ;
  assign n11254 = n3571 ^ x155 ^ 1'b0 ;
  assign n11255 = n5521 | n11254 ;
  assign n11256 = n2747 | n7613 ;
  assign n11257 = n10481 ^ n6653 ^ 1'b0 ;
  assign n11258 = n944 | n1981 ;
  assign n11259 = n11258 ^ n1880 ^ 1'b0 ;
  assign n11260 = n6864 & n11259 ;
  assign n11261 = n3864 ^ n1290 ^ 1'b0 ;
  assign n11262 = n10404 & n11261 ;
  assign n11263 = n4384 ^ n3762 ^ 1'b0 ;
  assign n11264 = n11263 ^ n2564 ^ 1'b0 ;
  assign n11265 = x143 & n2159 ;
  assign n11266 = n5783 & ~n11265 ;
  assign n11267 = n1809 & n11266 ;
  assign n11268 = n11267 ^ n3724 ^ 1'b0 ;
  assign n11269 = n11268 ^ n7631 ^ 1'b0 ;
  assign n11273 = n9721 ^ x9 ^ 1'b0 ;
  assign n11274 = n4869 | n11273 ;
  assign n11270 = ( n413 & n2418 ) | ( n413 & n4803 ) | ( n2418 & n4803 ) ;
  assign n11271 = n11270 ^ n2589 ^ 1'b0 ;
  assign n11272 = n11271 ^ n9284 ^ n7370 ;
  assign n11275 = n11274 ^ n11272 ^ 1'b0 ;
  assign n11276 = ~n3034 & n6564 ;
  assign n11277 = ( x120 & ~n420 ) | ( x120 & n1276 ) | ( ~n420 & n1276 ) ;
  assign n11278 = n4576 ^ n631 ^ 1'b0 ;
  assign n11279 = n7798 & n11278 ;
  assign n11280 = n11094 ^ n7831 ^ n796 ;
  assign n11283 = n3073 ^ n1336 ^ 1'b0 ;
  assign n11281 = n4553 ^ n3670 ^ 1'b0 ;
  assign n11282 = n500 | n11281 ;
  assign n11284 = n11283 ^ n11282 ^ 1'b0 ;
  assign n11285 = n8993 ^ n432 ^ 1'b0 ;
  assign n11286 = n11285 ^ n3325 ^ 1'b0 ;
  assign n11287 = n3405 & n11286 ;
  assign n11288 = ( ~n4204 & n4970 ) | ( ~n4204 & n9778 ) | ( n4970 & n9778 ) ;
  assign n11289 = ~n1301 & n7007 ;
  assign n11290 = n11289 ^ n10584 ^ 1'b0 ;
  assign n11291 = n11290 ^ n8358 ^ n3530 ;
  assign n11292 = n5061 ^ n1420 ^ 1'b0 ;
  assign n11294 = ~n5252 & n8855 ;
  assign n11295 = ~n1989 & n11294 ;
  assign n11293 = n3757 & n11040 ;
  assign n11296 = n11295 ^ n11293 ^ 1'b0 ;
  assign n11297 = n11296 ^ n7407 ^ 1'b0 ;
  assign n11298 = n11297 ^ n4837 ^ 1'b0 ;
  assign n11299 = n11292 & n11298 ;
  assign n11300 = n1735 & n6038 ;
  assign n11301 = n11300 ^ n6599 ^ 1'b0 ;
  assign n11302 = n11301 ^ n9853 ^ n7641 ;
  assign n11303 = n11302 ^ n289 ^ 1'b0 ;
  assign n11304 = n1447 | n1514 ;
  assign n11305 = n1447 & ~n11304 ;
  assign n11306 = n3966 & n7736 ;
  assign n11307 = ~n7736 & n11306 ;
  assign n11308 = n5087 | n11307 ;
  assign n11309 = n11307 & ~n11308 ;
  assign n11310 = n11305 | n11309 ;
  assign n11311 = n11303 | n11310 ;
  assign n11313 = n1157 & ~n2463 ;
  assign n11312 = n2592 & n4824 ;
  assign n11314 = n11313 ^ n11312 ^ 1'b0 ;
  assign n11315 = ~n483 & n1333 ;
  assign n11316 = n4499 & n11315 ;
  assign n11317 = n2061 | n11316 ;
  assign n11318 = n1989 | n11317 ;
  assign n11319 = ~n5722 & n11318 ;
  assign n11320 = n4537 ^ n858 ^ 1'b0 ;
  assign n11321 = n7723 ^ n1101 ^ 1'b0 ;
  assign n11322 = n4355 | n11321 ;
  assign n11323 = n11322 ^ n7130 ^ 1'b0 ;
  assign n11324 = n3613 & n11323 ;
  assign n11325 = n2259 ^ n1714 ^ 1'b0 ;
  assign n11326 = n9294 & ~n11325 ;
  assign n11327 = n1963 & ~n2191 ;
  assign n11328 = n8052 ^ n5786 ^ 1'b0 ;
  assign n11329 = n7368 ^ n2868 ^ 1'b0 ;
  assign n11330 = n2584 & n11329 ;
  assign n11331 = n1495 | n7742 ;
  assign n11332 = n4941 & n11331 ;
  assign n11333 = ~n9391 & n11332 ;
  assign n11334 = n7513 ^ n6755 ^ 1'b0 ;
  assign n11335 = n2098 & n3887 ;
  assign n11336 = ~n1832 & n11335 ;
  assign n11337 = n3106 | n8225 ;
  assign n11338 = n11337 ^ n1621 ^ 1'b0 ;
  assign n11339 = n3574 & ~n11338 ;
  assign n11340 = n11065 ^ n657 ^ 1'b0 ;
  assign n11341 = n3820 & ~n4293 ;
  assign n11342 = ~n2516 & n7794 ;
  assign n11343 = ~n1504 & n5596 ;
  assign n11344 = n11343 ^ n355 ^ 1'b0 ;
  assign n11345 = n11344 ^ n2210 ^ 1'b0 ;
  assign n11346 = n11342 & n11345 ;
  assign n11347 = x241 & ~n2497 ;
  assign n11348 = n6626 & ~n7763 ;
  assign n11349 = n595 & n3380 ;
  assign n11350 = n4867 | n11349 ;
  assign n11351 = n11348 | n11350 ;
  assign n11352 = ~n2474 & n2785 ;
  assign n11353 = ~n11351 & n11352 ;
  assign n11354 = n8011 ^ n1322 ^ 1'b0 ;
  assign n11355 = n11354 ^ n3041 ^ 1'b0 ;
  assign n11356 = n1045 ^ n888 ^ 1'b0 ;
  assign n11357 = n11356 ^ n2022 ^ n963 ;
  assign n11358 = n5627 ^ n1245 ^ 1'b0 ;
  assign n11359 = n7198 | n8822 ;
  assign n11360 = ~n1382 & n3007 ;
  assign n11361 = n11360 ^ n2208 ^ 1'b0 ;
  assign n11362 = n3114 | n10543 ;
  assign n11363 = n9289 & n11362 ;
  assign n11364 = n5700 & n11363 ;
  assign n11365 = ( ~n7827 & n8466 ) | ( ~n7827 & n11364 ) | ( n8466 & n11364 ) ;
  assign n11366 = n3213 ^ n3118 ^ 1'b0 ;
  assign n11367 = n4970 ^ n3967 ^ 1'b0 ;
  assign n11368 = n2929 & n11367 ;
  assign n11369 = n11366 & n11368 ;
  assign n11370 = ~n957 & n7732 ;
  assign n11371 = n11370 ^ n9218 ^ 1'b0 ;
  assign n11372 = n6315 | n11371 ;
  assign n11373 = n2983 | n8835 ;
  assign n11374 = ( ~n532 & n968 ) | ( ~n532 & n1023 ) | ( n968 & n1023 ) ;
  assign n11375 = ( n618 & ~n914 ) | ( n618 & n1684 ) | ( ~n914 & n1684 ) ;
  assign n11376 = ~n2311 & n6990 ;
  assign n11377 = n11375 & n11376 ;
  assign n11378 = ~n988 & n1018 ;
  assign n11379 = n11378 ^ n913 ^ 1'b0 ;
  assign n11380 = ~n2980 & n5078 ;
  assign n11381 = n11380 ^ n9644 ^ 1'b0 ;
  assign n11382 = n11381 ^ n7624 ^ 1'b0 ;
  assign n11383 = n8452 & ~n8724 ;
  assign n11384 = n8725 ^ x43 ^ 1'b0 ;
  assign n11385 = n10137 ^ n3007 ^ 1'b0 ;
  assign n11386 = ~n1871 & n11385 ;
  assign n11387 = n1579 & n11272 ;
  assign n11388 = n2355 & n11387 ;
  assign n11389 = n477 & ~n6360 ;
  assign n11390 = n9780 & ~n11389 ;
  assign n11391 = n6991 ^ x151 ^ 1'b0 ;
  assign n11392 = n6727 | n11391 ;
  assign n11393 = n1503 | n2354 ;
  assign n11394 = n11393 ^ n4698 ^ 1'b0 ;
  assign n11395 = n2703 | n11394 ;
  assign n11396 = n11395 ^ n7223 ^ 1'b0 ;
  assign n11397 = n3547 & n7971 ;
  assign n11398 = n11397 ^ n3231 ^ 1'b0 ;
  assign n11399 = n11398 ^ n8201 ^ 1'b0 ;
  assign n11400 = n6712 ^ n5840 ^ 1'b0 ;
  assign n11401 = n11400 ^ n268 ^ 1'b0 ;
  assign n11402 = n8683 ^ n8041 ^ 1'b0 ;
  assign n11403 = n6627 & ~n9438 ;
  assign n11404 = n5208 & n11403 ;
  assign n11405 = n11404 ^ n9360 ^ 1'b0 ;
  assign n11408 = n434 & ~n4718 ;
  assign n11409 = n11408 ^ n7490 ^ 1'b0 ;
  assign n11406 = n6260 ^ n5089 ^ 1'b0 ;
  assign n11407 = n10946 & ~n11406 ;
  assign n11410 = n11409 ^ n11407 ^ 1'b0 ;
  assign n11411 = n8532 & n11410 ;
  assign n11414 = n3731 | n4679 ;
  assign n11413 = ( n2688 & ~n7532 ) | ( n2688 & n7671 ) | ( ~n7532 & n7671 ) ;
  assign n11412 = n8087 ^ n1419 ^ 1'b0 ;
  assign n11415 = n11414 ^ n11413 ^ n11412 ;
  assign n11416 = n8466 ^ n5857 ^ n1649 ;
  assign n11425 = ~n677 & n1810 ;
  assign n11426 = n677 & n11425 ;
  assign n11427 = n11426 ^ n4327 ^ 1'b0 ;
  assign n11417 = ~n1437 & n1980 ;
  assign n11418 = n1437 & n11417 ;
  assign n11419 = n10356 | n11418 ;
  assign n11420 = n10356 & ~n11419 ;
  assign n11421 = n6895 | n11420 ;
  assign n11422 = n6895 & ~n11421 ;
  assign n11423 = ( n3535 & n7358 ) | ( n3535 & n9253 ) | ( n7358 & n9253 ) ;
  assign n11424 = ~n11422 & n11423 ;
  assign n11428 = n11427 ^ n11424 ^ 1'b0 ;
  assign n11429 = n6179 ^ n3655 ^ n283 ;
  assign n11430 = ~n2764 & n4093 ;
  assign n11431 = n11429 & ~n11430 ;
  assign n11432 = n4563 ^ n2817 ^ 1'b0 ;
  assign n11433 = n346 | n11432 ;
  assign n11434 = n11433 ^ n913 ^ 1'b0 ;
  assign n11435 = n5937 & n11434 ;
  assign n11436 = n11435 ^ n5936 ^ 1'b0 ;
  assign n11437 = ~x198 & n11436 ;
  assign n11442 = ~n1491 & n2912 ;
  assign n11438 = n6689 ^ n5842 ^ 1'b0 ;
  assign n11439 = n5021 & ~n11438 ;
  assign n11440 = n9383 ^ n5913 ^ 1'b0 ;
  assign n11441 = n11439 & ~n11440 ;
  assign n11443 = n11442 ^ n11441 ^ 1'b0 ;
  assign n11444 = n8476 ^ n2496 ^ 1'b0 ;
  assign n11445 = ~n3023 & n6024 ;
  assign n11446 = ~n4335 & n11445 ;
  assign n11447 = n11446 ^ n9117 ^ 1'b0 ;
  assign n11449 = x162 & ~n2521 ;
  assign n11450 = n3025 & n11449 ;
  assign n11448 = n3429 & ~n5099 ;
  assign n11451 = n11450 ^ n11448 ^ 1'b0 ;
  assign n11452 = n2646 & ~n11451 ;
  assign n11454 = x155 & n8064 ;
  assign n11453 = n3302 & ~n10408 ;
  assign n11455 = n11454 ^ n11453 ^ 1'b0 ;
  assign n11456 = n6200 ^ n5767 ^ 1'b0 ;
  assign n11457 = ( n1103 & n7515 ) | ( n1103 & n11456 ) | ( n7515 & n11456 ) ;
  assign n11458 = x242 & n3508 ;
  assign n11459 = ~n1462 & n3683 ;
  assign n11460 = n2356 & n10336 ;
  assign n11461 = n7326 ^ n666 ^ 1'b0 ;
  assign n11462 = n5692 ^ n1125 ^ 1'b0 ;
  assign n11463 = ~n9835 & n11462 ;
  assign n11464 = ~n4567 & n11463 ;
  assign n11465 = n3105 | n9041 ;
  assign n11466 = n1931 & n11465 ;
  assign n11467 = ~x253 & n11466 ;
  assign n11468 = ~x132 & n3010 ;
  assign n11469 = n11344 ^ n523 ^ 1'b0 ;
  assign n11470 = n1069 ^ x209 ^ 1'b0 ;
  assign n11471 = n3198 | n11470 ;
  assign n11472 = x0 | n11471 ;
  assign n11473 = n6332 ^ x123 ^ 1'b0 ;
  assign n11474 = n11472 & n11473 ;
  assign n11475 = n11469 & n11474 ;
  assign n11476 = n11475 ^ n5837 ^ 1'b0 ;
  assign n11477 = n2738 ^ n1365 ^ 1'b0 ;
  assign n11478 = n3468 ^ n3351 ^ 1'b0 ;
  assign n11479 = n3180 | n11478 ;
  assign n11480 = n11479 ^ n8059 ^ 1'b0 ;
  assign n11481 = n11477 | n11480 ;
  assign n11482 = n2830 & ~n11481 ;
  assign n11483 = n6607 ^ n6604 ^ n5333 ;
  assign n11484 = n3142 & ~n7145 ;
  assign n11485 = ~n1316 & n11484 ;
  assign n11486 = n8941 | n11485 ;
  assign n11487 = n11486 ^ n11446 ^ 1'b0 ;
  assign n11488 = n3705 & n6994 ;
  assign n11489 = n11488 ^ n6510 ^ 1'b0 ;
  assign n11490 = n7173 | n11489 ;
  assign n11491 = n7495 | n11490 ;
  assign n11492 = n3850 & n11491 ;
  assign n11493 = n11492 ^ n8514 ^ 1'b0 ;
  assign n11494 = n5366 ^ n5119 ^ n2983 ;
  assign n11495 = n9397 ^ n8103 ^ 1'b0 ;
  assign n11496 = n11494 & ~n11495 ;
  assign n11497 = ( n1871 & ~n10878 ) | ( n1871 & n11496 ) | ( ~n10878 & n11496 ) ;
  assign n11498 = n11497 ^ n1250 ^ 1'b0 ;
  assign n11499 = n2202 ^ n858 ^ n423 ;
  assign n11500 = n3546 & n8347 ;
  assign n11501 = n11499 & ~n11500 ;
  assign n11502 = ~n11262 & n11501 ;
  assign n11503 = n11206 ^ n7743 ^ 1'b0 ;
  assign n11504 = n2739 | n11503 ;
  assign n11505 = n1228 & ~n9074 ;
  assign n11506 = ~n708 & n11505 ;
  assign n11510 = n3747 & ~n4946 ;
  assign n11511 = n11510 ^ n3253 ^ 1'b0 ;
  assign n11507 = n3308 ^ n908 ^ 1'b0 ;
  assign n11508 = n5050 | n11507 ;
  assign n11509 = n8334 | n11508 ;
  assign n11512 = n11511 ^ n11509 ^ 1'b0 ;
  assign n11513 = n4241 | n11512 ;
  assign n11514 = n3199 | n11513 ;
  assign n11515 = ( ~n4193 & n11506 ) | ( ~n4193 & n11514 ) | ( n11506 & n11514 ) ;
  assign n11516 = x204 & n4599 ;
  assign n11517 = n1346 & n11516 ;
  assign n11518 = n2006 & ~n4018 ;
  assign n11519 = n11518 ^ n4691 ^ 1'b0 ;
  assign n11520 = n6889 & n11519 ;
  assign n11521 = ~n11517 & n11520 ;
  assign n11522 = ~n323 & n2446 ;
  assign n11523 = ~n4995 & n11522 ;
  assign n11524 = n780 | n4748 ;
  assign n11525 = n1084 & ~n11524 ;
  assign n11526 = n11525 ^ n7298 ^ 1'b0 ;
  assign n11527 = n11526 ^ n4242 ^ 1'b0 ;
  assign n11528 = ~n11523 & n11527 ;
  assign n11529 = n11528 ^ n9446 ^ 1'b0 ;
  assign n11530 = n11521 | n11529 ;
  assign n11531 = n11530 ^ n2638 ^ 1'b0 ;
  assign n11532 = n1571 ^ x231 ^ 1'b0 ;
  assign n11533 = n6761 | n11532 ;
  assign n11534 = ( ~n4691 & n6875 ) | ( ~n4691 & n11533 ) | ( n6875 & n11533 ) ;
  assign n11535 = x74 & ~n2476 ;
  assign n11536 = ~n5531 & n11535 ;
  assign n11537 = ~n2725 & n11536 ;
  assign n11538 = n11537 ^ n2881 ^ 1'b0 ;
  assign n11539 = n4413 & n11538 ;
  assign n11540 = n11539 ^ n4053 ^ 1'b0 ;
  assign n11541 = n5142 | n11540 ;
  assign n11542 = x143 & n8592 ;
  assign n11543 = n5891 ^ n2945 ^ 1'b0 ;
  assign n11544 = n11542 & n11543 ;
  assign n11545 = n7555 & ~n11544 ;
  assign n11546 = n675 & ~n8072 ;
  assign n11547 = n11545 & n11546 ;
  assign n11548 = n1486 & n3171 ;
  assign n11549 = n5859 & n10240 ;
  assign n11550 = n3050 | n5873 ;
  assign n11551 = n11550 ^ n7809 ^ 1'b0 ;
  assign n11552 = n885 & ~n11551 ;
  assign n11553 = n954 & n10925 ;
  assign n11554 = n11553 ^ n6398 ^ 1'b0 ;
  assign n11555 = n11554 ^ n7109 ^ 1'b0 ;
  assign n11556 = n1085 & ~n11555 ;
  assign n11558 = n6069 ^ n3926 ^ 1'b0 ;
  assign n11557 = ( n8863 & ~n10541 ) | ( n8863 & n10938 ) | ( ~n10541 & n10938 ) ;
  assign n11559 = n11558 ^ n11557 ^ 1'b0 ;
  assign n11560 = n11556 & n11559 ;
  assign n11561 = ( n7375 & ~n9299 ) | ( n7375 & n11560 ) | ( ~n9299 & n11560 ) ;
  assign n11562 = n4940 ^ n3156 ^ 1'b0 ;
  assign n11563 = ~n579 & n11562 ;
  assign n11564 = n4400 & n11563 ;
  assign n11565 = n11564 ^ n274 ^ 1'b0 ;
  assign n11566 = ~n1725 & n11565 ;
  assign n11567 = ( n4555 & n7002 ) | ( n4555 & n11566 ) | ( n7002 & n11566 ) ;
  assign n11568 = n11567 ^ n8167 ^ 1'b0 ;
  assign n11569 = n540 & n7736 ;
  assign n11570 = ~n1167 & n11569 ;
  assign n11571 = n11570 ^ n5135 ^ 1'b0 ;
  assign n11572 = n5082 ^ n3423 ^ 1'b0 ;
  assign n11573 = n9267 ^ n2559 ^ 1'b0 ;
  assign n11574 = n11572 & ~n11573 ;
  assign n11575 = ~n4294 & n11574 ;
  assign n11576 = ~n11571 & n11575 ;
  assign n11579 = n4542 ^ n1025 ^ 1'b0 ;
  assign n11580 = n8121 | n11579 ;
  assign n11581 = n11580 ^ n3319 ^ 1'b0 ;
  assign n11577 = n709 | n1877 ;
  assign n11578 = n11577 ^ n5440 ^ 1'b0 ;
  assign n11582 = n11581 ^ n11578 ^ 1'b0 ;
  assign n11583 = n8733 | n11582 ;
  assign n11584 = n11583 ^ n957 ^ 1'b0 ;
  assign n11585 = ~n1570 & n11584 ;
  assign n11586 = n10609 ^ n7439 ^ 1'b0 ;
  assign n11587 = n6877 ^ n794 ^ 1'b0 ;
  assign n11588 = n2730 | n11587 ;
  assign n11589 = n11588 ^ x118 ^ 1'b0 ;
  assign n11590 = n11589 ^ n1532 ^ n1492 ;
  assign n11591 = n984 & n11590 ;
  assign n11592 = ~n11586 & n11591 ;
  assign n11593 = n5675 & ~n11355 ;
  assign n11594 = n8760 ^ n6456 ^ 1'b0 ;
  assign n11595 = n5163 & ~n9360 ;
  assign n11596 = n11595 ^ n10167 ^ 1'b0 ;
  assign n11597 = n8455 ^ n1585 ^ 1'b0 ;
  assign n11598 = ~n11159 & n11597 ;
  assign n11599 = n11598 ^ n8028 ^ 1'b0 ;
  assign n11600 = n11599 ^ n5041 ^ 1'b0 ;
  assign n11601 = n5009 ^ n1985 ^ 1'b0 ;
  assign n11602 = n11600 | n11601 ;
  assign n11603 = ( n5041 & ~n6797 ) | ( n5041 & n8729 ) | ( ~n6797 & n8729 ) ;
  assign n11604 = n1784 & n7015 ;
  assign n11605 = n11604 ^ n6116 ^ 1'b0 ;
  assign n11606 = ~n2896 & n11605 ;
  assign n11607 = ~n5522 & n9996 ;
  assign n11608 = n2534 & ~n3296 ;
  assign n11609 = n1220 | n1768 ;
  assign n11610 = n1851 ^ n1563 ^ 1'b0 ;
  assign n11611 = n2082 & n3844 ;
  assign n11612 = n11610 & n11611 ;
  assign n11613 = n11612 ^ n2319 ^ 1'b0 ;
  assign n11614 = n5425 ^ n3196 ^ 1'b0 ;
  assign n11615 = n2023 & ~n6572 ;
  assign n11616 = n10084 ^ n5695 ^ 1'b0 ;
  assign n11617 = x180 | n11616 ;
  assign n11618 = n11615 | n11617 ;
  assign n11619 = n11618 ^ n11043 ^ 1'b0 ;
  assign n11620 = n10942 ^ n3761 ^ 1'b0 ;
  assign n11621 = ~n618 & n11620 ;
  assign n11622 = n8455 ^ n416 ^ 1'b0 ;
  assign n11623 = n4437 ^ n2622 ^ 1'b0 ;
  assign n11624 = ( ~n1786 & n3293 ) | ( ~n1786 & n8087 ) | ( n3293 & n8087 ) ;
  assign n11625 = n9083 & n11624 ;
  assign n11626 = n9621 ^ n3840 ^ 1'b0 ;
  assign n11627 = ~n4693 & n7407 ;
  assign n11628 = n11626 & ~n11627 ;
  assign n11629 = n6723 | n11628 ;
  assign n11630 = n11629 ^ n5396 ^ 1'b0 ;
  assign n11631 = ~n4181 & n6271 ;
  assign n11632 = n11631 ^ n10270 ^ 1'b0 ;
  assign n11633 = ( n997 & ~n2506 ) | ( n997 & n4406 ) | ( ~n2506 & n4406 ) ;
  assign n11634 = ~n854 & n5830 ;
  assign n11635 = n1318 & ~n6338 ;
  assign n11636 = ~n11634 & n11635 ;
  assign n11637 = n8268 ^ n2554 ^ 1'b0 ;
  assign n11638 = n6241 | n11637 ;
  assign n11639 = n11638 ^ x91 ^ 1'b0 ;
  assign n11640 = n6464 & n11639 ;
  assign n11642 = ~n2710 & n5660 ;
  assign n11643 = ~n625 & n11642 ;
  assign n11644 = n5034 & ~n11643 ;
  assign n11641 = n2528 | n3432 ;
  assign n11645 = n11644 ^ n11641 ^ 1'b0 ;
  assign n11646 = n5462 ^ n1159 ^ 1'b0 ;
  assign n11647 = n1482 | n11646 ;
  assign n11648 = n5705 | n11647 ;
  assign n11649 = n11648 ^ n3704 ^ 1'b0 ;
  assign n11650 = ~n1778 & n11649 ;
  assign n11651 = ~n518 & n943 ;
  assign n11652 = n11651 ^ n11099 ^ 1'b0 ;
  assign n11653 = ~n6393 & n11652 ;
  assign n11654 = ~n2518 & n7504 ;
  assign n11655 = n11654 ^ n2083 ^ 1'b0 ;
  assign n11658 = n3913 | n9012 ;
  assign n11659 = n2795 | n11658 ;
  assign n11657 = n8612 ^ n2685 ^ 1'b0 ;
  assign n11656 = n5241 | n6465 ;
  assign n11660 = n11659 ^ n11657 ^ n11656 ;
  assign n11661 = n7594 ^ n1198 ^ 1'b0 ;
  assign n11662 = x104 & n11661 ;
  assign n11663 = n11662 ^ n8754 ^ 1'b0 ;
  assign n11664 = n10403 ^ n4775 ^ 1'b0 ;
  assign n11665 = n4948 | n11664 ;
  assign n11666 = ( ~n2082 & n2193 ) | ( ~n2082 & n7398 ) | ( n2193 & n7398 ) ;
  assign n11667 = n2986 & ~n3926 ;
  assign n11668 = n11667 ^ n2202 ^ 1'b0 ;
  assign n11669 = n10914 ^ n6943 ^ 1'b0 ;
  assign n11670 = ~n716 & n11669 ;
  assign n11671 = ~n11668 & n11670 ;
  assign n11672 = n5136 & n6412 ;
  assign n11673 = ~n10391 & n11672 ;
  assign n11674 = n776 & n11673 ;
  assign n11675 = n7256 & ~n7759 ;
  assign n11676 = n11675 ^ x218 ^ 1'b0 ;
  assign n11677 = ~n11412 & n11676 ;
  assign n11678 = n8230 & ~n11677 ;
  assign n11679 = n6511 ^ n983 ^ 1'b0 ;
  assign n11680 = n8163 & n11679 ;
  assign n11681 = n7749 & n11680 ;
  assign n11682 = n3496 & ~n4316 ;
  assign n11683 = ~n7723 & n11682 ;
  assign n11684 = ( n4985 & ~n8375 ) | ( n4985 & n11683 ) | ( ~n8375 & n11683 ) ;
  assign n11685 = ( n980 & n11681 ) | ( n980 & n11684 ) | ( n11681 & n11684 ) ;
  assign n11686 = n2308 & n4852 ;
  assign n11687 = n11686 ^ n9885 ^ 1'b0 ;
  assign n11688 = ~n2924 & n10670 ;
  assign n11689 = n11688 ^ n5986 ^ 1'b0 ;
  assign n11690 = ~n4131 & n4416 ;
  assign n11691 = n11690 ^ n11276 ^ 1'b0 ;
  assign n11692 = n8033 ^ n3258 ^ n1420 ;
  assign n11693 = n3149 & n11692 ;
  assign n11694 = n11693 ^ n5433 ^ 1'b0 ;
  assign n11695 = ( ~n2584 & n7970 ) | ( ~n2584 & n11694 ) | ( n7970 & n11694 ) ;
  assign n11696 = n11695 ^ n4869 ^ 1'b0 ;
  assign n11697 = n11696 ^ n8117 ^ 1'b0 ;
  assign n11698 = ~n8948 & n11697 ;
  assign n11699 = n1351 & n11698 ;
  assign n11700 = n2378 & ~n8778 ;
  assign n11701 = n4078 ^ n1093 ^ 1'b0 ;
  assign n11704 = n4366 ^ n2267 ^ 1'b0 ;
  assign n11705 = n1288 | n11704 ;
  assign n11706 = n2006 & n9549 ;
  assign n11707 = n11705 & n11706 ;
  assign n11708 = n11707 ^ n3249 ^ 1'b0 ;
  assign n11703 = ( n2162 & n7433 ) | ( n2162 & n8071 ) | ( n7433 & n8071 ) ;
  assign n11702 = n2297 ^ x69 ^ 1'b0 ;
  assign n11709 = n11708 ^ n11703 ^ n11702 ;
  assign n11710 = x0 & ~n7181 ;
  assign n11711 = x116 & ~n2491 ;
  assign n11712 = ~n11710 & n11711 ;
  assign n11713 = n3782 | n5139 ;
  assign n11714 = ( n2086 & ~n5557 ) | ( n2086 & n11713 ) | ( ~n5557 & n11713 ) ;
  assign n11715 = n9180 & ~n11714 ;
  assign n11716 = n2466 & n10985 ;
  assign n11717 = ~n632 & n11716 ;
  assign n11718 = n10612 | n11717 ;
  assign n11719 = n11715 | n11718 ;
  assign n11720 = n7951 ^ n4372 ^ 1'b0 ;
  assign n11721 = n8139 & ~n11720 ;
  assign n11722 = n4795 & ~n6464 ;
  assign n11723 = n9702 & ~n11042 ;
  assign n11724 = n10846 ^ n8406 ^ 1'b0 ;
  assign n11725 = n5402 | n11724 ;
  assign n11726 = n3250 & ~n7023 ;
  assign n11727 = n6059 & n11201 ;
  assign n11728 = ~n11726 & n11727 ;
  assign n11729 = n1828 & ~n11728 ;
  assign n11730 = ~n5932 & n11729 ;
  assign n11734 = ( n1023 & n4279 ) | ( n1023 & ~n9100 ) | ( n4279 & ~n9100 ) ;
  assign n11731 = n3042 | n5243 ;
  assign n11732 = n2783 & n11731 ;
  assign n11733 = ( ~n2284 & n8365 ) | ( ~n2284 & n11732 ) | ( n8365 & n11732 ) ;
  assign n11735 = n11734 ^ n11733 ^ 1'b0 ;
  assign n11736 = n407 & n5888 ;
  assign n11737 = n6627 & n11736 ;
  assign n11738 = ~n1932 & n6700 ;
  assign n11739 = n11738 ^ n3980 ^ 1'b0 ;
  assign n11740 = ~n11737 & n11739 ;
  assign n11741 = n11740 ^ n10248 ^ 1'b0 ;
  assign n11742 = n4718 & ~n10179 ;
  assign n11743 = n11742 ^ n2883 ^ 1'b0 ;
  assign n11744 = n4325 & n6912 ;
  assign n11745 = n7173 & n11744 ;
  assign n11746 = n749 & n3576 ;
  assign n11747 = n3763 & n11746 ;
  assign n11748 = n11747 ^ n817 ^ 1'b0 ;
  assign n11749 = n10289 & ~n11748 ;
  assign n11750 = n4929 ^ n1244 ^ x164 ;
  assign n11751 = n11750 ^ n6019 ^ 1'b0 ;
  assign n11752 = n11751 ^ n4864 ^ 1'b0 ;
  assign n11753 = n9464 & n11752 ;
  assign n11754 = n4715 | n11753 ;
  assign n11755 = ( n1001 & ~n4925 ) | ( n1001 & n7102 ) | ( ~n4925 & n7102 ) ;
  assign n11756 = n3415 ^ n359 ^ 1'b0 ;
  assign n11757 = n1900 | n11756 ;
  assign n11758 = n1581 | n11084 ;
  assign n11759 = ( ~x88 & n2232 ) | ( ~x88 & n8591 ) | ( n2232 & n8591 ) ;
  assign n11760 = n11759 ^ n2399 ^ 1'b0 ;
  assign n11761 = n728 & ~n3973 ;
  assign n11762 = n11761 ^ n3481 ^ 1'b0 ;
  assign n11763 = n11760 & n11762 ;
  assign n11764 = n4450 & ~n7120 ;
  assign n11765 = n1599 | n11764 ;
  assign n11766 = n7120 & n11765 ;
  assign n11767 = n9892 & ~n9916 ;
  assign n11768 = n5678 ^ n4366 ^ 1'b0 ;
  assign n11769 = n7089 & ~n11768 ;
  assign n11770 = n7135 & n8808 ;
  assign n11771 = n9816 & ~n11770 ;
  assign n11772 = n11771 ^ n7310 ^ 1'b0 ;
  assign n11773 = n2323 ^ n1451 ^ 1'b0 ;
  assign n11774 = n1543 & ~n3317 ;
  assign n11775 = n4169 & n11774 ;
  assign n11776 = n1936 & ~n3385 ;
  assign n11777 = n11776 ^ n5783 ^ 1'b0 ;
  assign n11778 = n9609 & ~n11777 ;
  assign n11779 = n7495 & n8421 ;
  assign n11780 = n3011 & n11779 ;
  assign n11781 = n2369 & ~n10306 ;
  assign n11782 = n11781 ^ n916 ^ 1'b0 ;
  assign n11784 = x65 | n3237 ;
  assign n11785 = ~n819 & n5883 ;
  assign n11786 = ~n11784 & n11785 ;
  assign n11787 = ~n3179 & n11786 ;
  assign n11783 = n3961 & n9527 ;
  assign n11788 = n11787 ^ n11783 ^ 1'b0 ;
  assign n11789 = n1099 ^ n809 ^ 1'b0 ;
  assign n11790 = ~n2215 & n11789 ;
  assign n11791 = n9540 & n11790 ;
  assign n11792 = n11791 ^ n611 ^ 1'b0 ;
  assign n11793 = ( n746 & ~n7932 ) | ( n746 & n11792 ) | ( ~n7932 & n11792 ) ;
  assign n11794 = n5100 | n5525 ;
  assign n11795 = ~n3952 & n4894 ;
  assign n11796 = n11794 | n11795 ;
  assign n11797 = n1129 & n6998 ;
  assign n11798 = ~n3776 & n11797 ;
  assign n11802 = n1473 & n5428 ;
  assign n11801 = n9569 ^ n6741 ^ n845 ;
  assign n11803 = n11802 ^ n11801 ^ 1'b0 ;
  assign n11799 = n1053 & n1252 ;
  assign n11800 = n9919 & n11799 ;
  assign n11804 = n11803 ^ n11800 ^ 1'b0 ;
  assign n11805 = n4425 | n5769 ;
  assign n11806 = n8734 & n9681 ;
  assign n11807 = n11806 ^ n663 ^ 1'b0 ;
  assign n11808 = n3413 ^ n789 ^ 1'b0 ;
  assign n11809 = n2354 ^ n1979 ^ 1'b0 ;
  assign n11810 = ~n8671 & n11809 ;
  assign n11811 = n11810 ^ n1030 ^ 1'b0 ;
  assign n11812 = ~n3179 & n4078 ;
  assign n11813 = n11812 ^ n3878 ^ 1'b0 ;
  assign n11814 = n3791 | n11813 ;
  assign n11815 = n6159 ^ n5745 ^ n5313 ;
  assign n11816 = n8525 ^ n7736 ^ 1'b0 ;
  assign n11817 = ~n6419 & n11816 ;
  assign n11818 = x212 & n3041 ;
  assign n11819 = n2407 | n11818 ;
  assign n11820 = ~n1936 & n11819 ;
  assign n11821 = n11820 ^ n10131 ^ 1'b0 ;
  assign n11822 = n888 & n9956 ;
  assign n11824 = n2598 ^ n525 ^ 1'b0 ;
  assign n11825 = n2004 & ~n11824 ;
  assign n11826 = n4109 & n11825 ;
  assign n11827 = n11826 ^ n1877 ^ 1'b0 ;
  assign n11828 = n3331 & n11827 ;
  assign n11829 = ~n1588 & n11828 ;
  assign n11823 = n8011 & ~n11816 ;
  assign n11830 = n11829 ^ n11823 ^ 1'b0 ;
  assign n11831 = n445 & n9992 ;
  assign n11832 = n11831 ^ n2697 ^ 1'b0 ;
  assign n11833 = n11830 & ~n11832 ;
  assign n11834 = n3446 ^ n2661 ^ 1'b0 ;
  assign n11835 = n2937 & n11834 ;
  assign n11836 = ( n8222 & n11833 ) | ( n8222 & n11835 ) | ( n11833 & n11835 ) ;
  assign n11839 = n1176 ^ x181 ^ x125 ;
  assign n11837 = n3926 ^ n433 ^ 1'b0 ;
  assign n11838 = n766 | n11837 ;
  assign n11840 = n11839 ^ n11838 ^ 1'b0 ;
  assign n11841 = n4042 ^ n1366 ^ 1'b0 ;
  assign n11842 = n11841 ^ n677 ^ 1'b0 ;
  assign n11843 = n10150 ^ n3663 ^ 1'b0 ;
  assign n11844 = n1169 & n5190 ;
  assign n11845 = ~n1169 & n11844 ;
  assign n11846 = n3088 ^ n289 ^ 1'b0 ;
  assign n11847 = n11846 ^ n2566 ^ 1'b0 ;
  assign n11848 = ~n11845 & n11847 ;
  assign n11849 = n10715 ^ n6836 ^ 1'b0 ;
  assign n11851 = n11025 ^ n1843 ^ 1'b0 ;
  assign n11852 = ~n5318 & n11851 ;
  assign n11850 = n8693 ^ n4648 ^ n2674 ;
  assign n11853 = n11852 ^ n11850 ^ 1'b0 ;
  assign n11854 = n2227 & n2685 ;
  assign n11855 = n3851 | n11854 ;
  assign n11856 = n11855 ^ n951 ^ 1'b0 ;
  assign n11857 = ~n1598 & n6851 ;
  assign n11858 = ~n3287 & n10246 ;
  assign n11859 = n9395 ^ n2164 ^ n1365 ;
  assign n11860 = n11859 ^ n4616 ^ 1'b0 ;
  assign n11861 = n1109 & ~n11860 ;
  assign n11862 = n9348 ^ n477 ^ x80 ;
  assign n11863 = ~n1153 & n11488 ;
  assign n11864 = ~n11862 & n11863 ;
  assign n11865 = n4512 | n7999 ;
  assign n11866 = n11865 ^ n2825 ^ 1'b0 ;
  assign n11867 = ~n4758 & n11866 ;
  assign n11868 = n3617 ^ n3370 ^ 1'b0 ;
  assign n11869 = n4177 | n11868 ;
  assign n11870 = n3596 | n11869 ;
  assign n11871 = n1084 ^ n618 ^ 1'b0 ;
  assign n11872 = n10100 & ~n11871 ;
  assign n11873 = n5915 & ~n9526 ;
  assign n11874 = n2378 ^ x153 ^ 1'b0 ;
  assign n11875 = ~n2846 & n11874 ;
  assign n11877 = ~n883 & n1147 ;
  assign n11878 = n933 & ~n11877 ;
  assign n11879 = n11878 ^ n725 ^ 1'b0 ;
  assign n11876 = x123 & ~n6187 ;
  assign n11880 = n11879 ^ n11876 ^ 1'b0 ;
  assign n11881 = n5888 ^ n3753 ^ 1'b0 ;
  assign n11882 = x121 & n11881 ;
  assign n11883 = n11880 & n11882 ;
  assign n11884 = n11749 ^ n3683 ^ 1'b0 ;
  assign n11885 = n11883 | n11884 ;
  assign n11886 = ( n894 & n5130 ) | ( n894 & ~n5746 ) | ( n5130 & ~n5746 ) ;
  assign n11887 = n11099 & ~n11886 ;
  assign n11888 = n3974 & ~n7126 ;
  assign n11889 = n2316 & n11888 ;
  assign n11890 = n2086 & ~n7310 ;
  assign n11891 = n11889 & n11890 ;
  assign n11894 = n1208 | n3337 ;
  assign n11895 = n7042 & ~n11894 ;
  assign n11896 = n6634 | n11895 ;
  assign n11897 = n11896 ^ n3615 ^ 1'b0 ;
  assign n11892 = n1020 ^ n737 ^ 1'b0 ;
  assign n11893 = n2668 & n11892 ;
  assign n11898 = n11897 ^ n11893 ^ 1'b0 ;
  assign n11899 = n3190 & n9601 ;
  assign n11900 = ~n3196 & n10514 ;
  assign n11901 = n11900 ^ n8092 ^ 1'b0 ;
  assign n11902 = n11901 ^ n2297 ^ 1'b0 ;
  assign n11903 = ~x170 & n3601 ;
  assign n11904 = n1982 & ~n11903 ;
  assign n11905 = n3910 & n11904 ;
  assign n11906 = ( n3305 & n3619 ) | ( n3305 & n11905 ) | ( n3619 & n11905 ) ;
  assign n11907 = ~n875 & n1369 ;
  assign n11908 = n11906 | n11907 ;
  assign n11909 = n11450 & ~n11908 ;
  assign n11910 = n3627 ^ n740 ^ 1'b0 ;
  assign n11911 = n4493 ^ n2712 ^ 1'b0 ;
  assign n11915 = n1914 & n3823 ;
  assign n11916 = n277 & n11915 ;
  assign n11912 = n1807 ^ n635 ^ 1'b0 ;
  assign n11913 = n6141 | n11912 ;
  assign n11914 = n4824 | n11913 ;
  assign n11917 = n11916 ^ n11914 ^ 1'b0 ;
  assign n11918 = n3396 & n7470 ;
  assign n11919 = n4678 & n11918 ;
  assign n11920 = n11919 ^ n6695 ^ 1'b0 ;
  assign n11921 = n4368 | n11920 ;
  assign n11922 = n11921 ^ n10812 ^ 1'b0 ;
  assign n11923 = n10276 & ~n11922 ;
  assign n11924 = n9079 ^ n3535 ^ 1'b0 ;
  assign n11925 = ~n8371 & n8763 ;
  assign n11926 = ~n9967 & n11925 ;
  assign n11927 = n7449 ^ n1094 ^ 1'b0 ;
  assign n11928 = n5842 ^ n1871 ^ 1'b0 ;
  assign n11929 = n10749 & n11928 ;
  assign n11930 = n10943 ^ n2810 ^ 1'b0 ;
  assign n11931 = n4827 & ~n11760 ;
  assign n11932 = ~n6786 & n11931 ;
  assign n11933 = n4161 & ~n11932 ;
  assign n11934 = n11802 ^ n7351 ^ 1'b0 ;
  assign n11935 = n3646 & ~n11175 ;
  assign n11936 = n6583 ^ n464 ^ 1'b0 ;
  assign n11937 = n10247 & ~n10942 ;
  assign n11938 = ~n10258 & n11937 ;
  assign n11939 = n11938 ^ n4053 ^ 1'b0 ;
  assign n11940 = n11877 ^ n2337 ^ 1'b0 ;
  assign n11941 = n2746 & n11940 ;
  assign n11942 = n6809 ^ n5697 ^ n4783 ;
  assign n11943 = n11941 & n11942 ;
  assign n11944 = n11943 ^ n7330 ^ 1'b0 ;
  assign n11945 = ~x20 & n11944 ;
  assign n11946 = n11945 ^ n7693 ^ 1'b0 ;
  assign n11947 = n11946 ^ n617 ^ 1'b0 ;
  assign n11948 = n2353 & n3059 ;
  assign n11949 = n3009 | n11948 ;
  assign n11950 = n11949 ^ n3641 ^ 1'b0 ;
  assign n11951 = n11950 ^ n4443 ^ n349 ;
  assign n11952 = n11951 ^ n9878 ^ 1'b0 ;
  assign n11953 = n2620 ^ n810 ^ 1'b0 ;
  assign n11954 = x147 & n11953 ;
  assign n11955 = ( n317 & n9900 ) | ( n317 & n11954 ) | ( n9900 & n11954 ) ;
  assign n11956 = ~n3277 & n3560 ;
  assign n11957 = n11956 ^ n11084 ^ 1'b0 ;
  assign n11960 = n3661 & n3942 ;
  assign n11961 = ~n5055 & n11960 ;
  assign n11962 = n1772 ^ n729 ^ 1'b0 ;
  assign n11963 = n11961 | n11962 ;
  assign n11959 = n8236 ^ n3603 ^ n1500 ;
  assign n11964 = n11963 ^ n11959 ^ 1'b0 ;
  assign n11958 = n6189 & ~n10422 ;
  assign n11965 = n11964 ^ n11958 ^ 1'b0 ;
  assign n11966 = n3110 ^ n614 ^ 1'b0 ;
  assign n11967 = n7558 | n11966 ;
  assign n11968 = n5962 | n11967 ;
  assign n11969 = n2149 & n4051 ;
  assign n11970 = n9766 | n11969 ;
  assign n11971 = n7918 & ~n11970 ;
  assign n11972 = n11971 ^ n6360 ^ 1'b0 ;
  assign n11973 = n11570 ^ n6700 ^ 1'b0 ;
  assign n11974 = ~n3171 & n11973 ;
  assign n11975 = ~n2047 & n11344 ;
  assign n11976 = n7635 ^ n2884 ^ 1'b0 ;
  assign n11977 = n7304 & ~n11976 ;
  assign n11978 = n11977 ^ n4186 ^ 1'b0 ;
  assign n11979 = n11978 ^ n10872 ^ 1'b0 ;
  assign n11980 = n5669 ^ n3410 ^ 1'b0 ;
  assign n11981 = n11980 ^ n5273 ^ x196 ;
  assign n11982 = n11981 ^ n8989 ^ 1'b0 ;
  assign n11983 = ( ~n3353 & n3685 ) | ( ~n3353 & n7401 ) | ( n3685 & n7401 ) ;
  assign n11984 = n3879 & n11983 ;
  assign n11985 = n2361 & n11984 ;
  assign n11986 = ~n619 & n1766 ;
  assign n11987 = n11986 ^ n6918 ^ 1'b0 ;
  assign n11988 = n5688 | n11987 ;
  assign n11989 = n3613 | n11676 ;
  assign n11990 = n11989 ^ n532 ^ 1'b0 ;
  assign n11991 = n3804 ^ n3408 ^ 1'b0 ;
  assign n11992 = ( n11988 & n11990 ) | ( n11988 & n11991 ) | ( n11990 & n11991 ) ;
  assign n11993 = n5733 | n11992 ;
  assign n11994 = n6341 | n11993 ;
  assign n11995 = ~n673 & n4150 ;
  assign n11996 = n2067 & n8723 ;
  assign n11997 = ~n2507 & n11996 ;
  assign n11998 = n10004 | n11997 ;
  assign n11999 = n10666 & ~n11998 ;
  assign n12000 = n3592 & ~n11999 ;
  assign n12001 = ~n6828 & n9012 ;
  assign n12002 = n10295 & n12001 ;
  assign n12003 = n4206 | n5450 ;
  assign n12004 = n1450 & ~n12003 ;
  assign n12005 = n4381 | n12004 ;
  assign n12006 = n6012 | n12005 ;
  assign n12007 = n2693 | n3848 ;
  assign n12008 = n6404 & ~n12007 ;
  assign n12012 = x168 & ~n1442 ;
  assign n12013 = ~n9273 & n12012 ;
  assign n12014 = n12013 ^ n10090 ^ x19 ;
  assign n12009 = x40 & ~n4277 ;
  assign n12010 = n8943 | n10211 ;
  assign n12011 = n12009 & ~n12010 ;
  assign n12015 = n12014 ^ n12011 ^ 1'b0 ;
  assign n12016 = n5930 ^ n2434 ^ 1'b0 ;
  assign n12017 = ~n2095 & n12016 ;
  assign n12018 = n6019 & ~n7716 ;
  assign n12019 = n9295 & n12018 ;
  assign n12020 = ~n10920 & n10950 ;
  assign n12021 = n4539 | n6560 ;
  assign n12022 = n12021 ^ n592 ^ 1'b0 ;
  assign n12023 = n9406 & ~n11231 ;
  assign n12024 = n12023 ^ n2741 ^ 1'b0 ;
  assign n12026 = n11850 ^ n509 ^ 1'b0 ;
  assign n12027 = n4619 & n12026 ;
  assign n12025 = n4286 & n11681 ;
  assign n12028 = n12027 ^ n12025 ^ 1'b0 ;
  assign n12029 = n1153 | n5201 ;
  assign n12030 = n705 & ~n2263 ;
  assign n12031 = n12030 ^ n5150 ^ 1'b0 ;
  assign n12032 = n8031 | n12031 ;
  assign n12033 = n6857 ^ n2939 ^ 1'b0 ;
  assign n12034 = n12032 | n12033 ;
  assign n12035 = ~n725 & n8186 ;
  assign n12036 = n12035 ^ n7867 ^ 1'b0 ;
  assign n12037 = n10685 ^ n8349 ^ 1'b0 ;
  assign n12038 = n12036 & n12037 ;
  assign n12039 = n466 | n10179 ;
  assign n12040 = n12039 ^ n11981 ^ 1'b0 ;
  assign n12041 = n9115 & n11911 ;
  assign n12043 = ~n552 & n4824 ;
  assign n12044 = n12043 ^ x178 ^ 1'b0 ;
  assign n12045 = n5416 ^ n3823 ^ 1'b0 ;
  assign n12046 = n12044 | n12045 ;
  assign n12047 = n12046 ^ n1064 ^ 1'b0 ;
  assign n12042 = n2407 & ~n4988 ;
  assign n12048 = n12047 ^ n12042 ^ 1'b0 ;
  assign n12049 = n1129 & n8996 ;
  assign n12050 = n5565 & n12049 ;
  assign n12051 = n3843 | n12050 ;
  assign n12052 = n12048 | n12051 ;
  assign n12053 = n9226 ^ n6950 ^ 1'b0 ;
  assign n12055 = n5707 ^ n509 ^ 1'b0 ;
  assign n12054 = n9262 ^ n564 ^ 1'b0 ;
  assign n12056 = n12055 ^ n12054 ^ 1'b0 ;
  assign n12057 = n1133 & n12056 ;
  assign n12058 = n3032 & n6453 ;
  assign n12059 = n9992 ^ n1251 ^ 1'b0 ;
  assign n12060 = ~n3178 & n4287 ;
  assign n12061 = n12060 ^ n2735 ^ 1'b0 ;
  assign n12062 = n12061 ^ n5988 ^ 1'b0 ;
  assign n12063 = x63 & n12062 ;
  assign n12065 = n4547 ^ n1708 ^ 1'b0 ;
  assign n12064 = n3985 & ~n4319 ;
  assign n12066 = n12065 ^ n12064 ^ 1'b0 ;
  assign n12067 = n12066 ^ n4084 ^ 1'b0 ;
  assign n12068 = ~n11809 & n12067 ;
  assign n12069 = n492 ^ x63 ^ 1'b0 ;
  assign n12070 = ~n2135 & n12069 ;
  assign n12071 = n12070 ^ n4799 ^ n2481 ;
  assign n12072 = n12071 ^ n5469 ^ n5420 ;
  assign n12073 = n7513 & ~n11536 ;
  assign n12074 = ~n12072 & n12073 ;
  assign n12075 = n12074 ^ n1799 ^ 1'b0 ;
  assign n12076 = n5626 ^ n2329 ^ 1'b0 ;
  assign n12077 = ~n4632 & n12076 ;
  assign n12078 = n3039 ^ n2740 ^ 1'b0 ;
  assign n12079 = n848 & ~n12078 ;
  assign n12080 = n9578 ^ n7502 ^ n5664 ;
  assign n12081 = n8140 ^ n3479 ^ 1'b0 ;
  assign n12082 = n12081 ^ n6336 ^ 1'b0 ;
  assign n12083 = x116 & ~n12082 ;
  assign n12084 = ~n2464 & n10219 ;
  assign n12085 = n12084 ^ n9725 ^ 1'b0 ;
  assign n12086 = ~n10877 & n12085 ;
  assign n12087 = ~n5364 & n12086 ;
  assign n12088 = ~n1874 & n4918 ;
  assign n12089 = n12088 ^ n6271 ^ 1'b0 ;
  assign n12090 = n2580 | n12089 ;
  assign n12091 = ~n2670 & n2942 ;
  assign n12092 = ~x190 & n12091 ;
  assign n12096 = n3021 & n3970 ;
  assign n12097 = ~n2801 & n12096 ;
  assign n12093 = n3889 & n5188 ;
  assign n12094 = ~n6624 & n12093 ;
  assign n12095 = n1985 & ~n12094 ;
  assign n12098 = n12097 ^ n12095 ^ 1'b0 ;
  assign n12099 = ~n12092 & n12098 ;
  assign n12100 = n711 | n11659 ;
  assign n12101 = n7731 ^ n6555 ^ n1477 ;
  assign n12102 = n12101 ^ n10608 ^ 1'b0 ;
  assign n12103 = n8459 ^ n2936 ^ 1'b0 ;
  assign n12104 = n1382 | n12103 ;
  assign n12105 = n12104 ^ n5625 ^ 1'b0 ;
  assign n12106 = ~n3673 & n11077 ;
  assign n12107 = n1509 | n5427 ;
  assign n12108 = n7163 ^ n4711 ^ 1'b0 ;
  assign n12109 = n12108 ^ n765 ^ 1'b0 ;
  assign n12110 = x40 & ~n485 ;
  assign n12111 = n12110 ^ n5082 ^ 1'b0 ;
  assign n12112 = n12111 ^ n8660 ^ 1'b0 ;
  assign n12113 = n2764 ^ n1259 ^ 1'b0 ;
  assign n12115 = ~n1404 & n4275 ;
  assign n12116 = ~n4949 & n12115 ;
  assign n12117 = n9078 ^ n7282 ^ 1'b0 ;
  assign n12118 = n12116 & ~n12117 ;
  assign n12114 = n1148 & ~n1874 ;
  assign n12119 = n12118 ^ n12114 ^ 1'b0 ;
  assign n12120 = ~n10306 & n11175 ;
  assign n12121 = n2182 & ~n3291 ;
  assign n12122 = n12121 ^ n4210 ^ 1'b0 ;
  assign n12123 = n12122 ^ n1030 ^ 1'b0 ;
  assign n12124 = n6033 ^ n1389 ^ 1'b0 ;
  assign n12125 = n12123 & n12124 ;
  assign n12126 = n12125 ^ n7932 ^ 1'b0 ;
  assign n12128 = ~n2122 & n4031 ;
  assign n12127 = ~n1844 & n2299 ;
  assign n12129 = n12128 ^ n12127 ^ 1'b0 ;
  assign n12130 = ~n535 & n3257 ;
  assign n12131 = n4275 & n12130 ;
  assign n12132 = n1419 | n10164 ;
  assign n12133 = n7164 & ~n12132 ;
  assign n12134 = n2317 & ~n9195 ;
  assign n12135 = n6169 | n8928 ;
  assign n12136 = n2331 | n12135 ;
  assign n12137 = n12136 ^ n2944 ^ 1'b0 ;
  assign n12138 = n12134 | n12137 ;
  assign n12139 = n2682 ^ x250 ^ 1'b0 ;
  assign n12140 = n9543 ^ n2752 ^ 1'b0 ;
  assign n12141 = n4447 ^ n329 ^ 1'b0 ;
  assign n12142 = n10211 | n12141 ;
  assign n12143 = n7939 ^ n4503 ^ n863 ;
  assign n12144 = n12143 ^ n7255 ^ 1'b0 ;
  assign n12145 = ~n12142 & n12144 ;
  assign n12146 = ~n5047 & n5307 ;
  assign n12147 = n11749 & n12146 ;
  assign n12148 = n12147 ^ n11193 ^ 1'b0 ;
  assign n12149 = n1848 & n4389 ;
  assign n12150 = ~x72 & n12149 ;
  assign n12151 = n12150 ^ n1856 ^ 1'b0 ;
  assign n12152 = n7141 & ~n12151 ;
  assign n12153 = n12152 ^ n5665 ^ n1098 ;
  assign n12154 = n10577 ^ n10216 ^ 1'b0 ;
  assign n12155 = n8147 | n12154 ;
  assign n12156 = n7925 & ~n8694 ;
  assign n12157 = ~n8862 & n12156 ;
  assign n12158 = n655 & ~n10957 ;
  assign n12159 = n12158 ^ x9 ^ 1'b0 ;
  assign n12160 = n4535 ^ n3011 ^ 1'b0 ;
  assign n12161 = ~n10901 & n12160 ;
  assign n12162 = ( n797 & n2330 ) | ( n797 & ~n2600 ) | ( n2330 & ~n2600 ) ;
  assign n12163 = n12162 ^ n4770 ^ n635 ;
  assign n12164 = n12163 ^ n996 ^ 1'b0 ;
  assign n12165 = n5052 | n12164 ;
  assign n12166 = ~n3307 & n9154 ;
  assign n12167 = ~n12165 & n12166 ;
  assign n12178 = n9458 ^ n938 ^ 1'b0 ;
  assign n12179 = n5384 & ~n12178 ;
  assign n12168 = n5379 ^ n3569 ^ n1568 ;
  assign n12169 = n2153 | n9362 ;
  assign n12170 = ~n3894 & n12169 ;
  assign n12171 = n4949 ^ n977 ^ 1'b0 ;
  assign n12172 = n8011 & n12171 ;
  assign n12173 = ~n4498 & n12172 ;
  assign n12174 = n12173 ^ n10827 ^ 1'b0 ;
  assign n12175 = n12170 & n12174 ;
  assign n12176 = n12175 ^ n2306 ^ 1'b0 ;
  assign n12177 = n12168 & n12176 ;
  assign n12180 = n12179 ^ n12177 ^ 1'b0 ;
  assign n12181 = ~n1430 & n5570 ;
  assign n12182 = n12181 ^ n4094 ^ 1'b0 ;
  assign n12183 = n5413 ^ n1500 ^ x246 ;
  assign n12184 = n8295 ^ n6564 ^ 1'b0 ;
  assign n12185 = n5387 | n12184 ;
  assign n12186 = n8917 | n12185 ;
  assign n12187 = n4607 ^ n4198 ^ n1766 ;
  assign n12188 = n6199 & n8658 ;
  assign n12189 = n12188 ^ n9172 ^ 1'b0 ;
  assign n12190 = n12187 & ~n12189 ;
  assign n12191 = n4230 ^ n3260 ^ n1453 ;
  assign n12192 = ~n4038 & n12191 ;
  assign n12193 = n1176 | n1935 ;
  assign n12194 = n8360 ^ n1589 ^ 1'b0 ;
  assign n12195 = n9878 & ~n12194 ;
  assign n12196 = n2167 & n12195 ;
  assign n12197 = ~x64 & n12196 ;
  assign n12198 = n6151 ^ n2001 ^ 1'b0 ;
  assign n12199 = ~n1364 & n12198 ;
  assign n12200 = n12199 ^ n7815 ^ 1'b0 ;
  assign n12201 = n8180 ^ n5959 ^ 1'b0 ;
  assign n12202 = n1286 | n4741 ;
  assign n12203 = n3622 & ~n12202 ;
  assign n12204 = n6481 & ~n12203 ;
  assign n12205 = n5452 ^ n3942 ^ 1'b0 ;
  assign n12206 = ~n5650 & n9746 ;
  assign n12207 = ~n3023 & n12206 ;
  assign n12208 = n8883 | n12207 ;
  assign n12209 = n12208 ^ n10354 ^ 1'b0 ;
  assign n12210 = n5310 | n12209 ;
  assign n12211 = n4966 & n5488 ;
  assign n12212 = ~n2935 & n12211 ;
  assign n12213 = x249 & ~n287 ;
  assign n12214 = ~x159 & n12213 ;
  assign n12215 = n943 & ~n7035 ;
  assign n12216 = ~n657 & n9487 ;
  assign n12217 = n12215 | n12216 ;
  assign n12218 = n4610 & ~n4795 ;
  assign n12219 = n3246 ^ n1489 ^ 1'b0 ;
  assign n12220 = n12218 | n12219 ;
  assign n12223 = n1220 & n2721 ;
  assign n12224 = n12223 ^ n518 ^ 1'b0 ;
  assign n12221 = n1154 & ~n4512 ;
  assign n12222 = n12221 ^ n2790 ^ 1'b0 ;
  assign n12225 = n12224 ^ n12222 ^ 1'b0 ;
  assign n12226 = n1004 & ~n5038 ;
  assign n12227 = n2957 | n12226 ;
  assign n12228 = n12227 ^ n11674 ^ 1'b0 ;
  assign n12229 = n8336 ^ n7796 ^ n4953 ;
  assign n12230 = n12229 ^ n3588 ^ 1'b0 ;
  assign n12231 = n12230 ^ n5344 ^ 1'b0 ;
  assign n12232 = n12231 ^ n7555 ^ 1'b0 ;
  assign n12233 = n6106 ^ n3419 ^ x21 ;
  assign n12234 = n12233 ^ n7944 ^ 1'b0 ;
  assign n12235 = n1182 & ~n3769 ;
  assign n12236 = n12235 ^ n6187 ^ 1'b0 ;
  assign n12237 = n3663 ^ n3573 ^ 1'b0 ;
  assign n12238 = n389 & ~n12237 ;
  assign n12239 = n8639 & n12238 ;
  assign n12240 = n12239 ^ n9778 ^ 1'b0 ;
  assign n12241 = n3508 ^ n3146 ^ n810 ;
  assign n12242 = n2530 & ~n7825 ;
  assign n12243 = ~n1051 & n12242 ;
  assign n12244 = n7247 & n12243 ;
  assign n12245 = n11557 | n12244 ;
  assign n12246 = n10789 ^ n5671 ^ 1'b0 ;
  assign n12247 = n6490 ^ n5958 ^ 1'b0 ;
  assign n12248 = n12247 ^ n1824 ^ 1'b0 ;
  assign n12249 = ~n2301 & n12248 ;
  assign n12250 = ( n5773 & n9465 ) | ( n5773 & ~n12249 ) | ( n9465 & ~n12249 ) ;
  assign n12251 = n7825 | n12250 ;
  assign n12252 = n12251 ^ n5529 ^ 1'b0 ;
  assign n12253 = ~n4940 & n12252 ;
  assign n12254 = n3233 | n5330 ;
  assign n12255 = n7070 ^ n395 ^ 1'b0 ;
  assign n12256 = ~n6639 & n12255 ;
  assign n12257 = ~n6363 & n7245 ;
  assign n12258 = n12257 ^ n7421 ^ 1'b0 ;
  assign n12259 = n12258 ^ n10445 ^ 1'b0 ;
  assign n12260 = ~n6707 & n9198 ;
  assign n12261 = ~n5619 & n9204 ;
  assign n12262 = n12260 & n12261 ;
  assign n12263 = n2951 ^ n2948 ^ n1114 ;
  assign n12264 = n12263 ^ n1885 ^ 1'b0 ;
  assign n12265 = n6329 ^ n1550 ^ 1'b0 ;
  assign n12266 = ~n12264 & n12265 ;
  assign n12267 = n3663 ^ n3557 ^ 1'b0 ;
  assign n12268 = n3326 ^ n2646 ^ 1'b0 ;
  assign n12269 = ( ~n2464 & n4765 ) | ( ~n2464 & n12268 ) | ( n4765 & n12268 ) ;
  assign n12270 = ~n3581 & n12269 ;
  assign n12271 = n12270 ^ n2256 ^ 1'b0 ;
  assign n12272 = n7674 ^ n384 ^ 1'b0 ;
  assign n12273 = n7202 & n12272 ;
  assign n12274 = ( n5366 & n5748 ) | ( n5366 & n12273 ) | ( n5748 & n12273 ) ;
  assign n12275 = ~n2383 & n4865 ;
  assign n12276 = n1599 & n3777 ;
  assign n12277 = ~n10110 & n12276 ;
  assign n12278 = ~n12275 & n12277 ;
  assign n12279 = ~n7707 & n9824 ;
  assign n12280 = ~n5887 & n12279 ;
  assign n12281 = ( n1366 & n2240 ) | ( n1366 & ~n6313 ) | ( n2240 & ~n6313 ) ;
  assign n12282 = n6611 & n12281 ;
  assign n12283 = ~n10361 & n12282 ;
  assign n12284 = n10653 ^ n2629 ^ 1'b0 ;
  assign n12285 = n1964 & ~n12284 ;
  assign n12286 = ~n830 & n12285 ;
  assign n12287 = n7821 & n12286 ;
  assign n12288 = n5276 ^ n908 ^ n270 ;
  assign n12289 = n2165 ^ n302 ^ 1'b0 ;
  assign n12290 = n3333 | n12289 ;
  assign n12291 = ~n3039 & n4580 ;
  assign n12292 = n11617 & n12291 ;
  assign n12293 = ~n2590 & n5592 ;
  assign n12294 = n5410 ^ n4547 ^ n3805 ;
  assign n12295 = n12293 & ~n12294 ;
  assign n12296 = n445 & n4986 ;
  assign n12297 = n12296 ^ n4290 ^ 1'b0 ;
  assign n12298 = n8133 & ~n11891 ;
  assign n12300 = n7602 ^ n6118 ^ 1'b0 ;
  assign n12299 = n2415 & ~n3316 ;
  assign n12301 = n12300 ^ n12299 ^ n11995 ;
  assign n12302 = n3572 & n7319 ;
  assign n12303 = ~n10426 & n12302 ;
  assign n12304 = n847 & n10390 ;
  assign n12305 = ~n5317 & n12304 ;
  assign n12306 = ~n12303 & n12305 ;
  assign n12307 = n6620 ^ n1853 ^ 1'b0 ;
  assign n12308 = ~n6352 & n12307 ;
  assign n12309 = n5539 ^ n4794 ^ 1'b0 ;
  assign n12310 = n7375 ^ n6393 ^ 1'b0 ;
  assign n12311 = n2659 | n6826 ;
  assign n12312 = n6696 | n12311 ;
  assign n12313 = n11229 ^ n587 ^ 1'b0 ;
  assign n12314 = n3657 | n12313 ;
  assign n12315 = n12314 ^ n1234 ^ 1'b0 ;
  assign n12316 = n9699 & ~n12315 ;
  assign n12317 = n2858 ^ n370 ^ 1'b0 ;
  assign n12318 = n2942 & ~n12317 ;
  assign n12319 = n12318 ^ n6077 ^ 1'b0 ;
  assign n12320 = n2448 & n4871 ;
  assign n12321 = n9250 & n12320 ;
  assign n12322 = n12321 ^ n5481 ^ 1'b0 ;
  assign n12323 = ~n11640 & n12322 ;
  assign n12324 = n4227 | n6749 ;
  assign n12325 = n6689 | n12324 ;
  assign n12326 = n12325 ^ n4521 ^ 1'b0 ;
  assign n12327 = n12326 ^ n2371 ^ 1'b0 ;
  assign n12328 = n1284 | n12327 ;
  assign n12329 = n2821 & n12328 ;
  assign n12330 = n7827 ^ n4578 ^ 1'b0 ;
  assign n12331 = n8994 & n12330 ;
  assign n12332 = ~n11234 & n12331 ;
  assign n12333 = n9130 ^ n2163 ^ 1'b0 ;
  assign n12334 = n2269 & ~n6123 ;
  assign n12335 = n12334 ^ n4813 ^ 1'b0 ;
  assign n12336 = n3116 ^ n1079 ^ 1'b0 ;
  assign n12337 = n6129 & ~n12336 ;
  assign n12338 = n2037 ^ n1887 ^ 1'b0 ;
  assign n12339 = n3074 | n4672 ;
  assign n12340 = n12339 ^ n2433 ^ 1'b0 ;
  assign n12341 = n10487 & n12340 ;
  assign n12342 = n12341 ^ n7518 ^ 1'b0 ;
  assign n12343 = n1799 ^ n1695 ^ 1'b0 ;
  assign n12344 = n3277 | n12343 ;
  assign n12345 = n12344 ^ n4031 ^ 1'b0 ;
  assign n12346 = ~n2229 & n12345 ;
  assign n12347 = n8819 ^ n1174 ^ 1'b0 ;
  assign n12348 = n10625 & n12347 ;
  assign n12349 = ~n4170 & n12348 ;
  assign n12350 = n3990 | n8446 ;
  assign n12351 = n11930 & ~n12350 ;
  assign n12352 = n12349 & n12351 ;
  assign n12353 = n4568 ^ n1756 ^ 1'b0 ;
  assign n12354 = ~n1185 & n12353 ;
  assign n12355 = n6524 ^ n2047 ^ 1'b0 ;
  assign n12356 = n6340 & ~n12355 ;
  assign n12357 = n8488 & ~n12356 ;
  assign n12358 = n2634 & n7912 ;
  assign n12359 = ~n4787 & n12358 ;
  assign n12360 = n11684 & ~n12359 ;
  assign n12361 = n12360 ^ n2332 ^ 1'b0 ;
  assign n12362 = n7804 ^ n1249 ^ 1'b0 ;
  assign n12363 = n5595 & n12362 ;
  assign n12364 = n11151 ^ n617 ^ 1'b0 ;
  assign n12365 = n3018 & n4335 ;
  assign n12366 = n2934 & n12365 ;
  assign n12367 = ( n6585 & n8799 ) | ( n6585 & ~n12366 ) | ( n8799 & ~n12366 ) ;
  assign n12368 = n12058 ^ n10698 ^ 1'b0 ;
  assign n12369 = n2332 & ~n12368 ;
  assign n12370 = n8806 ^ n1846 ^ 1'b0 ;
  assign n12371 = ~n3277 & n12370 ;
  assign n12372 = x231 & ~n5209 ;
  assign n12373 = n1833 & ~n10395 ;
  assign n12374 = n12373 ^ n10866 ^ 1'b0 ;
  assign n12375 = n5223 | n12374 ;
  assign n12376 = n916 & ~n8319 ;
  assign n12377 = n12376 ^ n3837 ^ 1'b0 ;
  assign n12378 = x149 & n12377 ;
  assign n12379 = n9093 & n12378 ;
  assign n12380 = n2008 & n4313 ;
  assign n12381 = n4010 & ~n12380 ;
  assign n12382 = n9262 & n12381 ;
  assign n12383 = ~n7295 & n12382 ;
  assign n12384 = n12383 ^ n2104 ^ 1'b0 ;
  assign n12385 = n1862 & ~n1925 ;
  assign n12386 = ~n4364 & n12385 ;
  assign n12387 = n4363 & n7853 ;
  assign n12388 = n8253 & n12387 ;
  assign n12389 = ~n1503 & n6311 ;
  assign n12390 = n12389 ^ n2560 ^ 1'b0 ;
  assign n12391 = ~n1200 & n12390 ;
  assign n12392 = ~n8164 & n12391 ;
  assign n12393 = ~n2984 & n12392 ;
  assign n12394 = n11007 ^ n6957 ^ 1'b0 ;
  assign n12395 = n4736 ^ n3869 ^ 1'b0 ;
  assign n12396 = ~n5353 & n8996 ;
  assign n12397 = ~n8066 & n12396 ;
  assign n12398 = n271 | n12215 ;
  assign n12399 = n2078 | n6146 ;
  assign n12400 = ( n2304 & ~n4876 ) | ( n2304 & n12399 ) | ( ~n4876 & n12399 ) ;
  assign n12408 = n4258 & ~n10998 ;
  assign n12409 = n12408 ^ n4514 ^ 1'b0 ;
  assign n12401 = n1319 & ~n1328 ;
  assign n12402 = ~n1319 & n12401 ;
  assign n12403 = n3478 | n12402 ;
  assign n12404 = n3478 & ~n12403 ;
  assign n12405 = n5408 | n12404 ;
  assign n12406 = n12404 & ~n12405 ;
  assign n12407 = n8418 & ~n12406 ;
  assign n12410 = n12409 ^ n12407 ^ 1'b0 ;
  assign n12411 = n825 ^ x150 ^ 1'b0 ;
  assign n12412 = ~n4867 & n12411 ;
  assign n12413 = x250 & n12412 ;
  assign n12414 = n6453 ^ n1977 ^ 1'b0 ;
  assign n12415 = ~n1085 & n12414 ;
  assign n12416 = n10775 & ~n12415 ;
  assign n12417 = n12416 ^ n4619 ^ 1'b0 ;
  assign n12418 = n1177 ^ n862 ^ n380 ;
  assign n12419 = n12418 ^ n1848 ^ n591 ;
  assign n12420 = n7059 ^ n5229 ^ 1'b0 ;
  assign n12421 = n12419 & ~n12420 ;
  assign n12422 = n1853 & ~n7456 ;
  assign n12423 = n3576 ^ n1200 ^ 1'b0 ;
  assign n12424 = n9216 & ~n12423 ;
  assign n12425 = n1416 ^ n1196 ^ 1'b0 ;
  assign n12426 = n2677 & n12425 ;
  assign n12427 = n12424 & ~n12426 ;
  assign n12428 = n12427 ^ n2062 ^ 1'b0 ;
  assign n12429 = n5936 & n8462 ;
  assign n12431 = ~n8347 & n8684 ;
  assign n12432 = n8347 & n12431 ;
  assign n12433 = n12432 ^ n5621 ^ 1'b0 ;
  assign n12430 = n9074 & n11367 ;
  assign n12434 = n12433 ^ n12430 ^ 1'b0 ;
  assign n12435 = n6189 & n12434 ;
  assign n12437 = n6532 ^ n6442 ^ 1'b0 ;
  assign n12438 = ~n4530 & n12437 ;
  assign n12436 = n4020 & n10937 ;
  assign n12439 = n12438 ^ n12436 ^ 1'b0 ;
  assign n12440 = n3749 | n8413 ;
  assign n12441 = n4347 | n12440 ;
  assign n12442 = ( n2468 & n2550 ) | ( n2468 & ~n6292 ) | ( n2550 & ~n6292 ) ;
  assign n12443 = n6119 | n12442 ;
  assign n12444 = n10664 & ~n12443 ;
  assign n12445 = n6518 ^ n6421 ^ 1'b0 ;
  assign n12446 = ~n267 & n1591 ;
  assign n12447 = ~n2668 & n12446 ;
  assign n12448 = n1065 | n4426 ;
  assign n12449 = n12266 ^ n9866 ^ 1'b0 ;
  assign n12450 = n5767 ^ n5596 ^ 1'b0 ;
  assign n12451 = n5827 & ~n10172 ;
  assign n12454 = n266 & ~n3393 ;
  assign n12455 = n12454 ^ n4876 ^ 1'b0 ;
  assign n12456 = n9076 & n12455 ;
  assign n12457 = n12456 ^ n2276 ^ 1'b0 ;
  assign n12458 = n3590 | n5745 ;
  assign n12459 = n12457 & ~n12458 ;
  assign n12460 = n9311 & n12459 ;
  assign n12452 = n1311 & ~n2741 ;
  assign n12453 = ~n6602 & n12452 ;
  assign n12461 = n12460 ^ n12453 ^ 1'b0 ;
  assign n12462 = ~n5769 & n8236 ;
  assign n12463 = n3144 ^ n1225 ^ 1'b0 ;
  assign n12464 = n11392 | n12463 ;
  assign n12465 = n10909 ^ n2349 ^ 1'b0 ;
  assign n12466 = ( x32 & n5119 ) | ( x32 & ~n7470 ) | ( n5119 & ~n7470 ) ;
  assign n12467 = n5855 ^ n2516 ^ 1'b0 ;
  assign n12468 = n3174 & ~n12467 ;
  assign n12469 = ( ~n7398 & n12466 ) | ( ~n7398 & n12468 ) | ( n12466 & n12468 ) ;
  assign n12470 = n7300 ^ n3845 ^ 1'b0 ;
  assign n12471 = ~n12469 & n12470 ;
  assign n12472 = x243 & ~n4998 ;
  assign n12473 = n12472 ^ n9239 ^ 1'b0 ;
  assign n12474 = n2999 ^ n1730 ^ 1'b0 ;
  assign n12475 = n5254 & n5660 ;
  assign n12476 = n12474 & n12475 ;
  assign n12477 = n6690 ^ n4391 ^ n1174 ;
  assign n12478 = n1589 & n3601 ;
  assign n12479 = ~n12477 & n12478 ;
  assign n12480 = n426 & ~n1917 ;
  assign n12481 = n1727 | n1992 ;
  assign n12482 = n12481 ^ n2301 ^ 1'b0 ;
  assign n12483 = ~n7600 & n12482 ;
  assign n12484 = n1508 & n12483 ;
  assign n12485 = n12484 ^ n3007 ^ 1'b0 ;
  assign n12486 = n12485 ^ n11201 ^ n913 ;
  assign n12487 = ~n12480 & n12486 ;
  assign n12488 = n12487 ^ n3753 ^ 1'b0 ;
  assign n12489 = n5022 ^ n4657 ^ 1'b0 ;
  assign n12490 = n10938 & n12489 ;
  assign n12491 = n2567 | n11196 ;
  assign n12492 = n12491 ^ n9340 ^ 1'b0 ;
  assign n12493 = ~n6276 & n12492 ;
  assign n12494 = n2500 & ~n10958 ;
  assign n12495 = ~n12493 & n12494 ;
  assign n12496 = n5243 & n5949 ;
  assign n12497 = n12496 ^ n3785 ^ 1'b0 ;
  assign n12498 = n7726 ^ n5333 ^ 1'b0 ;
  assign n12499 = n12497 & ~n12498 ;
  assign n12500 = ~n7274 & n12499 ;
  assign n12501 = ~n375 & n12500 ;
  assign n12502 = n9397 ^ n5315 ^ 1'b0 ;
  assign n12503 = n12501 & n12502 ;
  assign n12504 = ~n908 & n8079 ;
  assign n12505 = n12504 ^ n988 ^ 1'b0 ;
  assign n12506 = n665 | n1928 ;
  assign n12507 = n1118 | n12506 ;
  assign n12508 = n7909 & ~n12507 ;
  assign n12509 = ~n12505 & n12508 ;
  assign n12510 = n3825 & ~n7902 ;
  assign n12511 = n12510 ^ n10425 ^ 1'b0 ;
  assign n12512 = n2702 ^ n1487 ^ 1'b0 ;
  assign n12513 = n5484 & n12512 ;
  assign n12514 = ~n5859 & n12513 ;
  assign n12515 = n467 ^ x45 ^ 1'b0 ;
  assign n12516 = ~n4933 & n12515 ;
  assign n12517 = n12516 ^ n5186 ^ 1'b0 ;
  assign n12518 = n12517 ^ n11403 ^ 1'b0 ;
  assign n12519 = ~n2075 & n12518 ;
  assign n12520 = n12519 ^ x146 ^ 1'b0 ;
  assign n12521 = n4708 & n7567 ;
  assign n12522 = n12521 ^ n7285 ^ 1'b0 ;
  assign n12523 = ~n4441 & n4730 ;
  assign n12524 = n12523 ^ n2631 ^ 1'b0 ;
  assign n12525 = n12524 ^ n10053 ^ 1'b0 ;
  assign n12526 = ~n9734 & n12525 ;
  assign n12527 = ~n834 & n6979 ;
  assign n12528 = ~n2697 & n12527 ;
  assign n12529 = n1017 | n3076 ;
  assign n12530 = n10405 | n12529 ;
  assign n12531 = ~x99 & n4921 ;
  assign n12532 = ~n7110 & n10735 ;
  assign n12533 = n12532 ^ n9063 ^ 1'b0 ;
  assign n12534 = n8483 ^ n5831 ^ 1'b0 ;
  assign n12535 = n3944 ^ n2697 ^ 1'b0 ;
  assign n12536 = n10846 ^ n3397 ^ 1'b0 ;
  assign n12537 = ~n4934 & n12536 ;
  assign n12538 = n4824 ^ n3064 ^ 1'b0 ;
  assign n12539 = n513 & n4406 ;
  assign n12540 = n2506 | n7771 ;
  assign n12541 = n12539 & ~n12540 ;
  assign n12542 = n556 | n12541 ;
  assign n12543 = ~n12538 & n12542 ;
  assign n12544 = ~n4311 & n12543 ;
  assign n12547 = n2613 & n8668 ;
  assign n12545 = ~n3670 & n7504 ;
  assign n12546 = n12545 ^ n1318 ^ 1'b0 ;
  assign n12548 = n12547 ^ n12546 ^ n2513 ;
  assign n12549 = n1958 | n12548 ;
  assign n12550 = n12538 ^ n9710 ^ n8838 ;
  assign n12551 = ~n3690 & n7273 ;
  assign n12552 = n2439 & ~n12551 ;
  assign n12553 = n1032 & ~n2464 ;
  assign n12554 = ~n6414 & n7218 ;
  assign n12555 = n6452 & n6910 ;
  assign n12556 = n12555 ^ n6004 ^ 1'b0 ;
  assign n12557 = n11472 ^ n9824 ^ 1'b0 ;
  assign n12558 = n9615 & n12557 ;
  assign n12559 = n12556 & n12558 ;
  assign n12560 = n11680 ^ n3704 ^ 1'b0 ;
  assign n12561 = n3653 | n7904 ;
  assign n12562 = n9725 & ~n12561 ;
  assign n12563 = n1820 | n9953 ;
  assign n12564 = n12562 & ~n12563 ;
  assign n12565 = ( n6177 & n12560 ) | ( n6177 & ~n12564 ) | ( n12560 & ~n12564 ) ;
  assign n12566 = n4733 & n7418 ;
  assign n12567 = ~n3420 & n12566 ;
  assign n12568 = n1039 & n1245 ;
  assign n12569 = n12568 ^ n4050 ^ 1'b0 ;
  assign n12570 = n12569 ^ n3477 ^ 1'b0 ;
  assign n12571 = n4696 & ~n12570 ;
  assign n12572 = n11094 & n12571 ;
  assign n12573 = n12572 ^ n6786 ^ 1'b0 ;
  assign n12574 = n12573 ^ n9819 ^ 1'b0 ;
  assign n12575 = n4824 ^ n4251 ^ n2139 ;
  assign n12576 = n4565 & ~n12575 ;
  assign n12577 = n9614 ^ n4400 ^ 1'b0 ;
  assign n12578 = n12576 | n12577 ;
  assign n12579 = n3085 | n6086 ;
  assign n12580 = n7086 | n12579 ;
  assign n12581 = n451 | n535 ;
  assign n12582 = ( n2741 & n4239 ) | ( n2741 & ~n12581 ) | ( n4239 & ~n12581 ) ;
  assign n12583 = n4059 & n12582 ;
  assign n12584 = n2533 ^ n709 ^ 1'b0 ;
  assign n12585 = n5169 & ~n12584 ;
  assign n12586 = n3001 & ~n4747 ;
  assign n12587 = ~x162 & n9959 ;
  assign n12588 = n12587 ^ n2229 ^ 1'b0 ;
  assign n12589 = ~n4302 & n7495 ;
  assign n12590 = n12588 & n12589 ;
  assign n12591 = n1977 & n12590 ;
  assign n12592 = n2788 & ~n5206 ;
  assign n12593 = n9874 ^ n2589 ^ 1'b0 ;
  assign n12594 = n5905 | n12593 ;
  assign n12595 = n1971 | n12594 ;
  assign n12596 = n12595 ^ n2661 ^ n1880 ;
  assign n12597 = n2789 | n4039 ;
  assign n12598 = ( ~n1626 & n2051 ) | ( ~n1626 & n11544 ) | ( n2051 & n11544 ) ;
  assign n12599 = n12598 ^ n3114 ^ 1'b0 ;
  assign n12600 = ~n9266 & n12057 ;
  assign n12601 = n12600 ^ n8863 ^ 1'b0 ;
  assign n12604 = ( ~x253 & n862 ) | ( ~x253 & n2990 ) | ( n862 & n2990 ) ;
  assign n12602 = n7377 ^ n2613 ^ 1'b0 ;
  assign n12603 = x158 & n12602 ;
  assign n12605 = n12604 ^ n12603 ^ 1'b0 ;
  assign n12606 = n11504 & ~n12605 ;
  assign n12607 = n1276 & n12606 ;
  assign n12608 = n9091 ^ n7275 ^ n2529 ;
  assign n12609 = n7383 ^ n7183 ^ 1'b0 ;
  assign n12610 = n7184 ^ n3626 ^ 1'b0 ;
  assign n12611 = ~n7252 & n8935 ;
  assign n12612 = n7594 ^ n3022 ^ 1'b0 ;
  assign n12613 = n10584 ^ n2345 ^ 1'b0 ;
  assign n12614 = n12612 & n12613 ;
  assign n12615 = n6155 ^ n943 ^ 1'b0 ;
  assign n12616 = n842 & n12615 ;
  assign n12617 = n8572 & n12616 ;
  assign n12618 = n8524 & n8857 ;
  assign n12619 = ~n6131 & n12618 ;
  assign n12620 = n3628 ^ n564 ^ 1'b0 ;
  assign n12621 = n8000 & n12620 ;
  assign n12622 = n12621 ^ n3785 ^ n2394 ;
  assign n12623 = ~n5218 & n12465 ;
  assign n12624 = n7188 ^ n2596 ^ 1'b0 ;
  assign n12625 = x92 & ~n12624 ;
  assign n12626 = n8799 ^ n3898 ^ 1'b0 ;
  assign n12627 = n12625 & ~n12626 ;
  assign n12628 = n12627 ^ n2968 ^ 1'b0 ;
  assign n12629 = n6022 & n10529 ;
  assign n12630 = n12629 ^ n5570 ^ 1'b0 ;
  assign n12631 = n3670 & ~n12630 ;
  assign n12632 = n12231 ^ n10759 ^ 1'b0 ;
  assign n12633 = n12632 ^ n5410 ^ x3 ;
  assign n12634 = n8784 ^ n8663 ^ 1'b0 ;
  assign n12635 = n7492 & ~n11406 ;
  assign n12636 = n12635 ^ n3311 ^ 1'b0 ;
  assign n12638 = n5915 ^ n3011 ^ 1'b0 ;
  assign n12637 = n2369 & n9215 ;
  assign n12639 = n12638 ^ n12637 ^ 1'b0 ;
  assign n12640 = n540 & n8286 ;
  assign n12641 = ~x3 & n12640 ;
  assign n12645 = n1138 & ~n6961 ;
  assign n12646 = n12645 ^ n2401 ^ 1'b0 ;
  assign n12647 = x118 & ~n12646 ;
  assign n12643 = n5390 | n6559 ;
  assign n12644 = n3563 | n12643 ;
  assign n12648 = n12647 ^ n12644 ^ 1'b0 ;
  assign n12649 = n872 & n12648 ;
  assign n12650 = n3984 & ~n12649 ;
  assign n12642 = n1389 & n2282 ;
  assign n12651 = n12650 ^ n12642 ^ n4100 ;
  assign n12652 = n8300 ^ n497 ^ 1'b0 ;
  assign n12653 = n2076 & n12652 ;
  assign n12654 = n4588 ^ n2634 ^ 1'b0 ;
  assign n12655 = n12653 & ~n12654 ;
  assign n12656 = n5554 | n5837 ;
  assign n12657 = ~n2877 & n6959 ;
  assign n12658 = x188 & n12657 ;
  assign n12659 = n11119 & n12658 ;
  assign n12660 = ( ~n2585 & n2936 ) | ( ~n2585 & n6602 ) | ( n2936 & n6602 ) ;
  assign n12661 = ~n1480 & n5182 ;
  assign n12662 = n4335 ^ n3619 ^ 1'b0 ;
  assign n12663 = n1055 & n12662 ;
  assign n12666 = ( n3768 & ~n7132 ) | ( n3768 & n10206 ) | ( ~n7132 & n10206 ) ;
  assign n12664 = n6027 & ~n10479 ;
  assign n12665 = ( n1049 & n10068 ) | ( n1049 & ~n12664 ) | ( n10068 & ~n12664 ) ;
  assign n12667 = n12666 ^ n12665 ^ 1'b0 ;
  assign n12668 = ~n1613 & n5660 ;
  assign n12669 = n12668 ^ n1780 ^ 1'b0 ;
  assign n12672 = n5606 & n11983 ;
  assign n12670 = n9955 ^ n1351 ^ 1'b0 ;
  assign n12671 = n9161 | n12670 ;
  assign n12673 = n12672 ^ n12671 ^ 1'b0 ;
  assign n12674 = ( n2472 & ~n7697 ) | ( n2472 & n9256 ) | ( ~n7697 & n9256 ) ;
  assign n12675 = n2176 ^ n543 ^ 1'b0 ;
  assign n12676 = x101 & ~n12675 ;
  assign n12677 = n5421 & n12676 ;
  assign n12678 = ~n1712 & n3383 ;
  assign n12679 = n12678 ^ n4610 ^ 1'b0 ;
  assign n12680 = n4315 ^ n1294 ^ n518 ;
  assign n12681 = n12679 | n12680 ;
  assign n12682 = n3535 | n12681 ;
  assign n12683 = n12677 | n12682 ;
  assign n12684 = n12138 ^ n7371 ^ 1'b0 ;
  assign n12685 = ~n716 & n2735 ;
  assign n12686 = n12685 ^ n9955 ^ 1'b0 ;
  assign n12687 = ~n4361 & n6338 ;
  assign n12688 = n9448 ^ n2946 ^ 1'b0 ;
  assign n12689 = n12688 ^ n8177 ^ 1'b0 ;
  assign n12690 = n12079 | n12689 ;
  assign n12691 = n3346 ^ n1321 ^ 1'b0 ;
  assign n12692 = ~n2809 & n12691 ;
  assign n12695 = ~n3007 & n7015 ;
  assign n12696 = n3900 & n12695 ;
  assign n12693 = ~n1220 & n8781 ;
  assign n12694 = n1665 & n12693 ;
  assign n12697 = n12696 ^ n12694 ^ n3892 ;
  assign n12698 = n9788 ^ n4462 ^ 1'b0 ;
  assign n12699 = n12698 ^ n8276 ^ 1'b0 ;
  assign n12700 = ~n1923 & n3684 ;
  assign n12701 = n3039 ^ n2668 ^ 1'b0 ;
  assign n12702 = n12700 & ~n12701 ;
  assign n12703 = n6303 ^ n1088 ^ 1'b0 ;
  assign n12704 = n12702 & n12703 ;
  assign n12705 = ~n1159 & n11615 ;
  assign n12706 = n1990 ^ n854 ^ 1'b0 ;
  assign n12707 = n7689 ^ n6847 ^ 1'b0 ;
  assign n12708 = n8678 | n12707 ;
  assign n12709 = n10124 ^ n7075 ^ 1'b0 ;
  assign n12710 = n8545 & ~n12680 ;
  assign n12711 = n12710 ^ n9856 ^ 1'b0 ;
  assign n12712 = ~n4202 & n9429 ;
  assign n12713 = ( n951 & ~n3702 ) | ( n951 & n7323 ) | ( ~n3702 & n7323 ) ;
  assign n12714 = ( n436 & n6525 ) | ( n436 & ~n12713 ) | ( n6525 & ~n12713 ) ;
  assign n12715 = ~n3168 & n12714 ;
  assign n12716 = n2940 & n12715 ;
  assign n12717 = ~n5330 & n10932 ;
  assign n12718 = n3022 & n12717 ;
  assign n12719 = n1867 | n3077 ;
  assign n12720 = n12719 ^ n9564 ^ n367 ;
  assign n12721 = n9603 | n10949 ;
  assign n12722 = ( x110 & n4803 ) | ( x110 & ~n12721 ) | ( n4803 & ~n12721 ) ;
  assign n12723 = n11358 ^ n2141 ^ 1'b0 ;
  assign n12724 = x19 & ~n12723 ;
  assign n12725 = n6884 & n12724 ;
  assign n12726 = n8174 ^ n992 ^ 1'b0 ;
  assign n12727 = n4688 | n12726 ;
  assign n12728 = n8877 ^ n3202 ^ 1'b0 ;
  assign n12729 = n12727 | n12728 ;
  assign n12730 = n12729 ^ n12036 ^ 1'b0 ;
  assign n12731 = x162 & n4510 ;
  assign n12732 = n12731 ^ n6561 ^ 1'b0 ;
  assign n12733 = ~n8945 & n9099 ;
  assign n12734 = n4779 ^ n4465 ^ 1'b0 ;
  assign n12735 = n12734 ^ n12597 ^ 1'b0 ;
  assign n12736 = n317 | n12735 ;
  assign n12737 = n2426 & ~n3034 ;
  assign n12738 = n8434 ^ n7850 ^ 1'b0 ;
  assign n12739 = n12738 ^ n716 ^ 1'b0 ;
  assign n12740 = n12737 & n12739 ;
  assign n12741 = n12740 ^ n1079 ^ 1'b0 ;
  assign n12742 = n5823 | n9549 ;
  assign n12743 = n9496 | n12064 ;
  assign n12744 = n12743 ^ n847 ^ 1'b0 ;
  assign n12745 = n9582 ^ n7387 ^ 1'b0 ;
  assign n12746 = n3396 ^ n3193 ^ n264 ;
  assign n12747 = ~n5492 & n12746 ;
  assign n12748 = n12747 ^ n6229 ^ 1'b0 ;
  assign n12749 = n12748 ^ n10368 ^ 1'b0 ;
  assign n12750 = n12323 & n12749 ;
  assign n12751 = n12564 & n12750 ;
  assign n12752 = n8315 & ~n10350 ;
  assign n12753 = n365 | n9049 ;
  assign n12754 = n12753 ^ n1125 ^ 1'b0 ;
  assign n12755 = ~n7644 & n12754 ;
  assign n12756 = n12755 ^ n2724 ^ 1'b0 ;
  assign n12757 = n6113 & n12756 ;
  assign n12758 = n12757 ^ n6879 ^ 1'b0 ;
  assign n12759 = n7831 ^ x165 ^ 1'b0 ;
  assign n12760 = n9368 & n12759 ;
  assign n12761 = n12245 ^ n3620 ^ 1'b0 ;
  assign n12762 = n12760 & ~n12761 ;
  assign n12763 = ~n4605 & n8401 ;
  assign n12764 = ( ~n420 & n2674 ) | ( ~n420 & n12763 ) | ( n2674 & n12763 ) ;
  assign n12765 = ( ~x148 & n1689 ) | ( ~x148 & n2672 ) | ( n1689 & n2672 ) ;
  assign n12766 = n1186 | n12765 ;
  assign n12767 = n12065 ^ n6452 ^ 1'b0 ;
  assign n12768 = n12767 ^ n7933 ^ 1'b0 ;
  assign n12769 = n12766 & n12768 ;
  assign n12770 = n10354 ^ n4515 ^ n3012 ;
  assign n12771 = n12770 ^ n11649 ^ 1'b0 ;
  assign n12772 = n10410 | n12581 ;
  assign n12773 = n12771 | n12772 ;
  assign n12774 = n970 & ~n10031 ;
  assign n12775 = n560 & n12774 ;
  assign n12777 = n11838 ^ n1223 ^ 1'b0 ;
  assign n12776 = n3546 & ~n6481 ;
  assign n12778 = n12777 ^ n12776 ^ 1'b0 ;
  assign n12779 = x24 & ~n655 ;
  assign n12780 = ~n9526 & n12779 ;
  assign n12781 = n12780 ^ n909 ^ 1'b0 ;
  assign n12782 = ~n9041 & n10540 ;
  assign n12783 = ( n767 & n7025 ) | ( n767 & n9722 ) | ( n7025 & n9722 ) ;
  assign n12784 = n6242 & ~n7173 ;
  assign n12785 = n12784 ^ n8591 ^ 1'b0 ;
  assign n12786 = n757 & ~n12785 ;
  assign n12787 = ~n7289 & n9816 ;
  assign n12788 = n11360 ^ n1137 ^ 1'b0 ;
  assign n12789 = ~n7806 & n12788 ;
  assign n12790 = ~n12217 & n12789 ;
  assign n12791 = ~n12787 & n12790 ;
  assign n12792 = n488 | n550 ;
  assign n12793 = ( n7242 & ~n7601 ) | ( n7242 & n12792 ) | ( ~n7601 & n12792 ) ;
  assign n12794 = ( n4037 & n4878 ) | ( n4037 & ~n8184 ) | ( n4878 & ~n8184 ) ;
  assign n12795 = n12794 ^ n2911 ^ 1'b0 ;
  assign n12796 = n12795 ^ n2409 ^ 1'b0 ;
  assign n12797 = n3042 | n12796 ;
  assign n12798 = x221 & ~n9350 ;
  assign n12799 = n12798 ^ n1997 ^ 1'b0 ;
  assign n12800 = n3543 & n12799 ;
  assign n12801 = n1311 & ~n4292 ;
  assign n12802 = n1554 & n12801 ;
  assign n12803 = n6060 | n12802 ;
  assign n12804 = n12803 ^ n6797 ^ 1'b0 ;
  assign n12805 = n2216 | n2743 ;
  assign n12806 = n12805 ^ n3193 ^ 1'b0 ;
  assign n12807 = n12528 ^ n11344 ^ 1'b0 ;
  assign n12808 = n7444 ^ n7251 ^ 1'b0 ;
  assign n12809 = n5324 & ~n12808 ;
  assign n12810 = n7173 | n12809 ;
  assign n12811 = x239 ^ x184 ^ 1'b0 ;
  assign n12812 = ~n780 & n12811 ;
  assign n12813 = n12812 ^ n4280 ^ 1'b0 ;
  assign n12815 = n5690 ^ n5554 ^ 1'b0 ;
  assign n12816 = n1556 | n12815 ;
  assign n12817 = n12816 ^ n1315 ^ 1'b0 ;
  assign n12814 = ~n8422 & n9709 ;
  assign n12818 = n12817 ^ n12814 ^ 1'b0 ;
  assign n12819 = ( ~n2789 & n3571 ) | ( ~n2789 & n9792 ) | ( n3571 & n9792 ) ;
  assign n12820 = ~n2715 & n12819 ;
  assign n12821 = n7083 & n10770 ;
  assign n12822 = n12821 ^ n1112 ^ 1'b0 ;
  assign n12828 = n946 & ~n3517 ;
  assign n12829 = ~n3490 & n12828 ;
  assign n12830 = n7257 & n12829 ;
  assign n12823 = ~n2272 & n7508 ;
  assign n12824 = ~n289 & n12823 ;
  assign n12825 = n5767 & ~n12824 ;
  assign n12826 = ~n10501 & n12825 ;
  assign n12827 = n7031 & ~n12826 ;
  assign n12831 = n12830 ^ n12827 ^ 1'b0 ;
  assign n12832 = ( n3291 & ~n9164 ) | ( n3291 & n9798 ) | ( ~n9164 & n9798 ) ;
  assign n12833 = ( n1931 & n7738 ) | ( n1931 & ~n7814 ) | ( n7738 & ~n7814 ) ;
  assign n12834 = n4937 & ~n6419 ;
  assign n12835 = n11406 & n12834 ;
  assign n12836 = ( ~n1346 & n2679 ) | ( ~n1346 & n12835 ) | ( n2679 & n12835 ) ;
  assign n12841 = n9693 ^ n7351 ^ n6269 ;
  assign n12837 = n4273 ^ n2390 ^ 1'b0 ;
  assign n12838 = n12837 ^ n4791 ^ 1'b0 ;
  assign n12839 = n10139 & n12838 ;
  assign n12840 = ~n9856 & n12839 ;
  assign n12842 = n12841 ^ n12840 ^ 1'b0 ;
  assign n12844 = n449 & ~n2357 ;
  assign n12845 = n4659 & n12844 ;
  assign n12843 = n6256 ^ n5408 ^ n4869 ;
  assign n12846 = n12845 ^ n12843 ^ n10267 ;
  assign n12847 = ~n2506 & n6978 ;
  assign n12848 = ~n6404 & n12847 ;
  assign n12849 = x34 & ~n12848 ;
  assign n12850 = n11583 & n12849 ;
  assign n12851 = n5732 ^ n2155 ^ 1'b0 ;
  assign n12852 = n3258 & ~n12851 ;
  assign n12853 = n12852 ^ n3281 ^ n1917 ;
  assign n12854 = ~n906 & n4315 ;
  assign n12855 = n7411 ^ n4175 ^ 1'b0 ;
  assign n12856 = n1156 & n9207 ;
  assign n12857 = n9844 ^ n7560 ^ 1'b0 ;
  assign n12858 = n12857 ^ n3904 ^ 1'b0 ;
  assign n12859 = n12856 | n12858 ;
  assign n12860 = n5316 ^ n1667 ^ 1'b0 ;
  assign n12861 = n970 | n12860 ;
  assign n12862 = n7783 & n12861 ;
  assign n12863 = n8196 ^ n2964 ^ 1'b0 ;
  assign n12864 = n11302 ^ n792 ^ 1'b0 ;
  assign n12865 = ~n810 & n6121 ;
  assign n12866 = n12864 & n12865 ;
  assign n12867 = n697 & n12866 ;
  assign n12870 = n9958 & ~n10394 ;
  assign n12869 = n3604 & n7162 ;
  assign n12871 = n12870 ^ n12869 ^ n4042 ;
  assign n12868 = ~n5452 & n7808 ;
  assign n12872 = n12871 ^ n12868 ^ 1'b0 ;
  assign n12874 = ( n1249 & n2016 ) | ( n1249 & ~n3831 ) | ( n2016 & ~n3831 ) ;
  assign n12873 = ~n7934 & n9526 ;
  assign n12875 = n12874 ^ n12873 ^ n1786 ;
  assign n12876 = n1720 | n5540 ;
  assign n12877 = x189 & ~n12876 ;
  assign n12878 = ( ~n3749 & n12551 ) | ( ~n3749 & n12877 ) | ( n12551 & n12877 ) ;
  assign n12879 = n10709 ^ n8366 ^ 1'b0 ;
  assign n12880 = n11605 ^ n6030 ^ 1'b0 ;
  assign n12881 = n12880 ^ n11917 ^ 1'b0 ;
  assign n12882 = n10180 & ~n12881 ;
  assign n12883 = n5438 & n12335 ;
  assign n12884 = ~n4754 & n12883 ;
  assign n12885 = n5786 ^ n3661 ^ 1'b0 ;
  assign n12886 = ~n8198 & n8845 ;
  assign n12887 = n12886 ^ x158 ^ 1'b0 ;
  assign n12888 = n5135 & ~n12887 ;
  assign n12889 = n12888 ^ n12721 ^ 1'b0 ;
  assign n12890 = ~n7022 & n12889 ;
  assign n12891 = n10283 ^ n1789 ^ 1'b0 ;
  assign n12892 = ( n4710 & n8198 ) | ( n4710 & ~n12891 ) | ( n8198 & ~n12891 ) ;
  assign n12895 = n3263 & ~n4204 ;
  assign n12896 = n12895 ^ n1765 ^ 1'b0 ;
  assign n12893 = n10639 ^ x113 ^ 1'b0 ;
  assign n12894 = n6934 | n12893 ;
  assign n12897 = n12896 ^ n12894 ^ 1'b0 ;
  assign n12898 = n1545 | n9853 ;
  assign n12902 = n5115 ^ n2158 ^ n817 ;
  assign n12903 = n9721 & ~n12902 ;
  assign n12899 = x225 & n10385 ;
  assign n12900 = n12899 ^ n8070 ^ 1'b0 ;
  assign n12901 = n2469 | n12900 ;
  assign n12904 = n12903 ^ n12901 ^ n4303 ;
  assign n12905 = n416 & ~n9470 ;
  assign n12906 = n8097 | n12905 ;
  assign n12907 = n10763 & ~n12906 ;
  assign n12908 = ~n2082 & n12300 ;
  assign n12909 = n12681 & n12908 ;
  assign n12910 = n12909 ^ n12605 ^ 1'b0 ;
  assign n12911 = ~n12907 & n12910 ;
  assign n12912 = x178 | n5315 ;
  assign n12913 = n12912 ^ n12386 ^ 1'b0 ;
  assign n12917 = n2582 & ~n9611 ;
  assign n12918 = ~n6819 & n12917 ;
  assign n12914 = n8182 ^ n7267 ^ 1'b0 ;
  assign n12915 = n5016 & n12914 ;
  assign n12916 = n8424 & n12915 ;
  assign n12919 = n12918 ^ n12916 ^ 1'b0 ;
  assign n12920 = n3105 | n6219 ;
  assign n12921 = n12920 ^ n3271 ^ 1'b0 ;
  assign n12922 = n12921 ^ n9703 ^ 1'b0 ;
  assign n12923 = ~n666 & n2964 ;
  assign n12924 = n6916 & n7704 ;
  assign n12925 = x131 & ~n996 ;
  assign n12926 = ~n1377 & n12925 ;
  assign n12927 = n10150 & ~n12926 ;
  assign n12928 = n927 & n12927 ;
  assign n12929 = n11178 & ~n11963 ;
  assign n12930 = n4595 ^ n872 ^ 1'b0 ;
  assign n12931 = n1956 & ~n12930 ;
  assign n12932 = n12931 ^ n11759 ^ 1'b0 ;
  assign n12933 = n12377 & ~n12932 ;
  assign n12937 = n2139 & ~n2788 ;
  assign n12934 = n8730 ^ n6008 ^ 1'b0 ;
  assign n12935 = n1342 | n12934 ;
  assign n12936 = ~n3291 & n12935 ;
  assign n12938 = n12937 ^ n12936 ^ 1'b0 ;
  assign n12939 = n2620 & ~n3302 ;
  assign n12940 = n6236 | n12939 ;
  assign n12941 = n5720 | n12940 ;
  assign n12942 = n10765 | n12941 ;
  assign n12943 = n10361 ^ n1504 ^ 1'b0 ;
  assign n12944 = ~n6023 & n8970 ;
  assign n12945 = n12943 | n12944 ;
  assign n12946 = n6017 | n8874 ;
  assign n12947 = n1828 | n12946 ;
  assign n12950 = n2472 ^ x119 ^ 1'b0 ;
  assign n12951 = n8281 & ~n12950 ;
  assign n12948 = n1591 & ~n2884 ;
  assign n12949 = ~n9916 & n12948 ;
  assign n12952 = n12951 ^ n12949 ^ 1'b0 ;
  assign n12962 = n7361 | n10187 ;
  assign n12963 = n12058 & ~n12962 ;
  assign n12953 = n2433 ^ n296 ^ 1'b0 ;
  assign n12954 = n1125 | n12953 ;
  assign n12955 = n12954 ^ n825 ^ 1'b0 ;
  assign n12957 = n1822 & n1880 ;
  assign n12958 = ~n5003 & n12957 ;
  assign n12959 = n7467 & n12958 ;
  assign n12956 = n5879 ^ n1069 ^ 1'b0 ;
  assign n12960 = n12959 ^ n12956 ^ 1'b0 ;
  assign n12961 = n12955 | n12960 ;
  assign n12964 = n12963 ^ n12961 ^ 1'b0 ;
  assign n12965 = n3508 & ~n12964 ;
  assign n12966 = n8744 & n12965 ;
  assign n12967 = n8583 ^ n4402 ^ n3527 ;
  assign n12968 = n3474 ^ n642 ^ 1'b0 ;
  assign n12969 = n1213 & n12968 ;
  assign n12970 = n12969 ^ n2900 ^ 1'b0 ;
  assign n12971 = n1878 & n10523 ;
  assign n12972 = n4608 ^ n1340 ^ 1'b0 ;
  assign n12973 = n12972 ^ n1430 ^ 1'b0 ;
  assign n12974 = n12971 & n12973 ;
  assign n12975 = n12342 ^ n8724 ^ 1'b0 ;
  assign n12976 = n5210 ^ n828 ^ 1'b0 ;
  assign n12977 = ~n5099 & n12976 ;
  assign n12978 = ( ~n3258 & n8454 ) | ( ~n3258 & n10014 ) | ( n8454 & n10014 ) ;
  assign n12979 = n12978 ^ n2622 ^ 1'b0 ;
  assign n12980 = ( ~n11124 & n12977 ) | ( ~n11124 & n12979 ) | ( n12977 & n12979 ) ;
  assign n12981 = n4374 | n7923 ;
  assign n12982 = n8330 ^ n1453 ^ 1'b0 ;
  assign n12983 = n7587 & ~n12982 ;
  assign n12984 = n1871 & n7757 ;
  assign n12985 = n7432 ^ n5231 ^ 1'b0 ;
  assign n12986 = ~n2062 & n2128 ;
  assign n12987 = ~n12985 & n12986 ;
  assign n12988 = n4739 ^ n2408 ^ 1'b0 ;
  assign n12989 = n1293 & ~n12988 ;
  assign n12990 = n12989 ^ n4595 ^ 1'b0 ;
  assign n12991 = ~n12987 & n12990 ;
  assign n12992 = n4345 | n4379 ;
  assign n12993 = n12992 ^ n6751 ^ 1'b0 ;
  assign n12994 = ~n1766 & n12993 ;
  assign n12995 = n12994 ^ n4920 ^ n2785 ;
  assign n12996 = n7093 ^ n4839 ^ x252 ;
  assign n12997 = n8210 & n10390 ;
  assign n12998 = ~n8573 & n12997 ;
  assign n13003 = n433 & n1770 ;
  assign n13004 = x253 & n13003 ;
  assign n12999 = n3633 ^ n389 ^ 1'b0 ;
  assign n13000 = ~n6211 & n12999 ;
  assign n13001 = n13000 ^ n4308 ^ 1'b0 ;
  assign n13002 = n6621 & n13001 ;
  assign n13005 = n13004 ^ n13002 ^ 1'b0 ;
  assign n13006 = n2219 | n12646 ;
  assign n13007 = n13006 ^ n6072 ^ 1'b0 ;
  assign n13008 = n453 & ~n13007 ;
  assign n13009 = n663 & ~n3712 ;
  assign n13010 = n3712 & n13009 ;
  assign n13012 = n10857 ^ n1439 ^ 1'b0 ;
  assign n13013 = ~n3133 & n13012 ;
  assign n13014 = n13013 ^ n562 ^ 1'b0 ;
  assign n13011 = n8042 ^ n3843 ^ 1'b0 ;
  assign n13015 = n13014 ^ n13011 ^ 1'b0 ;
  assign n13016 = n12331 & ~n13015 ;
  assign n13017 = ( n9527 & n13010 ) | ( n9527 & ~n13016 ) | ( n13010 & ~n13016 ) ;
  assign n13018 = n11040 & n11939 ;
  assign n13019 = n1628 | n5500 ;
  assign n13020 = n9264 ^ n6273 ^ 1'b0 ;
  assign n13021 = n267 | n13020 ;
  assign n13022 = n9063 | n13021 ;
  assign n13023 = n7314 ^ n5315 ^ 1'b0 ;
  assign n13024 = x159 | n2065 ;
  assign n13025 = n5014 & ~n13024 ;
  assign n13026 = n11178 & ~n13025 ;
  assign n13027 = n13023 | n13026 ;
  assign n13028 = n3722 ^ n2589 ^ x236 ;
  assign n13029 = n13028 ^ n2014 ^ 1'b0 ;
  assign n13030 = ~n8517 & n13029 ;
  assign n13031 = ( ~n1694 & n7809 ) | ( ~n1694 & n13030 ) | ( n7809 & n13030 ) ;
  assign n13032 = n11578 ^ n5919 ^ 1'b0 ;
  assign n13033 = n13031 & ~n13032 ;
  assign n13034 = n13033 ^ n3731 ^ 1'b0 ;
  assign n13035 = x51 & ~n9936 ;
  assign n13036 = n1172 | n2277 ;
  assign n13037 = n13036 ^ n7724 ^ 1'b0 ;
  assign n13038 = n3086 | n13037 ;
  assign n13039 = n1254 & ~n7814 ;
  assign n13040 = n5538 ^ n4718 ^ 1'b0 ;
  assign n13041 = ~n7617 & n13040 ;
  assign n13042 = n8109 ^ n7099 ^ 1'b0 ;
  assign n13043 = n10368 ^ n1523 ^ 1'b0 ;
  assign n13044 = ~n12476 & n13043 ;
  assign n13046 = n451 & n3871 ;
  assign n13047 = n6253 & n13046 ;
  assign n13045 = n5315 & ~n12795 ;
  assign n13048 = n13047 ^ n13045 ^ 1'b0 ;
  assign n13049 = n6159 ^ n2099 ^ 1'b0 ;
  assign n13050 = n10781 | n13049 ;
  assign n13051 = n11668 | n13050 ;
  assign n13052 = n13051 ^ n11243 ^ 1'b0 ;
  assign n13053 = n1244 | n13052 ;
  assign n13054 = ( ~n2268 & n6680 ) | ( ~n2268 & n8917 ) | ( n6680 & n8917 ) ;
  assign n13055 = n13054 ^ n3961 ^ 1'b0 ;
  assign n13056 = n3626 ^ n2557 ^ 1'b0 ;
  assign n13057 = ~n8025 & n13056 ;
  assign n13058 = ~x133 & n4472 ;
  assign n13059 = x175 & ~n13058 ;
  assign n13060 = n13059 ^ n12022 ^ 1'b0 ;
  assign n13061 = n5924 ^ n3826 ^ 1'b0 ;
  assign n13062 = n13061 ^ n11511 ^ 1'b0 ;
  assign n13063 = n4389 & ~n13062 ;
  assign n13064 = n1093 & n6781 ;
  assign n13065 = n2365 | n9551 ;
  assign n13066 = n7827 ^ n2685 ^ 1'b0 ;
  assign n13067 = x181 & n3685 ;
  assign n13068 = n13067 ^ n1001 ^ 1'b0 ;
  assign n13069 = n7160 & n13068 ;
  assign n13070 = ~n13066 & n13069 ;
  assign n13072 = n1839 & n9930 ;
  assign n13073 = ~n3371 & n13072 ;
  assign n13071 = ( x152 & n1053 ) | ( x152 & ~n2223 ) | ( n1053 & ~n2223 ) ;
  assign n13074 = n13073 ^ n13071 ^ 1'b0 ;
  assign n13075 = n5732 | n13074 ;
  assign n13076 = n421 & ~n3165 ;
  assign n13077 = n13076 ^ n944 ^ 1'b0 ;
  assign n13078 = n2378 & ~n13077 ;
  assign n13079 = x71 & n12353 ;
  assign n13080 = n13078 | n13079 ;
  assign n13081 = n12158 ^ n6218 ^ 1'b0 ;
  assign n13082 = n518 & n13081 ;
  assign n13083 = n12668 ^ n6533 ^ 1'b0 ;
  assign n13084 = n2668 & n4806 ;
  assign n13085 = n13084 ^ n779 ^ x76 ;
  assign n13086 = n6734 ^ n3025 ^ 1'b0 ;
  assign n13087 = n2307 & n13086 ;
  assign n13088 = n2988 & n13087 ;
  assign n13089 = n1416 | n8980 ;
  assign n13090 = ( n2231 & ~n6595 ) | ( n2231 & n8591 ) | ( ~n6595 & n8591 ) ;
  assign n13091 = n1535 & ~n2234 ;
  assign n13092 = n13091 ^ n3534 ^ 1'b0 ;
  assign n13093 = n11694 | n13092 ;
  assign n13094 = n2714 ^ n2433 ^ 1'b0 ;
  assign n13095 = ~n13093 & n13094 ;
  assign n13096 = ~n4910 & n13095 ;
  assign n13097 = ~n838 & n9816 ;
  assign n13098 = n2714 | n7864 ;
  assign n13099 = n13098 ^ n647 ^ 1'b0 ;
  assign n13100 = n2305 & ~n13099 ;
  assign n13101 = n1288 | n12612 ;
  assign n13102 = n13101 ^ n4959 ^ n4522 ;
  assign n13103 = ~n7518 & n13102 ;
  assign n13104 = ~n4932 & n13103 ;
  assign n13105 = n4840 | n11336 ;
  assign n13106 = n13105 ^ n11609 ^ 1'b0 ;
  assign n13107 = n8943 ^ n5879 ^ n1581 ;
  assign n13108 = x20 & ~x22 ;
  assign n13109 = n8104 | n8874 ;
  assign n13110 = n13109 ^ n3113 ^ 1'b0 ;
  assign n13111 = n1397 & ~n13110 ;
  assign n13112 = n8781 ^ n3461 ^ 1'b0 ;
  assign n13113 = n10837 | n13112 ;
  assign n13114 = n7107 & n13113 ;
  assign n13115 = n325 & ~n7271 ;
  assign n13116 = ~n5749 & n13115 ;
  assign n13117 = n6611 ^ n4091 ^ 1'b0 ;
  assign n13118 = n10272 | n13117 ;
  assign n13119 = n6582 ^ n5111 ^ 1'b0 ;
  assign n13120 = n9032 & ~n11485 ;
  assign n13121 = n13120 ^ n10356 ^ 1'b0 ;
  assign n13122 = n13121 ^ n1893 ^ 1'b0 ;
  assign n13123 = n10541 ^ n3496 ^ 1'b0 ;
  assign n13124 = ~n3186 & n13123 ;
  assign n13125 = ( n3115 & n7736 ) | ( n3115 & ~n13087 ) | ( n7736 & ~n13087 ) ;
  assign n13126 = n13125 ^ x227 ^ 1'b0 ;
  assign n13127 = ( n2715 & n7164 ) | ( n2715 & n13126 ) | ( n7164 & n13126 ) ;
  assign n13128 = n13127 ^ n7170 ^ 1'b0 ;
  assign n13129 = ~n813 & n13128 ;
  assign n13130 = n8000 & n13129 ;
  assign n13131 = ~n13124 & n13130 ;
  assign n13132 = n4449 & n9643 ;
  assign n13133 = n4940 & n13132 ;
  assign n13135 = n4059 & ~n8495 ;
  assign n13134 = n6301 | n7107 ;
  assign n13136 = n13135 ^ n13134 ^ 1'b0 ;
  assign n13137 = n2067 & ~n5798 ;
  assign n13138 = n3140 & n13137 ;
  assign n13139 = n7199 ^ n3355 ^ n815 ;
  assign n13140 = n4938 & n13139 ;
  assign n13141 = n13138 & n13140 ;
  assign n13142 = n3364 & n7968 ;
  assign n13143 = x203 | n8028 ;
  assign n13148 = n9260 ^ n5544 ^ 1'b0 ;
  assign n13149 = n3989 & n13148 ;
  assign n13144 = ~n571 & n7252 ;
  assign n13145 = n13144 ^ n10743 ^ 1'b0 ;
  assign n13146 = n889 | n13145 ;
  assign n13147 = n4562 & ~n13146 ;
  assign n13150 = n13149 ^ n13147 ^ 1'b0 ;
  assign n13151 = n13143 & n13150 ;
  assign n13152 = n13142 | n13151 ;
  assign n13153 = ~n3990 & n4686 ;
  assign n13154 = n13153 ^ n763 ^ 1'b0 ;
  assign n13155 = n13154 ^ n6514 ^ 1'b0 ;
  assign n13156 = n271 & n9026 ;
  assign n13157 = n2131 & n13156 ;
  assign n13158 = ( n7629 & n9516 ) | ( n7629 & ~n12173 ) | ( n9516 & ~n12173 ) ;
  assign n13159 = n13158 ^ n6284 ^ 1'b0 ;
  assign n13160 = n13157 | n13159 ;
  assign n13161 = n13160 ^ n1020 ^ 1'b0 ;
  assign n13162 = n13155 & ~n13161 ;
  assign n13163 = n5958 ^ n4642 ^ n1606 ;
  assign n13164 = x162 & ~n8495 ;
  assign n13165 = n13164 ^ n7066 ^ 1'b0 ;
  assign n13166 = n12890 ^ n8864 ^ 1'b0 ;
  assign n13167 = n9917 | n13166 ;
  assign n13168 = n4535 & ~n10424 ;
  assign n13169 = ~n6512 & n6616 ;
  assign n13170 = n13169 ^ n2813 ^ 1'b0 ;
  assign n13171 = ~n1593 & n10412 ;
  assign n13172 = n4434 & n10175 ;
  assign n13174 = n553 & n6824 ;
  assign n13175 = n13174 ^ n4730 ^ 1'b0 ;
  assign n13176 = n13175 ^ n510 ^ 1'b0 ;
  assign n13173 = ( n2569 & n3906 ) | ( n2569 & ~n5565 ) | ( n3906 & ~n5565 ) ;
  assign n13177 = n13176 ^ n13173 ^ n3256 ;
  assign n13178 = x2 & ~n11438 ;
  assign n13179 = n13178 ^ n1969 ^ 1'b0 ;
  assign n13180 = n9109 | n13116 ;
  assign n13181 = n1948 & ~n13180 ;
  assign n13182 = n2413 & ~n10730 ;
  assign n13183 = n6587 | n8217 ;
  assign n13184 = ~n673 & n12955 ;
  assign n13185 = n2460 & ~n13184 ;
  assign n13186 = n13183 & ~n13185 ;
  assign n13187 = n13186 ^ n8547 ^ 1'b0 ;
  assign n13190 = n11976 | n12848 ;
  assign n13191 = n12848 & ~n13190 ;
  assign n13188 = n11375 ^ n1867 ^ 1'b0 ;
  assign n13189 = n12285 & ~n13188 ;
  assign n13192 = n13191 ^ n13189 ^ n9481 ;
  assign n13193 = n3706 ^ n723 ^ 1'b0 ;
  assign n13194 = n13193 ^ n9609 ^ 1'b0 ;
  assign n13195 = ~n2853 & n13194 ;
  assign n13196 = ( n2170 & n4840 ) | ( n2170 & n13195 ) | ( n4840 & n13195 ) ;
  assign n13197 = n731 | n3589 ;
  assign n13198 = ~n5308 & n13197 ;
  assign n13199 = n4733 & n7693 ;
  assign n13200 = n13199 ^ n11833 ^ 1'b0 ;
  assign n13201 = n608 | n1096 ;
  assign n13202 = n1853 & ~n13201 ;
  assign n13203 = n5754 ^ n5616 ^ 1'b0 ;
  assign n13204 = n4347 & n13203 ;
  assign n13205 = ~n13202 & n13204 ;
  assign n13206 = n13205 ^ n6998 ^ 1'b0 ;
  assign n13207 = n13206 ^ n7130 ^ 1'b0 ;
  assign n13209 = ~n2054 & n3942 ;
  assign n13210 = ~n3942 & n13209 ;
  assign n13208 = n9100 & n10922 ;
  assign n13211 = n13210 ^ n13208 ^ 1'b0 ;
  assign n13212 = n6005 ^ n5022 ^ 1'b0 ;
  assign n13213 = n1662 & n13212 ;
  assign n13214 = ~n4400 & n13213 ;
  assign n13215 = n1757 & n5532 ;
  assign n13216 = n13215 ^ n2003 ^ 1'b0 ;
  assign n13217 = n7574 ^ n276 ^ 1'b0 ;
  assign n13218 = ( n6952 & ~n13216 ) | ( n6952 & n13217 ) | ( ~n13216 & n13217 ) ;
  assign n13219 = n13218 ^ n12929 ^ 1'b0 ;
  assign n13221 = n6653 & n10888 ;
  assign n13220 = n8536 & ~n12723 ;
  assign n13222 = n13221 ^ n13220 ^ 1'b0 ;
  assign n13223 = n5574 ^ n1981 ^ 1'b0 ;
  assign n13224 = n2259 & n13223 ;
  assign n13225 = n6015 ^ n3011 ^ 1'b0 ;
  assign n13226 = n12253 ^ n10158 ^ 1'b0 ;
  assign n13227 = ~n13225 & n13226 ;
  assign n13228 = n5432 ^ n3719 ^ 1'b0 ;
  assign n13229 = n13228 ^ n7050 ^ 1'b0 ;
  assign n13230 = n3608 | n10513 ;
  assign n13231 = n2402 | n11047 ;
  assign n13232 = ~n651 & n13231 ;
  assign n13233 = x165 & ~n1889 ;
  assign n13234 = n4036 & n5355 ;
  assign n13235 = n3037 & n13234 ;
  assign n13236 = n10455 & ~n13235 ;
  assign n13237 = n6684 ^ n2661 ^ 1'b0 ;
  assign n13238 = ~n4450 & n13237 ;
  assign n13239 = n13238 ^ n6688 ^ 1'b0 ;
  assign n13240 = ( n2110 & n2431 ) | ( n2110 & ~n10743 ) | ( n2431 & ~n10743 ) ;
  assign n13241 = n13240 ^ n1388 ^ 1'b0 ;
  assign n13242 = n7942 | n13241 ;
  assign n13243 = n13242 ^ x204 ^ 1'b0 ;
  assign n13244 = n3972 | n13243 ;
  assign n13245 = n3876 ^ n3102 ^ 1'b0 ;
  assign n13246 = n486 & n6102 ;
  assign n13247 = ~n860 & n13246 ;
  assign n13248 = n10208 & ~n13247 ;
  assign n13249 = n13248 ^ n3670 ^ 1'b0 ;
  assign n13250 = n13249 ^ n4588 ^ 1'b0 ;
  assign n13251 = n13245 | n13250 ;
  assign n13252 = n708 & n7251 ;
  assign n13253 = n1725 & n13252 ;
  assign n13254 = n13253 ^ n3154 ^ 1'b0 ;
  assign n13255 = n13254 ^ n7710 ^ n6184 ;
  assign n13256 = n9490 ^ n4402 ^ n3395 ;
  assign n13257 = n4290 ^ n2710 ^ 1'b0 ;
  assign n13258 = ~n13256 & n13257 ;
  assign n13259 = n2466 & n9111 ;
  assign n13260 = n5206 & ~n13259 ;
  assign n13261 = ~n7593 & n13260 ;
  assign n13262 = ~n4505 & n7630 ;
  assign n13263 = n3327 & n13262 ;
  assign n13264 = n13263 ^ n1504 ^ 1'b0 ;
  assign n13265 = n2668 & ~n4663 ;
  assign n13266 = ~n1387 & n13265 ;
  assign n13267 = x60 & n5168 ;
  assign n13268 = n10084 & ~n13267 ;
  assign n13271 = ~n3326 & n3876 ;
  assign n13272 = ~n6177 & n13271 ;
  assign n13269 = n9285 ^ n4545 ^ 1'b0 ;
  assign n13270 = n6412 & ~n13269 ;
  assign n13273 = n13272 ^ n13270 ^ 1'b0 ;
  assign n13274 = n1404 | n2321 ;
  assign n13275 = n6582 | n13274 ;
  assign n13276 = n13275 ^ n3714 ^ 1'b0 ;
  assign n13277 = n12048 & n13276 ;
  assign n13278 = n1272 & n5248 ;
  assign n13279 = n13278 ^ n12188 ^ n3686 ;
  assign n13280 = n8968 ^ n5352 ^ n1402 ;
  assign n13281 = n9340 & n13280 ;
  assign n13282 = n9541 ^ n9118 ^ 1'b0 ;
  assign n13283 = n4193 | n13282 ;
  assign n13284 = x222 & ~n4086 ;
  assign n13285 = n13284 ^ n357 ^ 1'b0 ;
  assign n13286 = n13285 ^ n772 ^ 1'b0 ;
  assign n13287 = n4824 ^ n1165 ^ 1'b0 ;
  assign n13288 = ~n1720 & n13287 ;
  assign n13289 = n1989 & ~n7242 ;
  assign n13290 = n1815 & n2948 ;
  assign n13291 = n13290 ^ n9109 ^ 1'b0 ;
  assign n13292 = n13291 ^ n7027 ^ 1'b0 ;
  assign n13293 = n11856 ^ n1481 ^ 1'b0 ;
  assign n13294 = ~n1720 & n10954 ;
  assign n13295 = n11978 ^ n2799 ^ 1'b0 ;
  assign n13296 = n8861 & n13295 ;
  assign n13297 = ( n2571 & n2982 ) | ( n2571 & ~n7248 ) | ( n2982 & ~n7248 ) ;
  assign n13298 = n262 & ~n13297 ;
  assign n13299 = n4856 & n13298 ;
  assign n13303 = n9964 ^ n446 ^ 1'b0 ;
  assign n13300 = n6619 & n8759 ;
  assign n13301 = n13300 ^ n6306 ^ 1'b0 ;
  assign n13302 = ~n963 & n13301 ;
  assign n13304 = n13303 ^ n13302 ^ 1'b0 ;
  assign n13305 = n1053 | n4214 ;
  assign n13308 = n7506 ^ n7361 ^ 1'b0 ;
  assign n13309 = n5309 | n13308 ;
  assign n13306 = n2095 ^ n1804 ^ 1'b0 ;
  assign n13307 = n2123 & n13306 ;
  assign n13310 = n13309 ^ n13307 ^ 1'b0 ;
  assign n13311 = n11533 & n13310 ;
  assign n13312 = n13311 ^ n7992 ^ n3893 ;
  assign n13313 = n7255 & ~n8951 ;
  assign n13314 = n13313 ^ n2701 ^ 1'b0 ;
  assign n13315 = n5031 | n13314 ;
  assign n13316 = ( n2566 & n7603 ) | ( n2566 & n7706 ) | ( n7603 & n7706 ) ;
  assign n13317 = n7378 ^ n2110 ^ 1'b0 ;
  assign n13318 = n13317 ^ n4085 ^ 1'b0 ;
  assign n13319 = n2198 | n5984 ;
  assign n13320 = x140 | n5865 ;
  assign n13321 = ~n6905 & n8815 ;
  assign n13322 = n882 & n13321 ;
  assign n13323 = x96 & ~n1728 ;
  assign n13324 = n13323 ^ n12235 ^ 1'b0 ;
  assign n13325 = n1605 | n13324 ;
  assign n13329 = ~n1657 & n12809 ;
  assign n13330 = n13329 ^ n6857 ^ 1'b0 ;
  assign n13326 = n5827 & n9100 ;
  assign n13327 = n13326 ^ n426 ^ 1'b0 ;
  assign n13328 = ~n10134 & n13327 ;
  assign n13331 = n13330 ^ n13328 ^ 1'b0 ;
  assign n13332 = n2069 & n7815 ;
  assign n13333 = ~n2069 & n13332 ;
  assign n13334 = ( n10242 & n12438 ) | ( n10242 & n13333 ) | ( n12438 & n13333 ) ;
  assign n13335 = n13334 ^ n11792 ^ 1'b0 ;
  assign n13337 = ~n2343 & n4263 ;
  assign n13338 = ~n5223 & n13337 ;
  assign n13336 = n4251 & n4970 ;
  assign n13339 = n13338 ^ n13336 ^ 1'b0 ;
  assign n13340 = n5177 ^ n1615 ^ 1'b0 ;
  assign n13341 = ~n2072 & n13340 ;
  assign n13342 = n6135 & n13341 ;
  assign n13343 = x110 & ~n13342 ;
  assign n13344 = n13343 ^ n2347 ^ 1'b0 ;
  assign n13345 = ~n12926 & n13344 ;
  assign n13348 = n9652 & n12249 ;
  assign n13349 = n3025 & n13348 ;
  assign n13346 = n1499 ^ x70 ^ 1'b0 ;
  assign n13347 = n13346 ^ n2282 ^ 1'b0 ;
  assign n13350 = n13349 ^ n13347 ^ 1'b0 ;
  assign n13351 = n781 & ~n13350 ;
  assign n13352 = n8933 ^ n8801 ^ 1'b0 ;
  assign n13354 = n4210 ^ n2367 ^ 1'b0 ;
  assign n13353 = n7746 ^ n2183 ^ x84 ;
  assign n13355 = n13354 ^ n13353 ^ 1'b0 ;
  assign n13356 = ( n387 & n9619 ) | ( n387 & n10629 ) | ( n9619 & n10629 ) ;
  assign n13357 = n9260 ^ n2641 ^ 1'b0 ;
  assign n13358 = n5018 | n13357 ;
  assign n13359 = n13356 & ~n13358 ;
  assign n13364 = n10398 ^ n8107 ^ n913 ;
  assign n13360 = n469 & n1570 ;
  assign n13361 = n5660 & ~n13360 ;
  assign n13362 = ~n3174 & n13361 ;
  assign n13363 = ~n3521 & n13362 ;
  assign n13365 = n13364 ^ n13363 ^ 1'b0 ;
  assign n13366 = n5915 & ~n6638 ;
  assign n13367 = n4360 | n10182 ;
  assign n13368 = n13367 ^ n6391 ^ 1'b0 ;
  assign n13372 = ~n3508 & n4425 ;
  assign n13370 = n4163 ^ n4004 ^ n3606 ;
  assign n13371 = n638 & n13370 ;
  assign n13373 = n13372 ^ n13371 ^ 1'b0 ;
  assign n13369 = n7507 | n13206 ;
  assign n13374 = n13373 ^ n13369 ^ 1'b0 ;
  assign n13375 = n2265 & ~n13374 ;
  assign n13376 = ~n2010 & n2544 ;
  assign n13377 = ~x33 & n13376 ;
  assign n13378 = n8358 & ~n13377 ;
  assign n13379 = n3890 & ~n11142 ;
  assign n13380 = n5509 ^ n1490 ^ n877 ;
  assign n13381 = ( ~n1837 & n10164 ) | ( ~n1837 & n10835 ) | ( n10164 & n10835 ) ;
  assign n13382 = n8352 ^ n7188 ^ 1'b0 ;
  assign n13383 = n9646 ^ n4665 ^ 1'b0 ;
  assign n13384 = ~n13382 & n13383 ;
  assign n13385 = n13384 ^ n4875 ^ n3777 ;
  assign n13389 = n10610 & n11943 ;
  assign n13390 = n13389 ^ n6042 ^ 1'b0 ;
  assign n13386 = n4044 | n8073 ;
  assign n13387 = n5772 | n13386 ;
  assign n13388 = ~n6260 & n13387 ;
  assign n13391 = n13390 ^ n13388 ^ 1'b0 ;
  assign n13392 = ~n4202 & n12896 ;
  assign n13393 = n13392 ^ n1432 ^ 1'b0 ;
  assign n13394 = n2782 | n13393 ;
  assign n13395 = x189 & ~n5347 ;
  assign n13396 = n13395 ^ n622 ^ 1'b0 ;
  assign n13397 = ~n10710 & n13396 ;
  assign n13398 = ~n4817 & n13397 ;
  assign n13399 = n13398 ^ n10897 ^ n2114 ;
  assign n13400 = n12264 ^ n10234 ^ 1'b0 ;
  assign n13401 = n6560 | n13400 ;
  assign n13402 = n3739 & ~n13401 ;
  assign n13403 = n12041 ^ n1822 ^ 1'b0 ;
  assign n13404 = n10454 & n13403 ;
  assign n13405 = n322 | n5953 ;
  assign n13407 = n12517 ^ n6395 ^ 1'b0 ;
  assign n13406 = ( n2593 & n5496 ) | ( n2593 & ~n8098 ) | ( n5496 & ~n8098 ) ;
  assign n13408 = n13407 ^ n13406 ^ 1'b0 ;
  assign n13409 = n1742 & n13408 ;
  assign n13410 = n10010 ^ n6781 ^ 1'b0 ;
  assign n13411 = n1945 & n8284 ;
  assign n13412 = ~n11776 & n13411 ;
  assign n13413 = n3271 & n4598 ;
  assign n13414 = ~n1213 & n13413 ;
  assign n13415 = n7019 ^ n3014 ^ 1'b0 ;
  assign n13416 = n13415 ^ n3637 ^ 1'b0 ;
  assign n13417 = n13414 | n13416 ;
  assign n13418 = n6037 ^ n4462 ^ n1553 ;
  assign n13420 = ~n6798 & n8897 ;
  assign n13419 = n11063 ^ n3186 ^ 1'b0 ;
  assign n13421 = n13420 ^ n13419 ^ 1'b0 ;
  assign n13422 = n13279 & ~n13421 ;
  assign n13423 = n13418 & n13422 ;
  assign n13424 = n6510 ^ n1593 ^ 1'b0 ;
  assign n13425 = n8730 ^ n6996 ^ n6397 ;
  assign n13426 = n13424 & n13425 ;
  assign n13427 = n7734 ^ n4848 ^ 1'b0 ;
  assign n13428 = n13427 ^ n3563 ^ 1'b0 ;
  assign n13429 = ~n8591 & n13428 ;
  assign n13430 = n13429 ^ x143 ^ 1'b0 ;
  assign n13431 = n13426 & ~n13430 ;
  assign n13437 = ( ~x125 & n1330 ) | ( ~x125 & n9437 ) | ( n1330 & n9437 ) ;
  assign n13438 = n6359 ^ n510 ^ 1'b0 ;
  assign n13439 = ( n12969 & n13437 ) | ( n12969 & ~n13438 ) | ( n13437 & ~n13438 ) ;
  assign n13432 = n4323 | n11580 ;
  assign n13433 = n3871 & ~n13432 ;
  assign n13434 = n12838 ^ n12359 ^ n5918 ;
  assign n13435 = n1545 & n13434 ;
  assign n13436 = ~n13433 & n13435 ;
  assign n13440 = n13439 ^ n13436 ^ 1'b0 ;
  assign n13441 = n4832 & n7338 ;
  assign n13442 = n3044 & n13441 ;
  assign n13443 = n1153 | n13442 ;
  assign n13444 = n11750 ^ n4305 ^ 1'b0 ;
  assign n13451 = n4447 ^ n2982 ^ 1'b0 ;
  assign n13447 = n3974 ^ n436 ^ 1'b0 ;
  assign n13448 = ~n1078 & n13447 ;
  assign n13445 = n3011 & n3016 ;
  assign n13446 = n8157 & n13445 ;
  assign n13449 = n13448 ^ n13446 ^ 1'b0 ;
  assign n13450 = n13449 ^ n3034 ^ 1'b0 ;
  assign n13452 = n13451 ^ n13450 ^ n4938 ;
  assign n13453 = n7830 & ~n9332 ;
  assign n13454 = ~n5118 & n13453 ;
  assign n13457 = ~n2061 & n8858 ;
  assign n13458 = ~n12455 & n13457 ;
  assign n13455 = ~n1557 & n11296 ;
  assign n13456 = n13455 ^ n11379 ^ 1'b0 ;
  assign n13459 = n13458 ^ n13456 ^ n4222 ;
  assign n13460 = n12162 ^ n9654 ^ 1'b0 ;
  assign n13461 = ~n8325 & n13460 ;
  assign n13462 = ~n3651 & n6954 ;
  assign n13463 = n6340 & n12586 ;
  assign n13464 = ~n622 & n2992 ;
  assign n13465 = n13464 ^ n12541 ^ n4673 ;
  assign n13466 = n8328 ^ x195 ^ 1'b0 ;
  assign n13467 = n10673 | n13466 ;
  assign n13468 = n5598 | n13467 ;
  assign n13469 = ~n3568 & n11094 ;
  assign n13470 = ( x68 & ~n3499 ) | ( x68 & n13469 ) | ( ~n3499 & n13469 ) ;
  assign n13471 = n11532 ^ x40 ^ 1'b0 ;
  assign n13472 = n7687 | n13471 ;
  assign n13473 = n13472 ^ n8580 ^ 1'b0 ;
  assign n13474 = n8138 | n13473 ;
  assign n13475 = ~n5602 & n10345 ;
  assign n13476 = n4867 & n13475 ;
  assign n13477 = n4254 | n5308 ;
  assign n13478 = n13477 ^ n2433 ^ 1'b0 ;
  assign n13479 = n3379 | n13478 ;
  assign n13480 = n4580 | n13479 ;
  assign n13481 = n1049 & n13480 ;
  assign n13482 = n6306 ^ n5571 ^ 1'b0 ;
  assign n13483 = ~n10172 & n13482 ;
  assign n13484 = n1073 | n13483 ;
  assign n13485 = n13484 ^ n9853 ^ 1'b0 ;
  assign n13486 = n9628 ^ n2274 ^ 1'b0 ;
  assign n13487 = n13486 ^ n4350 ^ 1'b0 ;
  assign n13488 = n11360 ^ n6157 ^ 1'b0 ;
  assign n13489 = n3294 & n13488 ;
  assign n13490 = n13489 ^ n2989 ^ 1'b0 ;
  assign n13491 = n13490 ^ n677 ^ 1'b0 ;
  assign n13493 = ( n4591 & ~n4723 ) | ( n4591 & n5957 ) | ( ~n4723 & n5957 ) ;
  assign n13492 = n2870 | n6462 ;
  assign n13494 = n13493 ^ n13492 ^ n12835 ;
  assign n13495 = n1878 & n9285 ;
  assign n13496 = n13495 ^ n9802 ^ 1'b0 ;
  assign n13498 = n4832 ^ n2883 ^ 1'b0 ;
  assign n13499 = n13498 ^ n1588 ^ 1'b0 ;
  assign n13500 = n5142 | n13499 ;
  assign n13497 = n6470 | n9017 ;
  assign n13501 = n13500 ^ n13497 ^ 1'b0 ;
  assign n13502 = n4357 & ~n13501 ;
  assign n13503 = n1177 ^ n359 ^ 1'b0 ;
  assign n13504 = n8693 ^ n7692 ^ 1'b0 ;
  assign n13505 = x128 & ~n2623 ;
  assign n13506 = n9365 | n13505 ;
  assign n13507 = n5076 ^ n3342 ^ 1'b0 ;
  assign n13508 = n6634 | n13507 ;
  assign n13509 = n13508 ^ n5001 ^ 1'b0 ;
  assign n13510 = n13509 ^ n7160 ^ 1'b0 ;
  assign n13511 = n8323 ^ n5569 ^ x229 ;
  assign n13512 = n5426 ^ n2954 ^ 1'b0 ;
  assign n13513 = n529 & ~n13512 ;
  assign n13514 = n8730 ^ n5028 ^ 1'b0 ;
  assign n13515 = n13513 & ~n13514 ;
  assign n13516 = n13515 ^ n4244 ^ 1'b0 ;
  assign n13517 = n5172 & n13516 ;
  assign n13518 = n7818 ^ n4097 ^ n2268 ;
  assign n13519 = n13518 ^ n3868 ^ 1'b0 ;
  assign n13520 = n13517 & n13519 ;
  assign n13521 = n11519 ^ n6342 ^ 1'b0 ;
  assign n13522 = n7677 ^ n4585 ^ 1'b0 ;
  assign n13523 = n5894 | n13522 ;
  assign n13524 = n9400 | n12481 ;
  assign n13525 = n779 & ~n2810 ;
  assign n13526 = ~n3600 & n9722 ;
  assign n13527 = ~n3092 & n13526 ;
  assign n13528 = n4534 ^ n2114 ^ 1'b0 ;
  assign n13529 = n8610 ^ n7635 ^ 1'b0 ;
  assign n13530 = n5274 ^ n4266 ^ n796 ;
  assign n13531 = n617 & ~n13530 ;
  assign n13532 = n5391 ^ n3215 ^ 1'b0 ;
  assign n13533 = n9355 ^ n2491 ^ 1'b0 ;
  assign n13534 = ~x137 & n12118 ;
  assign n13535 = n4222 ^ n2950 ^ 1'b0 ;
  assign n13536 = n6048 & ~n13535 ;
  assign n13537 = n13536 ^ n455 ^ 1'b0 ;
  assign n13538 = n9098 ^ n4220 ^ n1221 ;
  assign n13539 = ( ~n968 & n4209 ) | ( ~n968 & n9021 ) | ( n4209 & n9021 ) ;
  assign n13540 = ( x109 & n1758 ) | ( x109 & n1999 ) | ( n1758 & n1999 ) ;
  assign n13541 = ~n4360 & n13540 ;
  assign n13542 = ~x64 & n7736 ;
  assign n13543 = n13542 ^ n6460 ^ 1'b0 ;
  assign n13544 = n2011 & ~n13543 ;
  assign n13545 = ( n5611 & ~n8969 ) | ( n5611 & n10472 ) | ( ~n8969 & n10472 ) ;
  assign n13546 = n1602 & ~n3201 ;
  assign n13547 = n13546 ^ n10144 ^ 1'b0 ;
  assign n13549 = n6881 & ~n11972 ;
  assign n13548 = n5400 & n7972 ;
  assign n13550 = n13549 ^ n13548 ^ 1'b0 ;
  assign n13551 = n1284 | n2131 ;
  assign n13552 = n13551 ^ n7647 ^ 1'b0 ;
  assign n13553 = n1523 & n13552 ;
  assign n13554 = n9045 & n13553 ;
  assign n13555 = ~n2332 & n13554 ;
  assign n13556 = n7779 & n10630 ;
  assign n13557 = n13556 ^ n7018 ^ 1'b0 ;
  assign n13558 = n11558 & ~n13557 ;
  assign n13559 = n2868 | n9415 ;
  assign n13560 = n13559 ^ n1922 ^ 1'b0 ;
  assign n13561 = n3159 ^ n2775 ^ 1'b0 ;
  assign n13562 = n13560 & ~n13561 ;
  assign n13563 = n13562 ^ n6370 ^ n471 ;
  assign n13564 = n1503 ^ n1045 ^ 1'b0 ;
  assign n13565 = n13563 | n13564 ;
  assign n13566 = n13565 ^ n4229 ^ 1'b0 ;
  assign n13567 = n5949 & ~n13566 ;
  assign n13568 = n4868 ^ n1828 ^ 1'b0 ;
  assign n13569 = n6849 | n13568 ;
  assign n13570 = n9706 ^ n2576 ^ x119 ;
  assign n13571 = n3231 & n13570 ;
  assign n13572 = n2926 & n4995 ;
  assign n13573 = ~n4964 & n13572 ;
  assign n13574 = n3309 ^ n1295 ^ 1'b0 ;
  assign n13575 = ( ~n7360 & n13573 ) | ( ~n7360 & n13574 ) | ( n13573 & n13574 ) ;
  assign n13576 = ( ~x84 & n12152 ) | ( ~x84 & n13575 ) | ( n12152 & n13575 ) ;
  assign n13577 = n462 | n888 ;
  assign n13578 = n13577 ^ n6987 ^ 1'b0 ;
  assign n13582 = x148 & ~n2250 ;
  assign n13583 = ~n1210 & n13582 ;
  assign n13584 = n13583 ^ n11921 ^ 1'b0 ;
  assign n13579 = ( ~n676 & n3704 ) | ( ~n676 & n4995 ) | ( n3704 & n4995 ) ;
  assign n13580 = n11905 & n13579 ;
  assign n13581 = n2284 & n13580 ;
  assign n13585 = n13584 ^ n13581 ^ 1'b0 ;
  assign n13589 = n1866 & ~n11525 ;
  assign n13590 = ~n1866 & n13589 ;
  assign n13586 = n8119 ^ n3582 ^ 1'b0 ;
  assign n13587 = n6745 & n13586 ;
  assign n13588 = ~n13586 & n13587 ;
  assign n13591 = n13590 ^ n13588 ^ 1'b0 ;
  assign n13592 = n8853 & ~n13591 ;
  assign n13593 = ~n851 & n9511 ;
  assign n13594 = n13593 ^ n5685 ^ 1'b0 ;
  assign n13595 = n8169 ^ n3791 ^ 1'b0 ;
  assign n13596 = n3545 & ~n13595 ;
  assign n13597 = n13596 ^ n4540 ^ 1'b0 ;
  assign n13598 = ( ~n440 & n3019 ) | ( ~n440 & n13597 ) | ( n3019 & n13597 ) ;
  assign n13599 = ~n3425 & n7407 ;
  assign n13600 = n4085 & n13599 ;
  assign n13601 = ( n1186 & n5317 ) | ( n1186 & n13600 ) | ( n5317 & n13600 ) ;
  assign n13602 = ( n2928 & n3554 ) | ( n2928 & n7581 ) | ( n3554 & n7581 ) ;
  assign n13603 = n13602 ^ n9642 ^ 1'b0 ;
  assign n13604 = n10497 ^ n1276 ^ 1'b0 ;
  assign n13605 = n9237 & ~n13487 ;
  assign n13606 = n6604 & n13605 ;
  assign n13607 = n4675 ^ n2772 ^ 1'b0 ;
  assign n13608 = n13607 ^ n7961 ^ 1'b0 ;
  assign n13609 = n4350 & ~n11751 ;
  assign n13610 = n13609 ^ n4331 ^ 1'b0 ;
  assign n13611 = n7617 | n11817 ;
  assign n13613 = n2614 & ~n6437 ;
  assign n13612 = n449 & ~n9489 ;
  assign n13614 = n13613 ^ n13612 ^ 1'b0 ;
  assign n13615 = n8634 & n13614 ;
  assign n13616 = n11037 ^ n8382 ^ 1'b0 ;
  assign n13617 = n8145 ^ n2532 ^ 1'b0 ;
  assign n13618 = n13617 ^ n5384 ^ 1'b0 ;
  assign n13619 = n4910 ^ n2367 ^ 1'b0 ;
  assign n13620 = n4578 | n13619 ;
  assign n13621 = n9897 ^ n862 ^ 1'b0 ;
  assign n13622 = n13620 | n13621 ;
  assign n13623 = n13622 ^ n8752 ^ n1721 ;
  assign n13624 = n12108 ^ n4642 ^ 1'b0 ;
  assign n13625 = n13624 ^ n2622 ^ 1'b0 ;
  assign n13626 = n7375 & ~n13625 ;
  assign n13627 = n5595 & n13626 ;
  assign n13628 = n13623 & n13627 ;
  assign n13629 = ( ~n2587 & n3866 ) | ( ~n2587 & n4025 ) | ( n3866 & n4025 ) ;
  assign n13630 = n615 & ~n4310 ;
  assign n13631 = n5213 | n13630 ;
  assign n13632 = n13629 & ~n13631 ;
  assign n13633 = n3823 & n13632 ;
  assign n13634 = n9276 ^ n1490 ^ 1'b0 ;
  assign n13635 = n831 & ~n13634 ;
  assign n13636 = ( ~n5746 & n10756 ) | ( ~n5746 & n11497 ) | ( n10756 & n11497 ) ;
  assign n13637 = n10978 | n13636 ;
  assign n13638 = n13637 ^ n7495 ^ 1'b0 ;
  assign n13639 = n6348 | n8712 ;
  assign n13640 = n13639 ^ n2529 ^ 1'b0 ;
  assign n13641 = n1993 & n8717 ;
  assign n13642 = n2163 & n4213 ;
  assign n13643 = ~n13641 & n13642 ;
  assign n13644 = ( n3878 & ~n5280 ) | ( n3878 & n7920 ) | ( ~n5280 & n7920 ) ;
  assign n13645 = n13644 ^ n4821 ^ 1'b0 ;
  assign n13646 = n3412 & n13645 ;
  assign n13647 = ( n8083 & n13643 ) | ( n8083 & n13646 ) | ( n13643 & n13646 ) ;
  assign n13648 = n10268 ^ n4793 ^ 1'b0 ;
  assign n13649 = n6012 & n13648 ;
  assign n13650 = ( n1898 & ~n2245 ) | ( n1898 & n13649 ) | ( ~n2245 & n13649 ) ;
  assign n13651 = ~n946 & n1496 ;
  assign n13652 = n13651 ^ n9787 ^ 1'b0 ;
  assign n13653 = ~n5851 & n13652 ;
  assign n13654 = ( n10455 & n12574 ) | ( n10455 & n13653 ) | ( n12574 & n13653 ) ;
  assign n13656 = n2053 ^ n1124 ^ 1'b0 ;
  assign n13657 = n3841 & ~n13656 ;
  assign n13655 = n4375 & ~n7538 ;
  assign n13658 = n13657 ^ n13655 ^ 1'b0 ;
  assign n13659 = ~n865 & n3704 ;
  assign n13660 = n1589 & n13659 ;
  assign n13661 = n7685 & n13660 ;
  assign n13662 = n10155 ^ n6061 ^ 1'b0 ;
  assign n13663 = n1097 & n1919 ;
  assign n13664 = n13663 ^ n12765 ^ 1'b0 ;
  assign n13665 = n5998 ^ n5402 ^ 1'b0 ;
  assign n13666 = n13664 & n13665 ;
  assign n13667 = n6914 ^ n2735 ^ 1'b0 ;
  assign n13668 = n13666 & n13667 ;
  assign n13669 = n10131 & n13668 ;
  assign n13670 = ~n13662 & n13669 ;
  assign n13671 = n13670 ^ n10281 ^ 1'b0 ;
  assign n13672 = n6897 ^ n4837 ^ n2045 ;
  assign n13673 = n8663 | n13672 ;
  assign n13674 = n4954 & n10949 ;
  assign n13675 = ~n4976 & n13674 ;
  assign n13676 = n13675 ^ n5539 ^ 1'b0 ;
  assign n13677 = n3415 | n13676 ;
  assign n13678 = n2789 & ~n13677 ;
  assign n13679 = n6155 ^ n5488 ^ 1'b0 ;
  assign n13680 = n13679 ^ n10974 ^ 1'b0 ;
  assign n13681 = n12987 ^ n6120 ^ 1'b0 ;
  assign n13682 = n13680 & n13681 ;
  assign n13683 = ~n1985 & n4343 ;
  assign n13684 = ~n1215 & n5179 ;
  assign n13685 = n7738 & n13684 ;
  assign n13686 = n6741 ^ n1538 ^ 1'b0 ;
  assign n13687 = ~n9605 & n13686 ;
  assign n13688 = n1439 & n13687 ;
  assign n13689 = n436 & n640 ;
  assign n13690 = n4107 & ~n13689 ;
  assign n13691 = ~n4654 & n6596 ;
  assign n13692 = n11043 | n13691 ;
  assign n13693 = n342 & ~n11072 ;
  assign n13694 = n5313 & ~n5387 ;
  assign n13695 = ( n956 & ~n2556 ) | ( n956 & n13694 ) | ( ~n2556 & n13694 ) ;
  assign n13696 = n4094 | n13695 ;
  assign n13697 = n13693 | n13696 ;
  assign n13698 = n5818 ^ n3186 ^ 1'b0 ;
  assign n13699 = n4042 | n13698 ;
  assign n13700 = n9694 | n13699 ;
  assign n13701 = n810 | n1075 ;
  assign n13702 = n302 & n7315 ;
  assign n13703 = ~n302 & n13702 ;
  assign n13704 = n11264 | n13703 ;
  assign n13705 = n10606 & n13704 ;
  assign n13706 = n2554 ^ n520 ^ 1'b0 ;
  assign n13707 = n4511 ^ n2812 ^ 1'b0 ;
  assign n13708 = n2725 | n13707 ;
  assign n13709 = n518 & ~n13708 ;
  assign n13710 = ~n9204 & n13709 ;
  assign n13711 = n13710 ^ x125 ^ 1'b0 ;
  assign n13712 = n5983 | n13711 ;
  assign n13713 = n5205 & ~n13712 ;
  assign n13714 = n8660 ^ n4769 ^ n2593 ;
  assign n13715 = n7655 & ~n13714 ;
  assign n13716 = n13715 ^ n4180 ^ 1'b0 ;
  assign n13717 = n13716 ^ n872 ^ 1'b0 ;
  assign n13718 = ~n2828 & n13717 ;
  assign n13719 = n5767 & ~n13406 ;
  assign n13720 = n2726 & n10041 ;
  assign n13724 = n9068 ^ n5745 ^ 1'b0 ;
  assign n13725 = x73 & n13724 ;
  assign n13726 = n13725 ^ n10778 ^ 1'b0 ;
  assign n13721 = n1497 & n1611 ;
  assign n13722 = n13721 ^ n2877 ^ 1'b0 ;
  assign n13723 = ~n10169 & n13722 ;
  assign n13727 = n13726 ^ n13723 ^ 1'b0 ;
  assign n13728 = n1437 | n3683 ;
  assign n13729 = n7951 | n13728 ;
  assign n13730 = n13729 ^ n6903 ^ 1'b0 ;
  assign n13731 = n4678 ^ n789 ^ 1'b0 ;
  assign n13732 = n10843 & n13731 ;
  assign n13735 = n6352 & n10601 ;
  assign n13733 = n5976 & ~n13482 ;
  assign n13734 = ~n7228 & n13733 ;
  assign n13736 = n13735 ^ n13734 ^ 1'b0 ;
  assign n13737 = n5626 & n13736 ;
  assign n13738 = ~n3511 & n13737 ;
  assign n13739 = n3046 ^ n1019 ^ x214 ;
  assign n13740 = n13739 ^ n701 ^ 1'b0 ;
  assign n13741 = n13740 ^ n4195 ^ 1'b0 ;
  assign n13742 = n13741 ^ n1600 ^ 1'b0 ;
  assign n13743 = n13384 & n13742 ;
  assign n13744 = n2069 & ~n6723 ;
  assign n13745 = ~n2069 & n13744 ;
  assign n13746 = n8970 & n9804 ;
  assign n13747 = n3590 & n13746 ;
  assign n13749 = x59 & x148 ;
  assign n13750 = ~x59 & n13749 ;
  assign n13751 = n618 & n4480 ;
  assign n13752 = ~n618 & n13751 ;
  assign n13753 = n13750 & ~n13752 ;
  assign n13748 = n1364 | n5206 ;
  assign n13754 = n13753 ^ n13748 ^ 1'b0 ;
  assign n13755 = n13754 ^ n4316 ^ 1'b0 ;
  assign n13756 = n13747 | n13755 ;
  assign n13758 = n9549 & ~n11643 ;
  assign n13759 = n13758 ^ n2997 ^ 1'b0 ;
  assign n13757 = n891 & n6133 ;
  assign n13760 = n13759 ^ n13757 ^ 1'b0 ;
  assign n13761 = n4949 | n6120 ;
  assign n13762 = n13761 ^ n10480 ^ 1'b0 ;
  assign n13763 = ~n5029 & n13018 ;
  assign n13764 = ~n1873 & n1879 ;
  assign n13765 = n13764 ^ n10861 ^ 1'b0 ;
  assign n13766 = n9719 ^ n3674 ^ 1'b0 ;
  assign n13767 = n8927 ^ n3588 ^ 1'b0 ;
  assign n13768 = n2167 & n10374 ;
  assign n13769 = ~n3118 & n9815 ;
  assign n13772 = n3579 | n3749 ;
  assign n13773 = n13772 ^ n6949 ^ 1'b0 ;
  assign n13770 = n7647 & n10816 ;
  assign n13771 = ~n6918 & n13770 ;
  assign n13774 = n13773 ^ n13771 ^ 1'b0 ;
  assign n13775 = n2819 & n5248 ;
  assign n13776 = n13775 ^ n7996 ^ 1'b0 ;
  assign n13777 = ( n9451 & n13774 ) | ( n9451 & ~n13776 ) | ( n13774 & ~n13776 ) ;
  assign n13778 = ~n11857 & n12366 ;
  assign n13779 = ~n3805 & n5692 ;
  assign n13780 = ( n2287 & n3614 ) | ( n2287 & ~n13779 ) | ( n3614 & ~n13779 ) ;
  assign n13781 = n7543 & ~n10327 ;
  assign n13782 = n11068 ^ n3770 ^ 1'b0 ;
  assign n13783 = n12236 ^ n6693 ^ n6193 ;
  assign n13784 = ~n2867 & n2942 ;
  assign n13785 = n13784 ^ n5390 ^ 1'b0 ;
  assign n13786 = n13785 ^ n7872 ^ 1'b0 ;
  assign n13787 = ~n1215 & n13786 ;
  assign n13788 = n10281 ^ n3235 ^ 1'b0 ;
  assign n13789 = n1135 & ~n13788 ;
  assign n13790 = ~n3161 & n13789 ;
  assign n13791 = n10451 | n12798 ;
  assign n13792 = n13791 ^ n4542 ^ 1'b0 ;
  assign n13793 = n12937 & ~n13792 ;
  assign n13794 = n3966 & ~n9742 ;
  assign n13795 = n1775 | n3525 ;
  assign n13796 = ( n3704 & ~n13794 ) | ( n3704 & n13795 ) | ( ~n13794 & n13795 ) ;
  assign n13798 = n8104 ^ n2050 ^ 1'b0 ;
  assign n13799 = n13798 ^ n12835 ^ n1232 ;
  assign n13797 = n1020 | n7273 ;
  assign n13800 = n13799 ^ n13797 ^ 1'b0 ;
  assign n13801 = ~x94 & n8136 ;
  assign n13802 = ~n6424 & n9709 ;
  assign n13803 = ( n1276 & n5628 ) | ( n1276 & n9090 ) | ( n5628 & n9090 ) ;
  assign n13804 = n12001 ^ n10876 ^ 1'b0 ;
  assign n13805 = n13803 & n13804 ;
  assign n13806 = n13478 ^ n12436 ^ 1'b0 ;
  assign n13807 = n2228 & n6086 ;
  assign n13808 = n12322 ^ n3319 ^ 1'b0 ;
  assign n13809 = n5746 ^ n323 ^ 1'b0 ;
  assign n13810 = n11462 | n13809 ;
  assign n13811 = n5138 ^ n4109 ^ 1'b0 ;
  assign n13812 = n9754 | n13811 ;
  assign n13813 = ( n1696 & n2229 ) | ( n1696 & ~n4521 ) | ( n2229 & ~n4521 ) ;
  assign n13814 = n13813 ^ n6337 ^ 1'b0 ;
  assign n13815 = x144 & ~n4521 ;
  assign n13816 = n13815 ^ n3199 ^ 1'b0 ;
  assign n13817 = n13814 | n13816 ;
  assign n13818 = ~n8604 & n9704 ;
  assign n13819 = ~n3878 & n12017 ;
  assign n13820 = ~n12017 & n13819 ;
  assign n13821 = n540 & ~n12172 ;
  assign n13822 = n13820 | n13821 ;
  assign n13823 = n13820 & ~n13822 ;
  assign n13824 = n420 & ~n935 ;
  assign n13825 = n2877 | n3726 ;
  assign n13826 = n1338 & ~n2368 ;
  assign n13827 = ~n13825 & n13826 ;
  assign n13828 = n1167 & n13827 ;
  assign n13829 = n13824 & n13828 ;
  assign n13830 = n8548 | n13829 ;
  assign n13831 = n5488 ^ n1714 ^ 1'b0 ;
  assign n13832 = n327 | n6025 ;
  assign n13833 = n13832 ^ n10812 ^ 1'b0 ;
  assign n13834 = ~n13831 & n13833 ;
  assign n13835 = n12966 ^ n10433 ^ 1'b0 ;
  assign n13836 = n5058 ^ n889 ^ 1'b0 ;
  assign n13837 = ~n3169 & n8037 ;
  assign n13838 = n13837 ^ n1273 ^ 1'b0 ;
  assign n13839 = n13838 ^ n8691 ^ 1'b0 ;
  assign n13840 = n2609 & n5513 ;
  assign n13841 = n13840 ^ n8446 ^ 1'b0 ;
  assign n13842 = n13839 | n13841 ;
  assign n13843 = n2896 & ~n3650 ;
  assign n13844 = n13843 ^ n7266 ^ 1'b0 ;
  assign n13847 = n4035 & n4078 ;
  assign n13845 = n7368 ^ n3221 ^ 1'b0 ;
  assign n13846 = n13585 & ~n13845 ;
  assign n13848 = n13847 ^ n13846 ^ 1'b0 ;
  assign n13849 = n2287 & ~n3710 ;
  assign n13850 = n3600 & ~n9212 ;
  assign n13851 = n5743 & n13850 ;
  assign n13852 = n13851 ^ n3032 ^ 1'b0 ;
  assign n13853 = ~n12288 & n13852 ;
  assign n13854 = ~n2549 & n9643 ;
  assign n13855 = n8731 & n13854 ;
  assign n13856 = ~n1301 & n8150 ;
  assign n13857 = n13856 ^ n2016 ^ 1'b0 ;
  assign n13858 = n4610 ^ n444 ^ 1'b0 ;
  assign n13859 = n2196 | n13858 ;
  assign n13860 = n13859 ^ n8618 ^ 1'b0 ;
  assign n13861 = ( ~n2332 & n9803 ) | ( ~n2332 & n12466 ) | ( n9803 & n12466 ) ;
  assign n13862 = n13861 ^ n8547 ^ 1'b0 ;
  assign n13863 = n13679 ^ n2714 ^ 1'b0 ;
  assign n13864 = n7875 ^ n5458 ^ 1'b0 ;
  assign n13865 = x218 | n3161 ;
  assign n13866 = ~n13864 & n13865 ;
  assign n13867 = n7361 & n13866 ;
  assign n13868 = n9456 ^ n7038 ^ 1'b0 ;
  assign n13869 = n2312 & ~n13868 ;
  assign n13870 = ~n1114 & n2247 ;
  assign n13871 = ~n347 & n13629 ;
  assign n13872 = n5802 | n6753 ;
  assign n13873 = n13871 & ~n13872 ;
  assign n13874 = n10903 & ~n13873 ;
  assign n13875 = n13874 ^ n11010 ^ 1'b0 ;
  assign n13876 = n12553 & n13807 ;
  assign n13877 = n13876 ^ n4924 ^ 1'b0 ;
  assign n13878 = n10333 ^ n4222 ^ n3775 ;
  assign n13879 = n3978 & ~n5139 ;
  assign n13880 = n13878 & n13879 ;
  assign n13881 = ~n3255 & n4049 ;
  assign n13882 = n3481 & n13881 ;
  assign n13883 = n13882 ^ n6931 ^ n4149 ;
  assign n13884 = ~n5316 & n6553 ;
  assign n13885 = n13884 ^ n6263 ^ 1'b0 ;
  assign n13886 = n5237 ^ x55 ^ 1'b0 ;
  assign n13887 = ~n583 & n13886 ;
  assign n13888 = ~n8160 & n13887 ;
  assign n13889 = n13885 & n13888 ;
  assign n13890 = n7326 | n13794 ;
  assign n13891 = n13890 ^ n4144 ^ 1'b0 ;
  assign n13892 = n763 & n13891 ;
  assign n13893 = n4027 | n7294 ;
  assign n13894 = n13893 ^ n713 ^ 1'b0 ;
  assign n13895 = ( ~x23 & n9027 ) | ( ~x23 & n13894 ) | ( n9027 & n13894 ) ;
  assign n13896 = n13895 ^ n8325 ^ n1138 ;
  assign n13897 = n4125 & ~n12723 ;
  assign n13898 = ~n2394 & n9433 ;
  assign n13899 = n6345 & n13898 ;
  assign n13900 = n13508 & ~n13899 ;
  assign n13901 = n361 & ~n8704 ;
  assign n13902 = n8645 ^ n5187 ^ 1'b0 ;
  assign n13903 = n13901 & n13902 ;
  assign n13904 = n10038 ^ n6158 ^ 1'b0 ;
  assign n13905 = ~n4868 & n13904 ;
  assign n13906 = n9016 & n13905 ;
  assign n13907 = ~n5635 & n6898 ;
  assign n13908 = n13907 ^ n9290 ^ 1'b0 ;
  assign n13909 = ( n1254 & n13463 ) | ( n1254 & n13908 ) | ( n13463 & n13908 ) ;
  assign n13910 = n6987 | n13909 ;
  assign n13911 = n12704 | n13910 ;
  assign n13912 = n2881 ^ n537 ^ 1'b0 ;
  assign n13913 = n10085 & n13419 ;
  assign n13914 = n9402 ^ n6854 ^ 1'b0 ;
  assign n13916 = n3690 & n7923 ;
  assign n13917 = n13916 ^ n4679 ^ 1'b0 ;
  assign n13915 = x120 & ~n4395 ;
  assign n13918 = n13917 ^ n13915 ^ 1'b0 ;
  assign n13919 = n13914 & ~n13918 ;
  assign n13920 = n8822 ^ n3142 ^ 1'b0 ;
  assign n13921 = ~n12095 & n13920 ;
  assign n13922 = ~n1129 & n13921 ;
  assign n13923 = n9461 ^ n462 ^ 1'b0 ;
  assign n13924 = n3393 | n5292 ;
  assign n13925 = n13924 ^ n5737 ^ 1'b0 ;
  assign n13926 = n387 & ~n13925 ;
  assign n13927 = n7819 & n11795 ;
  assign n13928 = n13927 ^ n8815 ^ 1'b0 ;
  assign n13929 = n5051 & n13928 ;
  assign n13930 = ~n2199 & n13929 ;
  assign n13931 = n13930 ^ n9881 ^ 1'b0 ;
  assign n13932 = n13800 ^ n8048 ^ 1'b0 ;
  assign n13933 = n684 | n5373 ;
  assign n13934 = n3701 | n13933 ;
  assign n13935 = x155 & n13934 ;
  assign n13936 = n3768 & n13935 ;
  assign n13938 = n7630 ^ x141 ^ 1'b0 ;
  assign n13939 = ~n8968 & n13938 ;
  assign n13940 = n13939 ^ n7110 ^ 1'b0 ;
  assign n13937 = n1688 & n8604 ;
  assign n13941 = n13940 ^ n13937 ^ 1'b0 ;
  assign n13942 = n11089 & ~n13941 ;
  assign n13943 = n6903 ^ n2146 ^ 1'b0 ;
  assign n13944 = n6045 & n13943 ;
  assign n13945 = n13025 ^ n8604 ^ n4988 ;
  assign n13946 = n13944 & n13945 ;
  assign n13947 = n7162 ^ n4342 ^ 1'b0 ;
  assign n13949 = n7799 & n9484 ;
  assign n13948 = n1903 | n11818 ;
  assign n13950 = n13949 ^ n13948 ^ n9830 ;
  assign n13951 = n13950 ^ n13175 ^ 1'b0 ;
  assign n13952 = n9437 ^ n7028 ^ 1'b0 ;
  assign n13953 = n991 & n2499 ;
  assign n13954 = n13953 ^ n751 ^ 1'b0 ;
  assign n13955 = n8947 ^ n908 ^ 1'b0 ;
  assign n13956 = ~n5154 & n6138 ;
  assign n13957 = n5154 & n13956 ;
  assign n13958 = n7444 ^ n4724 ^ 1'b0 ;
  assign n13959 = n2228 & n13958 ;
  assign n13960 = n13959 ^ n2193 ^ 1'b0 ;
  assign n13961 = x76 & n9847 ;
  assign n13962 = n13961 ^ x236 ^ 1'b0 ;
  assign n13963 = n3364 & ~n13962 ;
  assign n13964 = ~n10449 & n13963 ;
  assign n13965 = n13405 ^ n7002 ^ 1'b0 ;
  assign n13966 = n13313 ^ n8967 ^ n3646 ;
  assign n13967 = n6474 | n11292 ;
  assign n13968 = n6496 & ~n13967 ;
  assign n13969 = n13968 ^ n2320 ^ 1'b0 ;
  assign n13970 = n5560 & n7402 ;
  assign n13971 = n13970 ^ n6339 ^ 1'b0 ;
  assign n13972 = n7371 & n13971 ;
  assign n13973 = ~n6345 & n13972 ;
  assign n13974 = n5912 | n6452 ;
  assign n13975 = n7502 ^ n5697 ^ 1'b0 ;
  assign n13976 = n5342 ^ n3858 ^ 1'b0 ;
  assign n13977 = n7059 ^ n1398 ^ 1'b0 ;
  assign n13978 = n13976 & ~n13977 ;
  assign n13979 = n566 & ~n13978 ;
  assign n13980 = n625 & n6425 ;
  assign n13981 = n542 & n13980 ;
  assign n13982 = ~n12547 & n13981 ;
  assign n13983 = n7385 | n13342 ;
  assign n13984 = n4361 & ~n13983 ;
  assign n13985 = n13984 ^ n3929 ^ 1'b0 ;
  assign n13986 = n2995 ^ n2443 ^ 1'b0 ;
  assign n13987 = n2334 & n4597 ;
  assign n13988 = n13987 ^ n11089 ^ 1'b0 ;
  assign n13989 = n13988 ^ n5390 ^ 1'b0 ;
  assign n13990 = n13986 & n13989 ;
  assign n13991 = ~n2622 & n5746 ;
  assign n13992 = n2178 & ~n13991 ;
  assign n13993 = n6059 ^ x130 ^ 1'b0 ;
  assign n13994 = n4124 & ~n13993 ;
  assign n13995 = ~n7643 & n13994 ;
  assign n13997 = n1366 & n6469 ;
  assign n13998 = ~n10298 & n13997 ;
  assign n13996 = ~n973 & n10072 ;
  assign n13999 = n13998 ^ n13996 ^ 1'b0 ;
  assign n14000 = ~x54 & n5456 ;
  assign n14001 = n10414 | n14000 ;
  assign n14002 = n1701 & ~n14001 ;
  assign n14003 = n13116 ^ n8125 ^ 1'b0 ;
  assign n14004 = n10781 ^ n3461 ^ 1'b0 ;
  assign n14005 = n1878 & n7949 ;
  assign n14006 = ~n1199 & n8314 ;
  assign n14007 = x144 & n5846 ;
  assign n14008 = n14006 | n14007 ;
  assign n14009 = n6808 ^ n4634 ^ 1'b0 ;
  assign n14010 = ~n9654 & n14009 ;
  assign n14011 = n1878 & ~n14010 ;
  assign n14012 = ~n14008 & n14011 ;
  assign n14013 = x40 & ~n7138 ;
  assign n14014 = ~n2155 & n14013 ;
  assign n14015 = n3925 ^ n1451 ^ 1'b0 ;
  assign n14016 = n14015 ^ n6797 ^ 1'b0 ;
  assign n14017 = n1999 ^ n572 ^ x141 ;
  assign n14018 = n3755 & n14017 ;
  assign n14019 = ~n14016 & n14018 ;
  assign n14020 = n8969 ^ n7275 ^ 1'b0 ;
  assign n14021 = n7727 ^ n5800 ^ 1'b0 ;
  assign n14022 = n3335 & ~n9425 ;
  assign n14023 = n8110 ^ n4114 ^ 1'b0 ;
  assign n14024 = ~n8594 & n10606 ;
  assign n14025 = ~n627 & n14024 ;
  assign n14026 = n14025 ^ n7601 ^ 1'b0 ;
  assign n14027 = n6412 & ~n14026 ;
  assign n14029 = ~n9654 & n10110 ;
  assign n14028 = n3823 & ~n12972 ;
  assign n14030 = n14029 ^ n14028 ^ 1'b0 ;
  assign n14031 = n6058 & n14030 ;
  assign n14032 = ~n14027 & n14031 ;
  assign n14033 = ~n11523 & n13693 ;
  assign n14034 = n14033 ^ n930 ^ 1'b0 ;
  assign n14035 = ~n634 & n8629 ;
  assign n14036 = n14034 & n14035 ;
  assign n14037 = ~n9354 & n11628 ;
  assign n14038 = n6152 ^ n2643 ^ 1'b0 ;
  assign n14039 = ~n3196 & n6769 ;
  assign n14040 = n14039 ^ n11206 ^ 1'b0 ;
  assign n14041 = ~n3880 & n14040 ;
  assign n14042 = n14041 ^ n1665 ^ 1'b0 ;
  assign n14043 = ~n1499 & n14042 ;
  assign n14044 = ~n14038 & n14043 ;
  assign n14045 = n5293 & ~n12826 ;
  assign n14046 = n1400 ^ n589 ^ 1'b0 ;
  assign n14047 = n949 & ~n14046 ;
  assign n14048 = n11323 & ~n14047 ;
  assign n14049 = ~n1288 & n7522 ;
  assign n14050 = n3362 & ~n7007 ;
  assign n14051 = n1045 & n14050 ;
  assign n14052 = ~n10625 & n14051 ;
  assign n14053 = n1950 & n3723 ;
  assign n14054 = n5416 | n8583 ;
  assign n14055 = n14054 ^ n12958 ^ 1'b0 ;
  assign n14056 = n772 & n1220 ;
  assign n14057 = ~n5005 & n14056 ;
  assign n14058 = n14055 | n14057 ;
  assign n14059 = n14053 | n14058 ;
  assign n14060 = n1328 | n2144 ;
  assign n14061 = n1170 & n6241 ;
  assign n14062 = n14061 ^ n3184 ^ 1'b0 ;
  assign n14063 = n9934 ^ n3677 ^ 1'b0 ;
  assign n14064 = x41 | n13474 ;
  assign n14065 = ( n614 & ~n808 ) | ( n614 & n1272 ) | ( ~n808 & n1272 ) ;
  assign n14066 = n14065 ^ n11430 ^ 1'b0 ;
  assign n14067 = n14066 ^ n3025 ^ 1'b0 ;
  assign n14068 = n12725 ^ n7418 ^ n6712 ;
  assign n14069 = n14067 & ~n14068 ;
  assign n14070 = n14069 ^ n2472 ^ 1'b0 ;
  assign n14071 = n2366 | n4172 ;
  assign n14072 = n14071 ^ n875 ^ 1'b0 ;
  assign n14073 = ( n1324 & ~n10350 ) | ( n1324 & n14072 ) | ( ~n10350 & n14072 ) ;
  assign n14074 = ~n3705 & n13807 ;
  assign n14075 = n4258 & n8981 ;
  assign n14076 = ~n6155 & n14075 ;
  assign n14077 = n4603 ^ n3186 ^ 1'b0 ;
  assign n14078 = n1356 & ~n14077 ;
  assign n14079 = n11483 & n14078 ;
  assign n14080 = n14079 ^ n4532 ^ 1'b0 ;
  assign n14081 = ( n11760 & n12108 ) | ( n11760 & ~n14080 ) | ( n12108 & ~n14080 ) ;
  assign n14082 = n917 & n6920 ;
  assign n14083 = n14082 ^ n11292 ^ 1'b0 ;
  assign n14084 = n3686 | n9809 ;
  assign n14085 = n2210 & n3677 ;
  assign n14086 = n14085 ^ n9967 ^ 1'b0 ;
  assign n14087 = n3145 ^ n2452 ^ 1'b0 ;
  assign n14088 = n14087 ^ n5857 ^ 1'b0 ;
  assign n14089 = ~n692 & n1445 ;
  assign n14090 = n14089 ^ n8058 ^ 1'b0 ;
  assign n14091 = n14090 ^ n3812 ^ 1'b0 ;
  assign n14092 = n11001 & n14091 ;
  assign n14093 = n6483 ^ n1630 ^ 1'b0 ;
  assign n14094 = ~n8658 & n14093 ;
  assign n14095 = n1333 & n14094 ;
  assign n14096 = n10089 & n14095 ;
  assign n14097 = ( n891 & ~n2252 ) | ( n891 & n4872 ) | ( ~n2252 & n4872 ) ;
  assign n14098 = ( n655 & n6273 ) | ( n655 & n7624 ) | ( n6273 & n7624 ) ;
  assign n14099 = ( n1125 & n4910 ) | ( n1125 & n7180 ) | ( n4910 & n7180 ) ;
  assign n14100 = n13340 ^ n4962 ^ 1'b0 ;
  assign n14101 = n9289 & ~n14100 ;
  assign n14102 = n1261 | n14101 ;
  assign n14103 = n14102 ^ n7516 ^ 1'b0 ;
  assign n14104 = n14099 & n14103 ;
  assign n14105 = n314 | n8185 ;
  assign n14106 = n10947 & ~n12036 ;
  assign n14107 = ~n2919 & n14106 ;
  assign n14108 = n11049 ^ n606 ^ 1'b0 ;
  assign n14109 = n10225 & ~n14108 ;
  assign n14110 = n1269 & n14109 ;
  assign n14111 = n14110 ^ n4632 ^ 1'b0 ;
  assign n14112 = n14107 & ~n14111 ;
  assign n14113 = n2408 & n12319 ;
  assign n14114 = ~n14112 & n14113 ;
  assign n14115 = n14114 ^ n1328 ^ n448 ;
  assign n14116 = n651 | n5034 ;
  assign n14117 = n14116 ^ n3641 ^ 1'b0 ;
  assign n14118 = n14117 ^ n6994 ^ 1'b0 ;
  assign n14119 = n1600 & ~n3449 ;
  assign n14120 = n3012 & n14119 ;
  assign n14121 = ( n765 & n12268 ) | ( n765 & ~n14120 ) | ( n12268 & ~n14120 ) ;
  assign n14122 = ~n10096 & n14121 ;
  assign n14123 = n9354 ^ n2294 ^ 1'b0 ;
  assign n14124 = n12972 | n14123 ;
  assign n14125 = ~n1124 & n7191 ;
  assign n14126 = ( x70 & x217 ) | ( x70 & ~n9705 ) | ( x217 & ~n9705 ) ;
  assign n14130 = n3121 ^ n932 ^ 1'b0 ;
  assign n14131 = ~n7326 & n14130 ;
  assign n14127 = ~n4913 & n4943 ;
  assign n14128 = n14127 ^ n1678 ^ 1'b0 ;
  assign n14129 = n4780 | n14128 ;
  assign n14132 = n14131 ^ n14129 ^ 1'b0 ;
  assign n14133 = n3018 ^ n2494 ^ 1'b0 ;
  assign n14134 = n2267 & ~n7231 ;
  assign n14135 = n4001 & n5163 ;
  assign n14136 = n7486 & n14135 ;
  assign n14137 = n1369 | n14136 ;
  assign n14138 = n14134 & ~n14137 ;
  assign n14139 = n9306 ^ n1992 ^ 1'b0 ;
  assign n14140 = n3719 ^ n2756 ^ 1'b0 ;
  assign n14141 = n7181 ^ n3271 ^ 1'b0 ;
  assign n14142 = n14141 ^ n8720 ^ 1'b0 ;
  assign n14143 = n7454 & n7553 ;
  assign n14146 = n3468 ^ n688 ^ 1'b0 ;
  assign n14144 = n3054 ^ n2529 ^ 1'b0 ;
  assign n14145 = n2073 | n14144 ;
  assign n14147 = n14146 ^ n14145 ^ 1'b0 ;
  assign n14148 = ( n464 & ~n6982 ) | ( n464 & n14147 ) | ( ~n6982 & n14147 ) ;
  assign n14149 = ~n3579 & n5625 ;
  assign n14150 = n14149 ^ n11170 ^ 1'b0 ;
  assign n14151 = ~n4426 & n14150 ;
  assign n14152 = n14151 ^ n2110 ^ 1'b0 ;
  assign n14153 = n6095 ^ n4209 ^ 1'b0 ;
  assign n14154 = n1937 | n3042 ;
  assign n14155 = n14154 ^ n10965 ^ 1'b0 ;
  assign n14156 = n11574 ^ n6923 ^ 1'b0 ;
  assign n14157 = n1521 & n10360 ;
  assign n14158 = n4892 & n14157 ;
  assign n14159 = x21 & ~n9204 ;
  assign n14160 = ( n6875 & n11433 ) | ( n6875 & ~n14159 ) | ( n11433 & ~n14159 ) ;
  assign n14161 = ~n4711 & n14160 ;
  assign n14162 = n8736 & n14161 ;
  assign n14163 = x142 & ~x234 ;
  assign n14164 = n11836 & n14163 ;
  assign n14165 = ( n1385 & ~n1948 ) | ( n1385 & n7501 ) | ( ~n1948 & n7501 ) ;
  assign n14166 = n14165 ^ n5786 ^ 1'b0 ;
  assign n14167 = n2167 ^ n1613 ^ n991 ;
  assign n14168 = n14167 ^ n6265 ^ 1'b0 ;
  assign n14169 = n886 & n3166 ;
  assign n14170 = ( ~x13 & n2230 ) | ( ~x13 & n14169 ) | ( n2230 & n14169 ) ;
  assign n14171 = n7350 & ~n10217 ;
  assign n14172 = n1718 | n14171 ;
  assign n14173 = n14172 ^ n7603 ^ 1'b0 ;
  assign n14174 = n2070 | n14173 ;
  assign n14175 = n6605 & ~n9749 ;
  assign n14176 = n8866 ^ n5821 ^ 1'b0 ;
  assign n14177 = n11549 | n14176 ;
  assign n14178 = n4739 ^ n2993 ^ n2936 ;
  assign n14179 = n6885 ^ n4708 ^ 1'b0 ;
  assign n14180 = n7161 ^ n3898 ^ 1'b0 ;
  assign n14181 = ~n4254 & n14180 ;
  assign n14182 = n8185 ^ n2436 ^ 1'b0 ;
  assign n14183 = ~n2799 & n14182 ;
  assign n14184 = n8842 & n14183 ;
  assign n14185 = n8504 & n14184 ;
  assign n14186 = ( n8725 & n13016 ) | ( n8725 & n14185 ) | ( n13016 & n14185 ) ;
  assign n14187 = n6794 & ~n6896 ;
  assign n14188 = ( ~n3265 & n5227 ) | ( ~n3265 & n12085 ) | ( n5227 & n12085 ) ;
  assign n14189 = n2653 & n14188 ;
  assign n14190 = n7999 & n14189 ;
  assign n14191 = ( ~n6589 & n9857 ) | ( ~n6589 & n14190 ) | ( n9857 & n14190 ) ;
  assign n14192 = n7846 & ~n11259 ;
  assign n14193 = n8352 ^ n6272 ^ n4251 ;
  assign n14194 = ~n2900 & n14193 ;
  assign n14195 = n1610 & ~n7447 ;
  assign n14196 = ~n7164 & n14195 ;
  assign n14197 = n8629 & ~n14196 ;
  assign n14198 = n11723 & n14197 ;
  assign n14199 = n8704 ^ n5837 ^ n3628 ;
  assign n14200 = n13978 ^ n4389 ^ 1'b0 ;
  assign n14201 = ~n11959 & n14200 ;
  assign n14202 = n11717 ^ n5122 ^ 1'b0 ;
  assign n14203 = n3412 ^ n2875 ^ 1'b0 ;
  assign n14204 = n2325 | n6682 ;
  assign n14205 = ~n2260 & n5579 ;
  assign n14206 = n4568 & n14205 ;
  assign n14207 = n9824 ^ n9371 ^ 1'b0 ;
  assign n14208 = n289 & n6642 ;
  assign n14209 = ~n14207 & n14208 ;
  assign n14210 = ~n14206 & n14209 ;
  assign n14211 = n4284 | n14210 ;
  assign n14212 = n14211 ^ n9086 ^ 1'b0 ;
  assign n14213 = n2872 | n5701 ;
  assign n14214 = n1262 & ~n2693 ;
  assign n14215 = n14214 ^ x11 ^ 1'b0 ;
  assign n14216 = ( n668 & n2589 ) | ( n668 & n14215 ) | ( n2589 & n14215 ) ;
  assign n14217 = x178 | n3297 ;
  assign n14218 = n4108 | n14217 ;
  assign n14219 = n3214 & ~n9850 ;
  assign n14220 = ~n14218 & n14219 ;
  assign n14221 = n2989 ^ n1508 ^ 1'b0 ;
  assign n14222 = n8070 & ~n14221 ;
  assign n14223 = ~n8116 & n8931 ;
  assign n14224 = ~n14222 & n14223 ;
  assign n14225 = n14224 ^ n5504 ^ 1'b0 ;
  assign n14226 = n14225 ^ n4844 ^ 1'b0 ;
  assign n14227 = n11672 & n14226 ;
  assign n14228 = n5849 & n7492 ;
  assign n14229 = n4279 & ~n13811 ;
  assign n14230 = ~n6497 & n14229 ;
  assign n14231 = n14230 ^ n12870 ^ 1'b0 ;
  assign n14232 = n5022 & n10648 ;
  assign n14236 = ( n419 & n3209 ) | ( n419 & ~n3749 ) | ( n3209 & ~n3749 ) ;
  assign n14233 = ~n6187 & n7791 ;
  assign n14234 = ~n3417 & n14233 ;
  assign n14235 = n14234 ^ n3047 ^ 1'b0 ;
  assign n14237 = n14236 ^ n14235 ^ 1'b0 ;
  assign n14238 = n13230 ^ n7271 ^ 1'b0 ;
  assign n14239 = n14237 | n14238 ;
  assign n14240 = ( ~n4004 & n4566 ) | ( ~n4004 & n11263 ) | ( n4566 & n11263 ) ;
  assign n14241 = n14240 ^ n10281 ^ n9571 ;
  assign n14242 = n14241 ^ n6660 ^ 1'b0 ;
  assign n14243 = n9853 ^ n8715 ^ 1'b0 ;
  assign n14244 = n14242 | n14243 ;
  assign n14245 = n1086 ^ x192 ^ 1'b0 ;
  assign n14246 = ~n3390 & n14245 ;
  assign n14247 = n11750 ^ n11626 ^ 1'b0 ;
  assign n14248 = n850 & ~n1244 ;
  assign n14249 = n1545 & n14248 ;
  assign n14250 = n9359 ^ n7539 ^ n1269 ;
  assign n14251 = n14249 | n14250 ;
  assign n14252 = n14251 ^ n5554 ^ 1'b0 ;
  assign n14253 = n11948 ^ x33 ^ 1'b0 ;
  assign n14254 = n9573 ^ n4752 ^ 1'b0 ;
  assign n14255 = n8513 ^ n7336 ^ 1'b0 ;
  assign n14256 = n6881 & ~n14255 ;
  assign n14257 = n14256 ^ n3105 ^ 1'b0 ;
  assign n14258 = x112 & ~n14257 ;
  assign n14259 = n1552 & ~n2343 ;
  assign n14260 = n8356 & n14104 ;
  assign n14261 = ~n14259 & n14260 ;
  assign n14262 = n6010 ^ n4757 ^ 1'b0 ;
  assign n14263 = n6842 ^ n2232 ^ 1'b0 ;
  assign n14264 = n14089 | n14263 ;
  assign n14265 = n14264 ^ n10034 ^ 1'b0 ;
  assign n14266 = n14265 ^ n7696 ^ 1'b0 ;
  assign n14267 = n14262 | n14266 ;
  assign n14268 = n2240 & n8612 ;
  assign n14269 = n14268 ^ n8745 ^ 1'b0 ;
  assign n14270 = ~n3319 & n5156 ;
  assign n14271 = ~n3973 & n11723 ;
  assign n14272 = n7379 ^ n1981 ^ 1'b0 ;
  assign n14275 = n2060 | n5688 ;
  assign n14276 = n14275 ^ n9368 ^ 1'b0 ;
  assign n14273 = n8735 ^ n7070 ^ 1'b0 ;
  assign n14274 = n6455 & n14273 ;
  assign n14277 = n14276 ^ n14274 ^ 1'b0 ;
  assign n14280 = n3509 | n9540 ;
  assign n14281 = n3147 & ~n14280 ;
  assign n14279 = n7724 | n9846 ;
  assign n14282 = n14281 ^ n14279 ^ n11185 ;
  assign n14278 = ~n7433 & n8760 ;
  assign n14283 = n14282 ^ n14278 ^ 1'b0 ;
  assign n14284 = n3957 ^ x54 ^ 1'b0 ;
  assign n14285 = ~x178 & n14284 ;
  assign n14286 = ~n3290 & n14285 ;
  assign n14287 = n14286 ^ n12197 ^ 1'b0 ;
  assign n14288 = n5221 ^ n3529 ^ 1'b0 ;
  assign n14289 = n2322 | n11458 ;
  assign n14290 = n751 | n14289 ;
  assign n14291 = n14290 ^ n8075 ^ 1'b0 ;
  assign n14292 = n8077 & n13382 ;
  assign n14293 = n2792 | n6555 ;
  assign n14294 = n14293 ^ n8781 ^ 1'b0 ;
  assign n14295 = n638 & n3782 ;
  assign n14296 = n10374 ^ n9187 ^ n1340 ;
  assign n14297 = n6825 | n14296 ;
  assign n14299 = n378 & n7160 ;
  assign n14300 = ~n12477 & n14299 ;
  assign n14298 = n13347 ^ n4335 ^ 1'b0 ;
  assign n14301 = n14300 ^ n14298 ^ n3435 ;
  assign n14302 = ~n2850 & n8740 ;
  assign n14303 = ( ~n2362 & n2598 ) | ( ~n2362 & n7819 ) | ( n2598 & n7819 ) ;
  assign n14304 = n2550 ^ n1002 ^ 1'b0 ;
  assign n14305 = ~n3217 & n9264 ;
  assign n14306 = n14304 & ~n14305 ;
  assign n14307 = x107 | n14306 ;
  assign n14308 = n8253 ^ n4410 ^ 1'b0 ;
  assign n14309 = n12956 ^ n1882 ^ 1'b0 ;
  assign n14310 = ~n9558 & n14309 ;
  assign n14311 = n4551 ^ n2448 ^ 1'b0 ;
  assign n14312 = ( n3856 & n5494 ) | ( n3856 & n14311 ) | ( n5494 & n14311 ) ;
  assign n14313 = n14312 ^ n5366 ^ 1'b0 ;
  assign n14314 = n445 & ~n1415 ;
  assign n14315 = ~n271 & n14314 ;
  assign n14316 = n671 & ~n14315 ;
  assign n14317 = n5525 & n14316 ;
  assign n14318 = ~n2020 & n14317 ;
  assign n14319 = n6360 | n11523 ;
  assign n14320 = n14319 ^ n1001 ^ 1'b0 ;
  assign n14321 = ~n4861 & n14320 ;
  assign n14322 = n2103 & ~n2297 ;
  assign n14323 = n2369 & n14322 ;
  assign n14324 = n1095 & n14323 ;
  assign n14325 = n13372 ^ n5170 ^ 1'b0 ;
  assign n14326 = n8224 ^ n5443 ^ 1'b0 ;
  assign n14327 = n12633 ^ n1813 ^ 1'b0 ;
  assign n14328 = ~n7177 & n7609 ;
  assign n14329 = n14328 ^ n3990 ^ 1'b0 ;
  assign n14330 = n14329 ^ n4476 ^ 1'b0 ;
  assign n14331 = n14222 ^ n5179 ^ 1'b0 ;
  assign n14334 = n1566 ^ n1508 ^ 1'b0 ;
  assign n14335 = n3515 | n14334 ;
  assign n14332 = n13217 ^ n12201 ^ 1'b0 ;
  assign n14333 = n11692 & ~n14332 ;
  assign n14336 = n14335 ^ n14333 ^ 1'b0 ;
  assign n14337 = n6421 ^ n1135 ^ 1'b0 ;
  assign n14338 = n8241 ^ x176 ^ 1'b0 ;
  assign n14339 = n14338 ^ n2249 ^ n694 ;
  assign n14340 = n1936 ^ n924 ^ 1'b0 ;
  assign n14341 = n6099 | n14340 ;
  assign n14342 = ( n2521 & n8755 ) | ( n2521 & n14341 ) | ( n8755 & n14341 ) ;
  assign n14344 = n1449 | n13014 ;
  assign n14345 = n14344 ^ n9363 ^ 1'b0 ;
  assign n14346 = n3198 | n14345 ;
  assign n14343 = ~n397 & n3569 ;
  assign n14347 = n14346 ^ n14343 ^ 1'b0 ;
  assign n14349 = n1742 & ~n2975 ;
  assign n14350 = ~n4465 & n14349 ;
  assign n14348 = n3928 & n8210 ;
  assign n14351 = n14350 ^ n14348 ^ 1'b0 ;
  assign n14352 = n12293 ^ n5818 ^ 1'b0 ;
  assign n14353 = n2685 ^ n1269 ^ 1'b0 ;
  assign n14354 = n14222 & n14353 ;
  assign n14355 = n14354 ^ n1579 ^ 1'b0 ;
  assign n14356 = ~n6612 & n13158 ;
  assign n14357 = n5242 & n14356 ;
  assign n14358 = n825 & ~n13263 ;
  assign n14359 = ( n497 & ~n5197 ) | ( n497 & n13708 ) | ( ~n5197 & n13708 ) ;
  assign n14360 = n14359 ^ n14067 ^ 1'b0 ;
  assign n14361 = n14360 ^ n9665 ^ 1'b0 ;
  assign n14362 = n8958 ^ n4238 ^ 1'b0 ;
  assign n14363 = n3646 & n14362 ;
  assign n14364 = n14363 ^ n13878 ^ n5812 ;
  assign n14365 = n14020 | n14364 ;
  assign n14366 = n2085 & ~n14365 ;
  assign n14367 = n2846 & ~n3627 ;
  assign n14368 = ~n3180 & n5626 ;
  assign n14369 = ~n7547 & n14368 ;
  assign n14370 = n545 & ~n14369 ;
  assign n14371 = ~n14367 & n14370 ;
  assign n14372 = n842 | n9271 ;
  assign n14373 = n12509 | n14372 ;
  assign n14374 = n1247 & n2394 ;
  assign n14375 = n9147 ^ n2467 ^ 1'b0 ;
  assign n14376 = n14375 ^ n6701 ^ 1'b0 ;
  assign n14377 = n6391 & ~n13680 ;
  assign n14378 = n6190 ^ n1165 ^ 1'b0 ;
  assign n14379 = n2208 & n14378 ;
  assign n14380 = ( n5043 & ~n7224 ) | ( n5043 & n14379 ) | ( ~n7224 & n14379 ) ;
  assign n14381 = ~n389 & n14380 ;
  assign n14382 = x61 & n4619 ;
  assign n14383 = n14382 ^ n3959 ^ 1'b0 ;
  assign n14384 = n14383 ^ n7848 ^ n2974 ;
  assign n14385 = n14381 & n14384 ;
  assign n14386 = ~n14381 & n14385 ;
  assign n14387 = n14386 ^ n11581 ^ n11529 ;
  assign n14390 = n4315 & n11563 ;
  assign n14391 = n14390 ^ n869 ^ 1'b0 ;
  assign n14388 = ~n1858 & n4368 ;
  assign n14389 = n5895 & n14388 ;
  assign n14392 = n14391 ^ n14389 ^ 1'b0 ;
  assign n14393 = n4479 & ~n5619 ;
  assign n14394 = ~n1796 & n14393 ;
  assign n14395 = n11031 | n14394 ;
  assign n14396 = n14392 | n14395 ;
  assign n14397 = ~n4055 & n9806 ;
  assign n14398 = ~n385 & n14397 ;
  assign n14399 = n14398 ^ n13692 ^ 1'b0 ;
  assign n14400 = n4635 & n8730 ;
  assign n14401 = n14400 ^ n2472 ^ 1'b0 ;
  assign n14402 = n14401 ^ n14015 ^ n8365 ;
  assign n14403 = ~n12578 & n14402 ;
  assign n14404 = n14403 ^ n2940 ^ 1'b0 ;
  assign n14405 = n3951 & n10527 ;
  assign n14406 = n7496 ^ n4273 ^ 1'b0 ;
  assign n14407 = n794 & n1734 ;
  assign n14408 = n14407 ^ n6450 ^ 1'b0 ;
  assign n14409 = n6058 & ~n6465 ;
  assign n14410 = n14409 ^ n1118 ^ 1'b0 ;
  assign n14413 = n2736 & ~n5769 ;
  assign n14414 = n14413 ^ n2615 ^ 1'b0 ;
  assign n14411 = n1338 & ~n2143 ;
  assign n14412 = ~x175 & n14411 ;
  assign n14415 = n14414 ^ n14412 ^ n3967 ;
  assign n14416 = n4673 | n5268 ;
  assign n14417 = n5005 & n14416 ;
  assign n14418 = ~n7199 & n9086 ;
  assign n14419 = n7583 & n14418 ;
  assign n14420 = n4107 & ~n5873 ;
  assign n14421 = ~n2785 & n4666 ;
  assign n14422 = n11416 & n14421 ;
  assign n14423 = ~n14420 & n14422 ;
  assign n14424 = n708 & n14423 ;
  assign n14425 = n8745 ^ n7294 ^ 1'b0 ;
  assign n14426 = n14425 ^ n6429 ^ 1'b0 ;
  assign n14427 = n12131 | n14426 ;
  assign n14428 = n11394 & ~n14427 ;
  assign n14429 = ( n9495 & ~n10016 ) | ( n9495 & n12044 ) | ( ~n10016 & n12044 ) ;
  assign n14430 = n14429 ^ n3926 ^ 1'b0 ;
  assign n14431 = n11956 ^ n2135 ^ 1'b0 ;
  assign n14432 = x17 & ~n1667 ;
  assign n14433 = ~n6424 & n14432 ;
  assign n14434 = ( n1611 & n11519 ) | ( n1611 & n14433 ) | ( n11519 & n14433 ) ;
  assign n14435 = n6400 ^ n346 ^ 1'b0 ;
  assign n14436 = n14434 & ~n14435 ;
  assign n14437 = ~n4545 & n9835 ;
  assign n14438 = n9093 & ~n14437 ;
  assign n14439 = n6921 ^ n889 ^ 1'b0 ;
  assign n14440 = x113 & n14439 ;
  assign n14441 = n14440 ^ n2281 ^ 1'b0 ;
  assign n14442 = n14438 | n14441 ;
  assign n14443 = n14436 & ~n14442 ;
  assign n14444 = ~n529 & n14443 ;
  assign n14445 = n12253 ^ n882 ^ 1'b0 ;
  assign n14446 = n2308 & n3796 ;
  assign n14447 = ~n10676 & n14446 ;
  assign n14448 = ( x82 & ~n3233 ) | ( x82 & n4269 ) | ( ~n3233 & n4269 ) ;
  assign n14449 = n1440 | n14448 ;
  assign n14450 = ~n11336 & n13372 ;
  assign n14451 = n9447 & n14450 ;
  assign n14452 = n2900 & n11038 ;
  assign n14453 = n14451 & n14452 ;
  assign n14454 = n1680 | n4908 ;
  assign n14455 = n14454 ^ n3157 ^ 1'b0 ;
  assign n14456 = n14455 ^ n558 ^ 1'b0 ;
  assign n14457 = n9026 ^ n3030 ^ 1'b0 ;
  assign n14458 = n1295 | n3656 ;
  assign n14459 = n14457 & n14458 ;
  assign n14460 = n3823 & n5605 ;
  assign n14462 = n1929 & n9536 ;
  assign n14461 = n7611 & ~n9292 ;
  assign n14463 = n14462 ^ n14461 ^ 1'b0 ;
  assign n14464 = ( n9014 & ~n9511 ) | ( n9014 & n14463 ) | ( ~n9511 & n14463 ) ;
  assign n14465 = n14071 ^ n7858 ^ 1'b0 ;
  assign n14466 = n11503 | n14465 ;
  assign n14467 = n8414 & ~n14466 ;
  assign n14468 = ~n3593 & n14467 ;
  assign n14469 = n14468 ^ n12411 ^ n591 ;
  assign n14470 = n11360 ^ x159 ^ 1'b0 ;
  assign n14471 = n5036 & n8841 ;
  assign n14472 = n14471 ^ n2942 ^ 1'b0 ;
  assign n14473 = ~n14470 & n14472 ;
  assign n14474 = n3030 | n4067 ;
  assign n14475 = n10271 & ~n14474 ;
  assign n14476 = n4056 & n12124 ;
  assign n14477 = n891 & ~n14476 ;
  assign n14478 = n14477 ^ n13476 ^ 1'b0 ;
  assign n14479 = n722 & n14478 ;
  assign n14480 = ~n1208 & n4288 ;
  assign n14481 = n6928 ^ n4793 ^ n3530 ;
  assign n14482 = n9649 ^ n3420 ^ 1'b0 ;
  assign n14483 = n6554 | n14482 ;
  assign n14484 = n14145 ^ n10713 ^ n9587 ;
  assign n14485 = n1839 & ~n9839 ;
  assign n14486 = x163 & n14485 ;
  assign n14487 = n14486 ^ n8928 ^ 1'b0 ;
  assign n14488 = n7053 ^ n2850 ^ n1979 ;
  assign n14489 = ~n3923 & n14488 ;
  assign n14490 = n2970 & n14489 ;
  assign n14491 = ( ~n4937 & n6073 ) | ( ~n4937 & n6080 ) | ( n6073 & n6080 ) ;
  assign n14492 = n12702 | n14491 ;
  assign n14493 = n13729 & n14492 ;
  assign n14494 = n10770 | n11130 ;
  assign n14495 = n2739 & n3666 ;
  assign n14496 = n14495 ^ n2748 ^ 1'b0 ;
  assign n14497 = n14496 ^ n5232 ^ 1'b0 ;
  assign n14498 = n2178 | n12212 ;
  assign n14499 = n14498 ^ n831 ^ 1'b0 ;
  assign n14500 = n6727 | n14499 ;
  assign n14501 = n11070 ^ n1606 ^ 1'b0 ;
  assign n14503 = ~n5839 & n7987 ;
  assign n14504 = n14503 ^ n5799 ^ 1'b0 ;
  assign n14502 = ~n10814 & n14025 ;
  assign n14505 = n14504 ^ n14502 ^ 1'b0 ;
  assign n14509 = ( ~n716 & n1884 ) | ( ~n716 & n4676 ) | ( n1884 & n4676 ) ;
  assign n14506 = ~n2061 & n3704 ;
  assign n14507 = ~n896 & n14506 ;
  assign n14508 = n4896 | n14507 ;
  assign n14510 = n14509 ^ n14508 ^ 1'b0 ;
  assign n14511 = n7193 ^ n1295 ^ 1'b0 ;
  assign n14512 = ~n874 & n1039 ;
  assign n14513 = n14512 ^ n7135 ^ 1'b0 ;
  assign n14514 = n6793 ^ n6276 ^ 1'b0 ;
  assign n14515 = n2357 | n5269 ;
  assign n14516 = n14514 & ~n14515 ;
  assign n14517 = n2051 & ~n14516 ;
  assign n14518 = n2489 & n14517 ;
  assign n14519 = n10931 ^ n8639 ^ 1'b0 ;
  assign n14520 = n501 & n5557 ;
  assign n14521 = n4282 & n14520 ;
  assign n14522 = n14521 ^ n6943 ^ 1'b0 ;
  assign n14523 = n9531 ^ n6698 ^ 1'b0 ;
  assign n14524 = n9495 ^ n2792 ^ 1'b0 ;
  assign n14525 = n3704 & n14524 ;
  assign n14526 = n1376 & n5047 ;
  assign n14527 = n14526 ^ n7667 ^ 1'b0 ;
  assign n14528 = n7914 & n14527 ;
  assign n14529 = n14528 ^ n13718 ^ 1'b0 ;
  assign n14531 = n3168 ^ n1894 ^ 1'b0 ;
  assign n14530 = ~n1797 & n2309 ;
  assign n14532 = n14531 ^ n14530 ^ 1'b0 ;
  assign n14533 = n7670 ^ n4614 ^ 1'b0 ;
  assign n14534 = n14533 ^ n10196 ^ 1'b0 ;
  assign n14535 = n10316 | n12079 ;
  assign n14536 = n8531 ^ n6166 ^ 1'b0 ;
  assign n14537 = n3838 & ~n11452 ;
  assign n14538 = n4872 & ~n9404 ;
  assign n14539 = n14538 ^ n8276 ^ n5965 ;
  assign n14540 = n9694 & n10596 ;
  assign n14541 = n8911 | n9373 ;
  assign n14542 = n14541 ^ x251 ^ 1'b0 ;
  assign n14543 = n14540 & n14542 ;
  assign n14544 = n7304 & n7353 ;
  assign n14545 = x216 & ~n2988 ;
  assign n14546 = ~n668 & n14545 ;
  assign n14547 = n4988 & n14546 ;
  assign n14548 = n2267 | n14547 ;
  assign n14549 = n535 | n14548 ;
  assign n14550 = n2891 ^ n331 ^ 1'b0 ;
  assign n14551 = n2047 | n14550 ;
  assign n14552 = n6883 ^ n1471 ^ 1'b0 ;
  assign n14553 = n2580 & ~n14552 ;
  assign n14554 = n14553 ^ n4439 ^ 1'b0 ;
  assign n14555 = n8962 | n14554 ;
  assign n14556 = n2627 & ~n4437 ;
  assign n14557 = n6020 ^ n4248 ^ n1070 ;
  assign n14563 = n6199 & ~n7626 ;
  assign n14564 = n5034 | n14563 ;
  assign n14565 = n10430 & ~n14564 ;
  assign n14566 = ~n2919 & n11881 ;
  assign n14567 = n14566 ^ x249 ^ 1'b0 ;
  assign n14568 = ( n485 & n1968 ) | ( n485 & ~n2070 ) | ( n1968 & ~n2070 ) ;
  assign n14569 = ( ~n11041 & n12007 ) | ( ~n11041 & n14568 ) | ( n12007 & n14568 ) ;
  assign n14570 = n14569 ^ n12638 ^ 1'b0 ;
  assign n14571 = n14567 & n14570 ;
  assign n14572 = ( n1534 & n5392 ) | ( n1534 & ~n8088 ) | ( n5392 & ~n8088 ) ;
  assign n14573 = n14572 ^ n10532 ^ n6644 ;
  assign n14574 = n14571 & ~n14573 ;
  assign n14575 = n14565 & n14574 ;
  assign n14561 = n1506 | n2562 ;
  assign n14562 = n14561 ^ n2584 ^ 1'b0 ;
  assign n14558 = n2900 | n5316 ;
  assign n14559 = ~n2323 & n14558 ;
  assign n14560 = n7421 & n14559 ;
  assign n14576 = n14575 ^ n14562 ^ n14560 ;
  assign n14577 = n1064 & ~n11612 ;
  assign n14578 = n1109 & n14577 ;
  assign n14579 = n14578 ^ n11680 ^ 1'b0 ;
  assign n14580 = n9357 & ~n14579 ;
  assign n14581 = n2051 | n4130 ;
  assign n14582 = n1379 | n14581 ;
  assign n14583 = n3871 & n14582 ;
  assign n14584 = n14583 ^ n5138 ^ 1'b0 ;
  assign n14585 = n7586 ^ n1647 ^ 1'b0 ;
  assign n14586 = ~n14584 & n14585 ;
  assign n14587 = n8490 & n14586 ;
  assign n14588 = ~n14580 & n14587 ;
  assign n14589 = n1841 & ~n5325 ;
  assign n14590 = n14589 ^ n3882 ^ 1'b0 ;
  assign n14591 = x100 | n14590 ;
  assign n14592 = n3710 & n9299 ;
  assign n14593 = n14591 & n14592 ;
  assign n14597 = n14090 ^ n6202 ^ 1'b0 ;
  assign n14594 = n4747 & ~n11643 ;
  assign n14595 = ~x248 & n14594 ;
  assign n14596 = n14595 ^ n12132 ^ 1'b0 ;
  assign n14598 = n14597 ^ n14596 ^ n12852 ;
  assign n14599 = n3022 ^ n1695 ^ n1315 ;
  assign n14600 = ~n2790 & n4470 ;
  assign n14601 = ~n1343 & n14600 ;
  assign n14602 = n1349 | n2286 ;
  assign n14603 = n14602 ^ n3596 ^ 1'b0 ;
  assign n14604 = ~n3961 & n14603 ;
  assign n14605 = n14601 & n14604 ;
  assign n14606 = n14599 & n14605 ;
  assign n14607 = n11735 ^ n8260 ^ 1'b0 ;
  assign n14608 = ( n9383 & n10072 ) | ( n9383 & n13575 ) | ( n10072 & n13575 ) ;
  assign n14609 = n14608 ^ n8052 ^ 1'b0 ;
  assign n14610 = ( n516 & n2949 ) | ( n516 & ~n6038 ) | ( n2949 & ~n6038 ) ;
  assign n14611 = n11902 | n14610 ;
  assign n14612 = n790 & ~n14611 ;
  assign n14613 = ( n4407 & ~n9735 ) | ( n4407 & n13807 ) | ( ~n9735 & n13807 ) ;
  assign n14614 = ~n3904 & n7856 ;
  assign n14615 = n14614 ^ n12783 ^ 1'b0 ;
  assign n14616 = n9557 & n14615 ;
  assign n14617 = n1519 & n2511 ;
  assign n14618 = n5231 | n13851 ;
  assign n14619 = n1744 | n1775 ;
  assign n14620 = x64 & n14619 ;
  assign n14622 = n4069 ^ n615 ^ n562 ;
  assign n14621 = n4244 & ~n11446 ;
  assign n14623 = n14622 ^ n14621 ^ 1'b0 ;
  assign n14624 = n3772 ^ n3595 ^ 1'b0 ;
  assign n14625 = ~n778 & n14624 ;
  assign n14626 = n14623 | n14625 ;
  assign n14627 = n6319 ^ n3028 ^ 1'b0 ;
  assign n14628 = n14396 | n14627 ;
  assign n14629 = ~n4970 & n5890 ;
  assign n14630 = n14629 ^ n13694 ^ 1'b0 ;
  assign n14631 = n14630 ^ n7101 ^ 1'b0 ;
  assign n14632 = n5625 ^ n3637 ^ 1'b0 ;
  assign n14633 = n5179 ^ n3659 ^ 1'b0 ;
  assign n14634 = x57 & n14633 ;
  assign n14635 = n4610 & n14634 ;
  assign n14639 = n7855 ^ n3539 ^ 1'b0 ;
  assign n14636 = n12415 ^ n5150 ^ 1'b0 ;
  assign n14637 = n10805 & ~n14636 ;
  assign n14638 = ~n7177 & n14637 ;
  assign n14640 = n14639 ^ n14638 ^ 1'b0 ;
  assign n14641 = n4432 & ~n14640 ;
  assign n14642 = ( n1465 & ~n10407 ) | ( n1465 & n14641 ) | ( ~n10407 & n14641 ) ;
  assign n14643 = n7757 ^ n3980 ^ 1'b0 ;
  assign n14644 = n7581 & ~n14643 ;
  assign n14645 = n14249 ^ n4115 ^ 1'b0 ;
  assign n14646 = ~n4869 & n14645 ;
  assign n14647 = n14646 ^ n4394 ^ 1'b0 ;
  assign n14648 = n2141 ^ n389 ^ 1'b0 ;
  assign n14649 = n3198 | n14648 ;
  assign n14650 = n1615 & n4597 ;
  assign n14651 = n11818 & n14650 ;
  assign n14652 = ~x211 & n2198 ;
  assign n14653 = ( n6604 & n10695 ) | ( n6604 & ~n14652 ) | ( n10695 & ~n14652 ) ;
  assign n14654 = n5130 ^ n1129 ^ 1'b0 ;
  assign n14655 = ~n14653 & n14654 ;
  assign n14656 = ~n3494 & n14516 ;
  assign n14657 = n1562 | n3037 ;
  assign n14658 = n451 | n14657 ;
  assign n14659 = ~n3843 & n14658 ;
  assign n14660 = ~n4900 & n14659 ;
  assign n14661 = ( n742 & n6640 ) | ( n742 & ~n7794 ) | ( n6640 & ~n7794 ) ;
  assign n14662 = n12852 ^ n9710 ^ n8241 ;
  assign n14663 = ~n7041 & n12874 ;
  assign n14664 = n14662 | n14663 ;
  assign n14665 = n3863 ^ n555 ^ 1'b0 ;
  assign n14666 = n12281 & ~n14665 ;
  assign n14667 = n7188 ^ n1099 ^ n737 ;
  assign n14668 = n8070 & ~n14667 ;
  assign n14669 = ~n14666 & n14668 ;
  assign n14670 = n4559 | n9862 ;
  assign n14671 = n2112 & ~n14670 ;
  assign n14672 = n14671 ^ n4227 ^ 1'b0 ;
  assign n14673 = ~n14669 & n14672 ;
  assign n14674 = n8512 ^ n2865 ^ n547 ;
  assign n14675 = n14674 ^ n8167 ^ 1'b0 ;
  assign n14676 = n3564 & ~n9291 ;
  assign n14677 = n14676 ^ n581 ^ 1'b0 ;
  assign n14678 = n14025 ^ n3825 ^ 1'b0 ;
  assign n14679 = n14677 | n14678 ;
  assign n14681 = ~n2730 & n13306 ;
  assign n14680 = ~n4165 & n9109 ;
  assign n14682 = n14681 ^ n14680 ^ 1'b0 ;
  assign n14683 = n1638 & ~n1968 ;
  assign n14684 = n1968 & n14683 ;
  assign n14685 = n5704 & ~n14684 ;
  assign n14686 = n7663 & ~n13423 ;
  assign n14687 = n14685 & n14686 ;
  assign n14688 = ( n1994 & ~n2018 ) | ( n1994 & n5497 ) | ( ~n2018 & n5497 ) ;
  assign n14689 = n1562 | n1654 ;
  assign n14690 = n4924 & ~n14689 ;
  assign n14691 = n14690 ^ n3458 ^ 1'b0 ;
  assign n14692 = n2978 & ~n14691 ;
  assign n14693 = n3922 ^ x100 ^ 1'b0 ;
  assign n14694 = ~n6803 & n12792 ;
  assign n14695 = n14693 & n14694 ;
  assign n14696 = n12574 ^ n2940 ^ 1'b0 ;
  assign n14697 = x237 & ~n5296 ;
  assign n14698 = n8564 | n10284 ;
  assign n14699 = n11496 ^ n11109 ^ 1'b0 ;
  assign n14702 = n5528 ^ n3646 ^ 1'b0 ;
  assign n14703 = n1915 & n14702 ;
  assign n14704 = n14703 ^ n10517 ^ 1'b0 ;
  assign n14705 = n13785 & ~n14704 ;
  assign n14700 = n8670 ^ n5412 ^ 1'b0 ;
  assign n14701 = ~n1718 & n14700 ;
  assign n14706 = n14705 ^ n14701 ^ n13693 ;
  assign n14707 = n10518 | n11531 ;
  assign n14708 = n10268 | n14707 ;
  assign n14709 = n1065 | n3805 ;
  assign n14710 = n1848 | n14709 ;
  assign n14711 = n9429 | n14710 ;
  assign n14715 = n8545 ^ n1382 ^ 1'b0 ;
  assign n14713 = ( ~n634 & n973 ) | ( ~n634 & n1867 ) | ( n973 & n1867 ) ;
  assign n14712 = n2532 & n9014 ;
  assign n14714 = n14713 ^ n14712 ^ 1'b0 ;
  assign n14716 = n14715 ^ n14714 ^ n8647 ;
  assign n14717 = n14716 ^ n2785 ^ 1'b0 ;
  assign n14718 = n7925 & ~n13796 ;
  assign n14719 = ~n14717 & n14718 ;
  assign n14720 = n4065 | n14614 ;
  assign n14721 = x115 & ~n3685 ;
  assign n14722 = n2804 & n14721 ;
  assign n14723 = ~n3256 & n3478 ;
  assign n14724 = n7251 ^ n4559 ^ 1'b0 ;
  assign n14725 = n14455 & n14724 ;
  assign n14726 = n14725 ^ n13496 ^ 1'b0 ;
  assign n14727 = n14723 | n14726 ;
  assign n14728 = ~n1933 & n6713 ;
  assign n14729 = n3462 & n14728 ;
  assign n14730 = n14729 ^ n7029 ^ 1'b0 ;
  assign n14731 = x213 & n14730 ;
  assign n14732 = n14727 & n14731 ;
  assign n14733 = n12115 ^ n5448 ^ 1'b0 ;
  assign n14734 = ~n11277 & n14733 ;
  assign n14735 = n14734 ^ n13840 ^ 1'b0 ;
  assign n14739 = n7113 ^ n419 ^ 1'b0 ;
  assign n14736 = n2428 & ~n3444 ;
  assign n14737 = n8072 | n9747 ;
  assign n14738 = n14736 | n14737 ;
  assign n14740 = n14739 ^ n14738 ^ 1'b0 ;
  assign n14741 = n7092 | n9920 ;
  assign n14742 = n5515 ^ n3806 ^ 1'b0 ;
  assign n14743 = n14742 ^ n10493 ^ 1'b0 ;
  assign n14744 = ~n11630 & n14743 ;
  assign n14745 = n1409 & n5671 ;
  assign n14746 = ~n9842 & n12222 ;
  assign n14747 = n14746 ^ n5578 ^ 1'b0 ;
  assign n14748 = n14160 ^ n12441 ^ 1'b0 ;
  assign n14749 = ~n14747 & n14748 ;
  assign n14750 = ~n4497 & n5455 ;
  assign n14751 = ~n779 & n3829 ;
  assign n14752 = n14751 ^ n830 ^ 1'b0 ;
  assign n14754 = n7201 ^ n6088 ^ 1'b0 ;
  assign n14753 = ~n2514 & n3769 ;
  assign n14755 = n14754 ^ n14753 ^ 1'b0 ;
  assign n14756 = n2049 & ~n10282 ;
  assign n14757 = ( n2335 & ~n14755 ) | ( n2335 & n14756 ) | ( ~n14755 & n14756 ) ;
  assign n14758 = n666 & n3576 ;
  assign n14759 = n14758 ^ n9662 ^ 1'b0 ;
  assign n14760 = n14757 & ~n14759 ;
  assign n14761 = n537 & ~n5315 ;
  assign n14762 = ~n3323 & n14761 ;
  assign n14763 = n1971 | n14762 ;
  assign n14765 = n3166 ^ n2431 ^ 1'b0 ;
  assign n14766 = ~n1306 & n14765 ;
  assign n14767 = ~n688 & n14766 ;
  assign n14768 = n834 | n14767 ;
  assign n14769 = n14768 ^ n9243 ^ 1'b0 ;
  assign n14764 = n6242 & n7349 ;
  assign n14770 = n14769 ^ n14764 ^ 1'b0 ;
  assign n14771 = n4919 & ~n14358 ;
  assign n14772 = n6661 & n8358 ;
  assign n14773 = x208 & n4964 ;
  assign n14774 = n14773 ^ n5973 ^ 1'b0 ;
  assign n14775 = n4295 ^ n3102 ^ 1'b0 ;
  assign n14776 = n328 & n6358 ;
  assign n14777 = n14776 ^ n3039 ^ 1'b0 ;
  assign n14778 = n14777 ^ n5839 ^ 1'b0 ;
  assign n14779 = n2644 & ~n14778 ;
  assign n14780 = n3856 & n14779 ;
  assign n14781 = n10069 & n14780 ;
  assign n14782 = n14781 ^ n3838 ^ 1'b0 ;
  assign n14783 = ~n14775 & n14782 ;
  assign n14784 = n14783 ^ n11492 ^ 1'b0 ;
  assign n14785 = n10207 & n12824 ;
  assign n14786 = n11351 & n12477 ;
  assign n14787 = n14786 ^ n8094 ^ 1'b0 ;
  assign n14788 = n1553 & n14787 ;
  assign n14791 = ~n2933 & n9296 ;
  assign n14792 = ~n5173 & n14791 ;
  assign n14789 = x159 & n2499 ;
  assign n14790 = x209 & n14789 ;
  assign n14793 = n14792 ^ n14790 ^ 1'b0 ;
  assign n14794 = n466 | n14793 ;
  assign n14795 = ~n14788 & n14794 ;
  assign n14796 = n14795 ^ n3255 ^ 1'b0 ;
  assign n14797 = n622 & n3323 ;
  assign n14798 = n14007 & n14797 ;
  assign n14799 = n14798 ^ n13143 ^ 1'b0 ;
  assign n14800 = n8103 ^ n6370 ^ 1'b0 ;
  assign n14801 = n14800 ^ n12260 ^ n389 ;
  assign n14802 = ~n1279 & n2812 ;
  assign n14803 = n1750 & n14802 ;
  assign n14804 = n11833 & ~n14803 ;
  assign n14805 = n14804 ^ n10484 ^ 1'b0 ;
  assign n14806 = ~n1557 & n14805 ;
  assign n14807 = n8724 & n14806 ;
  assign n14808 = n5031 | n11872 ;
  assign n14809 = n2366 | n3717 ;
  assign n14810 = n14809 ^ n8709 ^ 1'b0 ;
  assign n14811 = ~n3814 & n14810 ;
  assign n14812 = n14811 ^ n5576 ^ 1'b0 ;
  assign n14813 = n14812 ^ n5943 ^ 1'b0 ;
  assign n14814 = ~n11549 & n14813 ;
  assign n14815 = ~n5525 & n7681 ;
  assign n14816 = n14815 ^ n12058 ^ 1'b0 ;
  assign n14817 = n8341 & ~n14816 ;
  assign n14818 = n14817 ^ n2710 ^ 1'b0 ;
  assign n14819 = ~n1636 & n9744 ;
  assign n14820 = n14819 ^ n4267 ^ 1'b0 ;
  assign n14821 = n2554 | n11496 ;
  assign n14822 = n14821 ^ n9971 ^ 1'b0 ;
  assign n14823 = x12 & n14822 ;
  assign n14824 = n13748 ^ n5948 ^ n2245 ;
  assign n14825 = ~n12375 & n14824 ;
  assign n14826 = ~n6268 & n14825 ;
  assign n14827 = n10864 & n14826 ;
  assign n14828 = ~n3985 & n12575 ;
  assign n14829 = ~n2349 & n14828 ;
  assign n14830 = ( n1450 & ~n5197 ) | ( n1450 & n9310 ) | ( ~n5197 & n9310 ) ;
  assign n14831 = n14830 ^ n10596 ^ 1'b0 ;
  assign n14832 = n9619 ^ n5794 ^ n3392 ;
  assign n14833 = ~n14831 & n14832 ;
  assign n14834 = n4200 & n14833 ;
  assign n14835 = n14829 | n14834 ;
  assign n14836 = n14835 ^ x252 ^ 1'b0 ;
  assign n14837 = n3404 & n6781 ;
  assign n14838 = n14837 ^ n2829 ^ 1'b0 ;
  assign n14839 = n10126 & n14838 ;
  assign n14840 = n446 | n2219 ;
  assign n14841 = n14840 ^ x227 ^ 1'b0 ;
  assign n14842 = n4033 & n14841 ;
  assign n14843 = n8473 ^ n894 ^ 1'b0 ;
  assign n14844 = ~n14842 & n14843 ;
  assign n14845 = n14844 ^ n12758 ^ n7853 ;
  assign n14846 = n10885 & ~n14845 ;
  assign n14847 = ( ~n6750 & n7807 ) | ( ~n6750 & n14846 ) | ( n7807 & n14846 ) ;
  assign n14848 = n13073 ^ n4610 ^ 1'b0 ;
  assign n14849 = n2939 | n14848 ;
  assign n14850 = n14849 ^ n3747 ^ 1'b0 ;
  assign n14851 = n12372 | n14850 ;
  assign n14852 = n13080 | n14851 ;
  assign n14853 = n4830 & n11167 ;
  assign n14854 = n14853 ^ n7961 ^ 1'b0 ;
  assign n14855 = ( n1832 & n11403 ) | ( n1832 & n13271 ) | ( n11403 & n13271 ) ;
  assign n14856 = n5122 ^ n2258 ^ 1'b0 ;
  assign n14857 = n14856 ^ n4407 ^ 1'b0 ;
  assign n14858 = n6121 & ~n13809 ;
  assign n14859 = ~n3094 & n14858 ;
  assign n14860 = n6546 & n12862 ;
  assign n14861 = n9248 & n14860 ;
  assign n14862 = n5616 & ~n7941 ;
  assign n14863 = n5497 & n14862 ;
  assign n14864 = n14863 ^ n10586 ^ 1'b0 ;
  assign n14865 = n5181 ^ n2494 ^ 1'b0 ;
  assign n14866 = n5983 & n14865 ;
  assign n14869 = ( ~n5625 & n9540 ) | ( ~n5625 & n14218 ) | ( n9540 & n14218 ) ;
  assign n14867 = n1045 & ~n3542 ;
  assign n14868 = n5201 | n14867 ;
  assign n14870 = n14869 ^ n14868 ^ 1'b0 ;
  assign n14871 = n2936 & ~n5756 ;
  assign n14872 = ~n10070 & n14871 ;
  assign n14873 = ~n2579 & n3171 ;
  assign n14874 = ( n1170 & n8474 ) | ( n1170 & n14873 ) | ( n8474 & n14873 ) ;
  assign n14875 = n7444 ^ n5667 ^ 1'b0 ;
  assign n14876 = n4905 ^ n2258 ^ 1'b0 ;
  assign n14877 = n5364 & ~n14876 ;
  assign n14878 = ( n3230 & ~n4699 ) | ( n3230 & n6726 ) | ( ~n4699 & n6726 ) ;
  assign n14879 = n6261 ^ n449 ^ 1'b0 ;
  assign n14880 = n12819 & n14879 ;
  assign n14881 = n14878 & n14880 ;
  assign n14882 = n13646 ^ n1832 ^ 1'b0 ;
  assign n14883 = x213 & n14882 ;
  assign n14884 = ~n12815 & n14883 ;
  assign n14885 = n14881 & n14884 ;
  assign n14886 = n2966 ^ n1416 ^ 1'b0 ;
  assign n14887 = n5528 ^ n585 ^ 1'b0 ;
  assign n14888 = ~n3286 & n14887 ;
  assign n14889 = n14888 ^ n3221 ^ 1'b0 ;
  assign n14890 = ~n4302 & n4554 ;
  assign n14891 = n14890 ^ n8311 ^ 1'b0 ;
  assign n14892 = n10390 & ~n14885 ;
  assign n14893 = ~n5739 & n7737 ;
  assign n14894 = ~n8113 & n14893 ;
  assign n14895 = n3146 & ~n14894 ;
  assign n14896 = n3320 & n14895 ;
  assign n14897 = n14896 ^ n5003 ^ 1'b0 ;
  assign n14898 = ~n14608 & n14620 ;
  assign n14899 = n3115 & n3942 ;
  assign n14900 = n14899 ^ n4518 ^ 1'b0 ;
  assign n14901 = n1867 | n6902 ;
  assign n14902 = n14901 ^ n4703 ^ 1'b0 ;
  assign n14904 = n3114 & n5596 ;
  assign n14905 = n14904 ^ n3335 ^ 1'b0 ;
  assign n14903 = n858 & n10426 ;
  assign n14906 = n14905 ^ n14903 ^ 1'b0 ;
  assign n14908 = n1950 ^ n1142 ^ 1'b0 ;
  assign n14907 = ~n9973 & n11843 ;
  assign n14909 = n14908 ^ n14907 ^ 1'b0 ;
  assign n14910 = ~n2725 & n14560 ;
  assign n14911 = ~n3689 & n14910 ;
  assign n14912 = n6333 ^ n1486 ^ 1'b0 ;
  assign n14913 = n14912 ^ n2714 ^ 1'b0 ;
  assign n14914 = n8838 & ~n11154 ;
  assign n14915 = ~n12124 & n14914 ;
  assign n14916 = n14915 ^ n274 ^ 1'b0 ;
  assign n14917 = n8770 ^ n2544 ^ 1'b0 ;
  assign n14918 = n1045 & ~n14917 ;
  assign n14919 = ( n5018 & n7941 ) | ( n5018 & ~n10208 ) | ( n7941 & ~n10208 ) ;
  assign n14920 = n7939 & ~n14919 ;
  assign n14921 = n10545 & n14920 ;
  assign n14922 = n2284 & n2617 ;
  assign n14925 = n5977 ^ n1125 ^ 1'b0 ;
  assign n14926 = n4374 | n14925 ;
  assign n14923 = n7392 ^ x92 ^ 1'b0 ;
  assign n14924 = ~n2122 & n14923 ;
  assign n14927 = n14926 ^ n14924 ^ 1'b0 ;
  assign n14928 = n13442 ^ n1112 ^ 1'b0 ;
  assign n14929 = n5395 & ~n14928 ;
  assign n14930 = n2002 & ~n9067 ;
  assign n14931 = n14929 & n14930 ;
  assign n14932 = n4226 & n14931 ;
  assign n14933 = ~n473 & n14471 ;
  assign n14934 = n6524 | n10290 ;
  assign n14935 = n14000 & ~n14934 ;
  assign n14936 = ( n1475 & n3412 ) | ( n1475 & ~n4088 ) | ( n3412 & ~n4088 ) ;
  assign n14937 = n3154 & ~n14936 ;
  assign n14938 = n1078 | n14937 ;
  assign n14939 = n6369 & ~n14938 ;
  assign n14940 = n3307 | n14939 ;
  assign n14941 = n1473 | n14940 ;
  assign n14942 = ~n2883 & n10349 ;
  assign n14943 = n3032 & n14942 ;
  assign n14944 = n2797 | n14943 ;
  assign n14945 = n535 | n14944 ;
  assign n14946 = n1449 & ~n14945 ;
  assign n14947 = n14256 ^ n6850 ^ 1'b0 ;
  assign n14948 = ( n3706 & n6727 ) | ( n3706 & ~n14947 ) | ( n6727 & ~n14947 ) ;
  assign n14949 = n4511 ^ x195 ^ 1'b0 ;
  assign n14950 = ~n7838 & n14949 ;
  assign n14951 = n2542 & ~n4668 ;
  assign n14952 = n7968 & n14951 ;
  assign n14953 = n13538 & ~n14952 ;
  assign n14954 = n13472 & n14953 ;
  assign n14955 = n5698 & ~n11257 ;
  assign n14956 = n14955 ^ n4793 ^ 1'b0 ;
  assign n14957 = ~n4299 & n5961 ;
  assign n14958 = n9630 | n14957 ;
  assign n14959 = ~n4067 & n7097 ;
  assign n14960 = ~n7256 & n14959 ;
  assign n14961 = n14960 ^ n916 ^ 1'b0 ;
  assign n14962 = ( ~n10776 & n11130 ) | ( ~n10776 & n14961 ) | ( n11130 & n14961 ) ;
  assign n14963 = n14962 ^ n11777 ^ 1'b0 ;
  assign n14964 = n13023 ^ n2972 ^ n1373 ;
  assign n14965 = ( x207 & ~n3082 ) | ( x207 & n14964 ) | ( ~n3082 & n14964 ) ;
  assign n14966 = ~n322 & n4013 ;
  assign n14967 = ~n1231 & n14966 ;
  assign n14968 = ( ~n3532 & n3961 ) | ( ~n3532 & n14967 ) | ( n3961 & n14967 ) ;
  assign n14969 = n3704 & n4983 ;
  assign n14970 = ~n14968 & n14969 ;
  assign n14972 = n3634 ^ n1952 ^ 1'b0 ;
  assign n14973 = x240 & n14972 ;
  assign n14974 = ~n4537 & n14973 ;
  assign n14975 = n11472 | n14974 ;
  assign n14971 = n12961 ^ n9076 ^ 1'b0 ;
  assign n14976 = n14975 ^ n14971 ^ n3395 ;
  assign n14977 = n14976 ^ n6920 ^ 1'b0 ;
  assign n14978 = n11467 ^ n1750 ^ 1'b0 ;
  assign n14979 = ~n2375 & n13821 ;
  assign n14980 = n14366 | n14979 ;
  assign n14981 = n14980 ^ n5619 ^ 1'b0 ;
  assign n14982 = x54 & n5587 ;
  assign n14983 = n1867 & ~n7741 ;
  assign n14984 = n14983 ^ n7314 ^ 1'b0 ;
  assign n14985 = ( n10285 & ~n11170 ) | ( n10285 & n14984 ) | ( ~n11170 & n14984 ) ;
  assign n14986 = n14985 ^ n2775 ^ 1'b0 ;
  assign n14987 = n14982 & n14986 ;
  assign n14988 = n3028 & n14987 ;
  assign n14989 = n1741 | n9354 ;
  assign n14990 = n4437 | n14989 ;
  assign n14991 = ( n9973 & n13272 ) | ( n9973 & n14990 ) | ( n13272 & n14990 ) ;
  assign n14992 = ~n3279 & n8360 ;
  assign n14993 = n13327 ^ n7635 ^ 1'b0 ;
  assign n14994 = n9586 ^ x176 ^ 1'b0 ;
  assign n14995 = n14526 & n14994 ;
  assign n14996 = n14995 ^ n5915 ^ 1'b0 ;
  assign n14997 = n1726 | n13108 ;
  assign n14998 = n9371 ^ n7967 ^ 1'b0 ;
  assign n15001 = x56 & n2873 ;
  assign n14999 = n419 | n5785 ;
  assign n15000 = n5758 & ~n14999 ;
  assign n15002 = n15001 ^ n15000 ^ 1'b0 ;
  assign n15003 = n14998 | n15002 ;
  assign n15004 = n1681 & n1814 ;
  assign n15005 = ~n2203 & n6272 ;
  assign n15006 = ~n15004 & n15005 ;
  assign n15012 = n8907 ^ n1901 ^ 1'b0 ;
  assign n15007 = n3738 & ~n9938 ;
  assign n15008 = n15007 ^ n7283 ^ 1'b0 ;
  assign n15009 = n12845 ^ n5206 ^ 1'b0 ;
  assign n15010 = n4639 | n15009 ;
  assign n15011 = ( n10901 & ~n15008 ) | ( n10901 & n15010 ) | ( ~n15008 & n15010 ) ;
  assign n15013 = n15012 ^ n15011 ^ 1'b0 ;
  assign n15014 = n6632 | n15013 ;
  assign n15015 = n12616 ^ n2735 ^ 1'b0 ;
  assign n15016 = n9473 ^ n359 ^ 1'b0 ;
  assign n15017 = n15015 & n15016 ;
  assign n15018 = ~x192 & n8510 ;
  assign n15019 = n15018 ^ n12945 ^ 1'b0 ;
  assign n15020 = n4972 ^ n1075 ^ n420 ;
  assign n15021 = ~n765 & n1495 ;
  assign n15022 = ~n1885 & n15021 ;
  assign n15023 = n12835 | n15022 ;
  assign n15024 = n15023 ^ n11923 ^ 1'b0 ;
  assign n15025 = n2302 ^ n2103 ^ 1'b0 ;
  assign n15026 = n15025 ^ n14616 ^ 1'b0 ;
  assign n15027 = ( ~x219 & n2086 ) | ( ~x219 & n6015 ) | ( n2086 & n6015 ) ;
  assign n15028 = ( ~n3386 & n6851 ) | ( ~n3386 & n7672 ) | ( n6851 & n7672 ) ;
  assign n15029 = n3790 | n15028 ;
  assign n15030 = n9292 & ~n15029 ;
  assign n15031 = n15030 ^ n11795 ^ n7154 ;
  assign n15032 = n8553 | n10694 ;
  assign n15033 = n15032 ^ n7643 ^ 1'b0 ;
  assign n15034 = n13558 & n15033 ;
  assign n15035 = ~n1680 & n7936 ;
  assign n15036 = ~n5380 & n7184 ;
  assign n15037 = n5238 & n15036 ;
  assign n15038 = n12280 ^ n4260 ^ n1101 ;
  assign n15039 = n6550 ^ n4453 ^ 1'b0 ;
  assign n15040 = n4791 ^ n4415 ^ 1'b0 ;
  assign n15041 = ~n3838 & n15040 ;
  assign n15042 = ~n2807 & n15041 ;
  assign n15043 = n15042 ^ n4979 ^ 1'b0 ;
  assign n15044 = n11175 | n15043 ;
  assign n15045 = n11369 ^ n6864 ^ 1'b0 ;
  assign n15046 = n13834 & n15045 ;
  assign n15047 = n7873 | n12961 ;
  assign n15048 = n1330 | n15047 ;
  assign n15049 = n8915 & n11717 ;
  assign n15050 = n12344 ^ n3598 ^ 1'b0 ;
  assign n15051 = n13496 & n15050 ;
  assign n15052 = n5837 ^ n5201 ^ 1'b0 ;
  assign n15053 = n8336 & ~n15052 ;
  assign n15055 = n4519 ^ n296 ^ 1'b0 ;
  assign n15056 = ( n908 & n12569 ) | ( n908 & n15055 ) | ( n12569 & n15055 ) ;
  assign n15054 = ~n9769 & n10259 ;
  assign n15057 = n15056 ^ n15054 ^ 1'b0 ;
  assign n15058 = n3818 | n4909 ;
  assign n15059 = x251 | n15058 ;
  assign n15060 = n2856 & ~n15037 ;
  assign n15061 = n15060 ^ n9721 ^ 1'b0 ;
  assign n15062 = n5986 & n15061 ;
  assign n15063 = ~n15059 & n15062 ;
  assign n15064 = n10041 ^ x140 ^ 1'b0 ;
  assign n15065 = n6701 & n15064 ;
  assign n15066 = n4906 & n15065 ;
  assign n15067 = ~n446 & n15066 ;
  assign n15068 = n9281 ^ n5067 ^ 1'b0 ;
  assign n15069 = n5324 | n10847 ;
  assign n15070 = n5871 ^ n581 ^ 1'b0 ;
  assign n15071 = n15070 ^ n5276 ^ 1'b0 ;
  assign n15072 = n15071 ^ n3863 ^ 1'b0 ;
  assign n15073 = n15069 & ~n15072 ;
  assign n15074 = n7813 ^ n4014 ^ 1'b0 ;
  assign n15075 = n4122 & n12361 ;
  assign n15076 = n15075 ^ n2258 ^ 1'b0 ;
  assign n15077 = n5560 ^ n1554 ^ 1'b0 ;
  assign n15078 = n2904 & ~n15077 ;
  assign n15079 = ~n5232 & n15078 ;
  assign n15080 = ( ~n6378 & n10372 ) | ( ~n6378 & n12576 ) | ( n10372 & n12576 ) ;
  assign n15081 = n15080 ^ n9921 ^ 1'b0 ;
  assign n15082 = ~n4189 & n15081 ;
  assign n15083 = n8646 ^ n2262 ^ 1'b0 ;
  assign n15084 = n9622 | n15083 ;
  assign n15085 = n2533 & ~n13771 ;
  assign n15086 = n3069 & ~n5081 ;
  assign n15087 = n9450 ^ n5018 ^ 1'b0 ;
  assign n15088 = n15086 & n15087 ;
  assign n15089 = n11191 & n15088 ;
  assign n15090 = n6115 ^ n1215 ^ 1'b0 ;
  assign n15094 = n5465 ^ n1318 ^ 1'b0 ;
  assign n15091 = n10928 ^ n6933 ^ 1'b0 ;
  assign n15092 = n7490 | n15091 ;
  assign n15093 = n3272 & ~n15092 ;
  assign n15095 = n15094 ^ n15093 ^ n3054 ;
  assign n15096 = n1219 & n10827 ;
  assign n15097 = n15096 ^ n11578 ^ 1'b0 ;
  assign n15098 = n4575 | n15097 ;
  assign n15099 = n15098 ^ n12285 ^ 1'b0 ;
  assign n15100 = n10096 | n15099 ;
  assign n15101 = n3094 & n13615 ;
  assign n15102 = n2587 ^ n2192 ^ 1'b0 ;
  assign n15103 = n8822 & n15102 ;
  assign n15104 = n1532 & n15103 ;
  assign n15105 = n7577 | n15104 ;
  assign n15106 = n15105 ^ n3942 ^ 1'b0 ;
  assign n15107 = n4750 ^ n4360 ^ 1'b0 ;
  assign n15108 = n2018 & n15107 ;
  assign n15109 = n13288 & n15108 ;
  assign n15110 = ~n3635 & n12676 ;
  assign n15111 = n2062 & n15110 ;
  assign n15112 = n6409 | n11247 ;
  assign n15113 = ( n3131 & ~n10731 ) | ( n3131 & n10835 ) | ( ~n10731 & n10835 ) ;
  assign n15114 = x162 & ~n5238 ;
  assign n15115 = ~x48 & n15114 ;
  assign n15117 = n5942 & ~n8222 ;
  assign n15118 = n15117 ^ n7825 ^ 1'b0 ;
  assign n15119 = ~n627 & n15118 ;
  assign n15120 = ~n11001 & n15119 ;
  assign n15121 = n10737 | n15120 ;
  assign n15122 = n15121 ^ n10142 ^ 1'b0 ;
  assign n15116 = n3399 & ~n9998 ;
  assign n15123 = n15122 ^ n15116 ^ 1'b0 ;
  assign n15124 = n15123 ^ n5987 ^ 1'b0 ;
  assign n15125 = n4757 | n4997 ;
  assign n15126 = n15125 ^ n4074 ^ 1'b0 ;
  assign n15127 = n2487 ^ n631 ^ 1'b0 ;
  assign n15128 = n4132 & n15127 ;
  assign n15129 = n1887 & n15128 ;
  assign n15130 = x104 & ~n1932 ;
  assign n15131 = ~n15129 & n15130 ;
  assign n15132 = n4546 & ~n15131 ;
  assign n15133 = ~n10790 & n15132 ;
  assign n15134 = ~n5492 & n8295 ;
  assign n15135 = n15134 ^ n1133 ^ 1'b0 ;
  assign n15136 = n3736 | n7372 ;
  assign n15137 = n15136 ^ n9976 ^ 1'b0 ;
  assign n15138 = n2959 & n3765 ;
  assign n15139 = ~n5895 & n15138 ;
  assign n15140 = n11764 ^ n1473 ^ 1'b0 ;
  assign n15141 = n8578 ^ n2387 ^ n1566 ;
  assign n15142 = n3447 & n13038 ;
  assign n15143 = n15142 ^ n1835 ^ 1'b0 ;
  assign n15144 = n7266 ^ n1839 ^ 1'b0 ;
  assign n15145 = n7534 | n15144 ;
  assign n15146 = n3969 | n15145 ;
  assign n15147 = n8207 | n14724 ;
  assign n15148 = n3574 | n15147 ;
  assign n15149 = n15148 ^ n4267 ^ 1'b0 ;
  assign n15150 = n15146 | n15149 ;
  assign n15151 = n15150 ^ n2148 ^ 1'b0 ;
  assign n15152 = x57 & ~n11265 ;
  assign n15153 = ~n294 & n15152 ;
  assign n15154 = ( n917 & n3975 ) | ( n917 & ~n10253 ) | ( n3975 & ~n10253 ) ;
  assign n15155 = n9897 ^ n2859 ^ 1'b0 ;
  assign n15156 = n7426 & ~n8103 ;
  assign n15157 = n15156 ^ n10142 ^ 1'b0 ;
  assign n15158 = n3724 | n15157 ;
  assign n15159 = n599 ^ n315 ^ 1'b0 ;
  assign n15160 = n2123 & n15159 ;
  assign n15161 = n15160 ^ n9862 ^ n806 ;
  assign n15162 = ~n6243 & n15161 ;
  assign n15163 = n2323 & n7856 ;
  assign n15164 = n10061 ^ n3121 ^ 1'b0 ;
  assign n15165 = n2249 & n15164 ;
  assign n15166 = n6338 & n15165 ;
  assign n15167 = n4104 & ~n4370 ;
  assign n15168 = ~n4617 & n14445 ;
  assign n15169 = ~n15167 & n15168 ;
  assign n15170 = n3613 ^ n3308 ^ 1'b0 ;
  assign n15171 = ~n10391 & n15170 ;
  assign n15172 = n274 ^ x65 ^ 1'b0 ;
  assign n15173 = ~n6207 & n15172 ;
  assign n15174 = ~n3225 & n9652 ;
  assign n15175 = ~n2976 & n3098 ;
  assign n15176 = ~n15174 & n15175 ;
  assign n15177 = ~n7271 & n13658 ;
  assign n15178 = n10899 ^ n1101 ^ 1'b0 ;
  assign n15179 = ~n5425 & n7303 ;
  assign n15180 = n15179 ^ n12474 ^ 1'b0 ;
  assign n15181 = n15178 & ~n15180 ;
  assign n15182 = ~n4638 & n5986 ;
  assign n15183 = n15182 ^ n1557 ^ 1'b0 ;
  assign n15184 = n7457 | n10451 ;
  assign n15185 = n15184 ^ n3271 ^ 1'b0 ;
  assign n15186 = n2378 & n12123 ;
  assign n15187 = n15186 ^ n5481 ^ 1'b0 ;
  assign n15188 = n15187 ^ n13172 ^ 1'b0 ;
  assign n15189 = ~n851 & n10410 ;
  assign n15190 = n10527 & ~n15189 ;
  assign n15191 = ~n13079 & n15190 ;
  assign n15192 = n3440 | n15191 ;
  assign n15193 = ( n1189 & ~n7635 ) | ( n1189 & n11061 ) | ( ~n7635 & n11061 ) ;
  assign n15194 = ~n11549 & n15193 ;
  assign n15195 = n12840 & n15194 ;
  assign n15196 = n15195 ^ n7384 ^ 1'b0 ;
  assign n15197 = n15196 ^ n10959 ^ 1'b0 ;
  assign n15198 = n1975 & ~n13370 ;
  assign n15199 = ~n13399 & n15198 ;
  assign n15200 = n2688 ^ x157 ^ 1'b0 ;
  assign n15201 = n15199 & ~n15200 ;
  assign n15202 = n14381 ^ n7134 ^ 1'b0 ;
  assign n15206 = ~n1208 & n5515 ;
  assign n15207 = n15206 ^ n9571 ^ 1'b0 ;
  assign n15203 = ~n10895 & n12269 ;
  assign n15204 = n10767 & n15203 ;
  assign n15205 = n858 & ~n15204 ;
  assign n15208 = n15207 ^ n15205 ^ 1'b0 ;
  assign n15209 = n15208 ^ x225 ^ 1'b0 ;
  assign n15210 = n722 & n925 ;
  assign n15211 = n9440 & ~n11232 ;
  assign n15212 = ~n14694 & n15211 ;
  assign n15213 = n15212 ^ x192 ^ 1'b0 ;
  assign n15214 = ( ~n9672 & n15210 ) | ( ~n9672 & n15213 ) | ( n15210 & n15213 ) ;
  assign n15215 = n7351 & ~n15104 ;
  assign n15216 = n9291 ^ n3626 ^ 1'b0 ;
  assign n15217 = ~n2559 & n6358 ;
  assign n15218 = n11503 | n15217 ;
  assign n15219 = n5654 & ~n15218 ;
  assign n15220 = n10284 ^ n880 ^ 1'b0 ;
  assign n15221 = n3788 | n4791 ;
  assign n15222 = n8118 ^ n6864 ^ 1'b0 ;
  assign n15223 = n12445 ^ n12092 ^ 1'b0 ;
  assign n15224 = n15222 & n15223 ;
  assign n15225 = n2891 | n4423 ;
  assign n15226 = n7826 & n15225 ;
  assign n15227 = n13618 & n15226 ;
  assign n15228 = n5667 ^ n2167 ^ 1'b0 ;
  assign n15229 = n1757 & ~n9365 ;
  assign n15230 = ~n8577 & n15229 ;
  assign n15231 = n15230 ^ n10959 ^ 1'b0 ;
  assign n15232 = ~n1447 & n15231 ;
  assign n15235 = n436 & ~n6483 ;
  assign n15236 = ~n7670 & n15235 ;
  assign n15233 = n1342 & n14163 ;
  assign n15234 = ~n11905 & n15233 ;
  assign n15237 = n15236 ^ n15234 ^ 1'b0 ;
  assign n15238 = ~n10023 & n15237 ;
  assign n15239 = n11459 & n15238 ;
  assign n15240 = n6075 ^ n5066 ^ 1'b0 ;
  assign n15241 = n15240 ^ n991 ^ 1'b0 ;
  assign n15242 = n5909 ^ n3645 ^ 1'b0 ;
  assign n15243 = n3568 & n15242 ;
  assign n15244 = n5540 ^ n583 ^ 1'b0 ;
  assign n15245 = n15243 & ~n15244 ;
  assign n15246 = x186 & ~n15176 ;
  assign n15247 = n7040 & n15246 ;
  assign n15248 = x81 & n12538 ;
  assign n15249 = n2807 & ~n15248 ;
  assign n15250 = n3447 & ~n8460 ;
  assign n15251 = ~n15249 & n15250 ;
  assign n15252 = n444 | n1086 ;
  assign n15253 = n8921 & n15252 ;
  assign n15254 = n1116 | n1219 ;
  assign n15255 = n15254 ^ n13236 ^ 1'b0 ;
  assign n15256 = n12198 ^ n1200 ^ 1'b0 ;
  assign n15257 = ( n3886 & n10557 ) | ( n3886 & n10898 ) | ( n10557 & n10898 ) ;
  assign n15258 = n11063 ^ n9574 ^ 1'b0 ;
  assign n15259 = n10499 ^ n5069 ^ 1'b0 ;
  assign n15260 = ~n5619 & n8196 ;
  assign n15261 = n3508 | n15260 ;
  assign n15262 = ~n5195 & n15261 ;
  assign n15263 = n15259 & n15262 ;
  assign n15264 = n5651 & n6339 ;
  assign n15265 = n1486 & n1591 ;
  assign n15266 = ~n8423 & n15265 ;
  assign n15267 = n1261 | n11328 ;
  assign n15268 = n3490 & ~n15267 ;
  assign n15269 = n3977 & ~n15268 ;
  assign n15270 = n4861 | n10839 ;
  assign n15271 = n2992 | n15270 ;
  assign n15272 = n13607 ^ n2983 ^ 1'b0 ;
  assign n15273 = ~n2509 & n15272 ;
  assign n15274 = n5966 ^ n4494 ^ 1'b0 ;
  assign n15275 = ~n2103 & n15274 ;
  assign n15276 = n15275 ^ n4593 ^ 1'b0 ;
  assign n15277 = n5324 ^ x239 ^ 1'b0 ;
  assign n15278 = n15277 ^ n13526 ^ 1'b0 ;
  assign n15279 = n5767 & ~n15278 ;
  assign n15280 = n10687 & ~n15279 ;
  assign n15281 = n322 & n15280 ;
  assign n15282 = ~n2733 & n4153 ;
  assign n15283 = ( n6681 & n8718 ) | ( n6681 & ~n15282 ) | ( n8718 & ~n15282 ) ;
  assign n15284 = n4787 ^ x96 ^ 1'b0 ;
  assign n15285 = ~n11179 & n15284 ;
  assign n15286 = n2114 & ~n6639 ;
  assign n15287 = x42 & n4368 ;
  assign n15288 = ~n5722 & n15287 ;
  assign n15289 = n11199 ^ n7819 ^ n5848 ;
  assign n15290 = n8866 & ~n15289 ;
  assign n15291 = n5177 | n15290 ;
  assign n15292 = n15291 ^ n3596 ^ 1'b0 ;
  assign n15293 = n2378 ^ n1406 ^ 1'b0 ;
  assign n15294 = n13082 & n15293 ;
  assign n15295 = n5418 & n10055 ;
  assign n15296 = ~n12921 & n15295 ;
  assign n15297 = n12145 & n15296 ;
  assign n15298 = n2988 & ~n12802 ;
  assign n15299 = n5746 ^ n4285 ^ 1'b0 ;
  assign n15300 = n15299 ^ n4534 ^ 1'b0 ;
  assign n15301 = ~n9823 & n15300 ;
  assign n15302 = ~n9442 & n14335 ;
  assign n15303 = n15302 ^ n2378 ^ 1'b0 ;
  assign n15304 = n15303 ^ n4933 ^ 1'b0 ;
  assign n15305 = ( n1494 & n4788 ) | ( n1494 & ~n7329 ) | ( n4788 & ~n7329 ) ;
  assign n15306 = n8278 & n15305 ;
  assign n15307 = n15306 ^ n1393 ^ 1'b0 ;
  assign n15308 = n9573 ^ n4935 ^ 1'b0 ;
  assign n15309 = n3237 & ~n3926 ;
  assign n15310 = ( n3551 & ~n15308 ) | ( n3551 & n15309 ) | ( ~n15308 & n15309 ) ;
  assign n15311 = n1142 & ~n6158 ;
  assign n15312 = n15311 ^ n7092 ^ 1'b0 ;
  assign n15313 = n15312 ^ n12059 ^ n2007 ;
  assign n15314 = n15310 & n15313 ;
  assign n15315 = n558 & ~n2246 ;
  assign n15316 = n3864 & ~n15315 ;
  assign n15317 = n4752 ^ n1645 ^ 1'b0 ;
  assign n15318 = ~n3140 & n15317 ;
  assign n15319 = n15318 ^ n5632 ^ 1'b0 ;
  assign n15320 = n15319 ^ n6382 ^ n3109 ;
  assign n15321 = n9719 ^ n8022 ^ n7846 ;
  assign n15322 = ( n1994 & n8583 ) | ( n1994 & n15321 ) | ( n8583 & n15321 ) ;
  assign n15323 = n1854 & ~n5521 ;
  assign n15324 = n7810 & n15323 ;
  assign n15325 = n3386 | n15324 ;
  assign n15326 = n6448 ^ n547 ^ 1'b0 ;
  assign n15327 = ~n622 & n15326 ;
  assign n15328 = n13783 | n15327 ;
  assign n15329 = n4864 | n7856 ;
  assign n15330 = n15329 ^ n1956 ^ 1'b0 ;
  assign n15331 = n6886 & n15330 ;
  assign n15332 = n14591 ^ n1374 ^ 1'b0 ;
  assign n15333 = ( ~n957 & n2180 ) | ( ~n957 & n3844 ) | ( n2180 & n3844 ) ;
  assign n15334 = n3754 | n10203 ;
  assign n15335 = n10231 ^ n10146 ^ n6785 ;
  assign n15336 = n1093 & ~n11963 ;
  assign n15341 = n4074 ^ n2659 ^ 1'b0 ;
  assign n15337 = n5187 ^ n1344 ^ 1'b0 ;
  assign n15338 = ( ~n1550 & n2246 ) | ( ~n1550 & n15337 ) | ( n2246 & n15337 ) ;
  assign n15339 = n3481 | n4197 ;
  assign n15340 = n15338 & ~n15339 ;
  assign n15342 = n15341 ^ n15340 ^ 1'b0 ;
  assign n15343 = n2809 ^ n340 ^ 1'b0 ;
  assign n15344 = n938 | n9218 ;
  assign n15345 = n14089 & ~n15344 ;
  assign n15346 = n14010 & ~n15345 ;
  assign n15347 = n9004 ^ n3690 ^ 1'b0 ;
  assign n15348 = ( ~n1093 & n4432 ) | ( ~n1093 & n15347 ) | ( n4432 & n15347 ) ;
  assign n15349 = n11705 ^ n1775 ^ 1'b0 ;
  assign n15350 = n5874 ^ x185 ^ 1'b0 ;
  assign n15351 = n4256 & n15350 ;
  assign n15352 = ~n3351 & n15351 ;
  assign n15353 = ~n431 & n15352 ;
  assign n15354 = n14584 ^ n12936 ^ 1'b0 ;
  assign n15355 = n11681 ^ n3235 ^ 1'b0 ;
  assign n15356 = n13041 & n15355 ;
  assign n15357 = ~n6112 & n9060 ;
  assign n15358 = n2763 | n8746 ;
  assign n15359 = n15358 ^ n11369 ^ 1'b0 ;
  assign n15360 = n15357 | n15359 ;
  assign n15361 = n11012 | n12250 ;
  assign n15362 = n11461 & ~n12479 ;
  assign n15363 = n15362 ^ n10698 ^ 1'b0 ;
  assign n15364 = n15361 & ~n15363 ;
  assign n15365 = n15364 ^ n796 ^ 1'b0 ;
  assign n15366 = n4918 ^ n4547 ^ n3648 ;
  assign n15367 = x155 & ~n3481 ;
  assign n15368 = n15367 ^ n3183 ^ 1'b0 ;
  assign n15369 = n15366 | n15368 ;
  assign n15370 = n15369 ^ x79 ^ 1'b0 ;
  assign n15371 = ~n986 & n1553 ;
  assign n15372 = n15371 ^ n5160 ^ 1'b0 ;
  assign n15373 = n6655 & n6700 ;
  assign n15374 = n367 & ~n8233 ;
  assign n15375 = n15374 ^ n9872 ^ 1'b0 ;
  assign n15376 = n1651 ^ n1237 ^ 1'b0 ;
  assign n15377 = n2841 & n15376 ;
  assign n15378 = n4380 & n14159 ;
  assign n15379 = n5775 ^ n5205 ^ 1'b0 ;
  assign n15380 = ~n1409 & n15379 ;
  assign n15381 = n15380 ^ n3864 ^ 1'b0 ;
  assign n15382 = n5662 ^ n318 ^ 1'b0 ;
  assign n15383 = n9755 & ~n15382 ;
  assign n15384 = ~n7600 & n13511 ;
  assign n15385 = n1137 & n15384 ;
  assign n15386 = n5188 & n12081 ;
  assign n15387 = n2916 & n15386 ;
  assign n15388 = n1638 & n4976 ;
  assign n15389 = n15388 ^ n4282 ^ 1'b0 ;
  assign n15390 = n10256 & n15389 ;
  assign n15391 = n5969 ^ n2706 ^ 1'b0 ;
  assign n15392 = n1478 & ~n15391 ;
  assign n15393 = n15392 ^ n5187 ^ 1'b0 ;
  assign n15394 = ~n1442 & n15393 ;
  assign n15395 = n3378 & ~n10611 ;
  assign n15397 = n4837 & n4918 ;
  assign n15398 = n15397 ^ n4742 ^ 1'b0 ;
  assign n15396 = ~n11053 & n14929 ;
  assign n15399 = n15398 ^ n15396 ^ 1'b0 ;
  assign n15400 = n6465 ^ n2697 ^ n739 ;
  assign n15401 = ~n3395 & n15400 ;
  assign n15402 = n15401 ^ n2701 ^ 1'b0 ;
  assign n15403 = n6524 ^ n5234 ^ 1'b0 ;
  assign n15404 = ~n812 & n15403 ;
  assign n15405 = ( n4393 & n7770 ) | ( n4393 & n15404 ) | ( n7770 & n15404 ) ;
  assign n15406 = n15405 ^ n9747 ^ 1'b0 ;
  assign n15407 = n1153 & n14544 ;
  assign n15408 = n15406 & n15407 ;
  assign n15409 = n10529 & ~n13802 ;
  assign n15410 = n15409 ^ n12622 ^ 1'b0 ;
  assign n15411 = n860 | n7934 ;
  assign n15412 = n15411 ^ n7210 ^ 1'b0 ;
  assign n15413 = x158 & n15412 ;
  assign n15414 = ~n9755 & n15413 ;
  assign n15415 = n11112 ^ n7702 ^ 1'b0 ;
  assign n15416 = ~x118 & n15415 ;
  assign n15417 = ( n3845 & n6202 ) | ( n3845 & ~n15416 ) | ( n6202 & ~n15416 ) ;
  assign n15418 = n9824 ^ n8479 ^ 1'b0 ;
  assign n15419 = n15418 ^ n794 ^ 1'b0 ;
  assign n15420 = n3595 & n15419 ;
  assign n15421 = n8305 ^ n6341 ^ n2785 ;
  assign n15422 = ~n1809 & n15421 ;
  assign n15423 = n8300 & ~n15422 ;
  assign n15424 = ~n3138 & n4338 ;
  assign n15425 = n9340 & n15424 ;
  assign n15426 = n3542 & ~n6187 ;
  assign n15427 = n15426 ^ n1028 ^ 1'b0 ;
  assign n15428 = x55 | n15427 ;
  assign n15429 = x164 & n7452 ;
  assign n15430 = n8037 & n15429 ;
  assign n15431 = n11124 ^ x112 ^ 1'b0 ;
  assign n15432 = n2897 | n15431 ;
  assign n15433 = n5933 ^ n5350 ^ 1'b0 ;
  assign n15434 = n3205 & ~n3262 ;
  assign n15435 = ~n13359 & n15434 ;
  assign n15436 = n13845 & n15435 ;
  assign n15437 = n3010 ^ x154 ^ 1'b0 ;
  assign n15438 = n4730 | n15437 ;
  assign n15439 = ( n2204 & n8023 ) | ( n2204 & ~n9458 ) | ( n8023 & ~n9458 ) ;
  assign n15440 = n1600 & ~n14483 ;
  assign n15441 = ~n8607 & n15440 ;
  assign n15442 = n7903 ^ x139 ^ 1'b0 ;
  assign n15443 = n13658 & n15442 ;
  assign n15444 = n1208 | n8619 ;
  assign n15445 = n8827 & ~n15444 ;
  assign n15446 = ( n1669 & n4895 ) | ( n1669 & n15445 ) | ( n4895 & n15445 ) ;
  assign n15447 = n11498 & ~n14630 ;
  assign n15448 = n3237 & n15447 ;
  assign n15449 = n11386 & n15448 ;
  assign n15450 = n10164 & ~n15449 ;
  assign n15451 = ~n5704 & n15450 ;
  assign n15452 = ( ~n7198 & n15446 ) | ( ~n7198 & n15451 ) | ( n15446 & n15451 ) ;
  assign n15453 = n8849 & n9357 ;
  assign n15454 = n12349 ^ n8589 ^ 1'b0 ;
  assign n15455 = n15453 & n15454 ;
  assign n15459 = n7594 | n13666 ;
  assign n15460 = ( n640 & n8281 ) | ( n640 & ~n15459 ) | ( n8281 & ~n15459 ) ;
  assign n15456 = n3472 ^ n969 ^ n385 ;
  assign n15457 = n15456 ^ n14514 ^ 1'b0 ;
  assign n15458 = n11245 & ~n15457 ;
  assign n15461 = n15460 ^ n15458 ^ x3 ;
  assign n15462 = n5390 ^ n3332 ^ 1'b0 ;
  assign n15463 = ~n2244 & n15462 ;
  assign n15464 = ( n5428 & ~n10455 ) | ( n5428 & n15463 ) | ( ~n10455 & n15463 ) ;
  assign n15465 = ( n7579 & ~n7920 ) | ( n7579 & n11883 ) | ( ~n7920 & n11883 ) ;
  assign n15468 = n4018 | n9093 ;
  assign n15467 = n3214 & n6692 ;
  assign n15469 = n15468 ^ n15467 ^ 1'b0 ;
  assign n15466 = n7838 ^ n5425 ^ 1'b0 ;
  assign n15470 = n15469 ^ n15466 ^ 1'b0 ;
  assign n15471 = ~n15465 & n15470 ;
  assign n15472 = n5498 & n10735 ;
  assign n15473 = n9568 & ~n10914 ;
  assign n15474 = n15472 | n15473 ;
  assign n15475 = n12101 & ~n15474 ;
  assign n15476 = n15471 & ~n15475 ;
  assign n15477 = ~n10339 & n15476 ;
  assign n15478 = n8487 ^ n4345 ^ 1'b0 ;
  assign n15479 = n2674 & ~n15478 ;
  assign n15480 = n369 | n10905 ;
  assign n15481 = n15480 ^ n2919 ^ 1'b0 ;
  assign n15482 = x159 & ~n15481 ;
  assign n15483 = ~n15479 & n15482 ;
  assign n15484 = n1664 & ~n7331 ;
  assign n15485 = n10369 ^ n7383 ^ 1'b0 ;
  assign n15486 = n12575 ^ n8276 ^ n3075 ;
  assign n15487 = n15486 ^ n11921 ^ 1'b0 ;
  assign n15488 = n10024 ^ n6010 ^ 1'b0 ;
  assign n15489 = ( ~n2928 & n3421 ) | ( ~n2928 & n10949 ) | ( n3421 & n10949 ) ;
  assign n15490 = n860 & ~n15489 ;
  assign n15491 = ( n1126 & ~n15488 ) | ( n1126 & n15490 ) | ( ~n15488 & n15490 ) ;
  assign n15492 = ( n6093 & n6359 ) | ( n6093 & n15491 ) | ( n6359 & n15491 ) ;
  assign n15493 = ~n4649 & n9673 ;
  assign n15494 = ~n3105 & n7054 ;
  assign n15495 = ~n15493 & n15494 ;
  assign n15496 = n6847 ^ x232 ^ 1'b0 ;
  assign n15497 = n9347 & ~n15496 ;
  assign n15498 = ~n14829 & n15497 ;
  assign n15499 = n5739 ^ n3265 ^ 1'b0 ;
  assign n15500 = ~n579 & n15499 ;
  assign n15501 = n7329 & ~n15500 ;
  assign n15502 = n11105 ^ n5208 ^ 1'b0 ;
  assign n15503 = n12418 ^ n6712 ^ n1484 ;
  assign n15504 = n2343 | n15469 ;
  assign n15505 = n9142 & ~n15504 ;
  assign n15506 = ~n15503 & n15505 ;
  assign n15507 = ~n513 & n566 ;
  assign n15508 = n2681 ^ x231 ^ 1'b0 ;
  assign n15509 = n15507 & ~n15508 ;
  assign n15510 = n9655 & ~n15509 ;
  assign n15511 = n14496 ^ n13821 ^ n10064 ;
  assign n15512 = n1138 & ~n15511 ;
  assign n15513 = n10615 ^ n6576 ^ 1'b0 ;
  assign n15514 = n12347 & n15513 ;
  assign n15515 = n3104 ^ n1504 ^ 1'b0 ;
  assign n15516 = ( n12585 & n13668 ) | ( n12585 & ~n15515 ) | ( n13668 & ~n15515 ) ;
  assign n15517 = n1478 & n9225 ;
  assign n15518 = n15517 ^ n5364 ^ 1'b0 ;
  assign n15519 = n11619 | n15518 ;
  assign n15520 = n14878 & ~n15519 ;
  assign n15521 = ( n812 & n1273 ) | ( n812 & n12238 ) | ( n1273 & n12238 ) ;
  assign n15522 = ~n5315 & n8915 ;
  assign n15523 = n10589 & n15522 ;
  assign n15524 = n14990 & ~n15523 ;
  assign n15525 = n3238 ^ x89 ^ 1'b0 ;
  assign n15526 = n2275 & ~n15525 ;
  assign n15527 = ~n2771 & n5671 ;
  assign n15528 = n2771 & n15527 ;
  assign n15529 = n3747 & ~n15528 ;
  assign n15530 = ~n3747 & n15529 ;
  assign n15531 = n4498 | n15530 ;
  assign n15532 = n2794 & ~n15531 ;
  assign n15533 = n14222 ^ n12963 ^ 1'b0 ;
  assign n15534 = n4113 | n15533 ;
  assign n15535 = n8740 ^ n728 ^ 1'b0 ;
  assign n15536 = n10610 ^ n8087 ^ 1'b0 ;
  assign n15537 = ~n420 & n15536 ;
  assign n15538 = ~n3850 & n14035 ;
  assign n15539 = n2857 & ~n5255 ;
  assign n15540 = n676 & ~n1356 ;
  assign n15541 = ( n1206 & n8580 ) | ( n1206 & n10268 ) | ( n8580 & n10268 ) ;
  assign n15542 = n2556 & n8112 ;
  assign n15543 = ~n6383 & n15542 ;
  assign n15544 = ~n2554 & n9009 ;
  assign n15545 = ( n15541 & ~n15543 ) | ( n15541 & n15544 ) | ( ~n15543 & n15544 ) ;
  assign n15546 = n479 | n2477 ;
  assign n15547 = n15546 ^ n11570 ^ 1'b0 ;
  assign n15548 = n6737 & n15547 ;
  assign n15549 = n4806 & n15548 ;
  assign n15550 = n14964 ^ n1632 ^ 1'b0 ;
  assign n15551 = n15549 | n15550 ;
  assign n15552 = n5934 ^ n2308 ^ 1'b0 ;
  assign n15553 = ~n3007 & n15552 ;
  assign n15554 = n9841 & ~n12723 ;
  assign n15555 = ~n15553 & n15554 ;
  assign n15556 = n13971 ^ n3513 ^ 1'b0 ;
  assign n15557 = n4040 | n15556 ;
  assign n15558 = n357 & ~n14595 ;
  assign n15559 = n15557 & n15558 ;
  assign n15560 = n6346 ^ n2113 ^ 1'b0 ;
  assign n15561 = n15560 ^ n906 ^ 1'b0 ;
  assign n15562 = n6835 ^ n1947 ^ 1'b0 ;
  assign n15563 = n4506 & n15562 ;
  assign n15564 = n599 | n2748 ;
  assign n15565 = n9168 ^ n3481 ^ 1'b0 ;
  assign n15566 = n4576 ^ n813 ^ 1'b0 ;
  assign n15567 = n15565 | n15566 ;
  assign n15568 = ( n6947 & ~n15564 ) | ( n6947 & n15567 ) | ( ~n15564 & n15567 ) ;
  assign n15569 = n2287 | n6765 ;
  assign n15570 = n1276 & ~n15569 ;
  assign n15571 = n2719 & ~n3255 ;
  assign n15572 = n3690 | n8712 ;
  assign n15573 = ~n2174 & n15572 ;
  assign n15574 = n4093 ^ n2284 ^ 1'b0 ;
  assign n15575 = ( n801 & ~n8957 ) | ( n801 & n9807 ) | ( ~n8957 & n9807 ) ;
  assign n15576 = ~n7964 & n15575 ;
  assign n15577 = n15576 ^ n13539 ^ 1'b0 ;
  assign n15578 = n4411 & ~n10880 ;
  assign n15579 = n2911 ^ n1271 ^ 1'b0 ;
  assign n15580 = ~n7738 & n15579 ;
  assign n15581 = n15580 ^ n3588 ^ 1'b0 ;
  assign n15582 = n5416 | n15581 ;
  assign n15583 = n2928 ^ n2286 ^ 1'b0 ;
  assign n15584 = ~n986 & n12418 ;
  assign n15585 = ~n12418 & n15584 ;
  assign n15586 = n11002 | n15585 ;
  assign n15587 = n15583 & n15586 ;
  assign n15588 = x168 & ~n3133 ;
  assign n15589 = n3133 & n15588 ;
  assign n15590 = n4093 & n15589 ;
  assign n15591 = ~n15587 & n15590 ;
  assign n15592 = n15587 & n15591 ;
  assign n15593 = n5246 & n15592 ;
  assign n15594 = n4817 ^ n1735 ^ 1'b0 ;
  assign n15595 = ( n458 & ~n9284 ) | ( n458 & n15594 ) | ( ~n9284 & n15594 ) ;
  assign n15596 = ~n10570 & n15595 ;
  assign n15597 = n7833 ^ n5197 ^ 1'b0 ;
  assign n15598 = n4124 & ~n15597 ;
  assign n15599 = n12969 ^ n3513 ^ 1'b0 ;
  assign n15600 = n15598 & ~n15599 ;
  assign n15601 = ( n839 & ~n10068 ) | ( n839 & n15600 ) | ( ~n10068 & n15600 ) ;
  assign n15602 = ( n2445 & n7032 ) | ( n2445 & ~n8861 ) | ( n7032 & ~n8861 ) ;
  assign n15603 = n15601 | n15602 ;
  assign n15604 = ~n3622 & n4730 ;
  assign n15605 = n15604 ^ n11754 ^ 1'b0 ;
  assign n15606 = ~n9725 & n14434 ;
  assign n15607 = ~n5849 & n15606 ;
  assign n15608 = n9930 ^ n1255 ^ 1'b0 ;
  assign n15609 = n10333 | n15608 ;
  assign n15610 = n15607 | n15609 ;
  assign n15611 = n15605 & ~n15610 ;
  assign n15613 = ~n2506 & n9730 ;
  assign n15614 = n15613 ^ n11295 ^ 1'b0 ;
  assign n15612 = n5027 ^ n2568 ^ 1'b0 ;
  assign n15615 = n15614 ^ n15612 ^ n15169 ;
  assign n15616 = n14377 ^ n13502 ^ 1'b0 ;
  assign n15617 = n9051 ^ n3885 ^ 1'b0 ;
  assign n15618 = n9198 ^ n5317 ^ 1'b0 ;
  assign n15619 = n1028 & ~n15618 ;
  assign n15620 = n12264 ^ n9475 ^ 1'b0 ;
  assign n15621 = n15620 ^ n5012 ^ 1'b0 ;
  assign n15622 = n7846 & ~n15621 ;
  assign n15623 = n15622 ^ n3845 ^ 1'b0 ;
  assign n15624 = n15623 ^ x173 ^ 1'b0 ;
  assign n15625 = n5671 & n6298 ;
  assign n15626 = n867 & n15625 ;
  assign n15627 = n2611 & n15626 ;
  assign n15628 = n464 | n5745 ;
  assign n15629 = ( n8862 & n13152 ) | ( n8862 & n15628 ) | ( n13152 & n15628 ) ;
  assign n15630 = n13253 ^ n4269 ^ 1'b0 ;
  assign n15631 = n11581 ^ n6826 ^ 1'b0 ;
  assign n15632 = n5537 | n15631 ;
  assign n15633 = n15632 ^ n4122 ^ 1'b0 ;
  assign n15634 = ~n938 & n13586 ;
  assign n15635 = n15634 ^ n547 ^ 1'b0 ;
  assign n15636 = ~n3911 & n15635 ;
  assign n15637 = n15636 ^ n14228 ^ 1'b0 ;
  assign n15638 = ( n3966 & n5110 ) | ( n3966 & n13429 ) | ( n5110 & n13429 ) ;
  assign n15639 = n15638 ^ n1960 ^ 1'b0 ;
  assign n15640 = n11129 ^ n4132 ^ 1'b0 ;
  assign n15641 = n8551 & ~n14034 ;
  assign n15652 = n1404 ^ n953 ^ 1'b0 ;
  assign n15642 = n890 & ~n8347 ;
  assign n15643 = n15642 ^ n464 ^ 1'b0 ;
  assign n15644 = n15643 ^ n9634 ^ 1'b0 ;
  assign n15645 = n5278 ^ n3635 ^ 1'b0 ;
  assign n15646 = x39 & ~n15645 ;
  assign n15647 = ( n3956 & n9314 ) | ( n3956 & ~n15646 ) | ( n9314 & ~n15646 ) ;
  assign n15648 = n9961 ^ n3171 ^ n1768 ;
  assign n15649 = n15648 ^ n6907 ^ 1'b0 ;
  assign n15650 = ~n15647 & n15649 ;
  assign n15651 = n15644 & n15650 ;
  assign n15653 = n15652 ^ n15651 ^ 1'b0 ;
  assign n15654 = x3 & n1981 ;
  assign n15655 = n3619 & n6627 ;
  assign n15656 = n9706 | n15655 ;
  assign n15657 = n15654 & ~n15656 ;
  assign n15658 = n15657 ^ n13167 ^ 1'b0 ;
  assign n15659 = ~n1125 & n9552 ;
  assign n15660 = n15177 ^ n305 ^ 1'b0 ;
  assign n15661 = n3601 & n15660 ;
  assign n15662 = n10340 & ~n15661 ;
  assign n15663 = ~n2045 & n4985 ;
  assign n15664 = ~n9280 & n15663 ;
  assign n15665 = n7016 & n15664 ;
  assign n15666 = ~n10759 & n15665 ;
  assign n15667 = x48 & ~n1442 ;
  assign n15668 = ~n13798 & n15667 ;
  assign n15669 = n15668 ^ n2494 ^ 1'b0 ;
  assign n15670 = n6345 | n12409 ;
  assign n15671 = n15669 | n15670 ;
  assign n15672 = ~n5099 & n7496 ;
  assign n15673 = x8 & ~n11610 ;
  assign n15674 = ~n2918 & n15673 ;
  assign n15675 = ~n3034 & n15646 ;
  assign n15676 = n15674 & n15675 ;
  assign n15677 = n15676 ^ n8482 ^ 1'b0 ;
  assign n15678 = ~n11879 & n15677 ;
  assign n15679 = n464 & n6819 ;
  assign n15680 = n15679 ^ n8657 ^ 1'b0 ;
  assign n15681 = n15680 ^ n2091 ^ 1'b0 ;
  assign n15682 = x184 & n15681 ;
  assign n15683 = n15682 ^ n3747 ^ 1'b0 ;
  assign n15684 = n5713 ^ n4647 ^ n1404 ;
  assign n15685 = n992 | n13299 ;
  assign n15686 = n4754 | n15685 ;
  assign n15687 = n8157 & ~n14949 ;
  assign n15688 = ( ~n6739 & n9738 ) | ( ~n6739 & n11854 ) | ( n9738 & n11854 ) ;
  assign n15689 = ~n552 & n922 ;
  assign n15690 = n4637 | n4840 ;
  assign n15691 = n15689 | n15690 ;
  assign n15692 = ( n1006 & n2506 ) | ( n1006 & n4168 ) | ( n2506 & n4168 ) ;
  assign n15693 = ( n1851 & n9216 ) | ( n1851 & ~n15692 ) | ( n9216 & ~n15692 ) ;
  assign n15694 = n15693 ^ n14304 ^ 1'b0 ;
  assign n15695 = n5231 & n12638 ;
  assign n15696 = n15695 ^ n5525 ^ 1'b0 ;
  assign n15697 = n8145 & n15696 ;
  assign n15698 = n10615 & ~n12725 ;
  assign n15699 = ~n3796 & n4985 ;
  assign n15700 = n15699 ^ n4045 ^ 1'b0 ;
  assign n15701 = n1345 ^ x22 ^ 1'b0 ;
  assign n15706 = n7707 ^ n3942 ^ 1'b0 ;
  assign n15707 = n9397 | n15706 ;
  assign n15703 = n5720 ^ n2584 ^ 1'b0 ;
  assign n15702 = n4580 & n6661 ;
  assign n15704 = n15703 ^ n15702 ^ 1'b0 ;
  assign n15705 = n7455 & n15704 ;
  assign n15708 = n15707 ^ n15705 ^ 1'b0 ;
  assign n15709 = n2051 & n5107 ;
  assign n15710 = n3308 & ~n4512 ;
  assign n15711 = n1378 & n15710 ;
  assign n15712 = ~n2799 & n15711 ;
  assign n15713 = n9526 | n15712 ;
  assign n15714 = n7996 | n15713 ;
  assign n15715 = n2533 | n12694 ;
  assign n15716 = ~n10217 & n12347 ;
  assign n15717 = n891 & n14757 ;
  assign n15718 = ~n7822 & n15717 ;
  assign n15719 = ( ~x144 & n1426 ) | ( ~x144 & n7004 ) | ( n1426 & n7004 ) ;
  assign n15720 = n15719 ^ n7330 ^ 1'b0 ;
  assign n15721 = n6109 | n15720 ;
  assign n15722 = x96 & n15721 ;
  assign n15723 = n11268 ^ n3226 ^ 1'b0 ;
  assign n15724 = n6989 & ~n15723 ;
  assign n15725 = ~n5497 & n15724 ;
  assign n15726 = n2143 & ~n15050 ;
  assign n15727 = n4621 & ~n15726 ;
  assign n15728 = n15727 ^ n1510 ^ 1'b0 ;
  assign n15729 = ~n15725 & n15728 ;
  assign n15730 = n7178 ^ n3062 ^ 1'b0 ;
  assign n15731 = n3067 | n8084 ;
  assign n15732 = n15731 ^ n7000 ^ n4621 ;
  assign n15733 = n2297 | n11537 ;
  assign n15734 = x134 & ~n15733 ;
  assign n15735 = n9747 & n15734 ;
  assign n15736 = x90 & n10297 ;
  assign n15737 = n15736 ^ n8964 ^ 1'b0 ;
  assign n15738 = ~n2476 & n2870 ;
  assign n15739 = n4325 | n15738 ;
  assign n15740 = n9862 ^ n5232 ^ 1'b0 ;
  assign n15741 = ~n15739 & n15740 ;
  assign n15742 = n15741 ^ n5369 ^ 1'b0 ;
  assign n15743 = n15737 | n15742 ;
  assign n15746 = n1317 | n5891 ;
  assign n15747 = n10164 & ~n15746 ;
  assign n15744 = ~n7216 & n15128 ;
  assign n15745 = n15744 ^ n2831 ^ 1'b0 ;
  assign n15748 = n15747 ^ n15745 ^ 1'b0 ;
  assign n15749 = n11951 & ~n15748 ;
  assign n15750 = n550 | n4510 ;
  assign n15751 = ~n6520 & n11726 ;
  assign n15752 = n9719 & n15751 ;
  assign n15753 = n15752 ^ n7766 ^ 1'b0 ;
  assign n15754 = n724 | n15753 ;
  assign n15755 = n2654 & n9262 ;
  assign n15756 = n15755 ^ n5497 ^ 1'b0 ;
  assign n15757 = x140 & ~n7652 ;
  assign n15758 = n15757 ^ n13432 ^ 1'b0 ;
  assign n15759 = n8880 ^ x241 ^ 1'b0 ;
  assign n15760 = n3025 & n15759 ;
  assign n15761 = n15760 ^ n11973 ^ 1'b0 ;
  assign n15762 = ~n5079 & n11827 ;
  assign n15763 = n15762 ^ n6646 ^ 1'b0 ;
  assign n15764 = n7196 ^ n367 ^ 1'b0 ;
  assign n15765 = n2706 & n15764 ;
  assign n15766 = ~n3034 & n9383 ;
  assign n15768 = n6270 ^ n1032 ^ 1'b0 ;
  assign n15769 = n6991 & n15768 ;
  assign n15770 = n15769 ^ n8870 ^ 1'b0 ;
  assign n15767 = n923 | n10399 ;
  assign n15771 = n15770 ^ n15767 ^ 1'b0 ;
  assign n15772 = ~n7617 & n15771 ;
  assign n15773 = n2293 ^ n2167 ^ 1'b0 ;
  assign n15774 = n3504 & ~n15773 ;
  assign n15775 = n6088 ^ n4983 ^ n1245 ;
  assign n15776 = n1862 & n15775 ;
  assign n15777 = ~n2740 & n15776 ;
  assign n15778 = n9271 & ~n15777 ;
  assign n15779 = n15778 ^ n1199 ^ 1'b0 ;
  assign n15780 = n11323 ^ n897 ^ 1'b0 ;
  assign n15781 = n6985 & ~n15780 ;
  assign n15782 = n15779 & n15781 ;
  assign n15783 = n2711 & n15782 ;
  assign n15784 = ~x137 & n2232 ;
  assign n15785 = ~n12713 & n15784 ;
  assign n15786 = n15785 ^ n10589 ^ 1'b0 ;
  assign n15787 = ~n15783 & n15786 ;
  assign n15789 = n5446 & ~n11024 ;
  assign n15788 = n4635 & ~n12459 ;
  assign n15790 = n15789 ^ n15788 ^ 1'b0 ;
  assign n15791 = ~n15074 & n15790 ;
  assign n15792 = ~n11055 & n15791 ;
  assign n15793 = n4726 ^ n640 ^ 1'b0 ;
  assign n15794 = n7258 ^ n617 ^ 1'b0 ;
  assign n15795 = n5212 & ~n15794 ;
  assign n15796 = n5146 & ~n11630 ;
  assign n15797 = ~n15795 & n15796 ;
  assign n15798 = n5619 & ~n7712 ;
  assign n15799 = n15798 ^ n15466 ^ 1'b0 ;
  assign n15800 = n4679 & n15277 ;
  assign n15801 = n15800 ^ n12158 ^ 1'b0 ;
  assign n15802 = ~n1463 & n15801 ;
  assign n15803 = n10719 | n15802 ;
  assign n15804 = n6550 ^ n1695 ^ 1'b0 ;
  assign n15805 = n6745 & ~n8604 ;
  assign n15806 = n15805 ^ n12842 ^ 1'b0 ;
  assign n15807 = n15804 | n15806 ;
  assign n15808 = n10536 ^ n2096 ^ 1'b0 ;
  assign n15809 = n15807 | n15808 ;
  assign n15810 = n15809 ^ n2070 ^ 1'b0 ;
  assign n15811 = ~n3850 & n15810 ;
  assign n15812 = ~x48 & n9264 ;
  assign n15813 = n11976 | n13498 ;
  assign n15814 = n15813 ^ n14652 ^ 1'b0 ;
  assign n15815 = n14580 ^ n13056 ^ 1'b0 ;
  assign n15816 = n1121 & n15815 ;
  assign n15817 = n15816 ^ n5340 ^ 1'b0 ;
  assign n15818 = n12146 & n15817 ;
  assign n15819 = n11794 ^ n3521 ^ 1'b0 ;
  assign n15820 = n15819 ^ n5931 ^ 1'b0 ;
  assign n15823 = n4257 | n15804 ;
  assign n15824 = n15823 ^ n3593 ^ 1'b0 ;
  assign n15821 = n3257 & ~n5812 ;
  assign n15822 = n6746 | n15821 ;
  assign n15825 = n15824 ^ n15822 ^ 1'b0 ;
  assign n15826 = n9027 ^ n8668 ^ 1'b0 ;
  assign n15827 = n5189 ^ n4938 ^ 1'b0 ;
  assign n15828 = ~n8506 & n15827 ;
  assign n15829 = n15828 ^ n10172 ^ 1'b0 ;
  assign n15830 = n6278 | n15829 ;
  assign n15831 = n11605 & n14456 ;
  assign n15832 = n15831 ^ n3019 ^ 1'b0 ;
  assign n15835 = n9440 ^ n4149 ^ 1'b0 ;
  assign n15836 = n1036 & n15835 ;
  assign n15833 = n1417 & n8333 ;
  assign n15834 = ~n8577 & n15833 ;
  assign n15837 = n15836 ^ n15834 ^ 1'b0 ;
  assign n15838 = ~n419 & n4610 ;
  assign n15839 = ~n2144 & n15838 ;
  assign n15840 = n8219 | n13920 ;
  assign n15841 = n8845 & ~n15840 ;
  assign n15842 = n5502 & ~n13503 ;
  assign n15843 = x3 & n12989 ;
  assign n15844 = n954 & ~n2594 ;
  assign n15845 = ~n2287 & n15844 ;
  assign n15846 = n11963 ^ n7045 ^ 1'b0 ;
  assign n15847 = n15845 | n15846 ;
  assign n15848 = n271 & ~n6335 ;
  assign n15849 = n15847 & n15848 ;
  assign n15850 = n1589 & n1861 ;
  assign n15851 = n7248 ^ n921 ^ 1'b0 ;
  assign n15852 = n1614 & n15851 ;
  assign n15853 = ~n9456 & n15852 ;
  assign n15854 = ~n9080 & n15853 ;
  assign n15855 = n11532 & ~n15854 ;
  assign n15856 = ~n10911 & n15855 ;
  assign n15857 = ( n6670 & n15850 ) | ( n6670 & n15856 ) | ( n15850 & n15856 ) ;
  assign n15858 = n14815 ^ n11197 ^ 1'b0 ;
  assign n15860 = x212 & ~n11049 ;
  assign n15859 = ~n5749 & n11964 ;
  assign n15861 = n15860 ^ n15859 ^ 1'b0 ;
  assign n15862 = n5754 & ~n10420 ;
  assign n15863 = n15862 ^ n12649 ^ 1'b0 ;
  assign n15864 = n15861 & n15863 ;
  assign n15865 = n15864 ^ n4501 ^ 1'b0 ;
  assign n15866 = n5813 ^ n5169 ^ n473 ;
  assign n15867 = n537 & ~n15866 ;
  assign n15869 = ~n2263 & n3223 ;
  assign n15870 = n15869 ^ n3052 ^ 1'b0 ;
  assign n15871 = n15870 ^ n3518 ^ 1'b0 ;
  assign n15868 = n6225 | n14236 ;
  assign n15872 = n15871 ^ n15868 ^ n790 ;
  assign n15873 = n5749 & n10865 ;
  assign n15874 = n15873 ^ n3018 ^ 1'b0 ;
  assign n15875 = n6128 & n6293 ;
  assign n15876 = n7875 & n15816 ;
  assign n15877 = n15876 ^ n640 ^ 1'b0 ;
  assign n15878 = n7153 & n15877 ;
  assign n15879 = n11687 & n13354 ;
  assign n15880 = ~n13738 & n15879 ;
  assign n15881 = n7296 | n13699 ;
  assign n15882 = n10968 ^ n2174 ^ 1'b0 ;
  assign n15883 = n11483 ^ n6853 ^ 1'b0 ;
  assign n15884 = n6925 ^ n1859 ^ 1'b0 ;
  assign n15885 = n10028 & n15884 ;
  assign n15886 = n15885 ^ n11956 ^ 1'b0 ;
  assign n15887 = ~n6572 & n15886 ;
  assign n15888 = n4553 ^ n4119 ^ 1'b0 ;
  assign n15889 = n3041 | n15888 ;
  assign n15890 = n954 & ~n15889 ;
  assign n15891 = ~n12141 & n15890 ;
  assign n15892 = n9659 & n10800 ;
  assign n15893 = n4185 ^ n911 ^ 1'b0 ;
  assign n15894 = n13474 ^ n10855 ^ n453 ;
  assign n15907 = n11243 ^ n2465 ^ 1'b0 ;
  assign n15905 = x212 & ~n8216 ;
  assign n15899 = n13530 ^ n12046 ^ n2579 ;
  assign n15900 = n15899 ^ n12468 ^ n7426 ;
  assign n15901 = n3666 & ~n8432 ;
  assign n15902 = n15901 ^ n2937 ^ 1'b0 ;
  assign n15903 = ~n15900 & n15902 ;
  assign n15904 = ~n8007 & n15903 ;
  assign n15906 = n15905 ^ n15904 ^ 1'b0 ;
  assign n15908 = n15907 ^ n15906 ^ 1'b0 ;
  assign n15895 = ( n10522 & n12207 ) | ( n10522 & n15208 ) | ( n12207 & n15208 ) ;
  assign n15896 = n4867 | n15895 ;
  assign n15897 = n15896 ^ n15028 ^ 1'b0 ;
  assign n15898 = ~n5189 & n15897 ;
  assign n15909 = n15908 ^ n15898 ^ 1'b0 ;
  assign n15910 = n10472 ^ n7516 ^ n5610 ;
  assign n15911 = n15910 ^ n4003 ^ 1'b0 ;
  assign n15912 = ~n5698 & n7839 ;
  assign n15913 = n10908 & ~n15912 ;
  assign n15914 = n15913 ^ n9311 ^ 1'b0 ;
  assign n15915 = ~n6981 & n15086 ;
  assign n15916 = n10545 & n15915 ;
  assign n15917 = n1422 | n9611 ;
  assign n15918 = n3962 | n15917 ;
  assign n15919 = n11373 ^ n9428 ^ 1'b0 ;
  assign n15920 = n15918 & n15919 ;
  assign n15921 = n13630 & n15920 ;
  assign n15922 = n7810 | n8670 ;
  assign n15923 = n15922 ^ n12519 ^ 1'b0 ;
  assign n15924 = n8063 ^ n8005 ^ 1'b0 ;
  assign n15925 = n4941 ^ n3410 ^ 1'b0 ;
  assign n15926 = n15925 ^ n14760 ^ n2400 ;
  assign n15927 = n15324 ^ n13449 ^ 1'b0 ;
  assign n15928 = ~n12855 & n13155 ;
  assign n15929 = n671 & ~n6585 ;
  assign n15930 = n15929 ^ n13498 ^ n1828 ;
  assign n15931 = n15928 & ~n15930 ;
  assign n15932 = ~n2846 & n10922 ;
  assign n15934 = n8446 ^ x233 ^ 1'b0 ;
  assign n15935 = n1543 & ~n15934 ;
  assign n15936 = n15935 ^ n3683 ^ 1'b0 ;
  assign n15933 = x40 & n467 ;
  assign n15937 = n15936 ^ n15933 ^ 1'b0 ;
  assign n15938 = n4968 ^ x0 ^ 1'b0 ;
  assign n15939 = n1915 & ~n15938 ;
  assign n15940 = n15937 & n15939 ;
  assign n15941 = ~n14714 & n15940 ;
  assign n15942 = n15941 ^ x199 ^ 1'b0 ;
  assign n15943 = n15932 & n15942 ;
  assign n15944 = n13375 ^ n12632 ^ 1'b0 ;
  assign n15945 = n9557 & ~n15944 ;
  assign n15946 = ( ~x28 & n4047 ) | ( ~x28 & n5120 ) | ( n4047 & n5120 ) ;
  assign n15947 = n6187 | n15946 ;
  assign n15948 = n7351 & ~n15947 ;
  assign n15949 = n12828 | n15948 ;
  assign n15950 = n15949 ^ n15496 ^ 1'b0 ;
  assign n15951 = ~n928 & n3235 ;
  assign n15952 = n15951 ^ x70 ^ 1'b0 ;
  assign n15953 = ~n1467 & n15952 ;
  assign n15954 = n11659 ^ n7404 ^ 1'b0 ;
  assign n15955 = n1621 | n10111 ;
  assign n15956 = ~n9332 & n9836 ;
  assign n15957 = n14699 ^ n6281 ^ 1'b0 ;
  assign n15958 = n9457 ^ n8682 ^ n713 ;
  assign n15959 = n6442 & n7779 ;
  assign n15960 = n15959 ^ n11725 ^ 1'b0 ;
  assign n15961 = n12476 ^ n6689 ^ 1'b0 ;
  assign n15962 = n12455 ^ n4872 ^ 1'b0 ;
  assign n15963 = n9232 & n15962 ;
  assign n15964 = n15961 & n15963 ;
  assign n15965 = n7096 & n15663 ;
  assign n15966 = n15965 ^ n4985 ^ 1'b0 ;
  assign n15967 = ( n7594 & n14640 ) | ( n7594 & n15966 ) | ( n14640 & n15966 ) ;
  assign n15969 = n9501 ^ n2106 ^ 1'b0 ;
  assign n15968 = n7538 | n12131 ;
  assign n15970 = n15969 ^ n15968 ^ n13651 ;
  assign n15971 = n14276 ^ n12943 ^ n7876 ;
  assign n15972 = n6331 | n15971 ;
  assign n15973 = n15972 ^ n7702 ^ 1'b0 ;
  assign n15974 = n6921 | n11345 ;
  assign n15975 = n15974 ^ n6842 ^ 1'b0 ;
  assign n15976 = ( n2448 & n2647 ) | ( n2448 & n2747 ) | ( n2647 & n2747 ) ;
  assign n15977 = n15976 ^ n3298 ^ 1'b0 ;
  assign n15978 = ~n1424 & n3951 ;
  assign n15979 = n15978 ^ n6202 ^ 1'b0 ;
  assign n15980 = n15977 | n15979 ;
  assign n15981 = n12842 & ~n15980 ;
  assign n15982 = n11526 ^ n1383 ^ 1'b0 ;
  assign n15983 = n12022 & ~n15982 ;
  assign n15989 = ( n1725 & ~n1729 ) | ( n1725 & n1968 ) | ( ~n1729 & n1968 ) ;
  assign n15990 = n13095 & ~n15989 ;
  assign n15991 = n15990 ^ n6293 ^ 1'b0 ;
  assign n15984 = n2177 | n10827 ;
  assign n15985 = n8983 ^ n4144 ^ n4062 ;
  assign n15986 = n15187 & n15985 ;
  assign n15987 = n15984 & n15986 ;
  assign n15988 = n13579 & ~n15987 ;
  assign n15992 = n15991 ^ n15988 ^ 1'b0 ;
  assign n15993 = n15624 ^ n4142 ^ 1'b0 ;
  assign n15994 = ~n1912 & n7238 ;
  assign n15995 = ~n923 & n15994 ;
  assign n15996 = ~n2027 & n15995 ;
  assign n15997 = n15996 ^ n6421 ^ 1'b0 ;
  assign n15998 = n7393 & ~n15997 ;
  assign n15999 = ( ~n6433 & n14462 ) | ( ~n6433 & n15809 ) | ( n14462 & n15809 ) ;
  assign n16000 = n12394 ^ n7168 ^ 1'b0 ;
  assign n16001 = n12426 & n16000 ;
  assign n16002 = n4381 | n12719 ;
  assign n16003 = n3933 | n16002 ;
  assign n16004 = n4409 ^ n2143 ^ 1'b0 ;
  assign n16005 = n16003 & n16004 ;
  assign n16006 = ( n7623 & n13091 ) | ( n7623 & ~n16005 ) | ( n13091 & ~n16005 ) ;
  assign n16009 = n399 | n2521 ;
  assign n16010 = n1051 & ~n16009 ;
  assign n16007 = ~n4238 & n6012 ;
  assign n16008 = n16007 ^ n6358 ^ 1'b0 ;
  assign n16011 = n16010 ^ n16008 ^ 1'b0 ;
  assign n16012 = ~n13675 & n16011 ;
  assign n16013 = ~n5813 & n16012 ;
  assign n16014 = n16013 ^ n9511 ^ 1'b0 ;
  assign n16015 = n11035 | n14044 ;
  assign n16016 = n3904 & n9076 ;
  assign n16017 = n3956 | n8991 ;
  assign n16018 = n786 & n10345 ;
  assign n16032 = n6674 ^ n4521 ^ 1'b0 ;
  assign n16022 = n2817 & n10534 ;
  assign n16023 = n3561 ^ n1709 ^ 1'b0 ;
  assign n16024 = ~n1521 & n16023 ;
  assign n16025 = n16024 ^ n7013 ^ 1'b0 ;
  assign n16026 = n16025 ^ n3249 ^ 1'b0 ;
  assign n16027 = n10333 & n16026 ;
  assign n16028 = n7518 & n16027 ;
  assign n16029 = n16022 & ~n16028 ;
  assign n16030 = ~n8518 & n16029 ;
  assign n16019 = n7054 ^ n6912 ^ n1160 ;
  assign n16020 = n13433 & ~n16019 ;
  assign n16021 = n9594 & ~n16020 ;
  assign n16031 = n16030 ^ n16021 ^ 1'b0 ;
  assign n16033 = n16032 ^ n16031 ^ n8413 ;
  assign n16034 = n3603 ^ n1138 ^ 1'b0 ;
  assign n16035 = n6972 & ~n16034 ;
  assign n16036 = n5711 & ~n9783 ;
  assign n16037 = ~n16035 & n16036 ;
  assign n16041 = n3235 & ~n4388 ;
  assign n16042 = n16041 ^ n3959 ^ 1'b0 ;
  assign n16043 = n16042 ^ n8034 ^ 1'b0 ;
  assign n16044 = ~n5326 & n16043 ;
  assign n16038 = ( n3500 & n4380 ) | ( n3500 & ~n4589 ) | ( n4380 & ~n4589 ) ;
  assign n16039 = n16038 ^ n13363 ^ x106 ;
  assign n16040 = n9961 & ~n16039 ;
  assign n16045 = n16044 ^ n16040 ^ 1'b0 ;
  assign n16046 = n867 & ~n13297 ;
  assign n16047 = n16046 ^ n8200 ^ 1'b0 ;
  assign n16048 = ~n2525 & n11614 ;
  assign n16049 = n16048 ^ n3104 ^ 1'b0 ;
  assign n16052 = ~n589 & n10952 ;
  assign n16053 = n589 & n16052 ;
  assign n16054 = n941 | n16053 ;
  assign n16055 = n16053 & ~n16054 ;
  assign n16056 = n4027 & ~n16055 ;
  assign n16050 = ~n1969 & n13590 ;
  assign n16051 = ~n15809 & n16050 ;
  assign n16057 = n16056 ^ n16051 ^ 1'b0 ;
  assign n16058 = n3551 ^ n1208 ^ 1'b0 ;
  assign n16059 = n11512 & n16058 ;
  assign n16060 = ~n11285 & n16059 ;
  assign n16061 = n16060 ^ n10867 ^ 1'b0 ;
  assign n16062 = n6339 & n16061 ;
  assign n16069 = n4525 ^ n1395 ^ 1'b0 ;
  assign n16063 = n3001 & ~n7573 ;
  assign n16064 = ~x24 & n16063 ;
  assign n16065 = n6155 | n16064 ;
  assign n16066 = n507 & ~n16065 ;
  assign n16067 = n903 | n16066 ;
  assign n16068 = n276 & ~n16067 ;
  assign n16070 = n16069 ^ n16068 ^ 1'b0 ;
  assign n16071 = n5206 ^ n4516 ^ 1'b0 ;
  assign n16072 = n1208 ^ n1174 ^ 1'b0 ;
  assign n16073 = ( n3563 & n5043 ) | ( n3563 & ~n16072 ) | ( n5043 & ~n16072 ) ;
  assign n16074 = ( ~n1912 & n6446 ) | ( ~n1912 & n16073 ) | ( n6446 & n16073 ) ;
  assign n16075 = n1064 | n7828 ;
  assign n16076 = n4375 | n16075 ;
  assign n16077 = n16074 & ~n16076 ;
  assign n16078 = n8280 ^ n5406 ^ 1'b0 ;
  assign n16079 = n6177 & n7560 ;
  assign n16080 = n5160 & n11230 ;
  assign n16081 = ( n5855 & n8809 ) | ( n5855 & ~n16080 ) | ( n8809 & ~n16080 ) ;
  assign n16082 = n7679 & n16081 ;
  assign n16086 = n8501 | n10991 ;
  assign n16087 = n4316 & ~n16086 ;
  assign n16088 = n4720 & ~n16087 ;
  assign n16083 = ( n3598 & n4497 ) | ( n3598 & n8070 ) | ( n4497 & n8070 ) ;
  assign n16084 = n16083 ^ n3137 ^ 1'b0 ;
  assign n16085 = n2686 & n16084 ;
  assign n16089 = n16088 ^ n16085 ^ 1'b0 ;
  assign n16090 = n11360 | n16089 ;
  assign n16092 = n10391 ^ n5893 ^ 1'b0 ;
  assign n16091 = n13821 ^ n2091 ^ 1'b0 ;
  assign n16093 = n16092 ^ n16091 ^ n8814 ;
  assign n16094 = n12228 ^ n7623 ^ 1'b0 ;
  assign n16095 = n9209 & ~n16094 ;
  assign n16096 = n16095 ^ n15688 ^ 1'b0 ;
  assign n16097 = n4117 ^ n2003 ^ 1'b0 ;
  assign n16098 = ~n2809 & n16097 ;
  assign n16099 = ~n3335 & n3378 ;
  assign n16100 = n3657 & n16099 ;
  assign n16101 = n16100 ^ n6090 ^ n4826 ;
  assign n16102 = n1922 | n14327 ;
  assign n16103 = n3479 & n10331 ;
  assign n16104 = n16103 ^ n5461 ^ 1'b0 ;
  assign n16105 = n3368 & ~n10687 ;
  assign n16106 = n16104 & ~n16105 ;
  assign n16107 = n2681 | n5957 ;
  assign n16108 = n5560 | n16107 ;
  assign n16109 = ~n9293 & n16108 ;
  assign n16110 = n3823 & ~n8072 ;
  assign n16111 = n10277 & n16110 ;
  assign n16112 = n16111 ^ n11730 ^ 1'b0 ;
  assign n16113 = n2320 | n2741 ;
  assign n16114 = ~n8843 & n16113 ;
  assign n16115 = n4078 ^ n3323 ^ 1'b0 ;
  assign n16116 = n16114 & n16115 ;
  assign n16117 = n9350 ^ n2728 ^ 1'b0 ;
  assign n16118 = n11450 & n16117 ;
  assign n16119 = ~n7175 & n7490 ;
  assign n16120 = n16119 ^ n1729 ^ 1'b0 ;
  assign n16121 = n16118 & n16120 ;
  assign n16122 = n16121 ^ n13800 ^ 1'b0 ;
  assign n16123 = n2964 ^ n407 ^ 1'b0 ;
  assign n16124 = n4931 & n16123 ;
  assign n16125 = n8784 & n16124 ;
  assign n16126 = n6797 & ~n15744 ;
  assign n16127 = n4029 ^ n614 ^ 1'b0 ;
  assign n16128 = ~n6295 & n16127 ;
  assign n16129 = n16128 ^ n1001 ^ 1'b0 ;
  assign n16130 = n7222 & ~n16129 ;
  assign n16131 = n16130 ^ n4520 ^ 1'b0 ;
  assign n16132 = n6271 & n13845 ;
  assign n16133 = n12940 ^ n4865 ^ 1'b0 ;
  assign n16134 = n5063 | n16133 ;
  assign n16135 = n990 & n7242 ;
  assign n16136 = n1830 & ~n16135 ;
  assign n16137 = ~n8582 & n16136 ;
  assign n16138 = n15801 & ~n16137 ;
  assign n16139 = n13090 ^ n4234 ^ n274 ;
  assign n16140 = n359 & ~n908 ;
  assign n16141 = ( n13343 & ~n15858 ) | ( n13343 & n16140 ) | ( ~n15858 & n16140 ) ;
  assign n16142 = n4861 ^ n2073 ^ 1'b0 ;
  assign n16144 = n4402 ^ n689 ^ 1'b0 ;
  assign n16145 = n12111 | n16144 ;
  assign n16143 = ~n10112 & n12552 ;
  assign n16146 = n16145 ^ n16143 ^ 1'b0 ;
  assign n16147 = n1085 & ~n7340 ;
  assign n16148 = n16147 ^ n5895 ^ 1'b0 ;
  assign n16149 = ~n2191 & n8762 ;
  assign n16150 = x89 | n8751 ;
  assign n16151 = n14787 & n16150 ;
  assign n16152 = ~n4108 & n16151 ;
  assign n16153 = n8386 ^ n2873 ^ 1'b0 ;
  assign n16154 = n16153 ^ n3558 ^ 1'b0 ;
  assign n16155 = n13019 ^ n9846 ^ 1'b0 ;
  assign n16156 = ~n7722 & n16155 ;
  assign n16157 = n5232 ^ n2837 ^ 1'b0 ;
  assign n16158 = n10552 & ~n16157 ;
  assign n16159 = n14235 ^ n5475 ^ 1'b0 ;
  assign n16160 = n2735 | n16159 ;
  assign n16161 = n13193 ^ n12677 ^ 1'b0 ;
  assign n16162 = ~n872 & n16161 ;
  assign n16163 = n13404 ^ n2514 ^ 1'b0 ;
  assign n16164 = ~n3022 & n16163 ;
  assign n16165 = n9352 & ~n12569 ;
  assign n16166 = ~n4360 & n6106 ;
  assign n16167 = n16166 ^ n11608 ^ 1'b0 ;
  assign n16168 = ~n2653 & n9063 ;
  assign n16169 = ~n8034 & n12314 ;
  assign n16170 = n10971 & n16169 ;
  assign n16171 = ~n5571 & n14283 ;
  assign n16172 = ~n3895 & n10619 ;
  assign n16173 = n4014 & n4964 ;
  assign n16174 = n4534 & n16173 ;
  assign n16175 = n366 & ~n16174 ;
  assign n16176 = n16175 ^ n6920 ^ 1'b0 ;
  assign n16177 = n16176 ^ n14136 ^ 1'b0 ;
  assign n16178 = n16153 | n16177 ;
  assign n16179 = n2332 & ~n4074 ;
  assign n16180 = ~n5459 & n16179 ;
  assign n16181 = ~n532 & n13366 ;
  assign n16182 = n12842 ^ n2703 ^ 1'b0 ;
  assign n16183 = n9976 & n16182 ;
  assign n16184 = n11776 | n13423 ;
  assign n16185 = n941 & ~n5054 ;
  assign n16186 = n2817 & ~n6386 ;
  assign n16187 = ~n5922 & n16186 ;
  assign n16188 = n4650 | n7263 ;
  assign n16189 = n466 | n16188 ;
  assign n16190 = n5316 | n7521 ;
  assign n16191 = n16189 | n16190 ;
  assign n16192 = n13689 ^ n10827 ^ 1'b0 ;
  assign n16193 = n9992 | n16192 ;
  assign n16194 = n16193 ^ n2655 ^ 1'b0 ;
  assign n16195 = n16191 & ~n16194 ;
  assign n16196 = n8999 & ~n16195 ;
  assign n16197 = n7224 ^ n4276 ^ 1'b0 ;
  assign n16198 = ~n13867 & n16197 ;
  assign n16199 = n12789 & n13969 ;
  assign n16200 = n16199 ^ n890 ^ 1'b0 ;
  assign n16204 = n14572 ^ n9285 ^ 1'b0 ;
  assign n16201 = n784 & n2369 ;
  assign n16202 = n16201 ^ n5812 ^ 1'b0 ;
  assign n16203 = n15767 & ~n16202 ;
  assign n16205 = n16204 ^ n16203 ^ 1'b0 ;
  assign n16206 = n12451 & n16205 ;
  assign n16207 = ~n4405 & n16206 ;
  assign n16208 = n16207 ^ n6348 ^ 1'b0 ;
  assign n16209 = n1309 ^ n328 ^ 1'b0 ;
  assign n16211 = n3062 & n13740 ;
  assign n16212 = ~n2827 & n16211 ;
  assign n16210 = n863 & ~n5284 ;
  assign n16213 = n16212 ^ n16210 ^ n2227 ;
  assign n16214 = x83 & ~n7566 ;
  assign n16215 = n12240 & n16214 ;
  assign n16216 = n14120 ^ n2130 ^ n796 ;
  assign n16220 = ~n384 & n7748 ;
  assign n16221 = ~n11542 & n16220 ;
  assign n16217 = n12680 ^ n4821 ^ n3614 ;
  assign n16218 = n2154 & ~n16217 ;
  assign n16219 = ~n10485 & n16218 ;
  assign n16222 = n16221 ^ n16219 ^ 1'b0 ;
  assign n16223 = n16222 ^ n5876 ^ 1'b0 ;
  assign n16227 = n15941 ^ n3753 ^ 1'b0 ;
  assign n16224 = n709 & n14117 ;
  assign n16225 = n16224 ^ n4357 ^ 1'b0 ;
  assign n16226 = n3678 | n16225 ;
  assign n16228 = n16227 ^ n16226 ^ 1'b0 ;
  assign n16229 = n14097 ^ n11245 ^ 1'b0 ;
  assign n16230 = n13083 | n16229 ;
  assign n16231 = x159 | n2098 ;
  assign n16232 = n2306 | n16231 ;
  assign n16233 = n16232 ^ n13452 ^ 1'b0 ;
  assign n16234 = n1757 ^ n1393 ^ 1'b0 ;
  assign n16235 = n14936 & n16234 ;
  assign n16236 = ( n2946 & n11590 ) | ( n2946 & n16235 ) | ( n11590 & n16235 ) ;
  assign n16237 = n5675 ^ n3904 ^ 1'b0 ;
  assign n16238 = n2114 & ~n5264 ;
  assign n16239 = n12038 & n16238 ;
  assign n16240 = n3165 & n16239 ;
  assign n16241 = n16237 & ~n16240 ;
  assign n16242 = n6666 ^ n1045 ^ 1'b0 ;
  assign n16243 = x203 & ~n16242 ;
  assign n16244 = ~n264 & n16243 ;
  assign n16245 = x207 & n3903 ;
  assign n16246 = n3724 & n16245 ;
  assign n16247 = n16246 ^ n10503 ^ x43 ;
  assign n16248 = n10554 ^ n3957 ^ 1'b0 ;
  assign n16249 = n7024 & n9375 ;
  assign n16250 = n7813 | n16249 ;
  assign n16251 = n14705 & ~n16250 ;
  assign n16252 = n13917 & n16251 ;
  assign n16253 = ~n3111 & n14618 ;
  assign n16254 = ~n10557 & n16253 ;
  assign n16256 = n6294 & ~n8668 ;
  assign n16255 = n9420 ^ n4903 ^ n3601 ;
  assign n16257 = n16256 ^ n16255 ^ n11818 ;
  assign n16258 = n15319 ^ n7441 ^ 1'b0 ;
  assign n16259 = n16257 & ~n16258 ;
  assign n16260 = ( ~n2592 & n3861 ) | ( ~n2592 & n16259 ) | ( n3861 & n16259 ) ;
  assign n16261 = n14968 ^ n2706 ^ 1'b0 ;
  assign n16262 = n9944 & ~n16261 ;
  assign n16263 = n4985 & n16262 ;
  assign n16264 = ~n7083 & n16263 ;
  assign n16265 = n16264 ^ n15391 ^ 1'b0 ;
  assign n16266 = n2433 | n16265 ;
  assign n16267 = ( n6524 & ~n7629 ) | ( n6524 & n8322 ) | ( ~n7629 & n8322 ) ;
  assign n16268 = n4325 & ~n16267 ;
  assign n16269 = n5639 & n16268 ;
  assign n16270 = ~n3419 & n9280 ;
  assign n16271 = n16270 ^ n15145 ^ 1'b0 ;
  assign n16272 = n5621 & n16271 ;
  assign n16273 = n16272 ^ n5080 ^ 1'b0 ;
  assign n16274 = ~n5404 & n16273 ;
  assign n16275 = n752 & n16274 ;
  assign n16276 = n11774 & ~n16140 ;
  assign n16277 = n3216 ^ n596 ^ 1'b0 ;
  assign n16278 = n1812 ^ n1417 ^ 1'b0 ;
  assign n16279 = n8559 & ~n16278 ;
  assign n16280 = n16279 ^ n11372 ^ 1'b0 ;
  assign n16281 = n5642 ^ n4896 ^ 1'b0 ;
  assign n16282 = n3151 | n4510 ;
  assign n16283 = n16282 ^ n6067 ^ 1'b0 ;
  assign n16284 = ( n1813 & n9976 ) | ( n1813 & n11858 ) | ( n9976 & n11858 ) ;
  assign n16285 = n4546 ^ n2131 ^ x129 ;
  assign n16286 = n16285 ^ n9471 ^ 1'b0 ;
  assign n16287 = n684 | n3449 ;
  assign n16288 = n16287 ^ n1021 ^ 1'b0 ;
  assign n16289 = n5409 & ~n16288 ;
  assign n16290 = n6694 & n16289 ;
  assign n16291 = n16290 ^ n1298 ^ 1'b0 ;
  assign n16292 = n6336 | n16291 ;
  assign n16293 = n1659 | n16292 ;
  assign n16294 = n16293 ^ n1948 ^ 1'b0 ;
  assign n16295 = n6619 & ~n16294 ;
  assign n16296 = n9367 ^ n1602 ^ 1'b0 ;
  assign n16297 = n16296 ^ n15798 ^ 1'b0 ;
  assign n16298 = ~n6327 & n8417 ;
  assign n16299 = ~n3643 & n16298 ;
  assign n16300 = n15366 ^ n3670 ^ 1'b0 ;
  assign n16301 = n1435 & ~n6657 ;
  assign n16302 = n5406 & ~n8067 ;
  assign n16303 = n16302 ^ n6439 ^ 1'b0 ;
  assign n16304 = ~n9149 & n16303 ;
  assign n16305 = n11749 ^ n10036 ^ n6005 ;
  assign n16306 = n1084 | n3165 ;
  assign n16307 = n16306 ^ n1536 ^ 1'b0 ;
  assign n16308 = ~n11414 & n16307 ;
  assign n16309 = n14276 ^ x112 ^ 1'b0 ;
  assign n16310 = ~n12161 & n13743 ;
  assign n16311 = ~n2110 & n16310 ;
  assign n16312 = n3380 & ~n10692 ;
  assign n16313 = n1404 & n16312 ;
  assign n16317 = n14458 ^ n9986 ^ 1'b0 ;
  assign n16318 = n6325 & n16317 ;
  assign n16314 = n1286 | n8083 ;
  assign n16315 = n16314 ^ n14851 ^ 1'b0 ;
  assign n16316 = x136 & n16315 ;
  assign n16319 = n16318 ^ n16316 ^ 1'b0 ;
  assign n16320 = n12869 ^ n8536 ^ 1'b0 ;
  assign n16321 = n1846 | n3899 ;
  assign n16322 = n13545 ^ n294 ^ 1'b0 ;
  assign n16323 = n13291 ^ n4078 ^ 1'b0 ;
  assign n16324 = ~n4737 & n16323 ;
  assign n16325 = n7407 & n11361 ;
  assign n16326 = n16325 ^ n5932 ^ 1'b0 ;
  assign n16327 = n15819 ^ n9673 ^ n2161 ;
  assign n16328 = n2949 ^ n2308 ^ 1'b0 ;
  assign n16329 = n2148 & n16328 ;
  assign n16330 = n2855 & ~n9243 ;
  assign n16331 = ~n7058 & n16330 ;
  assign n16332 = ~n16074 & n16331 ;
  assign n16333 = n9683 ^ n589 ^ 1'b0 ;
  assign n16334 = n16333 ^ n16166 ^ 1'b0 ;
  assign n16338 = n1154 & ~n7428 ;
  assign n16339 = ~n13193 & n16338 ;
  assign n16340 = ( n12542 & n16137 ) | ( n12542 & n16339 ) | ( n16137 & n16339 ) ;
  assign n16335 = ~n9621 & n13429 ;
  assign n16336 = ~n12557 & n16335 ;
  assign n16337 = x110 & ~n16336 ;
  assign n16341 = n16340 ^ n16337 ^ 1'b0 ;
  assign n16342 = n2326 ^ x147 ^ 1'b0 ;
  assign n16343 = n5948 ^ n4270 ^ 1'b0 ;
  assign n16344 = n12515 ^ n6091 ^ 1'b0 ;
  assign n16345 = ( n8632 & n8751 ) | ( n8632 & ~n9228 ) | ( n8751 & ~n9228 ) ;
  assign n16346 = x135 & ~n16345 ;
  assign n16347 = n2404 & n2668 ;
  assign n16348 = n1203 & n16347 ;
  assign n16349 = n801 | n16348 ;
  assign n16350 = n2679 | n16349 ;
  assign n16351 = ~n3455 & n16350 ;
  assign n16352 = ~n16346 & n16351 ;
  assign n16353 = n16352 ^ n11013 ^ 1'b0 ;
  assign n16354 = n3806 ^ n3745 ^ 1'b0 ;
  assign n16355 = n16353 | n16354 ;
  assign n16356 = n12979 ^ n12840 ^ 1'b0 ;
  assign n16357 = ~n5992 & n9569 ;
  assign n16358 = n16357 ^ n9343 ^ 1'b0 ;
  assign n16359 = ~n491 & n16358 ;
  assign n16360 = n16359 ^ n3863 ^ 1'b0 ;
  assign n16361 = n16360 ^ n13347 ^ 1'b0 ;
  assign n16362 = n6017 | n8495 ;
  assign n16363 = ~n2385 & n4374 ;
  assign n16364 = n4242 ^ n2471 ^ 1'b0 ;
  assign n16365 = n16363 & n16364 ;
  assign n16366 = n16365 ^ n8547 ^ 1'b0 ;
  assign n16367 = n7709 | n8075 ;
  assign n16368 = n7757 | n16367 ;
  assign n16369 = n2900 & n9357 ;
  assign n16370 = n16369 ^ n3465 ^ 1'b0 ;
  assign n16371 = n16370 ^ n13095 ^ 1'b0 ;
  assign n16372 = n3086 ^ n2192 ^ 1'b0 ;
  assign n16373 = n13362 ^ n6208 ^ 1'b0 ;
  assign n16374 = n13483 ^ n8886 ^ n5392 ;
  assign n16375 = n16374 ^ n2120 ^ 1'b0 ;
  assign n16376 = n4269 ^ x13 ^ 1'b0 ;
  assign n16377 = n2116 & n16376 ;
  assign n16378 = n5664 & n16377 ;
  assign n16379 = n4906 & n16378 ;
  assign n16380 = n10700 ^ n8268 ^ 1'b0 ;
  assign n16382 = n7470 ^ n5637 ^ 1'b0 ;
  assign n16383 = n6030 | n16382 ;
  assign n16384 = ( n1742 & ~n3421 ) | ( n1742 & n10523 ) | ( ~n3421 & n10523 ) ;
  assign n16385 = n16383 | n16384 ;
  assign n16381 = n4679 & ~n8651 ;
  assign n16386 = n16385 ^ n16381 ^ 1'b0 ;
  assign n16387 = ~n1426 & n8557 ;
  assign n16388 = ~n15160 & n16387 ;
  assign n16389 = n8700 | n9883 ;
  assign n16390 = n16389 ^ n4520 ^ 1'b0 ;
  assign n16391 = n2728 & n4313 ;
  assign n16392 = n16391 ^ n14926 ^ 1'b0 ;
  assign n16393 = n799 | n16392 ;
  assign n16394 = n2203 | n15406 ;
  assign n16395 = n2951 | n16394 ;
  assign n16396 = ~n4264 & n11834 ;
  assign n16397 = n274 | n3830 ;
  assign n16398 = n16396 | n16397 ;
  assign n16399 = n2961 | n4388 ;
  assign n16400 = n16398 & ~n16399 ;
  assign n16401 = n16400 ^ n8664 ^ 1'b0 ;
  assign n16402 = n1931 & ~n13905 ;
  assign n16403 = n2743 | n16402 ;
  assign n16404 = ~n1521 & n7545 ;
  assign n16405 = ~n580 & n1138 ;
  assign n16406 = ~n4175 & n16405 ;
  assign n16407 = n16406 ^ n6664 ^ 1'b0 ;
  assign n16408 = n7851 ^ n1838 ^ 1'b0 ;
  assign n16409 = n8668 & n16408 ;
  assign n16410 = ~n11680 & n16409 ;
  assign n16411 = n14787 & ~n16410 ;
  assign n16412 = n16411 ^ n10157 ^ 1'b0 ;
  assign n16415 = n8079 ^ n1921 ^ 1'b0 ;
  assign n16413 = ( n7038 & ~n8315 ) | ( n7038 & n9600 ) | ( ~n8315 & n9600 ) ;
  assign n16414 = ~n5018 & n16413 ;
  assign n16416 = n16415 ^ n16414 ^ 1'b0 ;
  assign n16417 = n3431 & ~n6118 ;
  assign n16418 = n4202 | n16417 ;
  assign n16419 = n16418 ^ n7032 ^ 1'b0 ;
  assign n16420 = n6324 ^ n810 ^ 1'b0 ;
  assign n16421 = n14281 ^ n5840 ^ n5511 ;
  assign n16422 = n1820 & n7321 ;
  assign n16423 = n16422 ^ n882 ^ 1'b0 ;
  assign n16424 = n5039 ^ n692 ^ 1'b0 ;
  assign n16425 = n16424 ^ n2240 ^ 1'b0 ;
  assign n16429 = n407 & ~n2228 ;
  assign n16426 = n661 | n3913 ;
  assign n16427 = n5986 | n16426 ;
  assign n16428 = n16427 ^ n7904 ^ 1'b0 ;
  assign n16430 = n16429 ^ n16428 ^ n5273 ;
  assign n16431 = n7448 & ~n9507 ;
  assign n16432 = n7119 | n16431 ;
  assign n16433 = n16432 ^ n903 ^ 1'b0 ;
  assign n16434 = n3231 ^ n393 ^ 1'b0 ;
  assign n16435 = ~n16433 & n16434 ;
  assign n16436 = n3986 | n14514 ;
  assign n16437 = n2570 & ~n3688 ;
  assign n16438 = n2001 & n16437 ;
  assign n16439 = n10041 & ~n16438 ;
  assign n16440 = ( n1931 & n13231 ) | ( n1931 & n16439 ) | ( n13231 & n16439 ) ;
  assign n16441 = n4119 | n9552 ;
  assign n16442 = n7197 & n16441 ;
  assign n16443 = n9582 | n15631 ;
  assign n16444 = n3232 & n15204 ;
  assign n16445 = ( ~n13480 & n16443 ) | ( ~n13480 & n16444 ) | ( n16443 & n16444 ) ;
  assign n16446 = n9267 ^ n2178 ^ n1979 ;
  assign n16447 = n16446 ^ n5298 ^ 1'b0 ;
  assign n16449 = n4844 | n10470 ;
  assign n16448 = n3959 & n6469 ;
  assign n16450 = n16449 ^ n16448 ^ 1'b0 ;
  assign n16451 = x169 & ~n3397 ;
  assign n16452 = ~n13352 & n16451 ;
  assign n16453 = n4134 & ~n16452 ;
  assign n16454 = ~n8455 & n9224 ;
  assign n16455 = ~n10034 & n16454 ;
  assign n16456 = n7229 ^ n1258 ^ 1'b0 ;
  assign n16457 = n15290 ^ n3154 ^ 1'b0 ;
  assign n16458 = n2297 ^ n1563 ^ 1'b0 ;
  assign n16459 = n2507 & ~n16458 ;
  assign n16460 = n15638 & n16459 ;
  assign n16461 = n7443 & n15500 ;
  assign n16462 = n10520 & n16461 ;
  assign n16463 = n16462 ^ n2722 ^ 1'b0 ;
  assign n16464 = n466 | n987 ;
  assign n16465 = n5479 & n7349 ;
  assign n16466 = n16464 & n16465 ;
  assign n16467 = n2418 & ~n4649 ;
  assign n16468 = n908 & n3264 ;
  assign n16469 = n16468 ^ n9273 ^ 1'b0 ;
  assign n16470 = n16467 & n16469 ;
  assign n16471 = n16470 ^ n14703 ^ 1'b0 ;
  assign n16472 = n13976 & n15080 ;
  assign n16473 = n16471 & n16472 ;
  assign n16474 = n16473 ^ n3293 ^ 1'b0 ;
  assign n16475 = ( n3372 & n5659 ) | ( n3372 & ~n6607 ) | ( n5659 & ~n6607 ) ;
  assign n16476 = n3340 ^ n338 ^ 1'b0 ;
  assign n16477 = n3160 & n16476 ;
  assign n16478 = n10730 ^ n7118 ^ 1'b0 ;
  assign n16479 = n7890 | n8780 ;
  assign n16480 = n5697 & n5797 ;
  assign n16481 = n5650 ^ n2043 ^ 1'b0 ;
  assign n16482 = n9793 & n16481 ;
  assign n16483 = ~n3678 & n16482 ;
  assign n16484 = n16483 ^ n4159 ^ 1'b0 ;
  assign n16485 = n16480 & n16484 ;
  assign n16486 = n6346 & n16485 ;
  assign n16488 = n4449 & n7511 ;
  assign n16489 = ~n3684 & n16488 ;
  assign n16487 = ~n393 & n5967 ;
  assign n16490 = n16489 ^ n16487 ^ n547 ;
  assign n16491 = n3151 & n4953 ;
  assign n16492 = ( n2568 & n8005 ) | ( n2568 & n16491 ) | ( n8005 & n16491 ) ;
  assign n16493 = n5596 & ~n6357 ;
  assign n16494 = n9704 & n10965 ;
  assign n16495 = n7072 ^ n3021 ^ 1'b0 ;
  assign n16496 = n16495 ^ n6826 ^ n2020 ;
  assign n16497 = n5668 & n16496 ;
  assign n16498 = n1219 & n7547 ;
  assign n16499 = ~n2538 & n16498 ;
  assign n16500 = n16499 ^ n8845 ^ 1'b0 ;
  assign n16501 = n11988 ^ n991 ^ 1'b0 ;
  assign n16502 = n738 & ~n16501 ;
  assign n16503 = n16502 ^ n1148 ^ 1'b0 ;
  assign n16504 = n915 & n16503 ;
  assign n16505 = n16504 ^ n16047 ^ 1'b0 ;
  assign n16506 = n258 & ~n9813 ;
  assign n16507 = n2911 | n16506 ;
  assign n16508 = n3007 & ~n16507 ;
  assign n16509 = n1249 & n16508 ;
  assign n16510 = n14373 ^ n9578 ^ 1'b0 ;
  assign n16511 = n3568 & n16510 ;
  assign n16512 = ~n6719 & n9466 ;
  assign n16513 = ~n1032 & n16512 ;
  assign n16514 = n1684 & n8011 ;
  assign n16515 = n16514 ^ n5479 ^ 1'b0 ;
  assign n16516 = n16515 ^ n1328 ^ 1'b0 ;
  assign n16517 = n16513 | n16516 ;
  assign n16520 = n2103 | n3751 ;
  assign n16521 = n16520 ^ x195 ^ 1'b0 ;
  assign n16518 = n1935 & n7392 ;
  assign n16519 = ~n14525 & n16518 ;
  assign n16522 = n16521 ^ n16519 ^ 1'b0 ;
  assign n16524 = n4186 ^ n3600 ^ 1'b0 ;
  assign n16523 = n4844 & ~n9386 ;
  assign n16525 = n16524 ^ n16523 ^ n9549 ;
  assign n16526 = ~x100 & n9903 ;
  assign n16527 = ( n2426 & ~n4521 ) | ( n2426 & n8591 ) | ( ~n4521 & n8591 ) ;
  assign n16528 = ( n14588 & n16526 ) | ( n14588 & n16527 ) | ( n16526 & n16527 ) ;
  assign n16529 = n3892 | n8598 ;
  assign n16530 = n5919 & ~n16529 ;
  assign n16531 = n4876 | n16530 ;
  assign n16535 = n310 & n14936 ;
  assign n16532 = n14890 ^ n9902 ^ 1'b0 ;
  assign n16533 = n2946 & n6585 ;
  assign n16534 = n16532 | n16533 ;
  assign n16536 = n16535 ^ n16534 ^ 1'b0 ;
  assign n16537 = n6008 | n16536 ;
  assign n16538 = ~n3022 & n10305 ;
  assign n16539 = n16538 ^ n15862 ^ 1'b0 ;
  assign n16540 = n8456 | n11412 ;
  assign n16541 = ~n1067 & n1899 ;
  assign n16542 = n1067 & n16541 ;
  assign n16544 = n5478 & ~n6655 ;
  assign n16545 = n16544 ^ n2070 ^ 1'b0 ;
  assign n16543 = n1496 & n6661 ;
  assign n16546 = n16545 ^ n16543 ^ 1'b0 ;
  assign n16547 = ~n6893 & n16546 ;
  assign n16548 = ~n6259 & n16547 ;
  assign n16549 = ~n14389 & n16548 ;
  assign n16562 = ( ~x188 & n1240 ) | ( ~x188 & n2172 ) | ( n1240 & n2172 ) ;
  assign n16550 = ~n276 & n3166 ;
  assign n16551 = ~n3166 & n16550 ;
  assign n16552 = n1255 | n16551 ;
  assign n16553 = n16551 & ~n16552 ;
  assign n16554 = n7537 | n16553 ;
  assign n16555 = n7537 & ~n16554 ;
  assign n16556 = n1891 | n16555 ;
  assign n16557 = n1891 & ~n16556 ;
  assign n16558 = n12556 ^ n6567 ^ 1'b0 ;
  assign n16559 = n7779 & n16558 ;
  assign n16560 = n16559 ^ n5594 ^ 1'b0 ;
  assign n16561 = n16557 | n16560 ;
  assign n16563 = n16562 ^ n16561 ^ 1'b0 ;
  assign n16564 = n1570 | n16563 ;
  assign n16565 = n7177 ^ n6737 ^ 1'b0 ;
  assign n16566 = n16565 ^ n1981 ^ x121 ;
  assign n16567 = n3115 & ~n16566 ;
  assign n16568 = ~n7124 & n11866 ;
  assign n16569 = ~n3639 & n12857 ;
  assign n16570 = ~x143 & n7624 ;
  assign n16571 = ~n16569 & n16570 ;
  assign n16572 = ~x137 & n12676 ;
  assign n16573 = n16571 & n16572 ;
  assign n16575 = n10089 ^ n4229 ^ 1'b0 ;
  assign n16574 = n1782 | n7745 ;
  assign n16576 = n16575 ^ n16574 ^ 1'b0 ;
  assign n16577 = n5205 | n16576 ;
  assign n16578 = n13557 & ~n16577 ;
  assign n16579 = n3753 & n11106 ;
  assign n16580 = n16579 ^ n4218 ^ 1'b0 ;
  assign n16581 = n3380 & ~n16580 ;
  assign n16582 = n16581 ^ n813 ^ 1'b0 ;
  assign n16583 = n16582 ^ n7390 ^ 1'b0 ;
  assign n16584 = ~n8380 & n16583 ;
  assign n16585 = n3850 & ~n15010 ;
  assign n16586 = ~n5213 & n16585 ;
  assign n16587 = n1221 & n15108 ;
  assign n16588 = ~n12380 & n16587 ;
  assign n16589 = n5664 & ~n14873 ;
  assign n16590 = n6374 & ~n16589 ;
  assign n16591 = ~n1958 & n4807 ;
  assign n16592 = ( n6983 & ~n9457 ) | ( n6983 & n16591 ) | ( ~n9457 & n16591 ) ;
  assign n16593 = n4598 | n15069 ;
  assign n16594 = n4501 ^ n1777 ^ 1'b0 ;
  assign n16595 = ~n6881 & n16594 ;
  assign n16596 = n14540 ^ n4296 ^ 1'b0 ;
  assign n16597 = n12297 & ~n16596 ;
  assign n16598 = n1779 & ~n13309 ;
  assign n16599 = ~n1101 & n16598 ;
  assign n16600 = n3195 | n16599 ;
  assign n16602 = ~n1952 & n8488 ;
  assign n16603 = ~n2073 & n16602 ;
  assign n16601 = n3235 & n8447 ;
  assign n16604 = n16603 ^ n16601 ^ 1'b0 ;
  assign n16605 = ~n2441 & n3936 ;
  assign n16606 = ~n7876 & n16605 ;
  assign n16607 = n14143 ^ n871 ^ 1'b0 ;
  assign n16608 = ~n16606 & n16607 ;
  assign n16609 = n3348 ^ n276 ^ 1'b0 ;
  assign n16610 = n5490 & n7554 ;
  assign n16611 = n2661 & n4214 ;
  assign n16612 = n12987 & ~n16611 ;
  assign n16613 = n5978 | n16612 ;
  assign n16614 = n7395 ^ n1588 ^ 1'b0 ;
  assign n16615 = ( n5511 & ~n9140 ) | ( n5511 & n10408 ) | ( ~n9140 & n10408 ) ;
  assign n16616 = n1389 ^ n1295 ^ 1'b0 ;
  assign n16617 = ~n14840 & n16616 ;
  assign n16618 = ( n8334 & ~n9339 ) | ( n8334 & n16617 ) | ( ~n9339 & n16617 ) ;
  assign n16619 = n14803 ^ n723 ^ 1'b0 ;
  assign n16620 = n4306 & n16619 ;
  assign n16621 = n16620 ^ n3933 ^ n3750 ;
  assign n16622 = n7118 & ~n9332 ;
  assign n16623 = n2476 | n8638 ;
  assign n16624 = ( n387 & n779 ) | ( n387 & n2571 ) | ( n779 & n2571 ) ;
  assign n16625 = n8592 & n16624 ;
  assign n16626 = ~n2169 & n16625 ;
  assign n16627 = ~n12773 & n16626 ;
  assign n16628 = n11456 ^ n9340 ^ n7766 ;
  assign n16629 = x192 | n16628 ;
  assign n16630 = n16629 ^ n6144 ^ 1'b0 ;
  assign n16631 = n1710 & ~n15425 ;
  assign n16632 = n11410 & n16631 ;
  assign n16633 = ( ~x180 & n1045 ) | ( ~x180 & n10609 ) | ( n1045 & n10609 ) ;
  assign n16634 = n16633 ^ n496 ^ 1'b0 ;
  assign n16635 = x107 | n4956 ;
  assign n16636 = n16635 ^ n1802 ^ 1'b0 ;
  assign n16637 = n16636 ^ n3922 ^ 1'b0 ;
  assign n16638 = n3019 ^ n2265 ^ 1'b0 ;
  assign n16639 = ~n1301 & n2087 ;
  assign n16640 = n16639 ^ n2420 ^ 1'b0 ;
  assign n16641 = n6996 | n16640 ;
  assign n16642 = n1748 | n16641 ;
  assign n16643 = n6331 & n15553 ;
  assign n16644 = n16643 ^ n3745 ^ 1'b0 ;
  assign n16645 = n16644 ^ n13448 ^ 1'b0 ;
  assign n16646 = ( n4001 & ~n7485 ) | ( n4001 & n8073 ) | ( ~n7485 & n8073 ) ;
  assign n16647 = n16646 ^ n14040 ^ 1'b0 ;
  assign n16648 = n3954 & n10768 ;
  assign n16649 = n16648 ^ n5063 ^ 1'b0 ;
  assign n16650 = n11586 ^ n8141 ^ 1'b0 ;
  assign n16651 = ~n2023 & n16650 ;
  assign n16652 = n16649 & n16651 ;
  assign n16653 = n16647 & n16652 ;
  assign n16654 = ~n2169 & n8933 ;
  assign n16655 = n14017 & n16654 ;
  assign n16659 = n6660 ^ n5864 ^ 1'b0 ;
  assign n16660 = n4817 & n16659 ;
  assign n16656 = n12133 ^ n5276 ^ 1'b0 ;
  assign n16657 = n5427 | n16656 ;
  assign n16658 = n6358 & ~n16657 ;
  assign n16661 = n16660 ^ n16658 ^ 1'b0 ;
  assign n16662 = n13895 ^ n3050 ^ 1'b0 ;
  assign n16663 = n7301 ^ n3568 ^ 1'b0 ;
  assign n16664 = ~n2828 & n16663 ;
  assign n16665 = n2918 ^ n2086 ^ 1'b0 ;
  assign n16666 = n3331 & n16665 ;
  assign n16667 = n16666 ^ n13654 ^ 1'b0 ;
  assign n16668 = ~n5195 & n16667 ;
  assign n16669 = x206 & ~n16668 ;
  assign n16670 = n10022 & n11999 ;
  assign n16671 = n389 & ~n16508 ;
  assign n16672 = n16671 ^ n14191 ^ 1'b0 ;
  assign n16673 = n5563 ^ n4918 ^ 1'b0 ;
  assign n16674 = n12009 ^ n5213 ^ 1'b0 ;
  assign n16675 = n7195 & ~n16674 ;
  assign n16676 = n4887 | n11745 ;
  assign n16677 = n16676 ^ n5484 ^ 1'b0 ;
  assign n16678 = n16675 & n16677 ;
  assign n16679 = n9496 & n13757 ;
  assign n16680 = ~n2815 & n16679 ;
  assign n16681 = n16680 ^ n1294 ^ 1'b0 ;
  assign n16682 = n14381 ^ x110 ^ 1'b0 ;
  assign n16683 = n16682 ^ n16231 ^ n11745 ;
  assign n16684 = n15442 ^ n7693 ^ 1'b0 ;
  assign n16685 = n3231 | n16684 ;
  assign n16686 = n2004 ^ x36 ^ 1'b0 ;
  assign n16687 = n16686 ^ n3412 ^ 1'b0 ;
  assign n16688 = n16687 ^ n16308 ^ 1'b0 ;
  assign n16689 = n5920 ^ n2715 ^ 1'b0 ;
  assign n16690 = ~n2783 & n16689 ;
  assign n16691 = n10467 | n16690 ;
  assign n16692 = n11144 | n15370 ;
  assign n16693 = n14246 | n16692 ;
  assign n16694 = ~n1078 & n3431 ;
  assign n16695 = n16694 ^ n7732 ^ 1'b0 ;
  assign n16696 = n3814 ^ x60 ^ 1'b0 ;
  assign n16697 = n8966 | n16696 ;
  assign n16698 = n14912 & ~n16697 ;
  assign n16699 = n16698 ^ n6781 ^ 1'b0 ;
  assign n16700 = n3731 | n10990 ;
  assign n16701 = n7506 ^ n4589 ^ 1'b0 ;
  assign n16702 = ~n13689 & n16701 ;
  assign n16703 = n16702 ^ n2443 ^ 1'b0 ;
  assign n16704 = n6972 & ~n16703 ;
  assign n16705 = n16704 ^ n4226 ^ 1'b0 ;
  assign n16706 = x221 & n4321 ;
  assign n16707 = ~x111 & n16706 ;
  assign n16708 = n14455 ^ n367 ^ 1'b0 ;
  assign n16709 = n4395 | n4679 ;
  assign n16710 = n10778 ^ n3121 ^ 1'b0 ;
  assign n16711 = ~n6169 & n16710 ;
  assign n16712 = n16709 & n16711 ;
  assign n16713 = n5459 ^ n4193 ^ 1'b0 ;
  assign n16714 = n4831 & ~n16713 ;
  assign n16715 = n10541 & n16714 ;
  assign n16716 = n16712 & n16715 ;
  assign n16717 = n9525 ^ n2248 ^ 1'b0 ;
  assign n16718 = n12216 | n16717 ;
  assign n16719 = n16177 ^ n7321 ^ 1'b0 ;
  assign n16722 = ( ~n2045 & n10706 ) | ( ~n2045 & n12913 ) | ( n10706 & n12913 ) ;
  assign n16720 = n5046 & ~n6682 ;
  assign n16721 = ~n8463 & n16720 ;
  assign n16723 = n16722 ^ n16721 ^ 1'b0 ;
  assign n16724 = n7858 ^ n4169 ^ 1'b0 ;
  assign n16725 = n359 | n10954 ;
  assign n16726 = n558 & ~n12889 ;
  assign n16727 = n16725 & n16726 ;
  assign n16728 = n3210 ^ n766 ^ 1'b0 ;
  assign n16734 = x195 & n3875 ;
  assign n16735 = n16734 ^ n3710 ^ 1'b0 ;
  assign n16729 = n1211 | n5374 ;
  assign n16730 = n3081 & ~n16729 ;
  assign n16731 = n16730 ^ n10170 ^ n6033 ;
  assign n16732 = n12581 & n16731 ;
  assign n16733 = x99 | n16732 ;
  assign n16736 = n16735 ^ n16733 ^ 1'b0 ;
  assign n16737 = ~n16728 & n16736 ;
  assign n16738 = n5284 ^ n3565 ^ 1'b0 ;
  assign n16739 = n16737 & ~n16738 ;
  assign n16740 = n5177 | n14236 ;
  assign n16741 = n9260 ^ n296 ^ 1'b0 ;
  assign n16742 = n7513 & ~n16741 ;
  assign n16743 = n16742 ^ n2224 ^ 1'b0 ;
  assign n16744 = n2666 | n2703 ;
  assign n16745 = n3723 & ~n16744 ;
  assign n16746 = ~n3670 & n16745 ;
  assign n16747 = n16746 ^ n4608 ^ 1'b0 ;
  assign n16748 = n15271 & ~n15342 ;
  assign n16749 = n10325 & n16748 ;
  assign n16750 = n2255 & n4333 ;
  assign n16751 = n16750 ^ n13692 ^ 1'b0 ;
  assign n16752 = n2183 & n3950 ;
  assign n16753 = n6518 & n16752 ;
  assign n16754 = n15299 & ~n16753 ;
  assign n16755 = ~n3716 & n16754 ;
  assign n16756 = ~n7662 & n16755 ;
  assign n16757 = n3216 ^ x40 ^ 1'b0 ;
  assign n16758 = n16757 ^ n9713 ^ 1'b0 ;
  assign n16759 = ( n13693 & n16756 ) | ( n13693 & ~n16758 ) | ( n16756 & ~n16758 ) ;
  assign n16760 = ~n2715 & n3758 ;
  assign n16761 = n2018 | n2936 ;
  assign n16762 = n16761 ^ n6791 ^ 1'b0 ;
  assign n16763 = n15937 & ~n16762 ;
  assign n16764 = ( ~n291 & n1925 ) | ( ~n291 & n4946 ) | ( n1925 & n4946 ) ;
  assign n16765 = n16763 & ~n16764 ;
  assign n16766 = ~n1802 & n16765 ;
  assign n16767 = n16766 ^ n6952 ^ 1'b0 ;
  assign n16768 = ~n9788 & n16005 ;
  assign n16769 = n4405 | n15821 ;
  assign n16770 = n16768 & ~n16769 ;
  assign n16771 = n5088 ^ n2345 ^ 1'b0 ;
  assign n16772 = n16771 ^ n6393 ^ 1'b0 ;
  assign n16773 = n3134 | n16772 ;
  assign n16774 = ~n3985 & n5259 ;
  assign n16775 = n16773 & n16774 ;
  assign n16776 = n14087 ^ n11683 ^ x116 ;
  assign n16777 = ( n5676 & n16775 ) | ( n5676 & n16776 ) | ( n16775 & n16776 ) ;
  assign n16778 = n15018 ^ n5846 ^ 1'b0 ;
  assign n16779 = n16778 ^ n4793 ^ 1'b0 ;
  assign n16780 = n5984 & n14596 ;
  assign n16781 = ~n8235 & n8353 ;
  assign n16782 = n4460 ^ n2400 ^ 1'b0 ;
  assign n16783 = n16781 | n16782 ;
  assign n16784 = n6246 | n14971 ;
  assign n16785 = n5917 & ~n11080 ;
  assign n16786 = n16785 ^ n643 ^ 1'b0 ;
  assign n16787 = n7013 ^ n1608 ^ 1'b0 ;
  assign n16788 = n16786 & n16787 ;
  assign n16789 = n5509 & n16788 ;
  assign n16790 = ~n5978 & n16789 ;
  assign n16791 = n5309 & ~n10915 ;
  assign n16792 = n13022 | n14829 ;
  assign n16793 = ~n619 & n3840 ;
  assign n16794 = n780 & n16793 ;
  assign n16795 = n2743 | n16794 ;
  assign n16796 = n2640 & ~n4023 ;
  assign n16797 = n16796 ^ n1048 ^ 1'b0 ;
  assign n16798 = n2305 & n12233 ;
  assign n16799 = n16798 ^ x70 ^ 1'b0 ;
  assign n16800 = n14308 & n16799 ;
  assign n16801 = ~n349 & n2684 ;
  assign n16802 = ~n1086 & n16801 ;
  assign n16803 = n16802 ^ n9663 ^ 1'b0 ;
  assign n16804 = n4460 ^ n1347 ^ 1'b0 ;
  assign n16805 = n16804 ^ n4596 ^ 1'b0 ;
  assign n16806 = x79 & n7683 ;
  assign n16807 = n16806 ^ n6557 ^ 1'b0 ;
  assign n16808 = n16807 ^ n2726 ^ 1'b0 ;
  assign n16809 = ( n4428 & n16805 ) | ( n4428 & ~n16808 ) | ( n16805 & ~n16808 ) ;
  assign n16810 = x82 & ~n4911 ;
  assign n16811 = n8654 ^ n378 ^ 1'b0 ;
  assign n16812 = ~n13088 & n16811 ;
  assign n16813 = n2577 & n15233 ;
  assign n16814 = n9075 ^ n6817 ^ 1'b0 ;
  assign n16815 = n7868 & ~n16814 ;
  assign n16816 = ~n6141 & n16815 ;
  assign n16817 = n16816 ^ n2999 ^ 1'b0 ;
  assign n16818 = ~n3639 & n14044 ;
  assign n16819 = n4938 & ~n16818 ;
  assign n16820 = n13650 ^ n7384 ^ n3680 ;
  assign n16821 = n4984 & ~n12457 ;
  assign n16822 = ~x122 & n16821 ;
  assign n16823 = n6111 | n16822 ;
  assign n16824 = n16823 ^ n10102 ^ 1'b0 ;
  assign n16825 = n1995 ^ n787 ^ 1'b0 ;
  assign n16826 = n15904 & ~n16825 ;
  assign n16828 = n302 & n2317 ;
  assign n16829 = n16828 ^ n1001 ^ 1'b0 ;
  assign n16827 = ~n2521 & n16453 ;
  assign n16830 = n16829 ^ n16827 ^ 1'b0 ;
  assign n16831 = n12655 & ~n14089 ;
  assign n16832 = n16831 ^ n15416 ^ 1'b0 ;
  assign n16833 = ~n3060 & n7736 ;
  assign n16834 = ~n2942 & n16833 ;
  assign n16835 = n8241 ^ n4493 ^ 1'b0 ;
  assign n16836 = ~n16834 & n16835 ;
  assign n16837 = ~n12040 & n12168 ;
  assign n16838 = ~n7696 & n16668 ;
  assign n16839 = n2428 ^ x92 ^ 1'b0 ;
  assign n16840 = ~n7743 & n16839 ;
  assign n16841 = n16840 ^ n14768 ^ 1'b0 ;
  assign n16842 = n11451 | n16841 ;
  assign n16843 = n6038 ^ n2787 ^ 1'b0 ;
  assign n16844 = n1196 | n16843 ;
  assign n16845 = n7524 & n16844 ;
  assign n16846 = n7662 | n9088 ;
  assign n16847 = n16845 | n16846 ;
  assign n16848 = n16847 ^ n14703 ^ 1'b0 ;
  assign n16851 = x248 & n611 ;
  assign n16852 = n16851 ^ n5238 ^ 1'b0 ;
  assign n16849 = ~n2966 & n14263 ;
  assign n16850 = ~n2458 & n16849 ;
  assign n16853 = n16852 ^ n16850 ^ 1'b0 ;
  assign n16854 = n16853 ^ n10604 ^ 1'b0 ;
  assign n16855 = ~n16463 & n16854 ;
  assign n16856 = n4919 & n9260 ;
  assign n16857 = n16856 ^ n462 ^ 1'b0 ;
  assign n16858 = ( n7596 & n14421 ) | ( n7596 & ~n16857 ) | ( n14421 & ~n16857 ) ;
  assign n16862 = ~n825 & n14420 ;
  assign n16863 = n16862 ^ n3514 ^ 1'b0 ;
  assign n16859 = ~x132 & x146 ;
  assign n16860 = ~n988 & n16859 ;
  assign n16861 = n3913 & n16860 ;
  assign n16864 = n16863 ^ n16861 ^ 1'b0 ;
  assign n16865 = n8594 & n13814 ;
  assign n16866 = n9798 & n14106 ;
  assign n16867 = n2348 | n6623 ;
  assign n16868 = n16867 ^ n3721 ^ 1'b0 ;
  assign n16869 = n14803 ^ n3223 ^ n572 ;
  assign n16870 = n4227 & n16869 ;
  assign n16871 = n10219 ^ n3760 ^ n3183 ;
  assign n16872 = n13365 & ~n16871 ;
  assign n16873 = n16872 ^ n6537 ^ 1'b0 ;
  assign n16874 = n16851 ^ n4360 ^ 1'b0 ;
  assign n16875 = ~n8633 & n9717 ;
  assign n16876 = n4793 | n15468 ;
  assign n16877 = n16876 ^ n2366 ^ 1'b0 ;
  assign n16878 = ~n13405 & n16877 ;
  assign n16879 = n4123 ^ n2685 ^ 1'b0 ;
  assign n16880 = n16879 ^ n12714 ^ 1'b0 ;
  assign n16881 = n6580 & ~n11920 ;
  assign n16882 = n7904 & n16881 ;
  assign n16883 = n16882 ^ n3855 ^ 1'b0 ;
  assign n16884 = n16880 & ~n16883 ;
  assign n16885 = ( n1217 & n1494 ) | ( n1217 & ~n1615 ) | ( n1494 & ~n1615 ) ;
  assign n16886 = n585 & n16885 ;
  assign n16887 = ( n391 & n4525 ) | ( n391 & n14072 ) | ( n4525 & n14072 ) ;
  assign n16888 = n12380 & n15381 ;
  assign n16889 = n1621 & ~n4014 ;
  assign n16890 = n9153 | n16889 ;
  assign n16891 = n1231 | n16890 ;
  assign n16892 = ~n8849 & n16891 ;
  assign n16893 = n16892 ^ n13643 ^ n11838 ;
  assign n16894 = n1018 & n10499 ;
  assign n16895 = n16894 ^ n2967 ^ 1'b0 ;
  assign n16896 = x116 & n9782 ;
  assign n16897 = ~n2165 & n16896 ;
  assign n16899 = ~n3705 & n7418 ;
  assign n16898 = ( n1458 & n8269 ) | ( n1458 & ~n14865 ) | ( n8269 & ~n14865 ) ;
  assign n16900 = n16899 ^ n16898 ^ 1'b0 ;
  assign n16901 = n1544 & ~n8957 ;
  assign n16902 = n6259 ^ n3446 ^ 1'b0 ;
  assign n16903 = n16902 ^ n3544 ^ 1'b0 ;
  assign n16904 = n16903 ^ n9973 ^ 1'b0 ;
  assign n16905 = n16901 & ~n16904 ;
  assign n16906 = n12664 & n13887 ;
  assign n16907 = n16906 ^ n5374 ^ n3674 ;
  assign n16908 = n10455 ^ n4736 ^ 1'b0 ;
  assign n16909 = n4130 | n16908 ;
  assign n16910 = n11423 & n16484 ;
  assign n16911 = n16909 & n16910 ;
  assign n16912 = n2518 | n12638 ;
  assign n16913 = n1259 & n4380 ;
  assign n16914 = n4527 & ~n9407 ;
  assign n16915 = ~n12438 & n16914 ;
  assign n16916 = x86 & ~n16915 ;
  assign n16917 = n12293 ^ n9870 ^ 1'b0 ;
  assign n16918 = ~n8289 & n16917 ;
  assign n16919 = n16916 & n16918 ;
  assign n16920 = n14207 ^ n5459 ^ n3594 ;
  assign n16921 = n14000 & ~n16920 ;
  assign n16926 = n1588 | n2772 ;
  assign n16922 = n8654 ^ n666 ^ 1'b0 ;
  assign n16923 = ~n12953 & n16922 ;
  assign n16924 = n10280 & n16923 ;
  assign n16925 = ~n15547 & n16924 ;
  assign n16927 = n16926 ^ n16925 ^ n13185 ;
  assign n16928 = n899 | n6773 ;
  assign n16929 = n16928 ^ n5859 ^ 1'b0 ;
  assign n16930 = n8009 & ~n13300 ;
  assign n16931 = n3604 & ~n3880 ;
  assign n16932 = n16931 ^ x17 ^ 1'b0 ;
  assign n16933 = x105 & ~n9383 ;
  assign n16934 = n16933 ^ n2533 ^ 1'b0 ;
  assign n16935 = ( n8803 & n16932 ) | ( n8803 & ~n16934 ) | ( n16932 & ~n16934 ) ;
  assign n16936 = n2006 & ~n5934 ;
  assign n16937 = n11093 ^ n10106 ^ 1'b0 ;
  assign n16938 = ( n5746 & ~n8432 ) | ( n5746 & n13000 ) | ( ~n8432 & n13000 ) ;
  assign n16939 = ( n473 & n3385 ) | ( n473 & ~n7448 ) | ( n3385 & ~n7448 ) ;
  assign n16940 = ~n10172 & n15050 ;
  assign n16945 = n7409 ^ n1142 ^ 1'b0 ;
  assign n16941 = n11528 ^ n10014 ^ 1'b0 ;
  assign n16942 = ~n11002 & n16941 ;
  assign n16943 = n16942 ^ n1112 ^ 1'b0 ;
  assign n16944 = n11939 | n16943 ;
  assign n16946 = n16945 ^ n16944 ^ 1'b0 ;
  assign n16947 = ~x44 & n16946 ;
  assign n16948 = n16262 ^ n8583 ^ 1'b0 ;
  assign n16949 = n13666 & n16948 ;
  assign n16950 = n13737 & ~n14948 ;
  assign n16951 = ~n6660 & n15148 ;
  assign n16952 = n16951 ^ n2065 ^ 1'b0 ;
  assign n16953 = n14965 ^ n314 ^ 1'b0 ;
  assign n16954 = n3233 ^ n2341 ^ 1'b0 ;
  assign n16955 = n1896 & n16954 ;
  assign n16956 = n4174 & n16955 ;
  assign n16957 = n3286 | n13711 ;
  assign n16958 = n16957 ^ n9721 ^ 1'b0 ;
  assign n16959 = ~n4603 & n12838 ;
  assign n16960 = ( n428 & n1098 ) | ( n428 & n16959 ) | ( n1098 & n16959 ) ;
  assign n16961 = ~n6322 & n13662 ;
  assign n16962 = n5639 & n14179 ;
  assign n16963 = n9758 ^ n1547 ^ 1'b0 ;
  assign n16964 = n3400 | n16963 ;
  assign n16965 = n10248 ^ n913 ^ 1'b0 ;
  assign n16966 = n2262 ^ n1157 ^ 1'b0 ;
  assign n16967 = n11805 ^ n8319 ^ 1'b0 ;
  assign n16968 = n16967 ^ n10043 ^ 1'b0 ;
  assign n16969 = n5579 ^ n2369 ^ 1'b0 ;
  assign n16970 = ( n3607 & ~n6129 ) | ( n3607 & n6514 ) | ( ~n6129 & n6514 ) ;
  assign n16971 = n9996 ^ n3018 ^ 1'b0 ;
  assign n16972 = n4983 & n16971 ;
  assign n16973 = n16972 ^ n14383 ^ 1'b0 ;
  assign n16974 = n4933 & ~n16973 ;
  assign n16975 = n3451 | n8105 ;
  assign n16976 = n3431 & n16975 ;
  assign n16977 = n11536 ^ n8957 ^ n6639 ;
  assign n16978 = ( x48 & n11585 ) | ( x48 & n16977 ) | ( n11585 & n16977 ) ;
  assign n16979 = n6203 ^ n5990 ^ 1'b0 ;
  assign n16980 = n6935 | n16979 ;
  assign n16981 = n16980 ^ n6058 ^ 1'b0 ;
  assign n16982 = n14423 | n16981 ;
  assign n16983 = n16982 ^ n2859 ^ 1'b0 ;
  assign n16984 = n7072 & ~n13202 ;
  assign n16985 = n2474 | n7201 ;
  assign n16986 = n5347 & ~n16985 ;
  assign n16987 = ( n7703 & n16984 ) | ( n7703 & ~n16986 ) | ( n16984 & ~n16986 ) ;
  assign n16988 = ( n1768 & n7579 ) | ( n1768 & ~n11450 ) | ( n7579 & ~n11450 ) ;
  assign n16989 = n13488 ^ n4728 ^ 1'b0 ;
  assign n16990 = n16989 ^ n2262 ^ n1681 ;
  assign n16991 = ~n8354 & n16990 ;
  assign n16992 = n2710 & n12876 ;
  assign n16993 = n844 & n4580 ;
  assign n16994 = ~n4580 & n16993 ;
  assign n16995 = x104 & n16994 ;
  assign n16996 = n16995 ^ n12132 ^ 1'b0 ;
  assign n16997 = ~n7274 & n16996 ;
  assign n16998 = n7274 & n16997 ;
  assign n16999 = n3670 & n13171 ;
  assign n17001 = ~n1599 & n10191 ;
  assign n17000 = n11263 | n12416 ;
  assign n17002 = n17001 ^ n17000 ^ 1'b0 ;
  assign n17003 = ~n1950 & n17002 ;
  assign n17004 = n3887 & ~n9412 ;
  assign n17005 = ~n17003 & n17004 ;
  assign n17006 = n16859 ^ n6655 ^ 1'b0 ;
  assign n17007 = n15549 | n17006 ;
  assign n17008 = ~n260 & n7679 ;
  assign n17009 = n8531 & n8625 ;
  assign n17010 = ( n17007 & n17008 ) | ( n17007 & n17009 ) | ( n17008 & n17009 ) ;
  assign n17011 = n1439 | n6447 ;
  assign n17012 = n744 & ~n17011 ;
  assign n17013 = ~n4247 & n10827 ;
  assign n17014 = ~n17012 & n17013 ;
  assign n17015 = n17014 ^ n2446 ^ 1'b0 ;
  assign n17016 = n13790 | n17015 ;
  assign n17017 = n17016 ^ n1513 ^ 1'b0 ;
  assign n17018 = n11388 ^ n11351 ^ 1'b0 ;
  assign n17019 = n12828 ^ n6627 ^ 1'b0 ;
  assign n17021 = n7538 ^ n3966 ^ 1'b0 ;
  assign n17020 = n1109 | n11734 ;
  assign n17022 = n17021 ^ n17020 ^ 1'b0 ;
  assign n17023 = ~n5136 & n17022 ;
  assign n17024 = n8228 & n13510 ;
  assign n17025 = n17024 ^ n11318 ^ 1'b0 ;
  assign n17026 = n927 | n2531 ;
  assign n17027 = n703 | n17026 ;
  assign n17028 = ( n1813 & n3683 ) | ( n1813 & n8449 ) | ( n3683 & n8449 ) ;
  assign n17029 = ~n1342 & n17028 ;
  assign n17030 = n17027 & n17029 ;
  assign n17031 = n17030 ^ n13608 ^ 1'b0 ;
  assign n17038 = n12536 ^ n854 ^ 1'b0 ;
  assign n17032 = n3513 ^ n268 ^ 1'b0 ;
  assign n17033 = ( ~n4684 & n8353 ) | ( ~n4684 & n17032 ) | ( n8353 & n17032 ) ;
  assign n17034 = n8381 | n17033 ;
  assign n17035 = n17034 ^ n14444 ^ 1'b0 ;
  assign n17036 = n1025 & ~n16612 ;
  assign n17037 = n17035 & n17036 ;
  assign n17039 = n17038 ^ n17037 ^ n2399 ;
  assign n17040 = n12585 ^ n851 ^ 1'b0 ;
  assign n17041 = n5802 ^ n2299 ^ 1'b0 ;
  assign n17042 = n16735 | n17041 ;
  assign n17043 = n17040 & ~n17042 ;
  assign n17044 = n7515 & n16955 ;
  assign n17045 = ~n5170 & n17044 ;
  assign n17046 = n3296 & n6572 ;
  assign n17047 = n17045 & n17046 ;
  assign n17048 = ~n8517 & n16675 ;
  assign n17049 = n17048 ^ n2096 ^ 1'b0 ;
  assign n17050 = x152 & n9652 ;
  assign n17051 = n1332 & n17050 ;
  assign n17052 = n327 & ~n17051 ;
  assign n17053 = ( ~n4226 & n5169 ) | ( ~n4226 & n9578 ) | ( n5169 & n9578 ) ;
  assign n17054 = ~n17052 & n17053 ;
  assign n17055 = n17054 ^ n10408 ^ 1'b0 ;
  assign n17056 = n5243 & n10100 ;
  assign n17057 = n10742 & ~n17056 ;
  assign n17058 = ~n12299 & n17057 ;
  assign n17060 = n3172 & n4213 ;
  assign n17061 = n716 & n17060 ;
  assign n17062 = n1822 & ~n17061 ;
  assign n17063 = n17062 ^ n2133 ^ 1'b0 ;
  assign n17064 = n4462 | n17063 ;
  assign n17065 = n5403 | n17064 ;
  assign n17066 = n1333 & n13552 ;
  assign n17067 = ~n10431 & n17066 ;
  assign n17068 = n17065 & ~n17067 ;
  assign n17069 = ~n6666 & n17068 ;
  assign n17059 = n7231 | n7738 ;
  assign n17070 = n17069 ^ n17059 ^ 1'b0 ;
  assign n17073 = ~n10625 & n13546 ;
  assign n17071 = ( x207 & n1636 ) | ( x207 & ~n6908 ) | ( n1636 & ~n6908 ) ;
  assign n17072 = n5704 & n17071 ;
  assign n17074 = n17073 ^ n17072 ^ 1'b0 ;
  assign n17075 = n5065 ^ n4449 ^ n825 ;
  assign n17076 = ~n12146 & n17075 ;
  assign n17077 = n17076 ^ n7028 ^ 1'b0 ;
  assign n17078 = n754 ^ n529 ^ 1'b0 ;
  assign n17079 = n17078 ^ n6554 ^ 1'b0 ;
  assign n17080 = n13054 ^ n3567 ^ n779 ;
  assign n17081 = n15192 ^ n5027 ^ n2651 ;
  assign n17082 = n17081 ^ n4934 ^ 1'b0 ;
  assign n17083 = ~n11000 & n11821 ;
  assign n17084 = n16653 & n17083 ;
  assign n17085 = n2014 & ~n5646 ;
  assign n17086 = n17085 ^ n14873 ^ 1'b0 ;
  assign n17087 = n6404 | n12524 ;
  assign n17090 = ~n2845 & n11990 ;
  assign n17091 = n17090 ^ n372 ^ 1'b0 ;
  assign n17092 = n9335 & n17091 ;
  assign n17088 = n4405 | n15459 ;
  assign n17089 = n4869 & ~n17088 ;
  assign n17093 = n17092 ^ n17089 ^ 1'b0 ;
  assign n17094 = n2015 | n10516 ;
  assign n17095 = n17094 ^ n4505 ^ 1'b0 ;
  assign n17097 = n865 & n4195 ;
  assign n17096 = ~n1426 & n7388 ;
  assign n17098 = n17097 ^ n17096 ^ 1'b0 ;
  assign n17099 = n7637 ^ n1114 ^ 1'b0 ;
  assign n17100 = n14402 & ~n17099 ;
  assign n17101 = n8050 & n17100 ;
  assign n17102 = n17101 ^ n789 ^ 1'b0 ;
  assign n17103 = n8272 & ~n13666 ;
  assign n17105 = ~n7274 & n8638 ;
  assign n17106 = ~n10376 & n17105 ;
  assign n17107 = n6865 & n7431 ;
  assign n17108 = ~n17106 & n17107 ;
  assign n17109 = n3171 & n17108 ;
  assign n17104 = n3114 & ~n3298 ;
  assign n17110 = n17109 ^ n17104 ^ 1'b0 ;
  assign n17111 = n15178 & n17110 ;
  assign n17112 = n16313 & n17111 ;
  assign n17113 = n6305 & ~n9153 ;
  assign n17114 = n2324 | n17113 ;
  assign n17115 = n17114 ^ n6024 ^ 1'b0 ;
  assign n17116 = n6770 & ~n17115 ;
  assign n17117 = n7848 & n10778 ;
  assign n17118 = ~n2479 & n17117 ;
  assign n17119 = ~n5352 & n12451 ;
  assign n17120 = ~n12187 & n17119 ;
  assign n17121 = ~n2986 & n3685 ;
  assign n17122 = n724 | n9301 ;
  assign n17123 = n5135 | n7990 ;
  assign n17124 = n17123 ^ n15166 ^ 1'b0 ;
  assign n17125 = n5066 ^ n509 ^ 1'b0 ;
  assign n17126 = x160 & ~n17125 ;
  assign n17127 = n17126 ^ n961 ^ 1'b0 ;
  assign n17128 = n17127 ^ n11514 ^ 1'b0 ;
  assign n17129 = ~n9456 & n17128 ;
  assign n17136 = n9652 | n11699 ;
  assign n17131 = n6474 ^ n5688 ^ 1'b0 ;
  assign n17130 = n4506 & n12340 ;
  assign n17132 = n17131 ^ n17130 ^ 1'b0 ;
  assign n17133 = n17132 ^ n3704 ^ 1'b0 ;
  assign n17134 = n3974 & n17133 ;
  assign n17135 = ~x107 & n17134 ;
  assign n17137 = n17136 ^ n17135 ^ 1'b0 ;
  assign n17138 = n3804 | n7523 ;
  assign n17139 = n17138 ^ n7432 ^ 1'b0 ;
  assign n17140 = n17139 ^ n325 ^ 1'b0 ;
  assign n17141 = ( n1069 & n1505 ) | ( n1069 & n14522 ) | ( n1505 & n14522 ) ;
  assign n17142 = n17141 ^ n7868 ^ 1'b0 ;
  assign n17143 = n16878 & ~n17142 ;
  assign n17144 = n5445 | n5948 ;
  assign n17145 = n17144 ^ n3564 ^ 1'b0 ;
  assign n17146 = n17145 ^ n5996 ^ 1'b0 ;
  assign n17147 = n11433 ^ n6612 ^ 1'b0 ;
  assign n17148 = n17147 ^ n7026 ^ n3780 ;
  assign n17149 = n6668 & n15775 ;
  assign n17150 = ( n6503 & ~n8523 ) | ( n6503 & n17149 ) | ( ~n8523 & n17149 ) ;
  assign n17151 = n12604 ^ n10929 ^ 1'b0 ;
  assign n17152 = ~n17150 & n17151 ;
  assign n17153 = n810 & n7576 ;
  assign n17161 = ( n3745 & n4286 ) | ( n3745 & n16807 ) | ( n4286 & n16807 ) ;
  assign n17154 = ( n363 & n6521 ) | ( n363 & ~n6681 ) | ( n6521 & ~n6681 ) ;
  assign n17155 = n10287 & ~n17154 ;
  assign n17156 = n6827 ^ n4911 ^ 1'b0 ;
  assign n17157 = ~n17155 & n17156 ;
  assign n17158 = ~n8530 & n17157 ;
  assign n17159 = n17158 ^ n4807 ^ 1'b0 ;
  assign n17160 = n7959 & ~n17159 ;
  assign n17162 = n17161 ^ n17160 ^ n2980 ;
  assign n17163 = n7972 ^ n1456 ^ x236 ;
  assign n17164 = ~n6591 & n17163 ;
  assign n17165 = n12900 ^ n1686 ^ 1'b0 ;
  assign n17166 = n1861 ^ n1196 ^ 1'b0 ;
  assign n17167 = n3962 & n17166 ;
  assign n17168 = n15202 ^ n11166 ^ 1'b0 ;
  assign n17169 = n10017 ^ n3568 ^ 1'b0 ;
  assign n17170 = n6115 | n17169 ;
  assign n17171 = n2041 & ~n8279 ;
  assign n17172 = n1459 ^ x59 ^ 1'b0 ;
  assign n17173 = n9311 ^ n6388 ^ 1'b0 ;
  assign n17174 = n756 & n17173 ;
  assign n17175 = ~n17172 & n17174 ;
  assign n17176 = ( n6678 & ~n7116 ) | ( n6678 & n12700 ) | ( ~n7116 & n12700 ) ;
  assign n17177 = n16214 ^ n15929 ^ 1'b0 ;
  assign n17178 = n3856 & n17177 ;
  assign n17179 = ( n3030 & n17176 ) | ( n3030 & n17178 ) | ( n17176 & n17178 ) ;
  assign n17180 = n5703 & ~n17179 ;
  assign n17181 = n3539 & n17180 ;
  assign n17182 = n1126 & n12664 ;
  assign n17183 = ~n7805 & n17182 ;
  assign n17184 = ( ~n7240 & n7724 ) | ( ~n7240 & n17183 ) | ( n7724 & n17183 ) ;
  assign n17185 = n1458 | n8087 ;
  assign n17186 = n17185 ^ n4770 ^ 1'b0 ;
  assign n17187 = n4010 & n17186 ;
  assign n17188 = ( n11170 & n11699 ) | ( n11170 & n17187 ) | ( n11699 & n17187 ) ;
  assign n17189 = n1499 | n17188 ;
  assign n17190 = n17189 ^ n13456 ^ 1'b0 ;
  assign n17191 = n3973 ^ n2857 ^ 1'b0 ;
  assign n17192 = n890 & ~n17191 ;
  assign n17193 = ( n274 & n7379 ) | ( n274 & ~n17192 ) | ( n7379 & ~n17192 ) ;
  assign n17194 = x220 & n11726 ;
  assign n17195 = n17194 ^ n7179 ^ 1'b0 ;
  assign n17196 = n9903 ^ n7040 ^ 1'b0 ;
  assign n17198 = n1759 ^ n1388 ^ 1'b0 ;
  assign n17197 = n1369 & ~n2034 ;
  assign n17199 = n17198 ^ n17197 ^ 1'b0 ;
  assign n17200 = ~n3137 & n17199 ;
  assign n17201 = ( n10079 & n11152 ) | ( n10079 & ~n17200 ) | ( n11152 & ~n17200 ) ;
  assign n17202 = n11369 ^ n2034 ^ 1'b0 ;
  assign n17209 = n1103 & n1768 ;
  assign n17210 = ~n1103 & n17209 ;
  assign n17211 = n944 | n17210 ;
  assign n17212 = n17210 & ~n17211 ;
  assign n17213 = ~n4426 & n4691 ;
  assign n17214 = n17212 & n17213 ;
  assign n17203 = n372 | n2976 ;
  assign n17204 = n372 & ~n17203 ;
  assign n17205 = n2183 & ~n17204 ;
  assign n17206 = ~n2183 & n17205 ;
  assign n17207 = n1441 & n17206 ;
  assign n17208 = n11701 & ~n17207 ;
  assign n17215 = n17214 ^ n17208 ^ 1'b0 ;
  assign n17216 = n17215 ^ n12000 ^ 1'b0 ;
  assign n17220 = n3425 ^ n2625 ^ n346 ;
  assign n17221 = ~n875 & n17220 ;
  assign n17217 = n8556 | n12902 ;
  assign n17218 = n17217 ^ n17187 ^ 1'b0 ;
  assign n17219 = ~n8083 & n17218 ;
  assign n17222 = n17221 ^ n17219 ^ 1'b0 ;
  assign n17223 = n15549 ^ n1495 ^ 1'b0 ;
  assign n17224 = ~n1577 & n16208 ;
  assign n17229 = n13680 ^ n2827 ^ 1'b0 ;
  assign n17225 = n1522 & n4235 ;
  assign n17226 = ~n7352 & n17225 ;
  assign n17227 = x0 & ~n17226 ;
  assign n17228 = ~n9172 & n17227 ;
  assign n17230 = n17229 ^ n17228 ^ 1'b0 ;
  assign n17231 = n10217 & n17230 ;
  assign n17232 = n2831 | n8403 ;
  assign n17233 = n12611 ^ n1402 ^ 1'b0 ;
  assign n17234 = n10261 & n15261 ;
  assign n17235 = ~n17233 & n17234 ;
  assign n17241 = n6201 & n14014 ;
  assign n17236 = ( n1298 & n4837 ) | ( n1298 & ~n10180 ) | ( n4837 & ~n10180 ) ;
  assign n17237 = n9930 & n17236 ;
  assign n17238 = ~n11839 & n17237 ;
  assign n17239 = n6415 ^ n4769 ^ 1'b0 ;
  assign n17240 = ~n17238 & n17239 ;
  assign n17242 = n17241 ^ n17240 ^ n1999 ;
  assign n17243 = ( n1864 & n6615 ) | ( n1864 & n16333 ) | ( n6615 & n16333 ) ;
  assign n17244 = n5458 & ~n14667 ;
  assign n17250 = n801 & ~n2900 ;
  assign n17245 = n4045 & ~n9940 ;
  assign n17246 = n2819 & ~n17245 ;
  assign n17247 = n15721 & n17246 ;
  assign n17248 = n16880 & ~n17247 ;
  assign n17249 = n17248 ^ n16291 ^ 1'b0 ;
  assign n17251 = n17250 ^ n17249 ^ 1'b0 ;
  assign n17252 = n4503 ^ n3938 ^ n3596 ;
  assign n17253 = n17252 ^ n9714 ^ 1'b0 ;
  assign n17254 = n4635 | n13574 ;
  assign n17255 = n9402 ^ n7609 ^ n3291 ;
  assign n17256 = n14505 | n17255 ;
  assign n17257 = n17256 ^ n9059 ^ 1'b0 ;
  assign n17258 = n8939 ^ n256 ^ 1'b0 ;
  assign n17259 = n17258 ^ n6639 ^ n6263 ;
  assign n17260 = n6983 & n10292 ;
  assign n17261 = n17259 | n17260 ;
  assign n17262 = n16467 ^ n3382 ^ n3034 ;
  assign n17263 = n6306 & n17262 ;
  assign n17264 = n16309 | n17263 ;
  assign n17265 = n6788 ^ n716 ^ 1'b0 ;
  assign n17266 = n3674 | n17265 ;
  assign n17267 = ( n9262 & n9667 ) | ( n9262 & ~n12588 ) | ( n9667 & ~n12588 ) ;
  assign n17268 = n2916 & n17267 ;
  assign n17269 = n17268 ^ n3305 ^ 1'b0 ;
  assign n17270 = n3036 & n8916 ;
  assign n17271 = n17270 ^ n13443 ^ 1'b0 ;
  assign n17273 = n14335 ^ n779 ^ 1'b0 ;
  assign n17274 = n17273 ^ n16032 ^ n13961 ;
  assign n17272 = n15653 ^ n13288 ^ 1'b0 ;
  assign n17275 = n17274 ^ n17272 ^ n5986 ;
  assign n17276 = n4230 & n11951 ;
  assign n17277 = n17276 ^ n14145 ^ 1'b0 ;
  assign n17278 = n642 | n8273 ;
  assign n17279 = ~n5726 & n12679 ;
  assign n17280 = n17279 ^ n3041 ^ 1'b0 ;
  assign n17281 = ~n6157 & n15948 ;
  assign n17282 = n17281 ^ n3705 ^ 1'b0 ;
  assign n17283 = n3491 & n17282 ;
  assign n17285 = x89 | n5581 ;
  assign n17284 = n2960 & n11558 ;
  assign n17286 = n17285 ^ n17284 ^ 1'b0 ;
  assign n17287 = n14087 & ~n17286 ;
  assign n17288 = ~n4177 & n11943 ;
  assign n17289 = n17288 ^ n8301 ^ 1'b0 ;
  assign n17293 = n3455 ^ n1213 ^ 1'b0 ;
  assign n17294 = n4099 | n17293 ;
  assign n17295 = n14526 | n17294 ;
  assign n17290 = n1123 | n3793 ;
  assign n17291 = n17290 ^ n4974 ^ 1'b0 ;
  assign n17292 = n15137 | n17291 ;
  assign n17296 = n17295 ^ n17292 ^ 1'b0 ;
  assign n17297 = n1879 & ~n6077 ;
  assign n17298 = ~n10913 & n17297 ;
  assign n17299 = n15578 & n17298 ;
  assign n17300 = n8034 ^ n2291 ^ 1'b0 ;
  assign n17301 = n9161 ^ n8534 ^ 1'b0 ;
  assign n17302 = n14376 ^ n6123 ^ n1494 ;
  assign n17303 = n1466 & ~n7220 ;
  assign n17304 = n15429 | n17303 ;
  assign n17306 = n2912 & n5488 ;
  assign n17307 = n3096 & ~n17306 ;
  assign n17308 = n17307 ^ n4037 ^ 1'b0 ;
  assign n17305 = n6335 & ~n9892 ;
  assign n17309 = n17308 ^ n17305 ^ 1'b0 ;
  assign n17310 = n10596 & ~n17309 ;
  assign n17311 = n2081 | n6122 ;
  assign n17312 = n17311 ^ n10077 ^ n1430 ;
  assign n17313 = n7325 ^ n1805 ^ 1'b0 ;
  assign n17314 = ~n14774 & n17313 ;
  assign n17315 = n17312 & n17314 ;
  assign n17316 = n17315 ^ n8756 ^ n7043 ;
  assign n17317 = ( n1997 & n5061 ) | ( n1997 & ~n11371 ) | ( n5061 & ~n11371 ) ;
  assign n17318 = n4931 & n15446 ;
  assign n17319 = n17318 ^ n3603 ^ 1'b0 ;
  assign n17320 = n4410 ^ n2326 ^ 1'b0 ;
  assign n17321 = n5104 & n17320 ;
  assign n17322 = n7678 | n8191 ;
  assign n17323 = n17321 | n17322 ;
  assign n17324 = n11853 ^ n3888 ^ 1'b0 ;
  assign n17325 = n1523 ^ n503 ^ 1'b0 ;
  assign n17326 = ~n3022 & n17325 ;
  assign n17327 = n17326 ^ n9457 ^ 1'b0 ;
  assign n17328 = n6036 & n17327 ;
  assign n17329 = x4 & n17328 ;
  assign n17330 = n17329 ^ n2936 ^ 1'b0 ;
  assign n17331 = n1004 | n7999 ;
  assign n17332 = n6220 ^ n3594 ^ 1'b0 ;
  assign n17333 = n10145 & ~n14009 ;
  assign n17334 = n5511 | n8246 ;
  assign n17335 = n3817 ^ n1185 ^ 1'b0 ;
  assign n17336 = n3034 | n17335 ;
  assign n17337 = ~n4672 & n8073 ;
  assign n17338 = n17336 & n17337 ;
  assign n17339 = n17338 ^ n12863 ^ n3966 ;
  assign n17340 = n5470 ^ x48 ^ 1'b0 ;
  assign n17343 = n16212 ^ n15466 ^ 1'b0 ;
  assign n17341 = n4843 ^ n915 ^ 1'b0 ;
  assign n17342 = ~n1336 & n17341 ;
  assign n17344 = n17343 ^ n17342 ^ 1'b0 ;
  assign n17345 = n6722 & n17344 ;
  assign n17346 = ~n2246 & n8064 ;
  assign n17347 = n17346 ^ n14701 ^ 1'b0 ;
  assign n17348 = n2130 & ~n5195 ;
  assign n17349 = ~n10239 & n17348 ;
  assign n17350 = n13787 ^ n5616 ^ n4498 ;
  assign n17351 = n12914 ^ n7365 ^ 1'b0 ;
  assign n17352 = n2497 | n17351 ;
  assign n17353 = n17352 ^ n17116 ^ 1'b0 ;
  assign n17354 = x33 & ~n1271 ;
  assign n17355 = ~n7137 & n17354 ;
  assign n17356 = n4510 | n9298 ;
  assign n17357 = n8802 & ~n17356 ;
  assign n17358 = n17355 | n17357 ;
  assign n17359 = n4877 & n11498 ;
  assign n17360 = n17359 ^ n5861 ^ 1'b0 ;
  assign n17361 = n15668 ^ n8785 ^ n3547 ;
  assign n17362 = n13412 & n13429 ;
  assign n17363 = n6580 ^ n2960 ^ 1'b0 ;
  assign n17364 = n17362 & ~n17363 ;
  assign n17365 = n5811 ^ n3876 ^ 1'b0 ;
  assign n17366 = n2580 & ~n17365 ;
  assign n17367 = n3134 | n15324 ;
  assign n17368 = n17366 | n17367 ;
  assign n17369 = n17364 & ~n17368 ;
  assign n17370 = n9041 & n14227 ;
  assign n17371 = n1921 & n2255 ;
  assign n17372 = n17371 ^ n6083 ^ 1'b0 ;
  assign n17373 = n2831 | n17372 ;
  assign n17374 = ~n3523 & n5530 ;
  assign n17375 = n17373 & ~n17374 ;
  assign n17376 = n6135 & n17375 ;
  assign n17377 = n3627 & ~n13025 ;
  assign n17378 = n17376 | n17377 ;
  assign n17379 = n17378 ^ n11981 ^ n3653 ;
  assign n17380 = n1504 | n17379 ;
  assign n17381 = n3936 ^ x106 ^ 1'b0 ;
  assign n17382 = ~n6101 & n17381 ;
  assign n17383 = n17382 ^ n3001 ^ 1'b0 ;
  assign n17384 = n16080 ^ n7545 ^ 1'b0 ;
  assign n17385 = n5777 ^ n2950 ^ 1'b0 ;
  assign n17386 = n4861 & ~n17385 ;
  assign n17387 = ~n4031 & n5749 ;
  assign n17388 = ~n9628 & n17387 ;
  assign n17389 = n17173 & n17388 ;
  assign n17390 = ~n17386 & n17389 ;
  assign n17391 = n3265 ^ x48 ^ 1'b0 ;
  assign n17392 = ~n7377 & n17391 ;
  assign n17393 = n17392 ^ n16527 ^ n11348 ;
  assign n17395 = n1283 | n4754 ;
  assign n17394 = n2929 & n4016 ;
  assign n17396 = n17395 ^ n17394 ^ 1'b0 ;
  assign n17397 = n558 & n9715 ;
  assign n17398 = ~n6040 & n7325 ;
  assign n17399 = n17398 ^ n11102 ^ n6526 ;
  assign n17400 = ~n7107 & n9168 ;
  assign n17401 = n17400 ^ n2466 ^ 1'b0 ;
  assign n17402 = n17401 ^ n1284 ^ 1'b0 ;
  assign n17403 = n13093 ^ n12737 ^ 1'b0 ;
  assign n17404 = n10715 ^ n7608 ^ 1'b0 ;
  assign n17405 = n11726 & n17404 ;
  assign n17406 = x232 | n1109 ;
  assign n17407 = ~n12859 & n17406 ;
  assign n17408 = ~n17405 & n17407 ;
  assign n17409 = ( n1315 & n4737 ) | ( n1315 & ~n13202 ) | ( n4737 & ~n13202 ) ;
  assign n17410 = n17409 ^ n13845 ^ n11465 ;
  assign n17411 = n17410 ^ n755 ^ 1'b0 ;
  assign n17412 = ~n7981 & n12680 ;
  assign n17413 = n9892 ^ n8001 ^ 1'b0 ;
  assign n17414 = n17413 ^ n4413 ^ 1'b0 ;
  assign n17415 = ( ~n1311 & n4452 ) | ( ~n1311 & n7519 ) | ( n4452 & n7519 ) ;
  assign n17416 = n4236 & ~n9992 ;
  assign n17417 = n17416 ^ n10169 ^ 1'b0 ;
  assign n17418 = n17415 & n17417 ;
  assign n17419 = n6527 & n17418 ;
  assign n17420 = ( ~x34 & x112 ) | ( ~x34 & n3370 ) | ( x112 & n3370 ) ;
  assign n17421 = n560 | n17420 ;
  assign n17422 = ~n5745 & n13236 ;
  assign n17423 = n6805 & n17422 ;
  assign n17425 = n13729 ^ n3704 ^ 1'b0 ;
  assign n17426 = n5749 & ~n17425 ;
  assign n17424 = ~n7990 & n14312 ;
  assign n17427 = n17426 ^ n17424 ^ 1'b0 ;
  assign n17428 = n14392 ^ n8293 ^ 1'b0 ;
  assign n17429 = n14976 ^ n9316 ^ n7435 ;
  assign n17430 = n7933 ^ n6475 ^ n5122 ;
  assign n17431 = n17430 ^ x225 ^ 1'b0 ;
  assign n17432 = n12040 ^ n7273 ^ 1'b0 ;
  assign n17433 = n5323 & ~n17432 ;
  assign n17434 = n16887 ^ n4791 ^ 1'b0 ;
  assign n17435 = n10663 ^ n2389 ^ 1'b0 ;
  assign n17436 = n2855 & ~n12366 ;
  assign n17437 = n17436 ^ n3296 ^ 1'b0 ;
  assign n17438 = n6639 | n14713 ;
  assign n17439 = ( n17376 & n17437 ) | ( n17376 & ~n17438 ) | ( n17437 & ~n17438 ) ;
  assign n17440 = n4649 | n14849 ;
  assign n17441 = n17440 ^ n15312 ^ 1'b0 ;
  assign n17442 = n2514 & n17441 ;
  assign n17443 = ( n1492 & n2983 ) | ( n1492 & ~n16753 ) | ( n2983 & ~n16753 ) ;
  assign n17444 = n4698 & n6364 ;
  assign n17445 = n15878 | n17444 ;
  assign n17446 = n17445 ^ n4712 ^ 1'b0 ;
  assign n17451 = ~n8321 & n10333 ;
  assign n17452 = n17451 ^ n6655 ^ 1'b0 ;
  assign n17447 = ~n708 & n6303 ;
  assign n17448 = n4648 | n6856 ;
  assign n17449 = n17448 ^ n11871 ^ n8900 ;
  assign n17450 = n17447 & ~n17449 ;
  assign n17453 = n17452 ^ n17450 ^ 1'b0 ;
  assign n17454 = n15721 | n16988 ;
  assign n17455 = ( n2964 & n8991 ) | ( n2964 & ~n10403 ) | ( n8991 & ~n10403 ) ;
  assign n17456 = n3085 & ~n17455 ;
  assign n17457 = ~n2782 & n11610 ;
  assign n17458 = n17456 | n17457 ;
  assign n17459 = n908 & ~n17458 ;
  assign n17460 = ( ~n2307 & n8280 ) | ( ~n2307 & n16283 ) | ( n8280 & n16283 ) ;
  assign n17461 = n5392 ^ n1303 ^ 1'b0 ;
  assign n17462 = ~n12481 & n17461 ;
  assign n17463 = n17462 ^ n3325 ^ 1'b0 ;
  assign n17464 = ~n825 & n17463 ;
  assign n17465 = n17464 ^ n12280 ^ 1'b0 ;
  assign n17466 = n6125 | n10724 ;
  assign n17467 = n5465 & ~n17466 ;
  assign n17468 = n5295 | n15559 ;
  assign n17469 = n4361 ^ n663 ^ 1'b0 ;
  assign n17470 = n5613 & ~n17469 ;
  assign n17471 = n17470 ^ n6923 ^ 1'b0 ;
  assign n17472 = n3156 | n9883 ;
  assign n17473 = n17471 & ~n17472 ;
  assign n17474 = n11692 & ~n17473 ;
  assign n17478 = n1097 & ~n1322 ;
  assign n17476 = n1379 | n16339 ;
  assign n17475 = n3249 & n5293 ;
  assign n17477 = n17476 ^ n17475 ^ 1'b0 ;
  assign n17479 = n17478 ^ n17477 ^ 1'b0 ;
  assign n17480 = n946 & ~n17479 ;
  assign n17481 = n6036 & ~n6679 ;
  assign n17482 = ~n17480 & n17481 ;
  assign n17483 = n13419 ^ n12891 ^ 1'b0 ;
  assign n17484 = ~n4842 & n7203 ;
  assign n17485 = x99 & n14099 ;
  assign n17486 = n4084 & n17485 ;
  assign n17487 = n789 & ~n2663 ;
  assign n17488 = n17487 ^ n11000 ^ 1'b0 ;
  assign n17489 = n10142 ^ n6179 ^ 1'b0 ;
  assign n17490 = ( n17486 & n17488 ) | ( n17486 & n17489 ) | ( n17488 & n17489 ) ;
  assign n17491 = n13410 ^ n8824 ^ 1'b0 ;
  assign n17492 = n1562 | n1801 ;
  assign n17493 = n17492 ^ n6219 ^ 1'b0 ;
  assign n17494 = ( n4488 & n17491 ) | ( n4488 & ~n17493 ) | ( n17491 & ~n17493 ) ;
  assign n17495 = n6748 ^ n344 ^ 1'b0 ;
  assign n17496 = x92 & n17495 ;
  assign n17497 = n2375 & n7232 ;
  assign n17498 = n3400 & ~n8015 ;
  assign n17499 = n17498 ^ n5637 ^ 1'b0 ;
  assign n17500 = n17499 ^ n12983 ^ 1'b0 ;
  assign n17501 = ~n5406 & n8344 ;
  assign n17502 = n3694 & n7417 ;
  assign n17503 = n8326 & n17502 ;
  assign n17504 = n2416 & ~n6964 ;
  assign n17505 = n17504 ^ n1500 ^ 1'b0 ;
  assign n17506 = n17505 ^ n10373 ^ 1'b0 ;
  assign n17507 = n17503 | n17506 ;
  assign n17508 = n1470 & n16807 ;
  assign n17509 = ~n3830 & n7873 ;
  assign n17510 = n17508 & ~n17509 ;
  assign n17511 = n17510 ^ n15899 ^ 1'b0 ;
  assign n17513 = n6098 & ~n8962 ;
  assign n17514 = n12226 & n17513 ;
  assign n17512 = n1332 & ~n7738 ;
  assign n17515 = n17514 ^ n17512 ^ 1'b0 ;
  assign n17519 = ~n473 & n4861 ;
  assign n17516 = n4327 & ~n4481 ;
  assign n17517 = n17516 ^ n2439 ^ 1'b0 ;
  assign n17518 = n17517 ^ n3571 ^ 1'b0 ;
  assign n17520 = n17519 ^ n17518 ^ 1'b0 ;
  assign n17521 = ( ~n772 & n4835 ) | ( ~n772 & n17520 ) | ( n4835 & n17520 ) ;
  assign n17522 = n13726 ^ n4144 ^ 1'b0 ;
  assign n17523 = n3042 | n8892 ;
  assign n17524 = n17523 ^ n10861 ^ 1'b0 ;
  assign n17525 = ~x49 & n11874 ;
  assign n17526 = n17525 ^ n11983 ^ n4361 ;
  assign n17527 = ~n2501 & n17526 ;
  assign n17528 = ~n7058 & n17527 ;
  assign n17530 = n7228 ^ n593 ^ 1'b0 ;
  assign n17531 = n2082 & n17530 ;
  assign n17532 = n417 & ~n15946 ;
  assign n17533 = ~n17531 & n17532 ;
  assign n17534 = n1132 & n7270 ;
  assign n17535 = n17533 & n17534 ;
  assign n17529 = n4514 & n7872 ;
  assign n17536 = n17535 ^ n17529 ^ 1'b0 ;
  assign n17537 = n5837 ^ n5266 ^ 1'b0 ;
  assign n17538 = n16429 ^ n14606 ^ 1'b0 ;
  assign n17539 = ~n1595 & n9819 ;
  assign n17540 = n4698 & n17539 ;
  assign n17541 = n10398 | n16471 ;
  assign n17542 = n9586 ^ n1682 ^ 1'b0 ;
  assign n17543 = n3903 & ~n17542 ;
  assign n17544 = n17543 ^ n2062 ^ 1'b0 ;
  assign n17545 = n15781 | n17544 ;
  assign n17546 = n3515 | n12556 ;
  assign n17547 = n1053 & n14603 ;
  assign n17548 = n17547 ^ n15870 ^ 1'b0 ;
  assign n17549 = n17546 | n17548 ;
  assign n17550 = n17549 ^ n14908 ^ 1'b0 ;
  assign n17551 = x127 & n3677 ;
  assign n17552 = n3325 | n5632 ;
  assign n17553 = n4409 | n17552 ;
  assign n17554 = n1473 & ~n12771 ;
  assign n17555 = n17554 ^ n16967 ^ 1'b0 ;
  assign n17556 = n13486 ^ n4750 ^ 1'b0 ;
  assign n17557 = n7674 ^ n7467 ^ 1'b0 ;
  assign n17558 = n8793 ^ n1010 ^ 1'b0 ;
  assign n17559 = n2191 & ~n11392 ;
  assign n17560 = n3818 & n17559 ;
  assign n17562 = n6238 & ~n12541 ;
  assign n17563 = n12947 ^ n7695 ^ 1'b0 ;
  assign n17564 = n17562 & n17563 ;
  assign n17561 = n9582 ^ n9492 ^ 1'b0 ;
  assign n17565 = n17564 ^ n17561 ^ n7175 ;
  assign n17566 = n7352 & n13139 ;
  assign n17567 = n1261 | n7964 ;
  assign n17568 = n4892 & n12225 ;
  assign n17569 = n15042 ^ n2062 ^ 1'b0 ;
  assign n17570 = n17569 ^ n14912 ^ 1'b0 ;
  assign n17571 = n1632 & n8921 ;
  assign n17572 = n3845 ^ n1078 ^ 1'b0 ;
  assign n17573 = n3163 & n17572 ;
  assign n17574 = n7872 & ~n13616 ;
  assign n17575 = n3474 & n6204 ;
  assign n17576 = ~n14532 & n16068 ;
  assign n17577 = n4026 & ~n6521 ;
  assign n17578 = ( n2942 & n8974 ) | ( n2942 & n17577 ) | ( n8974 & n17577 ) ;
  assign n17579 = n13255 ^ n9661 ^ 1'b0 ;
  assign n17580 = n5685 & n17579 ;
  assign n17581 = n15109 & n17580 ;
  assign n17582 = n17581 ^ n13054 ^ 1'b0 ;
  assign n17583 = n3106 | n17238 ;
  assign n17585 = n13486 & n16545 ;
  assign n17586 = ~n8656 & n17585 ;
  assign n17584 = n15904 & ~n16944 ;
  assign n17587 = n17586 ^ n17584 ^ 1'b0 ;
  assign n17588 = n10470 ^ n3515 ^ 1'b0 ;
  assign n17589 = n4921 & n15233 ;
  assign n17590 = ( n2789 & n4282 ) | ( n2789 & n17589 ) | ( n4282 & n17589 ) ;
  assign n17591 = n3131 & n5145 ;
  assign n17592 = n17591 ^ n1358 ^ 1'b0 ;
  assign n17593 = n17592 ^ n6591 ^ 1'b0 ;
  assign n17594 = ~n6828 & n17593 ;
  assign n17595 = ~n3082 & n17594 ;
  assign n17596 = n7771 & n17595 ;
  assign n17597 = ( n2659 & n6225 ) | ( n2659 & ~n9720 ) | ( n6225 & ~n9720 ) ;
  assign n17598 = n17597 ^ n4914 ^ 1'b0 ;
  assign n17599 = ~n17596 & n17598 ;
  assign n17600 = ~n686 & n1975 ;
  assign n17601 = x118 & n17600 ;
  assign n17602 = n10783 & ~n17601 ;
  assign n17603 = n6348 | n8297 ;
  assign n17604 = n9708 & ~n17603 ;
  assign n17605 = n17604 ^ n708 ^ 1'b0 ;
  assign n17606 = n5722 & ~n15261 ;
  assign n17607 = ~n5014 & n17606 ;
  assign n17608 = n5325 & ~n14715 ;
  assign n17609 = n17608 ^ n4294 ^ 1'b0 ;
  assign n17610 = ~n17607 & n17609 ;
  assign n17611 = n16178 ^ n7630 ^ n6604 ;
  assign n17612 = n8600 & n15928 ;
  assign n17613 = n16496 ^ n10092 ^ 1'b0 ;
  assign n17614 = n6106 & n13305 ;
  assign n17615 = n17614 ^ n6609 ^ 1'b0 ;
  assign n17616 = n769 & n17615 ;
  assign n17625 = n7734 & ~n13110 ;
  assign n17626 = n17625 ^ n14762 ^ 1'b0 ;
  assign n17620 = n3508 | n6559 ;
  assign n17621 = n17620 ^ n5029 ^ 1'b0 ;
  assign n17617 = n7205 ^ n5727 ^ 1'b0 ;
  assign n17618 = n17617 ^ n4428 ^ 1'b0 ;
  assign n17619 = n4119 | n17618 ;
  assign n17622 = n17621 ^ n17619 ^ 1'b0 ;
  assign n17623 = n1221 & n17622 ;
  assign n17624 = ~x62 & n17623 ;
  assign n17627 = n17626 ^ n17624 ^ 1'b0 ;
  assign n17628 = n15995 | n17627 ;
  assign n17629 = n4562 ^ n1900 ^ 1'b0 ;
  assign n17630 = n1039 & ~n17629 ;
  assign n17631 = n17630 ^ n2957 ^ 1'b0 ;
  assign n17632 = n10584 ^ n3778 ^ 1'b0 ;
  assign n17633 = ~n4855 & n17632 ;
  assign n17634 = n17633 ^ n1294 ^ 1'b0 ;
  assign n17635 = n17631 & n17634 ;
  assign n17636 = n13075 ^ n13016 ^ 1'b0 ;
  assign n17637 = n17636 ^ n11138 ^ 1'b0 ;
  assign n17638 = n16069 ^ n7116 ^ n3950 ;
  assign n17639 = n17638 ^ n9200 ^ n3929 ;
  assign n17641 = ( n4668 & n4706 ) | ( n4668 & ~n7110 ) | ( n4706 & ~n7110 ) ;
  assign n17640 = n10264 & ~n14514 ;
  assign n17642 = n17641 ^ n17640 ^ 1'b0 ;
  assign n17643 = n3151 & n4976 ;
  assign n17644 = n6110 ^ n3293 ^ 1'b0 ;
  assign n17645 = n11137 | n17644 ;
  assign n17646 = n14845 ^ n1347 ^ 1'b0 ;
  assign n17650 = x190 & ~n8956 ;
  assign n17651 = ( n1878 & n5054 ) | ( n1878 & n5921 ) | ( n5054 & n5921 ) ;
  assign n17652 = n8340 & ~n17651 ;
  assign n17653 = ~n17650 & n17652 ;
  assign n17654 = n17653 ^ n15950 ^ n608 ;
  assign n17647 = n15412 ^ n4832 ^ 1'b0 ;
  assign n17648 = ~n6218 & n17647 ;
  assign n17649 = n17648 ^ n2249 ^ 1'b0 ;
  assign n17655 = n17654 ^ n17649 ^ 1'b0 ;
  assign n17656 = n14975 ^ n8291 ^ 1'b0 ;
  assign n17657 = n13330 | n17656 ;
  assign n17660 = n7199 ^ n5769 ^ n5665 ;
  assign n17658 = n5059 ^ n3311 ^ 1'b0 ;
  assign n17659 = ~n4920 & n17658 ;
  assign n17661 = n17660 ^ n17659 ^ 1'b0 ;
  assign n17662 = x175 | n17661 ;
  assign n17663 = ~n17657 & n17662 ;
  assign n17664 = n7448 & ~n14723 ;
  assign n17665 = n631 & n17664 ;
  assign n17666 = n6908 & n17665 ;
  assign n17667 = n12647 ^ n4430 ^ 1'b0 ;
  assign n17668 = n17666 | n17667 ;
  assign n17669 = n8670 ^ x36 ^ 1'b0 ;
  assign n17670 = x30 & n13641 ;
  assign n17671 = n17669 & n17670 ;
  assign n17672 = n12590 & ~n17671 ;
  assign n17673 = n17672 ^ x18 ^ 1'b0 ;
  assign n17674 = n17651 ^ n880 ^ 1'b0 ;
  assign n17675 = n6780 & n15850 ;
  assign n17676 = n17675 ^ n1230 ^ 1'b0 ;
  assign n17677 = ~n7858 & n11431 ;
  assign n17678 = n13364 & n17677 ;
  assign n17679 = ~n17676 & n17678 ;
  assign n17682 = n12647 ^ n4465 ^ 1'b0 ;
  assign n17680 = n794 & ~n4352 ;
  assign n17681 = n7356 & n17680 ;
  assign n17683 = n17682 ^ n17681 ^ 1'b0 ;
  assign n17684 = n17679 & ~n17683 ;
  assign n17685 = ~n17674 & n17684 ;
  assign n17686 = n3521 & ~n6620 ;
  assign n17687 = n17686 ^ n11919 ^ 1'b0 ;
  assign n17690 = ~n980 & n6267 ;
  assign n17688 = n1779 & ~n8905 ;
  assign n17689 = n17688 ^ n2746 ^ 1'b0 ;
  assign n17691 = n17690 ^ n17689 ^ 1'b0 ;
  assign n17692 = ~n6981 & n17691 ;
  assign n17693 = n13498 ^ n2889 ^ n2055 ;
  assign n17694 = ( ~n3911 & n7667 ) | ( ~n3911 & n11450 ) | ( n7667 & n11450 ) ;
  assign n17695 = n17693 & n17694 ;
  assign n17696 = x86 & ~n17695 ;
  assign n17697 = n17696 ^ n13493 ^ 1'b0 ;
  assign n17698 = ~n15520 & n15998 ;
  assign n17699 = n17698 ^ n7848 ^ 1'b0 ;
  assign n17700 = n2326 & n5315 ;
  assign n17701 = n17700 ^ n5153 ^ 1'b0 ;
  assign n17702 = n1500 & n14078 ;
  assign n17703 = n8649 & n17702 ;
  assign n17704 = n2047 | n2065 ;
  assign n17705 = n15221 & ~n17704 ;
  assign n17706 = n4933 & n10398 ;
  assign n17707 = n17706 ^ n2341 ^ 1'b0 ;
  assign n17708 = n17707 ^ n11381 ^ n3433 ;
  assign n17709 = n17705 & n17708 ;
  assign n17710 = n16330 ^ n2740 ^ 1'b0 ;
  assign n17711 = ~n2482 & n4815 ;
  assign n17712 = n7306 | n17711 ;
  assign n17713 = n17712 ^ n4603 ^ 1'b0 ;
  assign n17714 = n1635 & ~n9529 ;
  assign n17715 = n17714 ^ n5786 ^ 1'b0 ;
  assign n17716 = ~n7463 & n17715 ;
  assign n17717 = n606 & n2372 ;
  assign n17718 = n17717 ^ n16290 ^ n3166 ;
  assign n17719 = ~n2936 & n5469 ;
  assign n17720 = n1486 & n2529 ;
  assign n17721 = n17720 ^ n1489 ^ 1'b0 ;
  assign n17722 = ~n6979 & n17721 ;
  assign n17723 = n15511 ^ n15069 ^ 1'b0 ;
  assign n17724 = n14645 & n15802 ;
  assign n17725 = n12850 & n17724 ;
  assign n17726 = n537 & n1437 ;
  assign n17727 = n5152 & ~n5912 ;
  assign n17728 = n17727 ^ n1879 ^ 1'b0 ;
  assign n17729 = n6433 & ~n17728 ;
  assign n17730 = n17729 ^ n3000 ^ 1'b0 ;
  assign n17731 = n15681 & n17730 ;
  assign n17732 = ~n8157 & n17731 ;
  assign n17733 = n9544 ^ n2930 ^ 1'b0 ;
  assign n17735 = x139 & ~n5266 ;
  assign n17736 = n17735 ^ n2681 ^ 1'b0 ;
  assign n17734 = n4025 | n5534 ;
  assign n17737 = n17736 ^ n17734 ^ 1'b0 ;
  assign n17738 = ( n6112 & n13809 ) | ( n6112 & n14141 ) | ( n13809 & n14141 ) ;
  assign n17739 = n3400 & ~n12680 ;
  assign n17740 = n3629 ^ n1912 ^ 1'b0 ;
  assign n17741 = n1757 & ~n17740 ;
  assign n17742 = n6862 ^ n1025 ^ 1'b0 ;
  assign n17743 = n6991 | n17742 ;
  assign n17744 = n3100 & ~n17743 ;
  assign n17745 = ~n17741 & n17744 ;
  assign n17746 = n294 & ~n4252 ;
  assign n17747 = n17746 ^ n15282 ^ 1'b0 ;
  assign n17748 = ( n8428 & n11462 ) | ( n8428 & n17747 ) | ( n11462 & n17747 ) ;
  assign n17749 = n395 & ~n13706 ;
  assign n17750 = n6075 & n17749 ;
  assign n17751 = n4042 | n4562 ;
  assign n17752 = n1519 ^ x177 ^ 1'b0 ;
  assign n17753 = ~n7381 & n17752 ;
  assign n17754 = n17753 ^ n11557 ^ 1'b0 ;
  assign n17755 = n5438 & ~n17754 ;
  assign n17756 = n15935 ^ n6802 ^ n5269 ;
  assign n17757 = ~n2013 & n14504 ;
  assign n17758 = n17756 & n17757 ;
  assign n17759 = n10009 ^ n7210 ^ 1'b0 ;
  assign n17760 = n14448 & n17759 ;
  assign n17761 = n17760 ^ n6996 ^ 1'b0 ;
  assign n17762 = ( n1605 & n4451 ) | ( n1605 & n6122 ) | ( n4451 & n6122 ) ;
  assign n17763 = n17762 ^ n334 ^ 1'b0 ;
  assign n17764 = n14957 & n17763 ;
  assign n17765 = n4624 ^ n4072 ^ 1'b0 ;
  assign n17766 = n5650 & ~n17765 ;
  assign n17767 = n13942 ^ n574 ^ 1'b0 ;
  assign n17768 = n15192 & ~n17767 ;
  assign n17769 = n2289 | n6602 ;
  assign n17770 = n4769 | n17769 ;
  assign n17771 = ( n2675 & ~n14992 ) | ( n2675 & n17770 ) | ( ~n14992 & n17770 ) ;
  assign n17772 = n12877 & ~n15224 ;
  assign n17773 = ~n1595 & n6529 ;
  assign n17774 = n10371 ^ n1914 ^ 1'b0 ;
  assign n17775 = n1720 & ~n17774 ;
  assign n17776 = n10797 | n14799 ;
  assign n17777 = n17776 ^ n6540 ^ 1'b0 ;
  assign n17778 = n10823 ^ n5835 ^ 1'b0 ;
  assign n17779 = n3780 ^ n1249 ^ x142 ;
  assign n17780 = n8782 & ~n17779 ;
  assign n17781 = n17780 ^ n12013 ^ 1'b0 ;
  assign n17782 = ~n10484 & n17781 ;
  assign n17783 = ( n14499 & n15268 ) | ( n14499 & ~n17782 ) | ( n15268 & ~n17782 ) ;
  assign n17784 = ~n5529 & n7665 ;
  assign n17785 = n1890 | n17784 ;
  assign n17787 = ~n2122 & n7822 ;
  assign n17786 = n7685 & ~n9649 ;
  assign n17788 = n17787 ^ n17786 ^ 1'b0 ;
  assign n17789 = n1163 ^ x40 ^ 1'b0 ;
  assign n17790 = n8717 & ~n17789 ;
  assign n17791 = n7875 ^ n2204 ^ 1'b0 ;
  assign n17792 = n17156 ^ n3641 ^ n3049 ;
  assign n17793 = ~n11053 & n17792 ;
  assign n17794 = n5313 & n5924 ;
  assign n17795 = ~n7303 & n17794 ;
  assign n17796 = n7586 & n17795 ;
  assign n17797 = n17796 ^ n4417 ^ 1'b0 ;
  assign n17798 = n2015 & n7492 ;
  assign n17799 = ~x197 & n17798 ;
  assign n17800 = n3795 & n4705 ;
  assign n17801 = n17799 & n17800 ;
  assign n17802 = n5783 ^ n2934 ^ 1'b0 ;
  assign n17803 = n17802 ^ n9505 ^ 1'b0 ;
  assign n17804 = n17801 | n17803 ;
  assign n17805 = n425 & ~n9729 ;
  assign n17806 = ~n4512 & n17805 ;
  assign n17807 = ~n8236 & n16331 ;
  assign n17808 = n17807 ^ n10897 ^ 1'b0 ;
  assign n17809 = ( ~n2235 & n2491 ) | ( ~n2235 & n17808 ) | ( n2491 & n17808 ) ;
  assign n17810 = n3557 ^ n1937 ^ 1'b0 ;
  assign n17811 = n12838 & ~n17810 ;
  assign n17812 = n7089 & n17811 ;
  assign n17813 = n4192 & ~n12192 ;
  assign n17814 = n466 & n9999 ;
  assign n17815 = n13643 ^ n9126 ^ 1'b0 ;
  assign n17816 = ~n812 & n14977 ;
  assign n17817 = n17815 & n17816 ;
  assign n17818 = n4420 ^ n3705 ^ 1'b0 ;
  assign n17819 = n9642 & n12108 ;
  assign n17820 = ~n17818 & n17819 ;
  assign n17821 = n5925 ^ n3828 ^ 1'b0 ;
  assign n17822 = n12767 & ~n13032 ;
  assign n17823 = ~n8366 & n17822 ;
  assign n17824 = n3385 | n6346 ;
  assign n17825 = n5094 ^ n4829 ^ 1'b0 ;
  assign n17826 = n11253 ^ n2420 ^ 1'b0 ;
  assign n17827 = n3874 & ~n6623 ;
  assign n17828 = n4315 & n11031 ;
  assign n17829 = n6337 ^ n2559 ^ 1'b0 ;
  assign n17830 = n11137 & ~n17829 ;
  assign n17831 = n1470 & n17830 ;
  assign n17832 = n17831 ^ n15991 ^ 1'b0 ;
  assign n17834 = n12481 | n15228 ;
  assign n17835 = n7678 & ~n17834 ;
  assign n17833 = n1388 ^ n858 ^ 1'b0 ;
  assign n17836 = n17835 ^ n17833 ^ 1'b0 ;
  assign n17837 = n8642 ^ x243 ^ 1'b0 ;
  assign n17838 = n3321 ^ n1645 ^ 1'b0 ;
  assign n17839 = n17837 & ~n17838 ;
  assign n17840 = n17839 ^ n9377 ^ 1'b0 ;
  assign n17841 = n2206 & n3447 ;
  assign n17842 = n9719 & n17841 ;
  assign n17843 = n17842 ^ n7379 ^ 1'b0 ;
  assign n17844 = n4600 ^ n272 ^ 1'b0 ;
  assign n17845 = n4748 & n5812 ;
  assign n17846 = n3183 & ~n17845 ;
  assign n17847 = ~n2735 & n15970 ;
  assign n17848 = n6851 | n14225 ;
  assign n17849 = n17848 ^ n1062 ^ 1'b0 ;
  assign n17850 = n8141 & n17849 ;
  assign n17851 = n3255 ^ n1833 ^ 1'b0 ;
  assign n17852 = n5209 | n17851 ;
  assign n17853 = n1161 & ~n17852 ;
  assign n17854 = n17853 ^ n8760 ^ 1'b0 ;
  assign n17855 = n12792 | n17854 ;
  assign n17856 = n11619 | n17855 ;
  assign n17857 = n1468 | n4924 ;
  assign n17858 = n17857 ^ n9113 ^ 1'b0 ;
  assign n17859 = n17858 ^ n13740 ^ 1'b0 ;
  assign n17860 = n453 & n8216 ;
  assign n17861 = n17860 ^ n14285 ^ 1'b0 ;
  assign n17862 = n17859 | n17861 ;
  assign n17863 = n17862 ^ n6434 ^ 1'b0 ;
  assign n17864 = n2925 ^ n2540 ^ 1'b0 ;
  assign n17865 = ( n3941 & ~n6121 ) | ( n3941 & n17864 ) | ( ~n6121 & n17864 ) ;
  assign n17866 = n16410 ^ n5392 ^ 1'b0 ;
  assign n17867 = n6414 | n15094 ;
  assign n17868 = n12044 & n17867 ;
  assign n17869 = n11853 ^ n2741 ^ 1'b0 ;
  assign n17870 = n17382 ^ n9540 ^ 1'b0 ;
  assign n17871 = n7646 | n17870 ;
  assign n17872 = n17871 ^ n2317 ^ 1'b0 ;
  assign n17873 = n1185 & n10655 ;
  assign n17874 = n10259 | n11237 ;
  assign n17875 = ~n6188 & n17874 ;
  assign n17876 = ~n9540 & n12134 ;
  assign n17877 = n4090 & n15739 ;
  assign n17878 = n5696 ^ n4222 ^ 1'b0 ;
  assign n17879 = ~n17877 & n17878 ;
  assign n17880 = n5186 ^ x26 ^ 1'b0 ;
  assign n17881 = n12524 & n17880 ;
  assign n17882 = n4642 ^ n2426 ^ 1'b0 ;
  assign n17883 = ~n6099 & n17882 ;
  assign n17884 = n17883 ^ n10416 ^ 1'b0 ;
  assign n17885 = n3996 ^ n3686 ^ 1'b0 ;
  assign n17886 = n5746 & n14509 ;
  assign n17887 = x244 | n1869 ;
  assign n17888 = n7644 ^ n5111 ^ 1'b0 ;
  assign n17889 = n6214 | n7000 ;
  assign n17890 = n17889 ^ n14181 ^ n6338 ;
  assign n17894 = n1926 & n9673 ;
  assign n17895 = n17894 ^ n4357 ^ 1'b0 ;
  assign n17891 = n4115 & n4539 ;
  assign n17892 = n2032 & n17891 ;
  assign n17893 = n13941 | n17892 ;
  assign n17896 = n17895 ^ n17893 ^ 1'b0 ;
  assign n17900 = ~n1417 & n6847 ;
  assign n17897 = n1048 | n11265 ;
  assign n17898 = n17897 ^ n9903 ^ 1'b0 ;
  assign n17899 = n17898 ^ n14285 ^ n6487 ;
  assign n17901 = n17900 ^ n17899 ^ 1'b0 ;
  assign n17902 = n7791 | n14849 ;
  assign n17904 = n485 ^ x101 ^ 1'b0 ;
  assign n17905 = n17357 | n17904 ;
  assign n17903 = x192 & ~n1312 ;
  assign n17906 = n17905 ^ n17903 ^ 1'b0 ;
  assign n17907 = n270 | n15001 ;
  assign n17908 = n11103 & n12926 ;
  assign n17909 = n5410 & ~n13811 ;
  assign n17910 = ~n591 & n17909 ;
  assign n17911 = ~n1813 & n7178 ;
  assign n17912 = n17911 ^ n17646 ^ 1'b0 ;
  assign n17913 = n2785 & n8280 ;
  assign n17914 = n17913 ^ n7263 ^ 1'b0 ;
  assign n17915 = n17661 ^ n16992 ^ 1'b0 ;
  assign n17916 = n10649 | n17915 ;
  assign n17917 = n4699 ^ x34 ^ 1'b0 ;
  assign n17918 = n16250 | n17917 ;
  assign n17919 = n17918 ^ n10968 ^ n6005 ;
  assign n17920 = n14310 & ~n17919 ;
  assign n17921 = ~n4787 & n17920 ;
  assign n17922 = n10279 ^ n4836 ^ n4578 ;
  assign n17923 = n8063 & ~n17922 ;
  assign n17924 = n15902 ^ n7672 ^ 1'b0 ;
  assign n17925 = n15874 | n17924 ;
  assign n17926 = n4249 ^ x39 ^ 1'b0 ;
  assign n17927 = n2678 & ~n3656 ;
  assign n17928 = n17927 ^ n1711 ^ 1'b0 ;
  assign n17929 = n469 | n7130 ;
  assign n17930 = n17928 | n17929 ;
  assign n17931 = n17930 ^ n3579 ^ 1'b0 ;
  assign n17932 = n10131 & n17931 ;
  assign n17933 = n1969 & n3939 ;
  assign n17934 = n3235 ^ n2296 ^ 1'b0 ;
  assign n17935 = n17933 | n17934 ;
  assign n17936 = n15428 ^ n10286 ^ 1'b0 ;
  assign n17937 = n3572 & ~n9823 ;
  assign n17938 = ~n10174 & n17937 ;
  assign n17939 = ~n1525 & n17938 ;
  assign n17940 = ~n6737 & n8265 ;
  assign n17941 = n11895 ^ n5371 ^ n1356 ;
  assign n17942 = n17940 & n17941 ;
  assign n17943 = ~n3804 & n7566 ;
  assign n17944 = n14102 & n17943 ;
  assign n17945 = n3057 | n5429 ;
  assign n17946 = n17945 ^ n10717 ^ 1'b0 ;
  assign n17948 = ~n2972 & n7005 ;
  assign n17949 = ~n7050 & n17948 ;
  assign n17947 = x126 & ~n3455 ;
  assign n17950 = n17949 ^ n17947 ^ 1'b0 ;
  assign n17951 = n11264 ^ n10321 ^ n9030 ;
  assign n17952 = n11961 ^ n1575 ^ 1'b0 ;
  assign n17953 = n15309 ^ n12207 ^ n9912 ;
  assign n17954 = n5301 & ~n9720 ;
  assign n17955 = n17954 ^ n6321 ^ 1'b0 ;
  assign n17956 = n11277 | n17955 ;
  assign n17957 = ~n6327 & n6357 ;
  assign n17958 = n12604 & ~n17957 ;
  assign n17959 = n15351 ^ n500 ^ 1'b0 ;
  assign n17960 = n12714 | n17959 ;
  assign n17961 = n5917 & ~n6508 ;
  assign n17962 = ~n17405 & n17961 ;
  assign n17963 = ( n17958 & ~n17960 ) | ( n17958 & n17962 ) | ( ~n17960 & n17962 ) ;
  assign n17964 = n1744 & ~n2739 ;
  assign n17965 = ( n1620 & ~n4115 ) | ( n1620 & n9457 ) | ( ~n4115 & n9457 ) ;
  assign n17966 = ~n6393 & n6592 ;
  assign n17967 = n17966 ^ n5124 ^ 1'b0 ;
  assign n17968 = n17967 ^ n6880 ^ n3393 ;
  assign n17969 = n4657 ^ n3496 ^ 1'b0 ;
  assign n17970 = n17968 | n17969 ;
  assign n17971 = n17965 | n17970 ;
  assign n17972 = n8746 & ~n17971 ;
  assign n17973 = n1638 & ~n12044 ;
  assign n17974 = ~n3444 & n17973 ;
  assign n17975 = n11590 ^ n2135 ^ 1'b0 ;
  assign n17976 = n17974 | n17975 ;
  assign n17977 = n1259 | n8746 ;
  assign n17978 = n5295 | n17977 ;
  assign n17979 = n17978 ^ n14442 ^ 1'b0 ;
  assign n17980 = n1328 | n2843 ;
  assign n17981 = n11042 & ~n17980 ;
  assign n17982 = n17372 ^ n2513 ^ 1'b0 ;
  assign n17983 = n3650 | n17982 ;
  assign n17984 = n5600 & ~n17983 ;
  assign n17985 = ~n4970 & n17984 ;
  assign n17986 = n15327 ^ n3822 ^ 1'b0 ;
  assign n17987 = n3738 ^ n1262 ^ 1'b0 ;
  assign n17988 = n15752 | n15832 ;
  assign n17989 = n13993 & ~n17988 ;
  assign n17990 = n17987 & ~n17989 ;
  assign n17991 = ~x163 & n17990 ;
  assign n17992 = n13312 & ~n13688 ;
  assign n17993 = n9495 ^ n2167 ^ 1'b0 ;
  assign n17994 = n5994 ^ n2312 ^ 1'b0 ;
  assign n17995 = n11369 ^ n1605 ^ 1'b0 ;
  assign n17996 = n17994 & n17995 ;
  assign n17997 = n890 & n12485 ;
  assign n17998 = n17997 ^ n3993 ^ 1'b0 ;
  assign n17999 = n1138 | n17998 ;
  assign n18000 = n17999 ^ n14749 ^ 1'b0 ;
  assign n18001 = n5315 ^ n550 ^ 1'b0 ;
  assign n18002 = n990 & n18001 ;
  assign n18003 = n1118 & ~n1943 ;
  assign n18004 = n16853 & ~n18003 ;
  assign n18005 = ~n18002 & n18004 ;
  assign n18006 = n710 | n6327 ;
  assign n18007 = n8175 | n18006 ;
  assign n18008 = n14765 | n18007 ;
  assign n18009 = n1140 | n18008 ;
  assign n18010 = n4899 ^ n1387 ^ 1'b0 ;
  assign n18011 = ~n1259 & n18010 ;
  assign n18012 = n18011 ^ n8751 ^ 1'b0 ;
  assign n18013 = ~n856 & n18012 ;
  assign n18014 = n10835 & n17531 ;
  assign n18015 = n1674 ^ n525 ^ 1'b0 ;
  assign n18016 = n8981 & ~n18015 ;
  assign n18017 = ( n11692 & n15777 ) | ( n11692 & n18016 ) | ( n15777 & n18016 ) ;
  assign n18018 = n12918 ^ n3619 ^ 1'b0 ;
  assign n18019 = n10857 ^ n7241 ^ 1'b0 ;
  assign n18020 = ( n1653 & ~n18018 ) | ( n1653 & n18019 ) | ( ~n18018 & n18019 ) ;
  assign n18021 = n4773 ^ n258 ^ 1'b0 ;
  assign n18022 = n15347 & ~n18021 ;
  assign n18023 = n318 & n3812 ;
  assign n18027 = n12638 ^ n9307 ^ n9057 ;
  assign n18024 = n8815 & n11166 ;
  assign n18025 = n16906 ^ n4368 ^ 1'b0 ;
  assign n18026 = ~n18024 & n18025 ;
  assign n18028 = n18027 ^ n18026 ^ 1'b0 ;
  assign n18029 = n4828 ^ n4659 ^ 1'b0 ;
  assign n18030 = n6931 | n18029 ;
  assign n18031 = n18030 ^ n4356 ^ 1'b0 ;
  assign n18032 = n4209 | n18031 ;
  assign n18033 = n18032 ^ n7028 ^ 1'b0 ;
  assign n18034 = n12556 ^ n10231 ^ 1'b0 ;
  assign n18035 = n4803 & ~n18034 ;
  assign n18036 = n6157 | n6416 ;
  assign n18037 = n18036 ^ n13596 ^ 1'b0 ;
  assign n18038 = n13569 & n14812 ;
  assign n18039 = n18038 ^ n9556 ^ 1'b0 ;
  assign n18040 = ~x191 & n4605 ;
  assign n18041 = n16492 ^ n4085 ^ 1'b0 ;
  assign n18042 = ~n8207 & n10148 ;
  assign n18043 = n3290 ^ n1023 ^ 1'b0 ;
  assign n18044 = n8425 | n10893 ;
  assign n18045 = n18044 ^ n3189 ^ 1'b0 ;
  assign n18046 = ( n6171 & ~n13494 ) | ( n6171 & n18045 ) | ( ~n13494 & n18045 ) ;
  assign n18047 = n18043 & n18046 ;
  assign n18048 = ~n18042 & n18047 ;
  assign n18049 = ~n766 & n15835 ;
  assign n18050 = n18049 ^ n6695 ^ 1'b0 ;
  assign n18051 = ~n13769 & n17684 ;
  assign n18052 = ~n11649 & n18051 ;
  assign n18053 = n7306 ^ n2928 ^ 1'b0 ;
  assign n18054 = n10407 ^ n9072 ^ 1'b0 ;
  assign n18055 = x13 & ~n7032 ;
  assign n18056 = n1333 | n12773 ;
  assign n18057 = n9572 & ~n18056 ;
  assign n18058 = n16491 ^ n6079 ^ 1'b0 ;
  assign n18059 = n6670 & n18058 ;
  assign n18060 = n18059 ^ n6243 ^ 1'b0 ;
  assign n18061 = n12269 & n18060 ;
  assign n18062 = n3809 & n18061 ;
  assign n18063 = n7765 & ~n18062 ;
  assign n18064 = n18063 ^ n6340 ^ 1'b0 ;
  assign n18065 = ( x192 & n13071 ) | ( x192 & ~n14805 ) | ( n13071 & ~n14805 ) ;
  assign n18066 = n7061 ^ n2011 ^ 1'b0 ;
  assign n18067 = ~n4210 & n18066 ;
  assign n18068 = n18067 ^ n7671 ^ 1'b0 ;
  assign n18069 = n16674 & ~n18068 ;
  assign n18070 = n18069 ^ n16849 ^ n258 ;
  assign n18071 = n10851 | n12723 ;
  assign n18072 = n256 | n4481 ;
  assign n18073 = ~n8311 & n14779 ;
  assign n18074 = ~n15097 & n18073 ;
  assign n18075 = n18074 ^ n13030 ^ 1'b0 ;
  assign n18076 = n18075 ^ n13964 ^ n11268 ;
  assign n18077 = n3734 & n15210 ;
  assign n18078 = n18077 ^ n4906 ^ 1'b0 ;
  assign n18079 = n14562 & ~n15037 ;
  assign n18080 = n1395 & ~n1750 ;
  assign n18081 = n18080 ^ n1690 ^ 1'b0 ;
  assign n18082 = n7710 & n18081 ;
  assign n18083 = ~n9252 & n18082 ;
  assign n18085 = ~n8597 & n12625 ;
  assign n18086 = n18085 ^ n7056 ^ 1'b0 ;
  assign n18087 = ~n9085 & n18086 ;
  assign n18084 = n7771 ^ n1527 ^ 1'b0 ;
  assign n18088 = n18087 ^ n18084 ^ n4234 ;
  assign n18089 = n10679 & ~n18088 ;
  assign n18097 = n6703 & ~n10164 ;
  assign n18098 = n18097 ^ n7298 ^ 1'b0 ;
  assign n18090 = ~n1813 & n7260 ;
  assign n18091 = n2171 | n6207 ;
  assign n18092 = n18090 | n18091 ;
  assign n18093 = n9459 & n13306 ;
  assign n18094 = n18093 ^ n6424 ^ 1'b0 ;
  assign n18095 = n5820 | n18094 ;
  assign n18096 = n18092 | n18095 ;
  assign n18099 = n18098 ^ n18096 ^ 1'b0 ;
  assign n18100 = n353 | n9777 ;
  assign n18101 = n3231 | n18100 ;
  assign n18102 = n18101 ^ n10284 ^ 1'b0 ;
  assign n18103 = n5248 & ~n17780 ;
  assign n18104 = n18103 ^ n17051 ^ 1'b0 ;
  assign n18105 = ~n18102 & n18104 ;
  assign n18106 = n18105 ^ n2143 ^ 1'b0 ;
  assign n18107 = n7482 | n11751 ;
  assign n18108 = n4678 ^ n1505 ^ 1'b0 ;
  assign n18109 = n2117 & n11017 ;
  assign n18110 = ~n18108 & n18109 ;
  assign n18111 = n5371 | n5538 ;
  assign n18112 = n4445 | n18111 ;
  assign n18113 = n809 | n2946 ;
  assign n18114 = n18113 ^ n8100 ^ 1'b0 ;
  assign n18115 = n874 & n2232 ;
  assign n18116 = n7506 & ~n18115 ;
  assign n18117 = n18116 ^ n5328 ^ 1'b0 ;
  assign n18118 = n18114 & n18117 ;
  assign n18122 = ( n1986 & n11482 ) | ( n1986 & n11659 ) | ( n11482 & n11659 ) ;
  assign n18123 = n13629 & n18122 ;
  assign n18119 = x201 & ~n867 ;
  assign n18120 = n18119 ^ n4099 ^ 1'b0 ;
  assign n18121 = ~n17397 & n18120 ;
  assign n18124 = n18123 ^ n18121 ^ 1'b0 ;
  assign n18132 = n3728 & ~n6406 ;
  assign n18133 = ~n3853 & n18132 ;
  assign n18134 = n1611 & ~n18133 ;
  assign n18135 = n18134 ^ n1175 ^ 1'b0 ;
  assign n18130 = ~n579 & n12483 ;
  assign n18131 = n18130 ^ n7590 ^ 1'b0 ;
  assign n18136 = n18135 ^ n18131 ^ n15752 ;
  assign n18127 = n7392 & n9327 ;
  assign n18128 = n18127 ^ n8380 ^ 1'b0 ;
  assign n18125 = ~n10039 & n11775 ;
  assign n18126 = n18125 ^ n7083 ^ 1'b0 ;
  assign n18129 = n18128 ^ n18126 ^ x128 ;
  assign n18137 = n18136 ^ n18129 ^ 1'b0 ;
  assign n18138 = n14895 ^ n2349 ^ 1'b0 ;
  assign n18140 = x1 & n14972 ;
  assign n18141 = n347 & n18140 ;
  assign n18139 = n9976 & ~n17477 ;
  assign n18142 = n18141 ^ n18139 ^ 1'b0 ;
  assign n18143 = n13664 ^ n1079 ^ 1'b0 ;
  assign n18144 = n14025 | n18143 ;
  assign n18145 = n12832 & ~n18144 ;
  assign n18146 = n10174 ^ n3488 ^ 1'b0 ;
  assign n18147 = n6741 ^ n4107 ^ 1'b0 ;
  assign n18148 = n18147 ^ n8103 ^ 1'b0 ;
  assign n18149 = n18146 & ~n18148 ;
  assign n18150 = n9970 | n18149 ;
  assign n18151 = n11920 ^ n2679 ^ 1'b0 ;
  assign n18152 = n18150 | n18151 ;
  assign n18153 = n4421 ^ n2893 ^ 1'b0 ;
  assign n18154 = n10777 & n18153 ;
  assign n18155 = ( n9904 & n14081 ) | ( n9904 & ~n18154 ) | ( n14081 & ~n18154 ) ;
  assign n18156 = ~n6444 & n15391 ;
  assign n18157 = ~n1611 & n18156 ;
  assign n18158 = n880 & n2133 ;
  assign n18159 = n1571 & n10178 ;
  assign n18160 = n5608 & n18159 ;
  assign n18161 = ( n4209 & n11193 ) | ( n4209 & ~n15964 ) | ( n11193 & ~n15964 ) ;
  assign n18162 = n18161 ^ n5625 ^ 1'b0 ;
  assign n18163 = n3850 & n4656 ;
  assign n18164 = n7814 & n10009 ;
  assign n18165 = n18164 ^ n673 ^ 1'b0 ;
  assign n18166 = n14425 | n18165 ;
  assign n18168 = n394 | n3300 ;
  assign n18167 = n2779 & n15320 ;
  assign n18169 = n18168 ^ n18167 ^ 1'b0 ;
  assign n18170 = n4666 ^ n4553 ^ 1'b0 ;
  assign n18171 = ~n5700 & n18170 ;
  assign n18172 = n13500 ^ n4686 ^ 1'b0 ;
  assign n18173 = n4185 | n18172 ;
  assign n18174 = n18173 ^ n10655 ^ 1'b0 ;
  assign n18181 = n4797 & n17415 ;
  assign n18182 = n9540 | n18181 ;
  assign n18176 = n5782 ^ n2357 ^ 1'b0 ;
  assign n18177 = n1628 | n18176 ;
  assign n18175 = ~n9774 & n16350 ;
  assign n18178 = n18177 ^ n18175 ^ 1'b0 ;
  assign n18179 = n5482 & n18178 ;
  assign n18180 = n18179 ^ n5754 ^ 1'b0 ;
  assign n18183 = n18182 ^ n18180 ^ 1'b0 ;
  assign n18184 = ~n10364 & n15760 ;
  assign n18185 = n6300 & n13077 ;
  assign n18186 = ~n1866 & n18185 ;
  assign n18187 = ~n6693 & n10900 ;
  assign n18188 = n18187 ^ x2 ^ 1'b0 ;
  assign n18189 = ~n606 & n3853 ;
  assign n18190 = n18189 ^ n5278 ^ 1'b0 ;
  assign n18191 = n18190 ^ n3240 ^ 1'b0 ;
  assign n18192 = n7381 & ~n18191 ;
  assign n18193 = ~n1114 & n2746 ;
  assign n18194 = n4958 & n18193 ;
  assign n18195 = n16471 ^ n4553 ^ 1'b0 ;
  assign n18196 = ( n2783 & n18194 ) | ( n2783 & n18195 ) | ( n18194 & n18195 ) ;
  assign n18197 = ~n13286 & n14166 ;
  assign n18198 = n18197 ^ n2442 ^ 1'b0 ;
  assign n18199 = n1045 & ~n4719 ;
  assign n18200 = ~n8270 & n18199 ;
  assign n18201 = n7298 & ~n18200 ;
  assign n18202 = ~n7298 & n18201 ;
  assign n18203 = x187 & ~n18202 ;
  assign n18204 = n18203 ^ n9964 ^ 1'b0 ;
  assign n18205 = ~n992 & n11585 ;
  assign n18206 = n8530 ^ n7042 ^ 1'b0 ;
  assign n18207 = n6920 & n18206 ;
  assign n18208 = n18207 ^ n956 ^ 1'b0 ;
  assign n18209 = n18208 ^ n7745 ^ 1'b0 ;
  assign n18210 = n16665 ^ n5618 ^ 1'b0 ;
  assign n18211 = ~n1071 & n18210 ;
  assign n18212 = n11290 ^ n10250 ^ 1'b0 ;
  assign n18213 = n5686 & n18212 ;
  assign n18214 = n6803 ^ n6464 ^ 1'b0 ;
  assign n18215 = n7920 & ~n18214 ;
  assign n18216 = n18213 & n18215 ;
  assign n18217 = ~n3864 & n18216 ;
  assign n18218 = n18217 ^ n16543 ^ 1'b0 ;
  assign n18219 = ~n5771 & n14511 ;
  assign n18220 = n17297 ^ n1566 ^ 1'b0 ;
  assign n18221 = n5881 & ~n18220 ;
  assign n18222 = ( n3590 & ~n11153 ) | ( n3590 & n18221 ) | ( ~n11153 & n18221 ) ;
  assign n18223 = n18222 ^ n12280 ^ 1'b0 ;
  assign n18225 = n18131 ^ n8360 ^ 1'b0 ;
  assign n18226 = n5827 & ~n18225 ;
  assign n18224 = n1208 | n10515 ;
  assign n18227 = n18226 ^ n18224 ^ 1'b0 ;
  assign n18228 = n17791 | n18227 ;
  assign n18229 = n3886 & n10650 ;
  assign n18230 = ~n6639 & n18229 ;
  assign n18231 = n16042 & n18230 ;
  assign n18232 = n15695 ^ n12009 ^ 1'b0 ;
  assign n18233 = n966 & n15745 ;
  assign n18234 = n9536 ^ n4023 ^ 1'b0 ;
  assign n18235 = n2725 | n18234 ;
  assign n18236 = n7659 & ~n18235 ;
  assign n18237 = n18236 ^ x32 ^ 1'b0 ;
  assign n18238 = ~n10988 & n12839 ;
  assign n18239 = n9109 & n18238 ;
  assign n18240 = n9002 & ~n13620 ;
  assign n18241 = n18240 ^ n9708 ^ n1389 ;
  assign n18242 = n15662 | n18241 ;
  assign n18243 = n15867 ^ n5021 ^ 1'b0 ;
  assign n18244 = n1389 ^ n604 ^ 1'b0 ;
  assign n18245 = ~n16845 & n17452 ;
  assign n18246 = n18245 ^ n6737 ^ 1'b0 ;
  assign n18247 = n7070 & n16195 ;
  assign n18248 = ~n12994 & n18247 ;
  assign n18249 = n18248 ^ n3235 ^ 1'b0 ;
  assign n18250 = n12576 | n18249 ;
  assign n18251 = n3372 & n11271 ;
  assign n18252 = ~n17526 & n18251 ;
  assign n18253 = n18252 ^ n15984 ^ 1'b0 ;
  assign n18254 = n17641 ^ n4367 ^ 1'b0 ;
  assign n18255 = n1190 & n5261 ;
  assign n18256 = n18255 ^ n9529 ^ 1'b0 ;
  assign n18257 = n13189 & n18256 ;
  assign n18258 = ~n315 & n7070 ;
  assign n18259 = ~n897 & n9353 ;
  assign n18260 = n18258 & ~n18259 ;
  assign n18261 = n18260 ^ n8759 ^ 1'b0 ;
  assign n18262 = ~n4807 & n7147 ;
  assign n18263 = n9532 & n18262 ;
  assign n18264 = ~n2506 & n4705 ;
  assign n18265 = n2082 & n18264 ;
  assign n18266 = n18265 ^ n16975 ^ 1'b0 ;
  assign n18267 = n16582 ^ n7691 ^ 1'b0 ;
  assign n18272 = n7195 ^ n2351 ^ 1'b0 ;
  assign n18273 = n4342 | n18272 ;
  assign n18274 = n860 | n18273 ;
  assign n18275 = n18274 ^ n3069 ^ 1'b0 ;
  assign n18268 = n9317 ^ n6317 ^ 1'b0 ;
  assign n18269 = n1612 & n18268 ;
  assign n18270 = n18269 ^ n15579 ^ 1'b0 ;
  assign n18271 = n4943 & ~n18270 ;
  assign n18276 = n18275 ^ n18271 ^ 1'b0 ;
  assign n18277 = n4767 & n5660 ;
  assign n18282 = n5879 & ~n15668 ;
  assign n18278 = n9982 | n13360 ;
  assign n18279 = n18278 ^ n1516 ^ n1392 ;
  assign n18280 = n16482 & n18279 ;
  assign n18281 = n18280 ^ n5225 ^ 1'b0 ;
  assign n18283 = n18282 ^ n18281 ^ 1'b0 ;
  assign n18284 = ~n15523 & n18283 ;
  assign n18286 = n6821 ^ n6547 ^ 1'b0 ;
  assign n18285 = n5502 ^ n1386 ^ 1'b0 ;
  assign n18287 = n18286 ^ n18285 ^ 1'b0 ;
  assign n18288 = n9516 ^ n5154 ^ 1'b0 ;
  assign n18289 = n18288 ^ n5894 ^ n3508 ;
  assign n18290 = n18289 ^ n13812 ^ 1'b0 ;
  assign n18291 = n13729 ^ n7238 ^ 1'b0 ;
  assign n18292 = n5208 & n18291 ;
  assign n18293 = n8508 & n18292 ;
  assign n18294 = n10215 ^ x237 ^ 1'b0 ;
  assign n18295 = ~n865 & n18294 ;
  assign n18296 = n15643 ^ n13952 ^ n7123 ;
  assign n18297 = n5465 ^ n1006 ^ 1'b0 ;
  assign n18298 = n18297 ^ n7002 ^ 1'b0 ;
  assign n18299 = n6456 | n7828 ;
  assign n18300 = n18298 | n18299 ;
  assign n18301 = ~n302 & n18300 ;
  assign n18302 = n18301 ^ n17638 ^ 1'b0 ;
  assign n18303 = n14106 ^ n2246 ^ 1'b0 ;
  assign n18305 = n2900 & ~n4430 ;
  assign n18306 = n6144 & n18305 ;
  assign n18304 = n1506 & n11379 ;
  assign n18307 = n18306 ^ n18304 ^ 1'b0 ;
  assign n18308 = n2370 ^ n2131 ^ 1'b0 ;
  assign n18309 = n18307 & ~n18308 ;
  assign n18310 = n14546 ^ n7887 ^ n3729 ;
  assign n18311 = n6479 ^ x192 ^ 1'b0 ;
  assign n18312 = n18310 & n18311 ;
  assign n18313 = ( ~n1169 & n1589 ) | ( ~n1169 & n5428 ) | ( n1589 & n5428 ) ;
  assign n18314 = n5219 ^ n4327 ^ n2035 ;
  assign n18315 = n18314 ^ n17156 ^ n13433 ;
  assign n18316 = ~n1695 & n11534 ;
  assign n18317 = n17919 & n18316 ;
  assign n18318 = n3915 & ~n8724 ;
  assign n18319 = ( n1255 & n7806 ) | ( n1255 & ~n12777 ) | ( n7806 & ~n12777 ) ;
  assign n18320 = n8815 ^ n5023 ^ 1'b0 ;
  assign n18321 = n5459 & ~n18320 ;
  assign n18322 = n3159 | n17957 ;
  assign n18323 = n17957 & ~n18322 ;
  assign n18324 = n7353 ^ n3508 ^ 1'b0 ;
  assign n18325 = ( n977 & n1148 ) | ( n977 & ~n7355 ) | ( n1148 & ~n7355 ) ;
  assign n18326 = n6583 ^ n2901 ^ 1'b0 ;
  assign n18327 = n18326 ^ n977 ^ 1'b0 ;
  assign n18328 = n6546 & ~n18327 ;
  assign n18329 = n18328 ^ n18146 ^ 1'b0 ;
  assign n18330 = n16730 | n18329 ;
  assign n18331 = ~n817 & n6350 ;
  assign n18333 = n9385 | n16491 ;
  assign n18334 = n18333 ^ n10577 ^ 1'b0 ;
  assign n18335 = n10442 & n18334 ;
  assign n18336 = n18335 ^ n2070 ^ 1'b0 ;
  assign n18337 = n12328 ^ n2466 ^ 1'b0 ;
  assign n18338 = n18336 & n18337 ;
  assign n18332 = n2281 | n11500 ;
  assign n18339 = n18338 ^ n18332 ^ 1'b0 ;
  assign n18340 = n18339 ^ n16237 ^ 1'b0 ;
  assign n18341 = n8513 | n16129 ;
  assign n18342 = n7910 & ~n11157 ;
  assign n18343 = n17854 & n18342 ;
  assign n18344 = n5291 & ~n18343 ;
  assign n18345 = n18344 ^ n6628 ^ 1'b0 ;
  assign n18346 = n1909 & n13793 ;
  assign n18347 = n6031 & ~n18346 ;
  assign n18348 = ~n12338 & n18347 ;
  assign n18349 = ~n5639 & n14456 ;
  assign n18350 = n18349 ^ n17619 ^ 1'b0 ;
  assign n18351 = n810 | n9844 ;
  assign n18352 = n18351 ^ n9957 ^ 1'b0 ;
  assign n18353 = n4733 & ~n18352 ;
  assign n18354 = ~n847 & n18353 ;
  assign n18355 = n5573 | n13078 ;
  assign n18356 = n16374 & ~n18355 ;
  assign n18357 = ~n4484 & n15712 ;
  assign n18358 = n1351 & n14590 ;
  assign n18359 = ~n6662 & n18358 ;
  assign n18360 = n18359 ^ n12879 ^ 1'b0 ;
  assign n18361 = n8395 ^ n3202 ^ n1165 ;
  assign n18362 = n5867 | n18361 ;
  assign n18363 = n16989 ^ n13978 ^ 1'b0 ;
  assign n18364 = n2002 & n18363 ;
  assign n18365 = n18362 & n18364 ;
  assign n18366 = n5070 & ~n13374 ;
  assign n18367 = ~n9076 & n18366 ;
  assign n18368 = n12660 ^ n4906 ^ 1'b0 ;
  assign n18369 = ~n12936 & n18368 ;
  assign n18370 = n1093 & n5532 ;
  assign n18371 = n18370 ^ n1956 ^ 1'b0 ;
  assign n18372 = n8002 & ~n18371 ;
  assign n18373 = n18371 & n18372 ;
  assign n18374 = n8740 & n14840 ;
  assign n18375 = ~n14840 & n18374 ;
  assign n18376 = n11347 & n18375 ;
  assign n18377 = n18376 ^ n6187 ^ 1'b0 ;
  assign n18378 = n18373 | n18377 ;
  assign n18379 = n2262 & n5621 ;
  assign n18380 = n18379 ^ n9924 ^ 1'b0 ;
  assign n18381 = ~n7736 & n10950 ;
  assign n18382 = n18381 ^ n12167 ^ 1'b0 ;
  assign n18383 = ~n12737 & n18382 ;
  assign n18384 = n3820 | n18383 ;
  assign n18385 = n4836 ^ n1336 ^ 1'b0 ;
  assign n18386 = n18385 ^ n15294 ^ 1'b0 ;
  assign n18387 = n11372 ^ n6629 ^ 1'b0 ;
  assign n18388 = n11394 ^ x64 ^ 1'b0 ;
  assign n18389 = n18388 ^ n6959 ^ 1'b0 ;
  assign n18390 = n18387 & ~n18389 ;
  assign n18391 = ~x55 & n11367 ;
  assign n18392 = n9080 ^ n6202 ^ 1'b0 ;
  assign n18393 = n2489 | n18392 ;
  assign n18394 = n13785 & ~n18393 ;
  assign n18395 = n18391 & n18394 ;
  assign n18396 = ~n6324 & n18395 ;
  assign n18397 = n15089 ^ n6073 ^ 1'b0 ;
  assign n18398 = n946 & n7364 ;
  assign n18399 = n8725 & n18398 ;
  assign n18400 = n5849 ^ n2056 ^ 1'b0 ;
  assign n18401 = n4134 | n18083 ;
  assign n18402 = n1725 | n9057 ;
  assign n18403 = n12809 & n17708 ;
  assign n18404 = ~n1217 & n18403 ;
  assign n18405 = n18404 ^ n826 ^ 1'b0 ;
  assign n18406 = n8380 | n18405 ;
  assign n18407 = n4374 & ~n18181 ;
  assign n18408 = n18407 ^ n7210 ^ n2504 ;
  assign n18409 = n7448 | n7689 ;
  assign n18410 = n5927 & ~n18409 ;
  assign n18411 = n8030 & ~n18410 ;
  assign n18412 = n6094 ^ n4986 ^ 1'b0 ;
  assign n18413 = n7476 & ~n18412 ;
  assign n18414 = n13297 & n18413 ;
  assign n18415 = n17662 ^ n5662 ^ 1'b0 ;
  assign n18416 = n9310 ^ n289 ^ 1'b0 ;
  assign n18417 = n11093 ^ n9654 ^ 1'b0 ;
  assign n18418 = n1098 | n2687 ;
  assign n18419 = n18417 | n18418 ;
  assign n18420 = n1088 & ~n1678 ;
  assign n18421 = n6397 ^ n4277 ^ 1'b0 ;
  assign n18422 = n18420 & ~n18421 ;
  assign n18423 = n17690 ^ n5075 ^ 1'b0 ;
  assign n18424 = n3025 & ~n4542 ;
  assign n18425 = n18424 ^ n10941 ^ 1'b0 ;
  assign n18426 = n18425 ^ n7547 ^ 1'b0 ;
  assign n18427 = n18426 ^ n16348 ^ n10564 ;
  assign n18428 = n18427 ^ n5523 ^ 1'b0 ;
  assign n18429 = n4066 ^ n1369 ^ 1'b0 ;
  assign n18430 = ~n14065 & n18429 ;
  assign n18431 = ~n5864 & n8081 ;
  assign n18432 = ~n3871 & n18431 ;
  assign n18433 = n4203 & ~n11451 ;
  assign n18434 = n6875 ^ n270 ^ 1'b0 ;
  assign n18438 = x137 & n1433 ;
  assign n18439 = ~x137 & n18438 ;
  assign n18435 = n1619 & ~n9456 ;
  assign n18436 = n18435 ^ n566 ^ 1'b0 ;
  assign n18437 = n8438 & ~n18436 ;
  assign n18440 = n18439 ^ n18437 ^ 1'b0 ;
  assign n18443 = n6638 & n12557 ;
  assign n18441 = n3258 & n14652 ;
  assign n18442 = n7321 & n18441 ;
  assign n18444 = n18443 ^ n18442 ^ 1'b0 ;
  assign n18445 = ( ~n7576 & n18440 ) | ( ~n7576 & n18444 ) | ( n18440 & n18444 ) ;
  assign n18446 = n18445 ^ n15754 ^ 1'b0 ;
  assign n18447 = n18434 & n18446 ;
  assign n18448 = n3416 & ~n14622 ;
  assign n18449 = n18448 ^ n9876 ^ 1'b0 ;
  assign n18452 = n7025 ^ n3174 ^ 1'b0 ;
  assign n18450 = n11443 ^ n4795 ^ n3614 ;
  assign n18451 = n13830 & n18450 ;
  assign n18453 = n18452 ^ n18451 ^ 1'b0 ;
  assign n18455 = n2998 & ~n13570 ;
  assign n18456 = n10766 | n18455 ;
  assign n18457 = n18456 ^ n1623 ^ 1'b0 ;
  assign n18454 = x220 & ~n3388 ;
  assign n18458 = n18457 ^ n18454 ^ 1'b0 ;
  assign n18459 = ~n6817 & n8694 ;
  assign n18460 = n6259 & ~n7964 ;
  assign n18461 = n18460 ^ n7266 ^ 1'b0 ;
  assign n18462 = n6166 | n18461 ;
  assign n18463 = x139 | n16775 ;
  assign n18464 = n4387 & n13343 ;
  assign n18465 = n18463 & n18464 ;
  assign n18466 = n4225 & ~n4805 ;
  assign n18467 = n1398 | n18466 ;
  assign n18468 = n1822 | n18467 ;
  assign n18469 = n1186 | n5067 ;
  assign n18470 = n8317 ^ n3911 ^ 1'b0 ;
  assign n18471 = ~n8658 & n18470 ;
  assign n18472 = ( ~n18468 & n18469 ) | ( ~n18468 & n18471 ) | ( n18469 & n18471 ) ;
  assign n18473 = n6315 ^ n3127 ^ 1'b0 ;
  assign n18474 = n6996 & n18473 ;
  assign n18475 = n13396 ^ n11226 ^ n1119 ;
  assign n18476 = n5559 ^ n3284 ^ 1'b0 ;
  assign n18477 = n18476 ^ n9270 ^ 1'b0 ;
  assign n18478 = n10998 ^ n1397 ^ 1'b0 ;
  assign n18479 = n16509 & ~n18478 ;
  assign n18480 = n3707 & ~n18479 ;
  assign n18481 = n18477 & n18480 ;
  assign n18482 = n9867 ^ n2472 ^ 1'b0 ;
  assign n18484 = n13540 ^ n5758 ^ 1'b0 ;
  assign n18485 = ~n8713 & n18484 ;
  assign n18483 = ~n2369 & n15924 ;
  assign n18486 = n18485 ^ n18483 ^ 1'b0 ;
  assign n18488 = n7804 & n8063 ;
  assign n18489 = n8226 & ~n18488 ;
  assign n18490 = ~n9186 & n18489 ;
  assign n18487 = n13666 & ~n16892 ;
  assign n18491 = n18490 ^ n18487 ^ 1'b0 ;
  assign n18492 = n7862 ^ n5667 ^ 1'b0 ;
  assign n18493 = n14749 & n18492 ;
  assign n18494 = n5238 & ~n13225 ;
  assign n18495 = n14239 & ~n18494 ;
  assign n18496 = n11174 ^ n1748 ^ 1'b0 ;
  assign n18497 = ~n9212 & n18496 ;
  assign n18498 = ~n16270 & n18497 ;
  assign n18499 = n18498 ^ n3255 ^ 1'b0 ;
  assign n18500 = n18499 ^ n1557 ^ 1'b0 ;
  assign n18501 = n1853 | n1937 ;
  assign n18502 = n4441 & ~n18501 ;
  assign n18503 = n18502 ^ n779 ^ 1'b0 ;
  assign n18504 = n11680 & n18503 ;
  assign n18505 = n2622 & n7822 ;
  assign n18506 = ~n1688 & n18505 ;
  assign n18507 = n18506 ^ n15422 ^ 1'b0 ;
  assign n18508 = n18507 ^ n2004 ^ 1'b0 ;
  assign n18509 = n18504 & n18508 ;
  assign n18510 = n6977 & n15106 ;
  assign n18511 = n6782 & n18510 ;
  assign n18513 = n6465 ^ n5287 ^ 1'b0 ;
  assign n18512 = n12476 | n15626 ;
  assign n18514 = n18513 ^ n18512 ^ 1'b0 ;
  assign n18515 = n17197 ^ n3223 ^ 1'b0 ;
  assign n18516 = n13385 & n17321 ;
  assign n18517 = ~n3962 & n18516 ;
  assign n18518 = n12263 | n18517 ;
  assign n18519 = n18518 ^ n11650 ^ 1'b0 ;
  assign n18520 = ~n16221 & n18519 ;
  assign n18521 = n8963 & ~n15319 ;
  assign n18524 = ~n825 & n1945 ;
  assign n18525 = n8033 & n18524 ;
  assign n18526 = n14322 ^ n5816 ^ 1'b0 ;
  assign n18527 = n18526 ^ n6347 ^ 1'b0 ;
  assign n18528 = n18525 | n18527 ;
  assign n18529 = n18528 ^ n17874 ^ n1672 ;
  assign n18522 = n1795 & n3494 ;
  assign n18523 = n18522 ^ n5671 ^ 1'b0 ;
  assign n18530 = n18529 ^ n18523 ^ n2192 ;
  assign n18531 = n16069 ^ n6140 ^ 1'b0 ;
  assign n18532 = n1547 & n18531 ;
  assign n18533 = ~n4310 & n18532 ;
  assign n18534 = n4730 & n5195 ;
  assign n18535 = ( n349 & ~n2243 ) | ( n349 & n8915 ) | ( ~n2243 & n8915 ) ;
  assign n18536 = n4509 | n13682 ;
  assign n18537 = n7061 & ~n16663 ;
  assign n18538 = n10053 & n18537 ;
  assign n18540 = n10134 ^ n920 ^ n774 ;
  assign n18541 = n4021 ^ n2211 ^ 1'b0 ;
  assign n18543 = n3012 | n3702 ;
  assign n18542 = n1645 & ~n4701 ;
  assign n18544 = n18543 ^ n18542 ^ 1'b0 ;
  assign n18545 = n10556 | n10622 ;
  assign n18546 = n18544 | n18545 ;
  assign n18547 = n18541 & n18546 ;
  assign n18548 = n18540 & n18547 ;
  assign n18549 = n1898 & ~n18548 ;
  assign n18539 = n8656 & n14777 ;
  assign n18550 = n18549 ^ n18539 ^ 1'b0 ;
  assign n18551 = n4399 | n9958 ;
  assign n18552 = n18551 ^ x61 ^ 1'b0 ;
  assign n18553 = n1317 | n1364 ;
  assign n18554 = n18553 ^ n10229 ^ 1'b0 ;
  assign n18555 = ~n5965 & n18554 ;
  assign n18556 = n1142 & n4677 ;
  assign n18557 = n18556 ^ n5089 ^ 1'b0 ;
  assign n18558 = n18557 ^ n5282 ^ 1'b0 ;
  assign n18568 = ( n671 & n2783 ) | ( n671 & ~n8322 ) | ( n2783 & ~n8322 ) ;
  assign n18569 = n18568 ^ n6331 ^ 1'b0 ;
  assign n18561 = n2986 ^ n1496 ^ 1'b0 ;
  assign n18562 = n5103 & n18561 ;
  assign n18563 = n2296 & n18562 ;
  assign n18564 = n3176 | n5252 ;
  assign n18565 = n1648 & ~n18564 ;
  assign n18566 = n18563 | n18565 ;
  assign n18567 = n18566 ^ n10698 ^ 1'b0 ;
  assign n18570 = n18569 ^ n18567 ^ 1'b0 ;
  assign n18571 = n466 | n18570 ;
  assign n18559 = ~n2520 & n10133 ;
  assign n18560 = n1220 & n18559 ;
  assign n18572 = n18571 ^ n18560 ^ 1'b0 ;
  assign n18573 = ~n2202 & n10077 ;
  assign n18574 = n18573 ^ n9407 ^ 1'b0 ;
  assign n18575 = n8865 & n11091 ;
  assign n18576 = ~n18574 & n18575 ;
  assign n18577 = n6177 & ~n9830 ;
  assign n18578 = n18577 ^ n1649 ^ 1'b0 ;
  assign n18579 = ~n1867 & n14918 ;
  assign n18580 = n18579 ^ n12361 ^ 1'b0 ;
  assign n18581 = n18580 ^ n2702 ^ 1'b0 ;
  assign n18582 = n18578 & n18581 ;
  assign n18583 = n988 | n15238 ;
  assign n18584 = n599 & ~n18583 ;
  assign n18586 = n18578 ^ n14867 ^ n3879 ;
  assign n18585 = ~n5225 & n8114 ;
  assign n18587 = n18586 ^ n18585 ^ 1'b0 ;
  assign n18588 = n8883 | n9889 ;
  assign n18589 = n1579 | n8352 ;
  assign n18590 = n18589 ^ n14456 ^ 1'b0 ;
  assign n18591 = n1664 | n18590 ;
  assign n18592 = n11601 & ~n18591 ;
  assign n18593 = n1980 & ~n6802 ;
  assign n18594 = n9377 & n18593 ;
  assign n18595 = ( ~n3541 & n10140 ) | ( ~n3541 & n18594 ) | ( n10140 & n18594 ) ;
  assign n18596 = ( n327 & ~n3518 ) | ( n327 & n16899 ) | ( ~n3518 & n16899 ) ;
  assign n18597 = n1147 | n2369 ;
  assign n18598 = n18597 ^ n13644 ^ 1'b0 ;
  assign n18599 = n18596 & n18598 ;
  assign n18600 = n7737 ^ n6200 ^ 1'b0 ;
  assign n18601 = ~n5642 & n18600 ;
  assign n18602 = ~n3152 & n18601 ;
  assign n18603 = n14825 & ~n18602 ;
  assign n18604 = ~n11710 & n18603 ;
  assign n18605 = n13537 & n17480 ;
  assign n18606 = n1147 & n18605 ;
  assign n18607 = n4888 & n15562 ;
  assign n18608 = n4242 & n18607 ;
  assign n18609 = n17962 | n18608 ;
  assign n18610 = n5402 | n18609 ;
  assign n18617 = n18443 ^ n8198 ^ 1'b0 ;
  assign n18618 = n7371 & ~n18617 ;
  assign n18619 = ~n756 & n18618 ;
  assign n18611 = ( n4295 & ~n7617 ) | ( n4295 & n9731 ) | ( ~n7617 & n9731 ) ;
  assign n18612 = ~n7675 & n18611 ;
  assign n18613 = ~n6964 & n18612 ;
  assign n18614 = n14774 ^ n14730 ^ 1'b0 ;
  assign n18615 = ~n5476 & n18614 ;
  assign n18616 = ~n18613 & n18615 ;
  assign n18620 = n18619 ^ n18616 ^ 1'b0 ;
  assign n18621 = ~n1766 & n6692 ;
  assign n18622 = ~n6692 & n18621 ;
  assign n18623 = ~n2983 & n3738 ;
  assign n18624 = n18622 & n18623 ;
  assign n18625 = n4757 | n18624 ;
  assign n18626 = n4757 & ~n18625 ;
  assign n18628 = x218 & ~n11274 ;
  assign n18627 = n6698 | n15120 ;
  assign n18629 = n18628 ^ n18627 ^ 1'b0 ;
  assign n18631 = ( n5786 & n6959 ) | ( n5786 & n9330 ) | ( n6959 & n9330 ) ;
  assign n18630 = n4944 | n13660 ;
  assign n18632 = n18631 ^ n18630 ^ 1'b0 ;
  assign n18633 = ~n12090 & n18632 ;
  assign n18634 = n14816 ^ n2204 ^ 1'b0 ;
  assign n18635 = n18633 & ~n18634 ;
  assign n18637 = ~n8671 & n18031 ;
  assign n18636 = n14937 ^ n6555 ^ 1'b0 ;
  assign n18638 = n18637 ^ n18636 ^ n7727 ;
  assign n18639 = ~x172 & n18468 ;
  assign n18640 = n18639 ^ n13573 ^ 1'b0 ;
  assign n18641 = n18640 ^ n7196 ^ 1'b0 ;
  assign n18642 = n15571 ^ n7947 ^ 1'b0 ;
  assign n18643 = ~n18641 & n18642 ;
  assign n18644 = x163 & n15046 ;
  assign n18645 = n18644 ^ n17240 ^ 1'b0 ;
  assign n18646 = n3217 & n12096 ;
  assign n18647 = n635 & n18646 ;
  assign n18648 = n18647 ^ n17392 ^ 1'b0 ;
  assign n18649 = n9773 | n18648 ;
  assign n18650 = n3515 ^ x113 ^ 1'b0 ;
  assign n18651 = n8581 & n18650 ;
  assign n18652 = ~n11955 & n18651 ;
  assign n18653 = n12163 ^ n3568 ^ 1'b0 ;
  assign n18654 = n18653 ^ n4938 ^ 1'b0 ;
  assign n18655 = ~n1516 & n18654 ;
  assign n18656 = n13718 & ~n18655 ;
  assign n18657 = n4519 & n8720 ;
  assign n18658 = n9607 & n18657 ;
  assign n18659 = ~n11906 & n15238 ;
  assign n18660 = n1490 | n2223 ;
  assign n18661 = ~n12100 & n18660 ;
  assign n18663 = n4038 ^ n897 ^ n310 ;
  assign n18662 = n7352 & ~n13110 ;
  assign n18664 = n18663 ^ n18662 ^ 1'b0 ;
  assign n18665 = n18664 ^ n6278 ^ 1'b0 ;
  assign n18666 = ~n18661 & n18665 ;
  assign n18667 = n18637 ^ n15979 ^ 1'b0 ;
  assign n18668 = n18645 & ~n18667 ;
  assign n18669 = ~n7929 & n8771 ;
  assign n18670 = ~n4173 & n18669 ;
  assign n18671 = n8110 | n9540 ;
  assign n18672 = n2681 & ~n6951 ;
  assign n18673 = n18672 ^ n13030 ^ n2518 ;
  assign n18674 = ~n4348 & n5983 ;
  assign n18675 = ( n13253 & n18673 ) | ( n13253 & n18674 ) | ( n18673 & n18674 ) ;
  assign n18676 = n3062 & n5746 ;
  assign n18677 = n18676 ^ n1211 ^ 1'b0 ;
  assign n18678 = x163 | n547 ;
  assign n18679 = n18678 ^ n1848 ^ 1'b0 ;
  assign n18680 = n13045 | n18679 ;
  assign n18681 = n10612 ^ n3686 ^ 1'b0 ;
  assign n18682 = n17389 & ~n18681 ;
  assign n18683 = n16885 ^ n9062 ^ 1'b0 ;
  assign n18684 = n15595 & ~n18683 ;
  assign n18685 = n12719 ^ n10928 ^ 1'b0 ;
  assign n18686 = n18684 & ~n18685 ;
  assign n18687 = ~n2799 & n6222 ;
  assign n18688 = ~n18686 & n18687 ;
  assign n18696 = n7232 ^ n5213 ^ 1'b0 ;
  assign n18692 = n4415 | n16575 ;
  assign n18693 = n18692 ^ n2148 ^ 1'b0 ;
  assign n18689 = n16928 ^ n1220 ^ 1'b0 ;
  assign n18690 = n724 & ~n18689 ;
  assign n18691 = n18310 & n18690 ;
  assign n18694 = n18693 ^ n18691 ^ 1'b0 ;
  assign n18695 = n1645 & ~n18694 ;
  assign n18697 = n18696 ^ n18695 ^ 1'b0 ;
  assign n18698 = n11341 & ~n18697 ;
  assign n18699 = x137 & ~n10580 ;
  assign n18700 = ~n6959 & n18699 ;
  assign n18701 = n18700 ^ n5270 ^ 1'b0 ;
  assign n18702 = ( n3873 & n13644 ) | ( n3873 & ~n18701 ) | ( n13644 & ~n18701 ) ;
  assign n18703 = n15941 ^ n10039 ^ n3159 ;
  assign n18704 = n14354 & ~n18703 ;
  assign n18705 = n3198 | n6411 ;
  assign n18706 = n287 & n18705 ;
  assign n18707 = n18706 ^ n3286 ^ 1'b0 ;
  assign n18708 = n18707 ^ n1154 ^ 1'b0 ;
  assign n18709 = n17733 ^ n4619 ^ 1'b0 ;
  assign n18710 = n18708 | n18709 ;
  assign n18711 = n4988 | n18710 ;
  assign n18712 = n18711 ^ n2369 ^ 1'b0 ;
  assign n18713 = n4230 | n6628 ;
  assign n18714 = n16594 ^ n15983 ^ 1'b0 ;
  assign n18715 = ~n18713 & n18714 ;
  assign n18716 = n5571 ^ n2445 ^ 1'b0 ;
  assign n18717 = n11272 & ~n18716 ;
  assign n18718 = n5115 & n18717 ;
  assign n18719 = n4721 & n18718 ;
  assign n18720 = n18719 ^ n12275 ^ 1'b0 ;
  assign n18721 = n16795 & ~n17340 ;
  assign n18722 = n18721 ^ n18619 ^ 1'b0 ;
  assign n18724 = ~x249 & n7723 ;
  assign n18725 = n18724 ^ n4405 ^ 1'b0 ;
  assign n18726 = n2557 & n18725 ;
  assign n18723 = n2675 & ~n9809 ;
  assign n18727 = n18726 ^ n18723 ^ n18692 ;
  assign n18728 = n5831 & ~n13276 ;
  assign n18729 = ~n5118 & n18728 ;
  assign n18730 = ~n11899 & n18729 ;
  assign n18731 = n9489 ^ n3147 ^ 1'b0 ;
  assign n18732 = n3309 & ~n12597 ;
  assign n18733 = n6826 ^ n634 ^ 1'b0 ;
  assign n18734 = n11053 & ~n18733 ;
  assign n18735 = n18732 & ~n18734 ;
  assign n18736 = n11710 ^ n2959 ^ 1'b0 ;
  assign n18737 = ~n4266 & n18736 ;
  assign n18738 = ~n11129 & n16879 ;
  assign n18739 = n14634 ^ n11475 ^ 1'b0 ;
  assign n18740 = n11061 & ~n11939 ;
  assign n18741 = n2903 ^ n1583 ^ 1'b0 ;
  assign n18742 = n688 | n8117 ;
  assign n18743 = n18742 ^ n5173 ^ 1'b0 ;
  assign n18744 = n18741 & ~n18743 ;
  assign n18745 = n780 | n2765 ;
  assign n18746 = n1828 | n18745 ;
  assign n18747 = n11321 | n18746 ;
  assign n18748 = ~n6654 & n7022 ;
  assign n18749 = n18748 ^ n1866 ^ 1'b0 ;
  assign n18750 = n4752 & ~n18749 ;
  assign n18751 = ~n4673 & n17482 ;
  assign n18752 = n6352 & ~n12101 ;
  assign n18753 = n6006 & n18752 ;
  assign n18754 = ( n8585 & n9938 ) | ( n8585 & n18753 ) | ( n9938 & n18753 ) ;
  assign n18755 = ~n13871 & n18754 ;
  assign n18756 = n18755 ^ n15820 ^ 1'b0 ;
  assign n18757 = n1146 ^ x162 ^ 1'b0 ;
  assign n18762 = n9853 & n10831 ;
  assign n18758 = ( x60 & n1620 ) | ( x60 & ~n13202 ) | ( n1620 & ~n13202 ) ;
  assign n18759 = n10398 & n18758 ;
  assign n18760 = n3551 & ~n15010 ;
  assign n18761 = ~n18759 & n18760 ;
  assign n18763 = n18762 ^ n18761 ^ n16851 ;
  assign n18764 = n4470 & ~n16565 ;
  assign n18765 = n5313 ^ n611 ^ 1'b0 ;
  assign n18766 = n18764 & ~n18765 ;
  assign n18767 = n5878 | n8256 ;
  assign n18768 = n5254 | n18767 ;
  assign n18769 = n18768 ^ n4708 ^ 1'b0 ;
  assign n18770 = n18766 & n18769 ;
  assign n18771 = ~n367 & n3464 ;
  assign n18772 = n18771 ^ n13631 ^ 1'b0 ;
  assign n18773 = n7877 & ~n18772 ;
  assign n18774 = n9227 ^ n8225 ^ n7869 ;
  assign n18775 = n8705 & ~n18774 ;
  assign n18776 = n2317 & n5148 ;
  assign n18777 = n18776 ^ n6268 ^ 1'b0 ;
  assign n18778 = n11633 & ~n18777 ;
  assign n18779 = n18775 & n18778 ;
  assign n18780 = n1643 & ~n18779 ;
  assign n18781 = n1079 & n18780 ;
  assign n18782 = ~n2634 & n9664 ;
  assign n18783 = n14760 ^ n5673 ^ 1'b0 ;
  assign n18784 = n14124 | n17437 ;
  assign n18785 = n18784 ^ x180 ^ 1'b0 ;
  assign n18786 = n8071 ^ n1439 ^ 1'b0 ;
  assign n18787 = n18786 ^ n8561 ^ 1'b0 ;
  assign n18788 = ~n12047 & n18787 ;
  assign n18789 = n14521 & n18788 ;
  assign n18790 = n5616 & n7101 ;
  assign n18791 = n18790 ^ n17229 ^ 1'b0 ;
  assign n18792 = n2569 | n18791 ;
  assign n18793 = ~x154 & n7300 ;
  assign n18794 = n4208 | n18793 ;
  assign n18795 = n18794 ^ n5481 ^ 1'b0 ;
  assign n18796 = n15759 & n18795 ;
  assign n18797 = n4119 | n18147 ;
  assign n18798 = n18797 ^ n389 ^ 1'b0 ;
  assign n18799 = n10070 & ~n10377 ;
  assign n18800 = n18799 ^ n13444 ^ 1'b0 ;
  assign n18801 = n16181 ^ n12112 ^ 1'b0 ;
  assign n18802 = ( n1589 & ~n10761 ) | ( n1589 & n12714 ) | ( ~n10761 & n12714 ) ;
  assign n18803 = n8574 & ~n18802 ;
  assign n18804 = ~n4867 & n18803 ;
  assign n18805 = n643 | n1784 ;
  assign n18806 = ~n7541 & n7797 ;
  assign n18807 = n18806 ^ n16305 ^ 1'b0 ;
  assign n18808 = n6020 & n10397 ;
  assign n18809 = n10342 ^ n6171 ^ 1'b0 ;
  assign n18810 = ~n9454 & n18809 ;
  assign n18811 = n3584 ^ n3151 ^ 1'b0 ;
  assign n18812 = n12870 & ~n18811 ;
  assign n18813 = n1416 & n18812 ;
  assign n18814 = ~n4563 & n9316 ;
  assign n18815 = n18814 ^ n3302 ^ 1'b0 ;
  assign n18816 = n6332 ^ n3342 ^ 1'b0 ;
  assign n18817 = n1589 & ~n1619 ;
  assign n18818 = n11697 ^ n1513 ^ 1'b0 ;
  assign n18819 = x203 & n18818 ;
  assign n18821 = ( n3915 & n4292 ) | ( n3915 & ~n4460 ) | ( n4292 & ~n4460 ) ;
  assign n18820 = n1726 & n2615 ;
  assign n18822 = n18821 ^ n18820 ^ 1'b0 ;
  assign n18823 = n2316 & n18822 ;
  assign n18824 = n4169 & n18823 ;
  assign n18825 = n4027 ^ n3734 ^ 1'b0 ;
  assign n18826 = n1458 & ~n18825 ;
  assign n18827 = n8408 ^ n4325 ^ 1'b0 ;
  assign n18828 = n5980 | n18827 ;
  assign n18829 = n10502 & ~n18828 ;
  assign n18830 = ( n2150 & n18826 ) | ( n2150 & n18829 ) | ( n18826 & n18829 ) ;
  assign n18831 = n3412 & n5961 ;
  assign n18832 = n18831 ^ n16399 ^ 1'b0 ;
  assign n18835 = n14754 ^ n3317 ^ 1'b0 ;
  assign n18836 = n15768 & ~n18835 ;
  assign n18837 = n13511 & ~n18836 ;
  assign n18833 = n2130 & n11765 ;
  assign n18834 = n15777 & n18833 ;
  assign n18838 = n18837 ^ n18834 ^ 1'b0 ;
  assign n18839 = ~n18237 & n18838 ;
  assign n18840 = ~n3761 & n9751 ;
  assign n18841 = ~n2479 & n18840 ;
  assign n18842 = n18841 ^ n4645 ^ 1'b0 ;
  assign n18843 = n2453 & n18842 ;
  assign n18844 = n18843 ^ n876 ^ 1'b0 ;
  assign n18845 = n18844 ^ n12502 ^ 1'b0 ;
  assign n18846 = ~n4400 & n18845 ;
  assign n18847 = n5335 & n8529 ;
  assign n18848 = ( n6019 & n11410 ) | ( n6019 & ~n12669 ) | ( n11410 & ~n12669 ) ;
  assign n18849 = n14987 ^ n13584 ^ 1'b0 ;
  assign n18850 = n13390 & n18849 ;
  assign n18851 = n14354 & ~n18850 ;
  assign n18852 = n18851 ^ n10731 ^ 1'b0 ;
  assign n18853 = n18852 ^ n6180 ^ 1'b0 ;
  assign n18854 = n7964 | n18853 ;
  assign n18855 = n8891 & n10750 ;
  assign n18856 = ~n9465 & n18855 ;
  assign n18857 = n18856 ^ n14619 ^ n6412 ;
  assign n18858 = n18857 ^ n1981 ^ 1'b0 ;
  assign n18859 = n9009 ^ n2286 ^ 1'b0 ;
  assign n18863 = n18029 ^ n4845 ^ 1'b0 ;
  assign n18864 = n8119 & ~n18863 ;
  assign n18860 = n8112 | n9181 ;
  assign n18861 = n8632 | n18860 ;
  assign n18862 = n13493 & ~n18861 ;
  assign n18865 = n18864 ^ n18862 ^ 1'b0 ;
  assign n18866 = ~n3543 & n5966 ;
  assign n18867 = n11291 ^ n8121 ^ 1'b0 ;
  assign n18868 = n18867 ^ n5118 ^ n3980 ;
  assign n18869 = n17684 & n18868 ;
  assign n18870 = n5538 ^ x163 ^ 1'b0 ;
  assign n18871 = n3039 | n18870 ;
  assign n18872 = n14215 ^ n825 ^ 1'b0 ;
  assign n18873 = ~n5749 & n18872 ;
  assign n18874 = ~n7741 & n8544 ;
  assign n18875 = n3563 & n18874 ;
  assign n18876 = n7501 & n18875 ;
  assign n18877 = n4662 ^ n4343 ^ 1'b0 ;
  assign n18878 = n3913 & ~n4360 ;
  assign n18879 = n18878 ^ n14341 ^ 1'b0 ;
  assign n18880 = n11121 & n17868 ;
  assign n18881 = n9897 | n18880 ;
  assign n18882 = n18881 ^ n13629 ^ 1'b0 ;
  assign n18883 = n14757 ^ n10158 ^ 1'b0 ;
  assign n18884 = ~n16282 & n18883 ;
  assign n18885 = n2870 & ~n10612 ;
  assign n18886 = n18885 ^ n378 ^ 1'b0 ;
  assign n18887 = n3628 | n7112 ;
  assign n18888 = n13859 ^ n4553 ^ n3670 ;
  assign n18889 = n3059 ^ n370 ^ 1'b0 ;
  assign n18890 = n18889 ^ n18819 ^ 1'b0 ;
  assign n18891 = ~n1778 & n18890 ;
  assign n18892 = n1820 & ~n3539 ;
  assign n18893 = n4875 | n8502 ;
  assign n18894 = n16217 & ~n18893 ;
  assign n18895 = ~n18892 & n18894 ;
  assign n18896 = ~n10318 & n13666 ;
  assign n18897 = ~n16545 & n18896 ;
  assign n18898 = n18897 ^ n1465 ^ 1'b0 ;
  assign n18899 = n4397 & n8783 ;
  assign n18900 = n9012 & n16487 ;
  assign n18901 = n18900 ^ n15596 ^ 1'b0 ;
  assign n18902 = n18899 & n18901 ;
  assign n18903 = n14603 ^ n7742 ^ 1'b0 ;
  assign n18904 = n4946 | n18903 ;
  assign n18905 = n18904 ^ n8246 ^ n7513 ;
  assign n18906 = n6907 ^ n6155 ^ 1'b0 ;
  assign n18907 = n18906 ^ n4567 ^ 1'b0 ;
  assign n18908 = n18905 | n18907 ;
  assign n18909 = n1639 | n11146 ;
  assign n18910 = n725 | n875 ;
  assign n18911 = ~n11108 & n18910 ;
  assign n18912 = n15137 ^ n8584 ^ 1'b0 ;
  assign n18913 = ~n18911 & n18912 ;
  assign n18916 = n2507 ^ n1935 ^ 1'b0 ;
  assign n18917 = n8782 & n18916 ;
  assign n18914 = n11627 ^ n9684 ^ 1'b0 ;
  assign n18915 = n11818 | n18914 ;
  assign n18918 = n18917 ^ n18915 ^ 1'b0 ;
  assign n18919 = ( n2559 & n10176 ) | ( n2559 & ~n11908 ) | ( n10176 & ~n11908 ) ;
  assign n18920 = ~n14867 & n18919 ;
  assign n18921 = n13678 & n18920 ;
  assign n18922 = n15282 ^ n9053 ^ 1'b0 ;
  assign n18923 = n6057 & n18922 ;
  assign n18924 = n858 & n18923 ;
  assign n18925 = x2 & n1242 ;
  assign n18926 = n18924 & n18925 ;
  assign n18927 = n18926 ^ n16236 ^ 1'b0 ;
  assign n18928 = ~n5646 & n14825 ;
  assign n18929 = n2306 | n10129 ;
  assign n18930 = n18928 & ~n18929 ;
  assign n18931 = n17231 ^ n13697 ^ 1'b0 ;
  assign n18932 = n1025 & n18931 ;
  assign n18933 = n7557 ^ n7452 ^ 1'b0 ;
  assign n18934 = n5206 & n18933 ;
  assign n18935 = ~n5139 & n6851 ;
  assign n18936 = n6966 | n18935 ;
  assign n18937 = ~n389 & n3766 ;
  assign n18938 = ~n8715 & n18937 ;
  assign n18939 = ~n18936 & n18938 ;
  assign n18940 = n11809 ^ n5585 ^ 1'b0 ;
  assign n18941 = n11065 & n18940 ;
  assign n18943 = n10940 & ~n15631 ;
  assign n18942 = n15779 & n16815 ;
  assign n18944 = n18943 ^ n18942 ^ 1'b0 ;
  assign n18945 = ~n293 & n1926 ;
  assign n18946 = ~n8592 & n18945 ;
  assign n18947 = n18946 ^ n7242 ^ 1'b0 ;
  assign n18948 = n991 & n18947 ;
  assign n18949 = n18948 ^ n17149 ^ n7122 ;
  assign n18950 = n18949 ^ n1752 ^ 1'b0 ;
  assign n18951 = n13757 ^ n12876 ^ 1'b0 ;
  assign n18952 = n13065 & n18951 ;
  assign n18953 = n10284 ^ n9206 ^ n5055 ;
  assign n18954 = n18953 ^ n12447 ^ 1'b0 ;
  assign n18955 = n3699 & ~n4003 ;
  assign n18956 = n10169 & ~n18955 ;
  assign n18957 = x169 & n18956 ;
  assign n18958 = n12930 ^ n2382 ^ 1'b0 ;
  assign n18959 = n13766 & n18958 ;
  assign n18960 = n17929 & n18959 ;
  assign n18961 = n18960 ^ n9022 ^ 1'b0 ;
  assign n18962 = n5134 & ~n6415 ;
  assign n18963 = n7710 & ~n18436 ;
  assign n18964 = n18963 ^ n10449 ^ 1'b0 ;
  assign n18965 = n3308 & ~n7252 ;
  assign n18966 = n12694 & n18965 ;
  assign n18967 = ( n673 & ~n4031 ) | ( n673 & n14364 ) | ( ~n4031 & n14364 ) ;
  assign n18968 = n12811 ^ n9343 ^ 1'b0 ;
  assign n18969 = n18967 & n18968 ;
  assign n18970 = ( ~n1081 & n9595 ) | ( ~n1081 & n10172 ) | ( n9595 & n10172 ) ;
  assign n18971 = ( n8241 & n12514 ) | ( n8241 & ~n13657 ) | ( n12514 & ~n13657 ) ;
  assign n18972 = n11885 ^ n3699 ^ 1'b0 ;
  assign n18973 = n12009 ^ n10430 ^ 1'b0 ;
  assign n18974 = n18972 & n18973 ;
  assign n18975 = n3634 ^ n1402 ^ 1'b0 ;
  assign n18976 = n6307 & ~n18975 ;
  assign n18977 = n13917 ^ n5323 ^ 1'b0 ;
  assign n18978 = n7061 & ~n18977 ;
  assign n18979 = x214 & x249 ;
  assign n18980 = ~x249 & n18979 ;
  assign n18981 = n12406 | n18980 ;
  assign n18982 = n12406 & ~n18981 ;
  assign n18983 = ~n771 & n4033 ;
  assign n18984 = n771 & n18983 ;
  assign n18985 = ~n11477 & n18984 ;
  assign n18986 = n2593 & n4327 ;
  assign n18987 = ~n4327 & n18986 ;
  assign n18988 = n3887 & ~n18987 ;
  assign n18989 = n3323 & n4603 ;
  assign n18990 = ~n4603 & n18989 ;
  assign n18991 = n18988 & ~n18990 ;
  assign n18992 = n18985 & n18991 ;
  assign n18993 = n18992 ^ n9747 ^ 1'b0 ;
  assign n18994 = n9226 & n18993 ;
  assign n18995 = n18982 & n18994 ;
  assign n18996 = ~n455 & n1129 ;
  assign n18997 = n455 & n18996 ;
  assign n18998 = ~n2131 & n18997 ;
  assign n18999 = ~n18995 & n18998 ;
  assign n19000 = n18995 & n18999 ;
  assign n19001 = n2329 | n19000 ;
  assign n19002 = ( n18976 & ~n18978 ) | ( n18976 & n19001 ) | ( ~n18978 & n19001 ) ;
  assign n19003 = n4619 & n14516 ;
  assign n19005 = n4113 ^ x229 ^ 1'b0 ;
  assign n19004 = n707 & ~n15738 ;
  assign n19006 = n19005 ^ n19004 ^ 1'b0 ;
  assign n19007 = ( ~n4899 & n19003 ) | ( ~n4899 & n19006 ) | ( n19003 & n19006 ) ;
  assign n19008 = n446 & n995 ;
  assign n19009 = n11522 ^ n1649 ^ 1'b0 ;
  assign n19010 = n19009 ^ n7719 ^ 1'b0 ;
  assign n19011 = n12095 ^ n1477 ^ 1'b0 ;
  assign n19012 = n6540 ^ n2934 ^ 1'b0 ;
  assign n19013 = n2881 ^ x45 ^ 1'b0 ;
  assign n19014 = n3335 | n4845 ;
  assign n19016 = n7384 | n12987 ;
  assign n19015 = x192 & ~n11776 ;
  assign n19017 = n19016 ^ n19015 ^ 1'b0 ;
  assign n19018 = ( n7263 & n13451 ) | ( n7263 & ~n13644 ) | ( n13451 & ~n13644 ) ;
  assign n19019 = n3823 & n6811 ;
  assign n19020 = n16932 ^ n688 ^ 1'b0 ;
  assign n19021 = ~n19019 & n19020 ;
  assign n19022 = n3304 | n12203 ;
  assign n19023 = n5300 & ~n19022 ;
  assign n19024 = ~n18578 & n19023 ;
  assign n19025 = ~n2904 & n7871 ;
  assign n19026 = n19025 ^ n6872 ^ 1'b0 ;
  assign n19027 = n19026 ^ n1322 ^ 1'b0 ;
  assign n19028 = ~n11229 & n19027 ;
  assign n19029 = n3431 & n15893 ;
  assign n19030 = n19029 ^ n3429 ^ 1'b0 ;
  assign n19031 = ( n1606 & ~n1689 ) | ( n1606 & n19030 ) | ( ~n1689 & n19030 ) ;
  assign n19032 = n4108 ^ x165 ^ 1'b0 ;
  assign n19033 = n1073 | n19032 ;
  assign n19034 = n9476 | n19033 ;
  assign n19035 = n9070 & n19034 ;
  assign n19036 = ~n4436 & n4657 ;
  assign n19038 = ~n6680 & n10075 ;
  assign n19037 = n675 | n774 ;
  assign n19039 = n19038 ^ n19037 ^ 1'b0 ;
  assign n19040 = n19036 & n19039 ;
  assign n19041 = n13796 ^ n4784 ^ 1'b0 ;
  assign n19042 = ~n5408 & n5708 ;
  assign n19043 = n5729 ^ x22 ^ 1'b0 ;
  assign n19044 = n11517 ^ n7555 ^ 1'b0 ;
  assign n19045 = ~n11229 & n19044 ;
  assign n19046 = n19045 ^ x252 ^ 1'b0 ;
  assign n19047 = n19046 ^ x40 ^ 1'b0 ;
  assign n19048 = n16198 & n19047 ;
  assign n19049 = ~n19043 & n19048 ;
  assign n19050 = n17573 ^ n8851 ^ 1'b0 ;
  assign n19051 = n7147 ^ n6235 ^ 1'b0 ;
  assign n19052 = ~n8694 & n19051 ;
  assign n19053 = ~n9239 & n17875 ;
  assign n19054 = n19053 ^ n9714 ^ 1'b0 ;
  assign n19055 = n3275 | n5266 ;
  assign n19056 = n19055 ^ n14861 ^ 1'b0 ;
  assign n19057 = n2771 | n19056 ;
  assign n19058 = n11033 ^ n908 ^ 1'b0 ;
  assign n19059 = n6502 | n19058 ;
  assign n19060 = n14007 & ~n19059 ;
  assign n19061 = n19060 ^ n11597 ^ 1'b0 ;
  assign n19062 = ~n9452 & n13944 ;
  assign n19063 = ~n12136 & n19062 ;
  assign n19064 = n19063 ^ n11138 ^ 1'b0 ;
  assign n19065 = n4931 & ~n19064 ;
  assign n19066 = ~n4723 & n5227 ;
  assign n19067 = n19066 ^ n2701 ^ 1'b0 ;
  assign n19068 = n1367 & ~n19067 ;
  assign n19069 = x46 & n2102 ;
  assign n19070 = n19068 & n19069 ;
  assign n19071 = n7109 & n19070 ;
  assign n19072 = ~n7266 & n7836 ;
  assign n19073 = n19072 ^ n18949 ^ 1'b0 ;
  assign n19074 = n10279 & ~n11406 ;
  assign n19075 = n7964 | n14526 ;
  assign n19076 = n4333 ^ n1220 ^ 1'b0 ;
  assign n19077 = n19075 & n19076 ;
  assign n19078 = n11127 & ~n15279 ;
  assign n19079 = n9823 ^ n6098 ^ 1'b0 ;
  assign n19080 = n12225 & ~n19079 ;
  assign n19081 = n483 & n7238 ;
  assign n19082 = n10051 & n19081 ;
  assign n19083 = n10416 | n19082 ;
  assign n19084 = ( ~n2144 & n3114 ) | ( ~n2144 & n10129 ) | ( n3114 & n10129 ) ;
  assign n19085 = ( n16256 & n19083 ) | ( n16256 & ~n19084 ) | ( n19083 & ~n19084 ) ;
  assign n19086 = x226 & n3560 ;
  assign n19087 = n13497 ^ n997 ^ 1'b0 ;
  assign n19088 = n3046 & n4938 ;
  assign n19089 = n19088 ^ n4910 ^ 1'b0 ;
  assign n19090 = n19089 ^ n18734 ^ n8139 ;
  assign n19091 = n2215 ^ n1123 ^ 1'b0 ;
  assign n19092 = n5387 | n19091 ;
  assign n19093 = n10872 | n19092 ;
  assign n19094 = n4130 | n6017 ;
  assign n19095 = n1154 & ~n19094 ;
  assign n19096 = n5594 & ~n19037 ;
  assign n19097 = n12828 ^ n3557 ^ 1'b0 ;
  assign n19098 = n17859 | n19097 ;
  assign n19099 = n4139 ^ n1377 ^ 1'b0 ;
  assign n19100 = n17883 & ~n19099 ;
  assign n19101 = n18042 & n19100 ;
  assign n19102 = n19101 ^ x178 ^ 1'b0 ;
  assign n19103 = n2911 ^ x122 ^ 1'b0 ;
  assign n19104 = ~n7657 & n19103 ;
  assign n19105 = n8793 & n19104 ;
  assign n19106 = n19102 & n19105 ;
  assign n19107 = ( n2301 & ~n19098 ) | ( n2301 & n19106 ) | ( ~n19098 & n19106 ) ;
  assign n19108 = n15193 & n19107 ;
  assign n19109 = n10950 ^ n3565 ^ 1'b0 ;
  assign n19110 = n1900 | n11863 ;
  assign n19111 = x49 & ~n19068 ;
  assign n19112 = n10655 ^ n8645 ^ 1'b0 ;
  assign n19113 = ~n12592 & n19112 ;
  assign n19114 = n19113 ^ n7107 ^ 1'b0 ;
  assign n19115 = x167 & n19114 ;
  assign n19116 = ~n3765 & n9477 ;
  assign n19117 = ~n1742 & n19116 ;
  assign n19118 = n6546 & n7045 ;
  assign n19119 = ~n6546 & n19118 ;
  assign n19120 = ~n2514 & n5682 ;
  assign n19121 = n11109 ^ n8388 ^ n7340 ;
  assign n19122 = n11151 ^ n3349 ^ n1588 ;
  assign n19123 = n16622 ^ n13504 ^ 1'b0 ;
  assign n19124 = n6982 ^ n6827 ^ 1'b0 ;
  assign n19125 = n19124 ^ n11362 ^ 1'b0 ;
  assign n19126 = n5651 & ~n19125 ;
  assign n19127 = n7660 ^ n3007 ^ 1'b0 ;
  assign n19128 = n882 | n19127 ;
  assign n19129 = ( n3868 & n14580 ) | ( n3868 & ~n19128 ) | ( n14580 & ~n19128 ) ;
  assign n19130 = n12138 | n19129 ;
  assign n19131 = n4148 & ~n13142 ;
  assign n19132 = n18466 ^ n12811 ^ 1'b0 ;
  assign n19133 = n11460 | n19132 ;
  assign n19134 = ~n4864 & n14131 ;
  assign n19135 = n4539 | n19134 ;
  assign n19136 = n13070 ^ n11006 ^ 1'b0 ;
  assign n19137 = n15837 ^ n3876 ^ 1'b0 ;
  assign n19138 = n1367 & ~n19137 ;
  assign n19139 = ( ~n6898 & n18812 ) | ( ~n6898 & n19138 ) | ( n18812 & n19138 ) ;
  assign n19140 = ~n1016 & n19139 ;
  assign n19141 = n1016 & n19140 ;
  assign n19142 = n10390 ^ n5734 ^ 1'b0 ;
  assign n19143 = n11684 & n14436 ;
  assign n19144 = n9031 ^ n4380 ^ x106 ;
  assign n19145 = n5614 & n19144 ;
  assign n19146 = n19145 ^ n18723 ^ 1'b0 ;
  assign n19147 = n13305 & n19146 ;
  assign n19148 = n10984 | n19147 ;
  assign n19149 = n14369 ^ n8155 ^ 1'b0 ;
  assign n19150 = n854 & ~n19149 ;
  assign n19151 = n2778 ^ n1109 ^ 1'b0 ;
  assign n19152 = ~n14964 & n19151 ;
  assign n19153 = n19152 ^ n8243 ^ 1'b0 ;
  assign n19154 = ~n4169 & n15181 ;
  assign n19155 = n2560 | n3329 ;
  assign n19157 = n2387 ^ n917 ^ 1'b0 ;
  assign n19158 = n19157 ^ n6508 ^ 1'b0 ;
  assign n19156 = n3202 & n3939 ;
  assign n19159 = n19158 ^ n19156 ^ 1'b0 ;
  assign n19160 = n17552 & ~n19159 ;
  assign n19161 = n8976 & n10405 ;
  assign n19162 = n19161 ^ x96 ^ 1'b0 ;
  assign n19163 = n3174 & n19162 ;
  assign n19164 = n19163 ^ n4914 ^ 1'b0 ;
  assign n19165 = n5522 ^ n3515 ^ 1'b0 ;
  assign n19166 = n11040 ^ n4976 ^ 1'b0 ;
  assign n19167 = n2912 | n19166 ;
  assign n19168 = n10515 | n10878 ;
  assign n19169 = n19168 ^ n2456 ^ 1'b0 ;
  assign n19170 = n8535 ^ n1278 ^ n579 ;
  assign n19171 = n14679 ^ n7193 ^ 1'b0 ;
  assign n19172 = n9525 ^ n4679 ^ 1'b0 ;
  assign n19173 = n14391 & ~n19172 ;
  assign n19174 = n6304 | n7378 ;
  assign n19175 = n8130 ^ n3326 ^ 1'b0 ;
  assign n19176 = n9046 | n19175 ;
  assign n19177 = n19174 & ~n19176 ;
  assign n19178 = n15578 ^ n11204 ^ n6872 ;
  assign n19179 = n8698 & ~n13335 ;
  assign n19180 = n7373 & n10801 ;
  assign n19181 = n19180 ^ n1315 ^ 1'b0 ;
  assign n19182 = n5101 & ~n10049 ;
  assign n19183 = n5333 ^ n3044 ^ 1'b0 ;
  assign n19184 = n3882 | n9365 ;
  assign n19185 = n16651 | n19184 ;
  assign n19186 = n3474 | n15971 ;
  assign n19187 = n19186 ^ n14838 ^ 1'b0 ;
  assign n19188 = n17382 & n19187 ;
  assign n19189 = n19188 ^ n13737 ^ n1530 ;
  assign n19190 = n2343 | n15555 ;
  assign n19191 = n3266 & ~n19190 ;
  assign n19192 = n4369 ^ n2670 ^ 1'b0 ;
  assign n19193 = n19192 ^ n2579 ^ 1'b0 ;
  assign n19194 = x229 & n3757 ;
  assign n19195 = n19194 ^ n5490 ^ 1'b0 ;
  assign n19196 = n19195 ^ x132 ^ 1'b0 ;
  assign n19197 = ~n10299 & n18279 ;
  assign n19198 = ~n6662 & n14949 ;
  assign n19199 = n11435 ^ n5311 ^ 1'b0 ;
  assign n19200 = ( n703 & ~n1682 ) | ( n703 & n2566 ) | ( ~n1682 & n2566 ) ;
  assign n19201 = ~n9627 & n19200 ;
  assign n19202 = n920 & ~n19201 ;
  assign n19203 = n3853 & n19202 ;
  assign n19204 = n19199 & n19203 ;
  assign n19206 = n14225 ^ n2020 ^ 1'b0 ;
  assign n19207 = n5779 & n19206 ;
  assign n19205 = n8895 & ~n16662 ;
  assign n19208 = n19207 ^ n19205 ^ 1'b0 ;
  assign n19209 = ( x72 & n3371 ) | ( x72 & ~n14733 ) | ( n3371 & ~n14733 ) ;
  assign n19210 = n4567 & n4572 ;
  assign n19211 = n19210 ^ n7204 ^ n2622 ;
  assign n19212 = n19211 ^ n10700 ^ 1'b0 ;
  assign n19213 = n10596 & ~n19212 ;
  assign n19214 = ~n15785 & n19213 ;
  assign n19215 = ~n1565 & n19214 ;
  assign n19216 = n4970 & ~n19215 ;
  assign n19217 = n19216 ^ n2029 ^ 1'b0 ;
  assign n19218 = n16307 ^ n8916 ^ 1'b0 ;
  assign n19219 = n19218 ^ n18292 ^ 1'b0 ;
  assign n19221 = ~n9287 & n12670 ;
  assign n19222 = n19221 ^ n15745 ^ 1'b0 ;
  assign n19220 = ~n6818 & n9814 ;
  assign n19223 = n19222 ^ n19220 ^ 1'b0 ;
  assign n19224 = n9609 ^ n6587 ^ n1884 ;
  assign n19225 = ( n6359 & n11862 ) | ( n6359 & n19224 ) | ( n11862 & n19224 ) ;
  assign n19226 = n10189 ^ n2112 ^ 1'b0 ;
  assign n19227 = ~n2951 & n19226 ;
  assign n19228 = n12773 ^ n4072 ^ 1'b0 ;
  assign n19229 = ~x124 & n628 ;
  assign n19230 = n19229 ^ n8155 ^ n7593 ;
  assign n19231 = n19230 ^ n8568 ^ 1'b0 ;
  assign n19232 = n1500 & ~n19231 ;
  assign n19233 = n2338 | n19232 ;
  assign n19234 = n7736 ^ n4212 ^ 1'b0 ;
  assign n19235 = ~n11251 & n19234 ;
  assign n19236 = n19235 ^ n17524 ^ 1'b0 ;
  assign n19239 = n3213 | n3582 ;
  assign n19240 = n19239 ^ n4139 ^ 1'b0 ;
  assign n19241 = n19240 ^ n6207 ^ 1'b0 ;
  assign n19237 = ~n9766 & n12464 ;
  assign n19238 = n1517 & n19237 ;
  assign n19242 = n19241 ^ n19238 ^ 1'b0 ;
  assign n19243 = n2611 | n7629 ;
  assign n19244 = n19243 ^ n2735 ^ 1'b0 ;
  assign n19245 = n1633 & ~n16603 ;
  assign n19246 = n836 & n2170 ;
  assign n19247 = n10506 ^ n9194 ^ 1'b0 ;
  assign n19248 = n19247 ^ n9961 ^ 1'b0 ;
  assign n19249 = n10814 ^ n4621 ^ 1'b0 ;
  assign n19250 = ~n4185 & n19249 ;
  assign n19251 = n13549 & n19250 ;
  assign n19252 = n19251 ^ n17609 ^ 1'b0 ;
  assign n19253 = n2934 | n5456 ;
  assign n19254 = ~n4610 & n12571 ;
  assign n19255 = n6854 ^ n3377 ^ 1'b0 ;
  assign n19256 = n19255 ^ n4909 ^ 1'b0 ;
  assign n19257 = ~n1636 & n19256 ;
  assign n19258 = n890 | n8475 ;
  assign n19259 = ( n1938 & n9429 ) | ( n1938 & ~n19258 ) | ( n9429 & ~n19258 ) ;
  assign n19260 = n1859 & ~n11608 ;
  assign n19261 = n19260 ^ n8067 ^ 1'b0 ;
  assign n19262 = ~n1276 & n19261 ;
  assign n19263 = n19262 ^ n15725 ^ 1'b0 ;
  assign n19264 = x26 & n2243 ;
  assign n19265 = n19264 ^ n14803 ^ 1'b0 ;
  assign n19266 = n7855 ^ n1311 ^ 1'b0 ;
  assign n19267 = n4424 & ~n19266 ;
  assign n19268 = n19267 ^ n17363 ^ 1'b0 ;
  assign n19269 = n16059 & n19268 ;
  assign n19270 = n18336 ^ n16834 ^ n11720 ;
  assign n19271 = n7801 ^ n4567 ^ 1'b0 ;
  assign n19274 = n10047 ^ n7460 ^ 1'b0 ;
  assign n19275 = x195 & n19274 ;
  assign n19272 = n5367 | n8954 ;
  assign n19273 = n7417 | n19272 ;
  assign n19276 = n19275 ^ n19273 ^ 1'b0 ;
  assign n19277 = n7002 & n19276 ;
  assign n19278 = ~n16421 & n19277 ;
  assign n19279 = n2242 | n4168 ;
  assign n19280 = n19279 ^ n5431 ^ 1'b0 ;
  assign n19281 = ~n5428 & n19280 ;
  assign n19283 = n8300 ^ n2721 ^ n1530 ;
  assign n19282 = n7247 | n9955 ;
  assign n19284 = n19283 ^ n19282 ^ 1'b0 ;
  assign n19285 = n446 & n12919 ;
  assign n19286 = n19284 | n19285 ;
  assign n19287 = ~n5485 & n5659 ;
  assign n19288 = n4605 ^ n4598 ^ n3594 ;
  assign n19289 = ~n1079 & n3309 ;
  assign n19290 = ~n2929 & n19289 ;
  assign n19291 = n1742 & n19290 ;
  assign n19292 = ~n17747 & n19291 ;
  assign n19293 = n564 ^ n384 ^ 1'b0 ;
  assign n19294 = ~n17717 & n19293 ;
  assign n19295 = n15078 ^ n4519 ^ 1'b0 ;
  assign n19296 = x55 & ~n11097 ;
  assign n19297 = ~n11755 & n19296 ;
  assign n19298 = n19297 ^ n2332 ^ n905 ;
  assign n19299 = ~n6746 & n7199 ;
  assign n19300 = n19299 ^ n10758 ^ 1'b0 ;
  assign n19301 = n19298 | n19300 ;
  assign n19302 = n15137 | n19301 ;
  assign n19303 = n1903 | n19302 ;
  assign n19304 = ( n6726 & ~n14985 ) | ( n6726 & n15594 ) | ( ~n14985 & n15594 ) ;
  assign n19307 = n5359 & n10625 ;
  assign n19305 = ~n2032 & n2257 ;
  assign n19306 = n19305 ^ n810 ^ 1'b0 ;
  assign n19308 = n19307 ^ n19306 ^ 1'b0 ;
  assign n19310 = n16350 ^ n5836 ^ 1'b0 ;
  assign n19309 = ~n3498 & n5187 ;
  assign n19311 = n19310 ^ n19309 ^ 1'b0 ;
  assign n19312 = n19308 | n19311 ;
  assign n19313 = n16989 ^ n7466 ^ 1'b0 ;
  assign n19314 = n19312 | n19313 ;
  assign n19315 = n3635 ^ x13 ^ 1'b0 ;
  assign n19316 = ~n3284 & n5713 ;
  assign n19317 = ~n19315 & n19316 ;
  assign n19318 = n19317 ^ n5047 ^ 1'b0 ;
  assign n19319 = n9901 & n13054 ;
  assign n19320 = n5745 & n19319 ;
  assign n19321 = n668 & ~n13462 ;
  assign n19322 = n19320 & n19321 ;
  assign n19323 = n825 | n11625 ;
  assign n19324 = n1335 & ~n2958 ;
  assign n19325 = n19324 ^ n8897 ^ 1'b0 ;
  assign n19326 = n19325 ^ n19011 ^ 1'b0 ;
  assign n19327 = n7800 ^ n4691 ^ 1'b0 ;
  assign n19328 = n11776 ^ n3654 ^ 1'b0 ;
  assign n19329 = n4740 & ~n19328 ;
  assign n19330 = n19329 ^ n7603 ^ 1'b0 ;
  assign n19331 = n1759 & ~n16429 ;
  assign n19332 = n16576 ^ n6563 ^ 1'b0 ;
  assign n19333 = n3396 ^ n3011 ^ 1'b0 ;
  assign n19334 = n293 | n15730 ;
  assign n19335 = n440 & ~n19334 ;
  assign n19336 = n11619 ^ n7183 ^ 1'b0 ;
  assign n19337 = ~n2307 & n8627 ;
  assign n19338 = n19336 & ~n19337 ;
  assign n19339 = n19335 & n19338 ;
  assign n19340 = n19339 ^ n16030 ^ 1'b0 ;
  assign n19341 = n7287 ^ n4288 ^ 1'b0 ;
  assign n19342 = n6500 | n19341 ;
  assign n19343 = n1070 & n11197 ;
  assign n19344 = n19342 & n19343 ;
  assign n19345 = n13540 ^ n708 ^ 1'b0 ;
  assign n19346 = n19344 | n19345 ;
  assign n19347 = n17689 | n19346 ;
  assign n19348 = ~n340 & n5153 ;
  assign n19349 = n3925 ^ n2537 ^ n320 ;
  assign n19350 = n17616 & ~n19349 ;
  assign n19351 = n1249 & n19350 ;
  assign n19352 = n19348 & n19351 ;
  assign n19353 = n2083 & ~n10420 ;
  assign n19354 = n19352 & n19353 ;
  assign n19355 = x75 & n3392 ;
  assign n19356 = n287 & n19355 ;
  assign n19357 = n19356 ^ n3594 ^ 1'b0 ;
  assign n19358 = ~n5683 & n19357 ;
  assign n19359 = n10374 ^ n6467 ^ 1'b0 ;
  assign n19360 = n15312 & n19359 ;
  assign n19361 = ( n6693 & n19358 ) | ( n6693 & n19360 ) | ( n19358 & n19360 ) ;
  assign n19362 = n7748 & ~n19361 ;
  assign n19363 = n9742 & ~n12681 ;
  assign n19364 = n19363 ^ n9693 ^ 1'b0 ;
  assign n19365 = n2040 & ~n12714 ;
  assign n19366 = n4794 | n19365 ;
  assign n19367 = n7065 | n11935 ;
  assign n19368 = n2529 | n19367 ;
  assign n19369 = n19368 ^ n14829 ^ 1'b0 ;
  assign n19370 = n4222 ^ n483 ^ n464 ;
  assign n19371 = n19370 ^ n16625 ^ 1'b0 ;
  assign n19374 = x208 & ~n3846 ;
  assign n19375 = n19374 ^ x100 ^ 1'b0 ;
  assign n19376 = n10807 | n19375 ;
  assign n19377 = n19376 ^ n8071 ^ 1'b0 ;
  assign n19378 = n19377 ^ n2070 ^ 1'b0 ;
  assign n19379 = n11255 | n19378 ;
  assign n19372 = ~n672 & n12030 ;
  assign n19373 = n19372 ^ n8819 ^ n6036 ;
  assign n19380 = n19379 ^ n19373 ^ n10272 ;
  assign n19381 = ~n1497 & n11784 ;
  assign n19382 = n2665 | n13245 ;
  assign n19383 = n19382 ^ n632 ^ 1'b0 ;
  assign n19384 = n19383 ^ n6073 ^ 1'b0 ;
  assign n19385 = n19381 & ~n19384 ;
  assign n19386 = n3939 & n10246 ;
  assign n19387 = x195 & n19386 ;
  assign n19388 = ~n7818 & n19387 ;
  assign n19389 = n19388 ^ n15046 ^ 1'b0 ;
  assign n19390 = n2798 | n9278 ;
  assign n19391 = n19390 ^ n17476 ^ 1'b0 ;
  assign n19392 = n5350 & n19391 ;
  assign n19393 = n16042 ^ n9938 ^ 1'b0 ;
  assign n19394 = ~n1815 & n19393 ;
  assign n19395 = n19394 ^ n6769 ^ 1'b0 ;
  assign n19396 = n18046 & ~n19395 ;
  assign n19397 = n19396 ^ n4235 ^ 1'b0 ;
  assign n19398 = n6154 ^ n5270 ^ 1'b0 ;
  assign n19399 = n2856 & n19398 ;
  assign n19400 = ~n13126 & n19399 ;
  assign n19401 = n8649 & n19400 ;
  assign n19402 = n3106 & n14509 ;
  assign n19403 = n12142 | n15704 ;
  assign n19404 = n8534 & ~n19403 ;
  assign n19405 = n19404 ^ n11146 ^ 1'b0 ;
  assign n19406 = x45 & n19405 ;
  assign n19407 = n15475 ^ n13300 ^ 1'b0 ;
  assign n19408 = n19406 & n19407 ;
  assign n19409 = n19201 ^ n16887 ^ 1'b0 ;
  assign n19410 = n13537 ^ n11272 ^ 1'b0 ;
  assign n19411 = ~n4563 & n19410 ;
  assign n19412 = n19411 ^ n618 ^ 1'b0 ;
  assign n19413 = ( n949 & ~n3368 ) | ( n949 & n6474 ) | ( ~n3368 & n6474 ) ;
  assign n19414 = n3796 & ~n19413 ;
  assign n19415 = n3234 & n19414 ;
  assign n19416 = n9573 | n19415 ;
  assign n19417 = ( n8293 & ~n9132 ) | ( n8293 & n19416 ) | ( ~n9132 & n19416 ) ;
  assign n19418 = n2655 & n19417 ;
  assign n19419 = ~n3796 & n19418 ;
  assign n19420 = n13479 ^ n8725 ^ n7836 ;
  assign n19421 = n9919 & n11950 ;
  assign n19422 = ~n1161 & n19421 ;
  assign n19423 = n3782 & n9271 ;
  assign n19424 = n19423 ^ n14694 ^ 1'b0 ;
  assign n19425 = n19422 | n19424 ;
  assign n19426 = n2407 & n11662 ;
  assign n19427 = n12698 & n19426 ;
  assign n19428 = ~n320 & n8902 ;
  assign n19429 = n12215 | n13962 ;
  assign n19430 = n19429 ^ n4391 ^ 1'b0 ;
  assign n19431 = n19430 ^ n15703 ^ 1'b0 ;
  assign n19432 = ~n16580 & n19431 ;
  assign n19433 = n2004 | n3997 ;
  assign n19438 = n7051 & ~n7145 ;
  assign n19439 = ~n9440 & n19438 ;
  assign n19436 = n7868 ^ n2845 ^ 1'b0 ;
  assign n19437 = n1854 & ~n19436 ;
  assign n19440 = n19439 ^ n19437 ^ n13895 ;
  assign n19434 = ~n4792 & n14790 ;
  assign n19435 = n19434 ^ n13263 ^ 1'b0 ;
  assign n19441 = n19440 ^ n19435 ^ 1'b0 ;
  assign n19442 = n638 & n1055 ;
  assign n19443 = n1705 & n19442 ;
  assign n19444 = n13766 | n19443 ;
  assign n19445 = n12915 | n19444 ;
  assign n19446 = n17896 & n19445 ;
  assign n19447 = ~n6650 & n19446 ;
  assign n19448 = ( n970 & n1995 ) | ( n970 & ~n2845 ) | ( n1995 & ~n2845 ) ;
  assign n19449 = ~n11723 & n19448 ;
  assign n19450 = n19449 ^ n17141 ^ 1'b0 ;
  assign n19451 = n7903 ^ n2237 ^ 1'b0 ;
  assign n19452 = n12308 & ~n19298 ;
  assign n19453 = n19452 ^ n18075 ^ 1'b0 ;
  assign n19456 = n363 & n8360 ;
  assign n19454 = ~n3889 & n9016 ;
  assign n19455 = n15510 | n19454 ;
  assign n19457 = n19456 ^ n19455 ^ 1'b0 ;
  assign n19458 = n19457 ^ n8365 ^ 1'b0 ;
  assign n19459 = n15335 ^ n4325 ^ 1'b0 ;
  assign n19460 = n7321 ^ n6627 ^ n2492 ;
  assign n19461 = n19460 ^ n6333 ^ 1'b0 ;
  assign n19462 = ~n5859 & n19461 ;
  assign n19463 = n18181 ^ n15468 ^ 1'b0 ;
  assign n19464 = ( n2210 & n6264 ) | ( n2210 & n6734 ) | ( n6264 & n6734 ) ;
  assign n19476 = n4267 | n9733 ;
  assign n19477 = n19476 ^ n7457 ^ 1'b0 ;
  assign n19465 = n4436 | n10729 ;
  assign n19466 = n14428 & n19465 ;
  assign n19467 = n1553 ^ n742 ^ 1'b0 ;
  assign n19471 = x148 & n998 ;
  assign n19468 = n10917 & n13806 ;
  assign n19469 = n19468 ^ n6990 ^ 1'b0 ;
  assign n19470 = n9230 | n19469 ;
  assign n19472 = n19471 ^ n19470 ^ 1'b0 ;
  assign n19473 = n9353 & n19472 ;
  assign n19474 = n19467 & ~n19473 ;
  assign n19475 = n19466 & n19474 ;
  assign n19478 = n19477 ^ n19475 ^ 1'b0 ;
  assign n19479 = n9674 | n19478 ;
  assign n19480 = ( ~n4301 & n6511 ) | ( ~n4301 & n15489 ) | ( n6511 & n15489 ) ;
  assign n19482 = n7396 ^ n1657 ^ 1'b0 ;
  assign n19481 = n10475 & n19045 ;
  assign n19483 = n19482 ^ n19481 ^ 1'b0 ;
  assign n19484 = n19483 ^ n4123 ^ 1'b0 ;
  assign n19485 = n19480 & n19484 ;
  assign n19486 = n1473 | n4023 ;
  assign n19487 = n583 | n1075 ;
  assign n19488 = n19487 ^ n16562 ^ 1'b0 ;
  assign n19489 = ( x214 & n7135 ) | ( x214 & n9973 ) | ( n7135 & n9973 ) ;
  assign n19490 = n19488 & ~n19489 ;
  assign n19491 = n19490 ^ x3 ^ 1'b0 ;
  assign n19492 = n19486 & ~n19491 ;
  assign n19493 = n3880 ^ n1797 ^ 1'b0 ;
  assign n19494 = ( n10129 & n15875 ) | ( n10129 & n19493 ) | ( n15875 & n19493 ) ;
  assign n19501 = ( n2358 & n12162 ) | ( n2358 & n12571 ) | ( n12162 & n12571 ) ;
  assign n19496 = n2873 ^ n2194 ^ 1'b0 ;
  assign n19497 = ( n378 & n2020 ) | ( n378 & n19496 ) | ( n2020 & n19496 ) ;
  assign n19495 = n6202 & n11945 ;
  assign n19498 = n19497 ^ n19495 ^ 1'b0 ;
  assign n19499 = n4991 & ~n8295 ;
  assign n19500 = n19498 & n19499 ;
  assign n19502 = n19501 ^ n19500 ^ n1506 ;
  assign n19503 = ( n4259 & n14964 ) | ( n4259 & n16072 ) | ( n14964 & n16072 ) ;
  assign n19504 = ( n14303 & ~n16989 ) | ( n14303 & n19503 ) | ( ~n16989 & n19503 ) ;
  assign n19505 = n8125 ^ n1565 ^ 1'b0 ;
  assign n19506 = n19504 | n19505 ;
  assign n19507 = n19506 ^ n13899 ^ n11617 ;
  assign n19508 = n6794 ^ n2199 ^ 1'b0 ;
  assign n19509 = n3011 | n19508 ;
  assign n19510 = n961 & ~n3898 ;
  assign n19511 = n3898 & n19510 ;
  assign n19512 = n16551 ^ n274 ^ 1'b0 ;
  assign n19513 = n19512 ^ n13493 ^ 1'b0 ;
  assign n19514 = n19511 | n19513 ;
  assign n19515 = n19514 ^ n6077 ^ n6072 ;
  assign n19516 = n19509 & n19515 ;
  assign n19517 = n1125 & n19516 ;
  assign n19518 = n7448 ^ n5815 ^ 1'b0 ;
  assign n19519 = n12632 | n19518 ;
  assign n19521 = n5595 ^ n4309 ^ 1'b0 ;
  assign n19520 = ~n1119 & n8666 ;
  assign n19522 = n19521 ^ n19520 ^ 1'b0 ;
  assign n19523 = ~n8555 & n19522 ;
  assign n19524 = n8162 ^ n4676 ^ 1'b0 ;
  assign n19525 = n14159 ^ n11674 ^ 1'b0 ;
  assign n19526 = n19524 & ~n19525 ;
  assign n19527 = n19526 ^ n7734 ^ 1'b0 ;
  assign n19528 = n10837 ^ n5685 ^ 1'b0 ;
  assign n19529 = n19283 & n19528 ;
  assign n19530 = n7846 ^ n5315 ^ n2608 ;
  assign n19531 = n5632 & ~n19530 ;
  assign n19532 = ~n19529 & n19531 ;
  assign n19533 = n6046 ^ n3776 ^ 1'b0 ;
  assign n19534 = n618 | n15929 ;
  assign n19535 = ~n3047 & n5987 ;
  assign n19536 = n19535 ^ n11237 ^ 1'b0 ;
  assign n19537 = n13554 | n19536 ;
  assign n19538 = n9360 & ~n19537 ;
  assign n19539 = n1599 & n5490 ;
  assign n19540 = x115 & n19539 ;
  assign n19541 = n19540 ^ n6109 ^ 1'b0 ;
  assign n19542 = ~n8625 & n19541 ;
  assign n19543 = ~n17753 & n19542 ;
  assign n19544 = n4169 | n17733 ;
  assign n19545 = n19544 ^ n15899 ^ 1'b0 ;
  assign n19546 = n1985 ^ n1982 ^ 1'b0 ;
  assign n19547 = n911 & n19546 ;
  assign n19548 = n14851 ^ n3628 ^ 1'b0 ;
  assign n19549 = n19350 ^ n3611 ^ 1'b0 ;
  assign n19550 = n2446 | n10914 ;
  assign n19551 = n4480 ^ n2785 ^ 1'b0 ;
  assign n19552 = ~n4400 & n19551 ;
  assign n19553 = n19550 | n19552 ;
  assign n19555 = ~n473 & n9735 ;
  assign n19554 = n8916 ^ n8844 ^ n2743 ;
  assign n19556 = n19555 ^ n19554 ^ n12809 ;
  assign n19557 = n19556 ^ n6613 ^ n2840 ;
  assign n19558 = ~n2897 & n19306 ;
  assign n19559 = ~n1369 & n18453 ;
  assign n19564 = n11063 ^ x86 ^ 1'b0 ;
  assign n19565 = n4514 & ~n19564 ;
  assign n19566 = n19565 ^ n4180 ^ 1'b0 ;
  assign n19567 = n19566 ^ n5540 ^ 1'b0 ;
  assign n19560 = n10232 ^ n4131 ^ 1'b0 ;
  assign n19561 = n1257 | n19560 ;
  assign n19562 = n4003 | n19561 ;
  assign n19563 = n12131 | n19562 ;
  assign n19568 = n19567 ^ n19563 ^ 1'b0 ;
  assign n19569 = n1509 | n5075 ;
  assign n19570 = ( n1405 & ~n8118 ) | ( n1405 & n18948 ) | ( ~n8118 & n18948 ) ;
  assign n19571 = n8052 & ~n19570 ;
  assign n19572 = ~n6907 & n7737 ;
  assign n19573 = n16386 ^ n9711 ^ 1'b0 ;
  assign n19574 = n4767 | n5856 ;
  assign n19575 = n14157 | n19574 ;
  assign n19576 = n2950 | n3775 ;
  assign n19577 = n19576 ^ n4046 ^ 1'b0 ;
  assign n19578 = n14030 & n19577 ;
  assign n19579 = n9587 ^ n4778 ^ 1'b0 ;
  assign n19580 = ~n2430 & n19579 ;
  assign n19581 = n19580 ^ n2827 ^ 1'b0 ;
  assign n19582 = n3163 & n6447 ;
  assign n19583 = n14068 | n18742 ;
  assign n19584 = n19583 ^ n12578 ^ 1'b0 ;
  assign n19585 = ~n19582 & n19584 ;
  assign n19586 = ~n7072 & n10295 ;
  assign n19587 = ~n7404 & n19586 ;
  assign n19588 = ( n603 & ~n2149 ) | ( n603 & n8547 ) | ( ~n2149 & n8547 ) ;
  assign n19589 = n19588 ^ n13851 ^ 1'b0 ;
  assign n19590 = n1899 & ~n8725 ;
  assign n19591 = n1632 & n19590 ;
  assign n19592 = n19591 ^ n6350 ^ 1'b0 ;
  assign n19593 = n19592 ^ n12443 ^ 1'b0 ;
  assign n19594 = n19589 & ~n19593 ;
  assign n19595 = n6516 | n12353 ;
  assign n19596 = n2978 & ~n14491 ;
  assign n19597 = n6817 & n19596 ;
  assign n19598 = n19595 | n19597 ;
  assign n19599 = n19598 ^ n5047 ^ 1'b0 ;
  assign n19600 = n12610 ^ n3467 ^ 1'b0 ;
  assign n19601 = ~n7399 & n14620 ;
  assign n19602 = n6155 & n19601 ;
  assign n19603 = n6341 & n19602 ;
  assign n19604 = n15279 ^ n9646 ^ 1'b0 ;
  assign n19605 = n1494 & n5678 ;
  assign n19606 = n4400 & n12032 ;
  assign n19609 = n15572 ^ n4877 ^ 1'b0 ;
  assign n19610 = n15636 & n19609 ;
  assign n19607 = ~n9536 & n10407 ;
  assign n19608 = n19607 ^ n6014 ^ 1'b0 ;
  assign n19611 = n19610 ^ n19608 ^ 1'b0 ;
  assign n19612 = n16903 & n19611 ;
  assign n19613 = n18070 & n18700 ;
  assign n19615 = n12617 ^ n11030 ^ 1'b0 ;
  assign n19616 = n15828 & ~n19615 ;
  assign n19614 = n8022 | n14090 ;
  assign n19617 = n19616 ^ n19614 ^ 1'b0 ;
  assign n19618 = x73 & ~n19593 ;
  assign n19619 = n12612 ^ n1775 ^ 1'b0 ;
  assign n19620 = n14869 ^ n4325 ^ 1'b0 ;
  assign n19621 = n2080 & n19620 ;
  assign n19622 = n19621 ^ n9180 ^ 1'b0 ;
  assign n19623 = n19619 & n19622 ;
  assign n19624 = n9582 ^ n8676 ^ 1'b0 ;
  assign n19625 = n17355 | n19624 ;
  assign n19626 = n2767 & ~n6593 ;
  assign n19627 = n11449 & ~n14775 ;
  assign n19628 = ~n2530 & n19627 ;
  assign n19629 = n10746 | n19628 ;
  assign n19630 = n634 & ~n19629 ;
  assign n19631 = n12222 & ~n14900 ;
  assign n19632 = n1896 & ~n12528 ;
  assign n19633 = n632 & n19632 ;
  assign n19634 = n11905 ^ n3837 ^ 1'b0 ;
  assign n19635 = n4993 & n13817 ;
  assign n19636 = n19635 ^ n2116 ^ 1'b0 ;
  assign n19637 = n6391 & n13212 ;
  assign n19638 = n466 & n7506 ;
  assign n19639 = n9123 & n19638 ;
  assign n19640 = n19637 | n19639 ;
  assign n19641 = ( n4100 & n7868 ) | ( n4100 & n19640 ) | ( n7868 & n19640 ) ;
  assign n19642 = n19641 ^ n11891 ^ 1'b0 ;
  assign n19643 = n12340 & n13807 ;
  assign n19644 = n19643 ^ n3988 ^ 1'b0 ;
  assign n19645 = n14816 ^ n9377 ^ 1'b0 ;
  assign n19646 = n15524 ^ n3806 ^ x242 ;
  assign n19647 = n8054 ^ n2347 ^ 1'b0 ;
  assign n19648 = n1416 & n19647 ;
  assign n19649 = n1371 | n8591 ;
  assign n19650 = n19649 ^ n10615 ^ 1'b0 ;
  assign n19651 = ( n4234 & n19648 ) | ( n4234 & n19650 ) | ( n19648 & n19650 ) ;
  assign n19652 = n2050 & ~n5475 ;
  assign n19653 = n19652 ^ n18461 ^ 1'b0 ;
  assign n19654 = n6229 & ~n8178 ;
  assign n19655 = n1859 & n14879 ;
  assign n19656 = n19655 ^ n6934 ^ 1'b0 ;
  assign n19657 = n19654 | n19656 ;
  assign n19658 = n15866 ^ n2008 ^ 1'b0 ;
  assign n19659 = n11251 | n11892 ;
  assign n19660 = x185 & ~n12811 ;
  assign n19661 = ( n2540 & n13297 ) | ( n2540 & n14747 ) | ( n13297 & n14747 ) ;
  assign n19662 = n19661 ^ n3665 ^ 1'b0 ;
  assign n19663 = n10395 ^ n4210 ^ 1'b0 ;
  assign n19664 = n10601 | n12751 ;
  assign n19665 = n19664 ^ n5665 ^ 1'b0 ;
  assign n19666 = n19665 ^ n10177 ^ 1'b0 ;
  assign n19667 = n9905 ^ n1402 ^ 1'b0 ;
  assign n19668 = n17392 & n19667 ;
  assign n19669 = n14111 & n19668 ;
  assign n19670 = n19669 ^ n12083 ^ 1'b0 ;
  assign n19671 = ( ~n4260 & n7432 ) | ( ~n4260 & n11303 ) | ( n7432 & n11303 ) ;
  assign n19672 = n8456 & n19671 ;
  assign n19673 = n19672 ^ n17491 ^ 1'b0 ;
  assign n19674 = n10268 & ~n19673 ;
  assign n19675 = ~x75 & n19674 ;
  assign n19676 = n3560 ^ n2919 ^ 1'b0 ;
  assign n19677 = ~n9009 & n19676 ;
  assign n19678 = n19677 ^ n16254 ^ 1'b0 ;
  assign n19679 = n19678 ^ n19409 ^ 1'b0 ;
  assign n19682 = n18776 ^ n10729 ^ 1'b0 ;
  assign n19680 = n8512 & ~n14998 ;
  assign n19681 = n19680 ^ n7846 ^ 1'b0 ;
  assign n19683 = n19682 ^ n19681 ^ 1'b0 ;
  assign n19684 = n842 & n19683 ;
  assign n19685 = n14433 & n19684 ;
  assign n19686 = n18244 ^ n16539 ^ 1'b0 ;
  assign n19687 = ~n776 & n2141 ;
  assign n19688 = n7057 & n19687 ;
  assign n19689 = n10203 | n19688 ;
  assign n19690 = n19689 ^ n7759 ^ 1'b0 ;
  assign n19691 = n8008 & ~n9463 ;
  assign n19692 = ( ~n854 & n19690 ) | ( ~n854 & n19691 ) | ( n19690 & n19691 ) ;
  assign n19693 = n15689 | n19692 ;
  assign n19694 = n3408 | n6972 ;
  assign n19695 = n432 | n8401 ;
  assign n19696 = n17355 & n19695 ;
  assign n19697 = n17326 ^ x89 ^ 1'b0 ;
  assign n19698 = n11978 & ~n19697 ;
  assign n19699 = n3910 ^ n2840 ^ 1'b0 ;
  assign n19700 = n3573 & ~n19699 ;
  assign n19701 = ~n2310 & n19700 ;
  assign n19702 = n2158 & n19701 ;
  assign n19703 = n5475 | n5830 ;
  assign n19704 = n19703 ^ n547 ^ 1'b0 ;
  assign n19705 = n19704 ^ n10373 ^ 1'b0 ;
  assign n19706 = ~n10498 & n19705 ;
  assign n19707 = n19706 ^ n10244 ^ 1'b0 ;
  assign n19708 = n6580 & n19707 ;
  assign n19709 = n19708 ^ n6788 ^ 1'b0 ;
  assign n19710 = n1952 & n8845 ;
  assign n19711 = n2799 & ~n4184 ;
  assign n19712 = n17796 & n18450 ;
  assign n19713 = ~n2901 & n6177 ;
  assign n19714 = n631 | n19713 ;
  assign n19715 = n19714 ^ n9876 ^ 1'b0 ;
  assign n19716 = n3300 ^ n2399 ^ n1376 ;
  assign n19717 = n2054 | n3251 ;
  assign n19718 = n19716 | n19717 ;
  assign n19719 = n19718 ^ n7929 ^ 1'b0 ;
  assign n19720 = n19719 ^ x221 ^ 1'b0 ;
  assign n19721 = ~n954 & n19720 ;
  assign n19722 = n923 & n7435 ;
  assign n19723 = ~n9835 & n19722 ;
  assign n19724 = n19723 ^ n7107 ^ 1'b0 ;
  assign n19725 = n7524 & ~n19724 ;
  assign n19726 = n908 | n8207 ;
  assign n19727 = n11813 & ~n19726 ;
  assign n19728 = n16885 ^ n1274 ^ 1'b0 ;
  assign n19729 = n4245 & n5696 ;
  assign n19730 = n14742 ^ n2371 ^ 1'b0 ;
  assign n19731 = ~n8172 & n19730 ;
  assign n19732 = ~n12647 & n19731 ;
  assign n19733 = n3255 & ~n9708 ;
  assign n19734 = n19733 ^ n14428 ^ n4638 ;
  assign n19735 = n19734 ^ n9691 ^ 1'b0 ;
  assign n19736 = n18836 ^ n9213 ^ 1'b0 ;
  assign n19737 = n3023 | n9724 ;
  assign n19738 = n19737 ^ n1739 ^ 1'b0 ;
  assign n19739 = n14565 ^ n11330 ^ 1'b0 ;
  assign n19740 = n13207 | n19739 ;
  assign n19741 = ( n2226 & ~n2693 ) | ( n2226 & n5192 ) | ( ~n2693 & n5192 ) ;
  assign n19742 = ~n17949 & n19741 ;
  assign n19743 = ~n16505 & n18462 ;
  assign n19744 = n6295 | n10599 ;
  assign n19745 = ( n2620 & n14797 ) | ( n2620 & ~n19744 ) | ( n14797 & ~n19744 ) ;
  assign n19746 = n14996 & n15561 ;
  assign n19747 = n19746 ^ n15658 ^ 1'b0 ;
  assign n19748 = x70 & n17738 ;
  assign n19749 = n15370 & n19748 ;
  assign n19750 = n2275 & n12677 ;
  assign n19751 = n19750 ^ n16975 ^ 1'b0 ;
  assign n19752 = n2749 ^ n875 ^ 1'b0 ;
  assign n19753 = n4236 & ~n5428 ;
  assign n19754 = ( n16531 & n19752 ) | ( n16531 & ~n19753 ) | ( n19752 & ~n19753 ) ;
  assign n19755 = n627 ^ n525 ^ 1'b0 ;
  assign n19756 = ~n1981 & n9218 ;
  assign n19758 = n2634 & ~n11375 ;
  assign n19757 = ~n13776 & n17448 ;
  assign n19759 = n19758 ^ n19757 ^ 1'b0 ;
  assign n19760 = ~n17914 & n19759 ;
  assign n19761 = ( ~n19755 & n19756 ) | ( ~n19755 & n19760 ) | ( n19756 & n19760 ) ;
  assign n19762 = x221 & n2334 ;
  assign n19763 = n19762 ^ n3838 ^ 1'b0 ;
  assign n19764 = n6851 ^ n2108 ^ 1'b0 ;
  assign n19765 = n9030 & n19764 ;
  assign n19766 = n19765 ^ n16083 ^ 1'b0 ;
  assign n19767 = n6309 | n19766 ;
  assign n19768 = n5734 & ~n6976 ;
  assign n19769 = ~n19767 & n19768 ;
  assign n19770 = n6104 ^ n3075 ^ x153 ;
  assign n19771 = n1528 & n7987 ;
  assign n19772 = ~n15503 & n19771 ;
  assign n19773 = n10057 ^ n6849 ^ 1'b0 ;
  assign n19774 = n4755 & ~n19773 ;
  assign n19775 = ~n17686 & n18972 ;
  assign n19776 = n19775 ^ n11981 ^ 1'b0 ;
  assign n19780 = n2011 & ~n2909 ;
  assign n19781 = n9227 & n19780 ;
  assign n19777 = n2799 ^ n1623 ^ 1'b0 ;
  assign n19778 = n18381 ^ n3598 ^ n3134 ;
  assign n19779 = n19777 | n19778 ;
  assign n19782 = n19781 ^ n19779 ^ 1'b0 ;
  assign n19783 = ~n1664 & n7411 ;
  assign n19784 = n19783 ^ n14134 ^ 1'b0 ;
  assign n19785 = n5207 ^ n2416 ^ n1928 ;
  assign n19786 = n14531 ^ n11772 ^ 1'b0 ;
  assign n19787 = n19785 | n19786 ;
  assign n19788 = n19787 ^ n4145 ^ 1'b0 ;
  assign n19789 = n19788 ^ n18045 ^ 1'b0 ;
  assign n19790 = n8104 ^ n2622 ^ 1'b0 ;
  assign n19791 = n6164 ^ n4885 ^ 1'b0 ;
  assign n19792 = n3665 & ~n19791 ;
  assign n19793 = n19792 ^ n1028 ^ 1'b0 ;
  assign n19794 = ~n2819 & n5420 ;
  assign n19795 = n3488 | n19794 ;
  assign n19796 = n19795 ^ n2875 ^ 1'b0 ;
  assign n19797 = n5954 ^ n789 ^ 1'b0 ;
  assign n19798 = n4840 ^ n2895 ^ 1'b0 ;
  assign n19799 = n8256 ^ n1492 ^ 1'b0 ;
  assign n19800 = n19798 & n19799 ;
  assign n19801 = n19797 & n19800 ;
  assign n19802 = n19801 ^ n19597 ^ 1'b0 ;
  assign n19803 = n13338 ^ n6199 ^ 1'b0 ;
  assign n19804 = n6616 & n7877 ;
  assign n19805 = n19804 ^ n9669 ^ 1'b0 ;
  assign n19806 = n13038 ^ n4508 ^ 1'b0 ;
  assign n19807 = n17486 | n19806 ;
  assign n19808 = n10437 & ~n14315 ;
  assign n19809 = n19808 ^ n5442 ^ 1'b0 ;
  assign n19810 = n5193 ^ n4626 ^ x146 ;
  assign n19811 = n12172 & ~n19810 ;
  assign n19812 = n4543 & ~n17958 ;
  assign n19813 = ~n2127 & n5962 ;
  assign n19814 = n7499 | n10957 ;
  assign n19815 = n479 & ~n19814 ;
  assign n19816 = n19815 ^ n5626 ^ 1'b0 ;
  assign n19817 = n19813 & ~n19816 ;
  assign n19818 = n15405 ^ n3251 ^ 1'b0 ;
  assign n19819 = ~x254 & n336 ;
  assign n19820 = n19819 ^ n17910 ^ 1'b0 ;
  assign n19821 = ~n8312 & n19820 ;
  assign n19822 = n5941 & ~n10139 ;
  assign n19823 = ~n3007 & n18758 ;
  assign n19824 = n19823 ^ n9995 ^ 1'b0 ;
  assign n19825 = ~n2951 & n5851 ;
  assign n19826 = n11429 ^ x135 ^ 1'b0 ;
  assign n19827 = n16929 | n19826 ;
  assign n19828 = n15533 & ~n19827 ;
  assign n19829 = n11766 ^ n8729 ^ 1'b0 ;
  assign n19830 = n5135 & ~n19829 ;
  assign n19831 = ~n19828 & n19830 ;
  assign n19832 = n19825 & n19831 ;
  assign n19833 = n19824 | n19832 ;
  assign n19834 = n19822 & ~n19833 ;
  assign n19835 = n7190 & n18000 ;
  assign n19836 = n19835 ^ n5264 ^ 1'b0 ;
  assign n19837 = n8110 ^ n6173 ^ 1'b0 ;
  assign n19838 = n8585 & ~n14827 ;
  assign n19839 = n19838 ^ n9988 ^ 1'b0 ;
  assign n19840 = ~n426 & n789 ;
  assign n19841 = n426 & n19840 ;
  assign n19842 = n759 & n3294 ;
  assign n19843 = ~n759 & n19842 ;
  assign n19844 = x99 & ~n1509 ;
  assign n19845 = ~x99 & n19844 ;
  assign n19846 = n466 & ~n19845 ;
  assign n19847 = n19843 & n19846 ;
  assign n19848 = n19841 & ~n19847 ;
  assign n19849 = n13650 ^ n4204 ^ 1'b0 ;
  assign n19850 = n19848 & n19849 ;
  assign n19851 = ~n1456 & n19850 ;
  assign n19852 = n12402 & n13158 ;
  assign n19853 = n1734 & ~n18114 ;
  assign n19854 = ~n1734 & n19853 ;
  assign n19855 = n16422 | n19854 ;
  assign n19856 = n19854 & ~n19855 ;
  assign n19857 = n19852 & ~n19856 ;
  assign n19858 = ~n19851 & n19857 ;
  assign n19859 = n10145 & n10540 ;
  assign n19860 = n13531 & ~n19859 ;
  assign n19861 = n18766 ^ n13949 ^ 1'b0 ;
  assign n19862 = n3211 & n9912 ;
  assign n19863 = n19862 ^ n10569 ^ 1'b0 ;
  assign n19864 = n8921 & n10070 ;
  assign n19865 = ~n7958 & n19864 ;
  assign n19866 = ~n2075 & n2544 ;
  assign n19867 = n19866 ^ n3493 ^ 1'b0 ;
  assign n19868 = n13954 ^ n3074 ^ 1'b0 ;
  assign n19869 = x249 | n19868 ;
  assign n19870 = n17968 ^ n9730 ^ 1'b0 ;
  assign n19871 = n1416 | n19870 ;
  assign n19872 = n6686 & n14584 ;
  assign n19873 = n3134 & n4173 ;
  assign n19874 = n10337 ^ n361 ^ 1'b0 ;
  assign n19875 = n5488 & n19874 ;
  assign n19876 = n17858 & n19875 ;
  assign n19877 = ~n9187 & n19876 ;
  assign n19878 = ~n5236 & n19098 ;
  assign n19879 = n16764 ^ n12074 ^ n2240 ;
  assign n19880 = n2903 & n19879 ;
  assign n19881 = n9156 | n16100 ;
  assign n19882 = n19881 ^ n7968 ^ n4432 ;
  assign n19883 = n19882 ^ n10403 ^ 1'b0 ;
  assign n19884 = n8404 ^ n8344 ^ 1'b0 ;
  assign n19885 = n2424 | n19884 ;
  assign n19886 = n19885 ^ n9976 ^ n4691 ;
  assign n19887 = n7013 & ~n17756 ;
  assign n19888 = ~n1671 & n19887 ;
  assign n19889 = n10445 | n19888 ;
  assign n19890 = ( ~n11360 & n17741 ) | ( ~n11360 & n19889 ) | ( n17741 & n19889 ) ;
  assign n19891 = ~n19886 & n19890 ;
  assign n19892 = n5320 & n19891 ;
  assign n19893 = n2192 | n10405 ;
  assign n19894 = n19893 ^ n6018 ^ 1'b0 ;
  assign n19895 = n1073 & n19894 ;
  assign n19896 = n740 ^ x77 ^ 1'b0 ;
  assign n19897 = ~n11864 & n19896 ;
  assign n19898 = ( n3565 & n16202 ) | ( n3565 & ~n19897 ) | ( n16202 & ~n19897 ) ;
  assign n19899 = ~n2799 & n5519 ;
  assign n19900 = n19899 ^ n7191 ^ n6759 ;
  assign n19901 = ~n948 & n2397 ;
  assign n19902 = n4197 | n7759 ;
  assign n19903 = n19902 ^ n14062 ^ 1'b0 ;
  assign n19904 = n3372 & ~n16473 ;
  assign n19905 = n19904 ^ n12696 ^ 1'b0 ;
  assign n19906 = ~n7157 & n16313 ;
  assign n19907 = n5355 & ~n11295 ;
  assign n19908 = ~n19906 & n19907 ;
  assign n19909 = ( n1774 & ~n1798 ) | ( n1774 & n16252 ) | ( ~n1798 & n16252 ) ;
  assign n19910 = ~n2970 & n14002 ;
  assign n19911 = n17433 & n18554 ;
  assign n19912 = n6884 & n15210 ;
  assign n19913 = n6061 & ~n19912 ;
  assign n19914 = n19913 ^ n8251 ^ 1'b0 ;
  assign n19915 = n8670 ^ n1111 ^ 1'b0 ;
  assign n19916 = n19915 ^ n12288 ^ 1'b0 ;
  assign n19917 = n3090 & ~n19916 ;
  assign n19918 = n4387 & n4417 ;
  assign n19919 = n19918 ^ n17903 ^ 1'b0 ;
  assign n19920 = n4929 & n6171 ;
  assign n19921 = n19920 ^ n1620 ^ 1'b0 ;
  assign n19922 = n7637 & ~n11743 ;
  assign n19923 = n19922 ^ n12513 ^ n2403 ;
  assign n19924 = n8276 | n11511 ;
  assign n19925 = n19466 & ~n19924 ;
  assign n19926 = n19925 ^ n2083 ^ 1'b0 ;
  assign n19927 = n8311 ^ n2130 ^ 1'b0 ;
  assign n19928 = n7951 & n17755 ;
  assign n19929 = n3993 & ~n14029 ;
  assign n19930 = n12297 ^ n10347 ^ 1'b0 ;
  assign n19931 = ~n10172 & n14639 ;
  assign n19932 = n19931 ^ n6350 ^ 1'b0 ;
  assign n19933 = n6626 & n7264 ;
  assign n19934 = n19933 ^ n11653 ^ 1'b0 ;
  assign n19935 = n6155 | n10689 ;
  assign n19936 = n19935 ^ n4260 ^ 1'b0 ;
  assign n19937 = n14765 ^ n13694 ^ 1'b0 ;
  assign n19938 = n10243 | n19937 ;
  assign n19939 = n19936 | n19938 ;
  assign n19940 = n17067 ^ n2001 ^ 1'b0 ;
  assign n19941 = n19940 ^ n16674 ^ 1'b0 ;
  assign n19942 = n8293 ^ n1293 ^ 1'b0 ;
  assign n19943 = n18641 | n19942 ;
  assign n19944 = n14436 & ~n17507 ;
  assign n19945 = n2123 & ~n13776 ;
  assign n19946 = n19945 ^ n5296 ^ 1'b0 ;
  assign n19947 = n16495 & ~n19946 ;
  assign n19948 = n12887 & n14040 ;
  assign n19949 = n16778 ^ n11041 ^ 1'b0 ;
  assign n19950 = n2950 & n19949 ;
  assign n19951 = n2041 & ~n6270 ;
  assign n19952 = n509 & n19951 ;
  assign n19953 = n19952 ^ n10903 ^ 1'b0 ;
  assign n19954 = n9615 & ~n14185 ;
  assign n19955 = n9747 & n17287 ;
  assign n19956 = n4254 & n6540 ;
  assign n19957 = n5578 & ~n5665 ;
  assign n19958 = n19957 ^ n7964 ^ 1'b0 ;
  assign n19959 = n18694 | n19958 ;
  assign n19960 = n845 & ~n19959 ;
  assign n19961 = n1915 | n3225 ;
  assign n19962 = n3659 ^ n2535 ^ 1'b0 ;
  assign n19963 = n1723 & n19962 ;
  assign n19964 = n9177 & ~n19963 ;
  assign n19965 = n14487 ^ x117 ^ 1'b0 ;
  assign n19966 = ~n4218 & n19965 ;
  assign n19967 = n19964 & n19966 ;
  assign n19968 = n387 & ~n10031 ;
  assign n19969 = n19968 ^ n11863 ^ 1'b0 ;
  assign n19970 = n8172 ^ n6122 ^ 1'b0 ;
  assign n19971 = n19970 ^ n19777 ^ 1'b0 ;
  assign n19972 = n4009 & ~n4253 ;
  assign n19973 = n19972 ^ n7134 ^ 1'b0 ;
  assign n19974 = n329 & ~n4450 ;
  assign n19975 = ~n11030 & n19974 ;
  assign n19976 = n6470 & n19975 ;
  assign n19977 = n19976 ^ n8792 ^ 1'b0 ;
  assign n19978 = n7291 & ~n12708 ;
  assign n19979 = n19978 ^ n6875 ^ 1'b0 ;
  assign n19980 = n11287 & n19979 ;
  assign n19981 = n17875 ^ n5307 ^ 1'b0 ;
  assign n19982 = ~n18384 & n19981 ;
  assign n19983 = n2925 | n10053 ;
  assign n19984 = n19983 ^ n10606 ^ 1'b0 ;
  assign n19985 = ~n4506 & n17808 ;
  assign n19986 = x47 & ~n1788 ;
  assign n19987 = ( n6495 & ~n8523 ) | ( n6495 & n19986 ) | ( ~n8523 & n19986 ) ;
  assign n19988 = ( x87 & ~n10239 ) | ( x87 & n15886 ) | ( ~n10239 & n15886 ) ;
  assign n19989 = ~n4508 & n18726 ;
  assign n19990 = n19989 ^ n1383 ^ 1'b0 ;
  assign n19991 = n10911 & ~n19990 ;
  assign n19992 = n19988 & n19991 ;
  assign n19993 = n8688 | n16686 ;
  assign n19994 = n1468 & ~n19993 ;
  assign n19995 = n16786 & ~n19994 ;
  assign n19996 = n14242 & n19995 ;
  assign n19997 = n3178 | n14007 ;
  assign n19998 = ~n6987 & n19997 ;
  assign n19999 = n15910 ^ n10847 ^ 1'b0 ;
  assign n20000 = ~n9213 & n19999 ;
  assign n20001 = n2465 & n20000 ;
  assign n20002 = n12124 & ~n14062 ;
  assign n20003 = ~n3451 & n15273 ;
  assign n20004 = n20002 & n20003 ;
  assign n20005 = n18022 ^ n11415 ^ 1'b0 ;
  assign n20006 = n20004 | n20005 ;
  assign n20007 = n1165 | n12094 ;
  assign n20008 = n20006 & ~n20007 ;
  assign n20009 = ~n3345 & n6271 ;
  assign n20010 = n20009 ^ n774 ^ 1'b0 ;
  assign n20011 = ~n3554 & n7659 ;
  assign n20012 = ~n20010 & n20011 ;
  assign n20013 = n20012 ^ n11084 ^ 1'b0 ;
  assign n20014 = ~n4222 & n20013 ;
  assign n20015 = n5296 & n11483 ;
  assign n20016 = n20014 & n20015 ;
  assign n20017 = x152 | n20016 ;
  assign n20018 = n10191 ^ n492 ^ 1'b0 ;
  assign n20019 = n16913 & n20018 ;
  assign n20020 = n18856 ^ n8639 ^ 1'b0 ;
  assign n20021 = n19599 ^ n10152 ^ 1'b0 ;
  assign n20022 = ~n4094 & n16329 ;
  assign n20023 = ~n16487 & n20022 ;
  assign n20024 = ( n11010 & ~n14240 ) | ( n11010 & n20023 ) | ( ~n14240 & n20023 ) ;
  assign n20025 = ~n11737 & n12786 ;
  assign n20026 = n12940 & n20025 ;
  assign n20027 = n14555 ^ n3898 ^ 1'b0 ;
  assign n20028 = ~n1204 & n20027 ;
  assign n20029 = n3012 | n7456 ;
  assign n20030 = n6638 | n20029 ;
  assign n20031 = n9905 & ~n15777 ;
  assign n20032 = ~n2167 & n20031 ;
  assign n20033 = n1853 & ~n15761 ;
  assign n20034 = ~n1779 & n12310 ;
  assign n20035 = ~n12962 & n17837 ;
  assign n20036 = n5235 & n20035 ;
  assign n20037 = n20036 ^ n2246 ^ n2024 ;
  assign n20038 = n15647 ^ n5544 ^ 1'b0 ;
  assign n20039 = n17533 & n19493 ;
  assign n20040 = n1354 | n20039 ;
  assign n20041 = n20040 ^ n6355 ^ 1'b0 ;
  assign n20042 = n6015 & n20041 ;
  assign n20043 = ~n1410 & n20042 ;
  assign n20044 = n4500 & ~n12301 ;
  assign n20045 = n10867 ^ n5010 ^ 1'b0 ;
  assign n20046 = n5160 | n20045 ;
  assign n20047 = n11777 & ~n20046 ;
  assign n20048 = n12841 & n20047 ;
  assign n20049 = n20048 ^ n2056 ^ 1'b0 ;
  assign n20050 = n1328 | n2846 ;
  assign n20051 = n20050 ^ n5602 ^ 1'b0 ;
  assign n20052 = ( ~n19317 & n20049 ) | ( ~n19317 & n20051 ) | ( n20049 & n20051 ) ;
  assign n20053 = n5492 | n15880 ;
  assign n20054 = n20053 ^ n16193 ^ 1'b0 ;
  assign n20055 = ( n4430 & n9270 ) | ( n4430 & n20054 ) | ( n9270 & n20054 ) ;
  assign n20056 = ( n1583 & n3571 ) | ( n1583 & ~n8104 ) | ( n3571 & ~n8104 ) ;
  assign n20057 = n2746 & ~n20056 ;
  assign n20058 = ~n14843 & n20057 ;
  assign n20059 = n10731 & ~n17308 ;
  assign n20060 = n16804 & n20059 ;
  assign n20062 = n5912 ^ n1968 ^ 1'b0 ;
  assign n20063 = n5474 & n20062 ;
  assign n20061 = n6359 | n6731 ;
  assign n20064 = n20063 ^ n20061 ^ 1'b0 ;
  assign n20067 = n12856 ^ n7606 ^ 1'b0 ;
  assign n20065 = n591 & n5848 ;
  assign n20066 = n10298 | n20065 ;
  assign n20068 = n20067 ^ n20066 ^ 1'b0 ;
  assign n20069 = n20068 ^ n10794 ^ 1'b0 ;
  assign n20070 = n15042 ^ n8855 ^ 1'b0 ;
  assign n20071 = n17933 | n20070 ;
  assign n20072 = n6999 | n8519 ;
  assign n20073 = n20072 ^ n8424 ^ 1'b0 ;
  assign n20074 = ~n6927 & n11819 ;
  assign n20075 = ~n19936 & n20074 ;
  assign n20076 = ( ~n5768 & n18268 ) | ( ~n5768 & n20075 ) | ( n18268 & n20075 ) ;
  assign n20077 = n2076 & ~n16240 ;
  assign n20078 = n20077 ^ n7877 ^ 1'b0 ;
  assign n20079 = n20076 | n20078 ;
  assign n20080 = n14542 ^ n14311 ^ 1'b0 ;
  assign n20081 = ~n20079 & n20080 ;
  assign n20082 = n20081 ^ n618 ^ 1'b0 ;
  assign n20083 = n20073 & ~n20082 ;
  assign n20084 = n3806 & ~n3929 ;
  assign n20085 = n20084 ^ n4348 ^ 1'b0 ;
  assign n20086 = n8222 | n20085 ;
  assign n20087 = n3420 & ~n11926 ;
  assign n20088 = ~n604 & n20087 ;
  assign n20089 = n10737 ^ n9659 ^ x70 ;
  assign n20090 = ~n1473 & n20089 ;
  assign n20091 = n8470 ^ n6723 ^ 1'b0 ;
  assign n20092 = n20091 ^ n5604 ^ 1'b0 ;
  assign n20093 = n10242 | n20092 ;
  assign n20094 = n16990 ^ n10545 ^ n5404 ;
  assign n20095 = n13836 | n19594 ;
  assign n20096 = n5049 & ~n7084 ;
  assign n20097 = n3411 & ~n20096 ;
  assign n20098 = n20097 ^ n10305 ^ 1'b0 ;
  assign n20099 = n13443 ^ n4966 ^ 1'b0 ;
  assign n20100 = n17631 & ~n20099 ;
  assign n20104 = n8823 ^ n3007 ^ x163 ;
  assign n20105 = n20104 ^ n12688 ^ 1'b0 ;
  assign n20101 = n4122 ^ n3012 ^ 1'b0 ;
  assign n20102 = n597 & n20101 ;
  assign n20103 = ~n1638 & n20102 ;
  assign n20106 = n20105 ^ n20103 ^ 1'b0 ;
  assign n20107 = n2697 | n15819 ;
  assign n20108 = n8487 ^ n4811 ^ 1'b0 ;
  assign n20109 = n1613 & n1698 ;
  assign n20110 = ~n20108 & n20109 ;
  assign n20111 = ( ~x154 & n2301 ) | ( ~x154 & n9400 ) | ( n2301 & n9400 ) ;
  assign n20112 = n3312 | n20111 ;
  assign n20113 = n17229 & ~n19102 ;
  assign n20114 = ( ~n7385 & n20112 ) | ( ~n7385 & n20113 ) | ( n20112 & n20113 ) ;
  assign n20115 = n15181 & ~n20114 ;
  assign n20116 = n14937 ^ n6730 ^ 1'b0 ;
  assign n20118 = n16360 ^ n7807 ^ 1'b0 ;
  assign n20117 = n14193 & n14363 ;
  assign n20119 = n20118 ^ n20117 ^ 1'b0 ;
  assign n20120 = n6030 | n11776 ;
  assign n20121 = ~n16241 & n20120 ;
  assign n20124 = n7839 & n10180 ;
  assign n20125 = n12719 & n20124 ;
  assign n20122 = n12596 ^ n11347 ^ 1'b0 ;
  assign n20123 = ~n3676 & n20122 ;
  assign n20126 = n20125 ^ n20123 ^ 1'b0 ;
  assign n20127 = n10280 ^ n9890 ^ 1'b0 ;
  assign n20128 = n9981 & ~n20127 ;
  assign n20129 = n18663 ^ n8968 ^ 1'b0 ;
  assign n20130 = n675 & n9072 ;
  assign n20131 = n1100 & ~n3806 ;
  assign n20132 = ~n2020 & n2200 ;
  assign n20133 = n20132 ^ n6605 ^ 1'b0 ;
  assign n20134 = n7134 | n20133 ;
  assign n20135 = n16627 ^ n13253 ^ n4527 ;
  assign n20136 = n20135 ^ x15 ^ 1'b0 ;
  assign n20137 = ( n661 & n3724 ) | ( n661 & n9695 ) | ( n3724 & n9695 ) ;
  assign n20138 = ~n1332 & n20137 ;
  assign n20139 = n12204 ^ n7053 ^ 1'b0 ;
  assign n20140 = ~n15459 & n20139 ;
  assign n20141 = n16095 ^ n14442 ^ 1'b0 ;
  assign n20142 = ~n6782 & n13101 ;
  assign n20143 = n20142 ^ n19200 ^ 1'b0 ;
  assign n20144 = ( n6483 & ~n10714 ) | ( n6483 & n11645 ) | ( ~n10714 & n11645 ) ;
  assign n20145 = n20144 ^ n5542 ^ x206 ;
  assign n20146 = n20145 ^ n9621 ^ 1'b0 ;
  assign n20147 = ~n14762 & n17763 ;
  assign n20148 = n4325 & n20147 ;
  assign n20149 = n20146 & ~n20148 ;
  assign n20150 = ~n5906 & n20149 ;
  assign n20151 = n20150 ^ n12830 ^ 1'b0 ;
  assign n20153 = n5551 & n6561 ;
  assign n20152 = ~n320 & n4792 ;
  assign n20154 = n20153 ^ n20152 ^ 1'b0 ;
  assign n20158 = n2919 ^ n496 ^ 1'b0 ;
  assign n20155 = n13649 & ~n15368 ;
  assign n20156 = n11871 & n20155 ;
  assign n20157 = n4758 | n20156 ;
  assign n20159 = n20158 ^ n20157 ^ 1'b0 ;
  assign n20160 = n19649 ^ n4424 ^ 1'b0 ;
  assign n20161 = n20160 ^ n18690 ^ 1'b0 ;
  assign n20162 = n4903 & n20161 ;
  assign n20163 = n2164 & ~n14209 ;
  assign n20164 = n20163 ^ x118 ^ 1'b0 ;
  assign n20165 = n20162 & n20164 ;
  assign n20166 = n12463 & ~n20165 ;
  assign n20167 = n1392 & ~n7241 ;
  assign n20168 = n20167 ^ n7521 ^ 1'b0 ;
  assign n20169 = ~n1630 & n20168 ;
  assign n20170 = ~n10694 & n12898 ;
  assign n20171 = n13521 & ~n16834 ;
  assign n20172 = n2627 & n20171 ;
  assign n20173 = n3588 & n10630 ;
  assign n20174 = n20173 ^ n16231 ^ 1'b0 ;
  assign n20175 = ~n7356 & n20174 ;
  assign n20176 = ~n8049 & n20175 ;
  assign n20177 = n4766 & n20176 ;
  assign n20178 = ~n13849 & n15185 ;
  assign n20179 = n13849 & n20178 ;
  assign n20180 = n5293 ^ n306 ^ 1'b0 ;
  assign n20181 = n8902 | n13620 ;
  assign n20182 = n12714 & n20181 ;
  assign n20183 = ~n1213 & n7295 ;
  assign n20184 = n20183 ^ n3917 ^ 1'b0 ;
  assign n20185 = n8308 & n9520 ;
  assign n20186 = n20185 ^ n4652 ^ 1'b0 ;
  assign n20187 = n16528 ^ n8951 ^ 1'b0 ;
  assign n20188 = n879 & n10615 ;
  assign n20189 = ~n2001 & n3817 ;
  assign n20190 = ~n8872 & n20189 ;
  assign n20191 = n12100 ^ n10305 ^ 1'b0 ;
  assign n20192 = ~n14234 & n20191 ;
  assign n20193 = n20192 ^ n10988 ^ 1'b0 ;
  assign n20195 = ( n2936 & ~n4956 ) | ( n2936 & n15037 ) | ( ~n4956 & n15037 ) ;
  assign n20196 = ~n5870 & n20195 ;
  assign n20194 = n1903 & ~n10004 ;
  assign n20197 = n20196 ^ n20194 ^ 1'b0 ;
  assign n20198 = n18184 ^ n2463 ^ 1'b0 ;
  assign n20199 = ~n2611 & n13912 ;
  assign n20200 = n1100 & n20199 ;
  assign n20201 = n611 & n4260 ;
  assign n20202 = n20201 ^ n9782 ^ n8671 ;
  assign n20203 = n8764 & ~n16105 ;
  assign n20204 = ( n2570 & n5177 ) | ( n2570 & ~n11403 ) | ( n5177 & ~n11403 ) ;
  assign n20205 = n9605 ^ n2348 ^ 1'b0 ;
  assign n20206 = n18326 & n20205 ;
  assign n20207 = ~n20204 & n20206 ;
  assign n20208 = n14273 & n20207 ;
  assign n20209 = ~n8305 & n20208 ;
  assign n20210 = n2092 & n20209 ;
  assign n20211 = ( n1073 & n7258 ) | ( n1073 & ~n9753 ) | ( n7258 & ~n9753 ) ;
  assign n20212 = n1525 | n2890 ;
  assign n20213 = n20212 ^ n6238 ^ 1'b0 ;
  assign n20214 = ~n3113 & n20213 ;
  assign n20215 = n9640 & ~n16224 ;
  assign n20216 = ~n20214 & n20215 ;
  assign n20217 = n8471 ^ n6441 ^ 1'b0 ;
  assign n20219 = ~n2337 & n3576 ;
  assign n20220 = n8827 & n20219 ;
  assign n20218 = n5813 | n13675 ;
  assign n20221 = n20220 ^ n20218 ^ 1'b0 ;
  assign n20222 = ~n6256 & n11323 ;
  assign n20223 = n8681 & n17711 ;
  assign n20224 = n5920 | n11483 ;
  assign n20225 = ~n13739 & n18468 ;
  assign n20226 = n20224 | n20225 ;
  assign n20227 = n17045 & ~n20226 ;
  assign n20228 = ~n9134 & n12414 ;
  assign n20229 = n6559 & n20228 ;
  assign n20230 = n7939 & ~n20229 ;
  assign n20231 = n6263 & n20230 ;
  assign n20240 = ~x89 & n11105 ;
  assign n20241 = n20240 ^ n6157 ^ 1'b0 ;
  assign n20242 = n16144 & ~n20241 ;
  assign n20232 = n7940 & ~n14756 ;
  assign n20233 = n20232 ^ n4095 ^ 1'b0 ;
  assign n20234 = n7308 ^ n4287 ^ 1'b0 ;
  assign n20235 = n12587 & n20234 ;
  assign n20236 = n3439 | n20235 ;
  assign n20237 = n20236 ^ n13011 ^ 1'b0 ;
  assign n20238 = n20233 | n20237 ;
  assign n20239 = n13305 & ~n20238 ;
  assign n20243 = n20242 ^ n20239 ^ 1'b0 ;
  assign n20244 = ~n1251 & n8622 ;
  assign n20245 = ( n10403 & n14737 ) | ( n10403 & ~n20244 ) | ( n14737 & ~n20244 ) ;
  assign n20246 = n9572 & ~n18814 ;
  assign n20247 = n20246 ^ n19470 ^ 1'b0 ;
  assign n20248 = n749 & ~n16025 ;
  assign n20249 = n20248 ^ n3364 ^ 1'b0 ;
  assign n20250 = n9347 ^ n7462 ^ 1'b0 ;
  assign n20251 = ( n4619 & n10530 ) | ( n4619 & n15674 ) | ( n10530 & n15674 ) ;
  assign n20252 = ~n8622 & n15889 ;
  assign n20253 = n4135 & ~n18597 ;
  assign n20255 = ~n1020 & n2073 ;
  assign n20256 = ~x253 & n20255 ;
  assign n20254 = ~x21 & n6023 ;
  assign n20257 = n20256 ^ n20254 ^ 1'b0 ;
  assign n20258 = n7526 & n20257 ;
  assign n20259 = n8116 ^ n2937 ^ 1'b0 ;
  assign n20260 = ( ~n17409 & n20258 ) | ( ~n17409 & n20259 ) | ( n20258 & n20259 ) ;
  assign n20261 = n577 | n14305 ;
  assign n20262 = n20261 ^ n8150 ^ n6483 ;
  assign n20263 = n17648 ^ n15543 ^ 1'b0 ;
  assign n20264 = n9885 | n20263 ;
  assign n20265 = n7038 & ~n7999 ;
  assign n20266 = n18733 ^ n17345 ^ 1'b0 ;
  assign n20267 = n12971 & ~n20266 ;
  assign n20268 = ~n6088 & n20267 ;
  assign n20269 = n20268 ^ n8414 ^ 1'b0 ;
  assign n20270 = n13986 ^ n3410 ^ 1'b0 ;
  assign n20271 = n19126 ^ n2718 ^ n1620 ;
  assign n20272 = n9721 ^ n8959 ^ 1'b0 ;
  assign n20273 = n11028 & ~n20272 ;
  assign n20274 = n6952 ^ n4923 ^ 1'b0 ;
  assign n20275 = ~n3549 & n20274 ;
  assign n20277 = n2950 ^ n903 ^ 1'b0 ;
  assign n20276 = ~n8244 & n18397 ;
  assign n20278 = n20277 ^ n20276 ^ 1'b0 ;
  assign n20280 = n13944 ^ n3498 ^ 1'b0 ;
  assign n20279 = ( n4654 & n9128 ) | ( n4654 & ~n13353 ) | ( n9128 & ~n13353 ) ;
  assign n20281 = n20280 ^ n20279 ^ n11345 ;
  assign n20282 = n12516 ^ n10177 ^ n2055 ;
  assign n20283 = n1931 | n20282 ;
  assign n20287 = n312 | n1989 ;
  assign n20286 = n1600 & ~n12939 ;
  assign n20288 = n20287 ^ n20286 ^ 1'b0 ;
  assign n20284 = n2866 & n3795 ;
  assign n20285 = n9505 & n20284 ;
  assign n20289 = n20288 ^ n20285 ^ n12719 ;
  assign n20290 = ~n3699 & n12146 ;
  assign n20291 = n20289 & n20290 ;
  assign n20292 = n2319 & n20291 ;
  assign n20293 = ( n4061 & n10387 ) | ( n4061 & ~n10675 ) | ( n10387 & ~n10675 ) ;
  assign n20294 = n9934 ^ n3614 ^ 1'b0 ;
  assign n20295 = n20293 & ~n20294 ;
  assign n20300 = n17333 ^ n7437 ^ 1'b0 ;
  assign n20301 = n16348 | n20300 ;
  assign n20296 = n4520 & ~n6348 ;
  assign n20297 = n20296 ^ n5190 ^ 1'b0 ;
  assign n20298 = n1509 & ~n3520 ;
  assign n20299 = n20297 & n20298 ;
  assign n20302 = n20301 ^ n20299 ^ 1'b0 ;
  assign n20303 = n2835 | n5509 ;
  assign n20304 = ~n6632 & n20303 ;
  assign n20305 = n2122 & n20304 ;
  assign n20306 = n20305 ^ n15662 ^ n8592 ;
  assign n20307 = n15080 ^ n4755 ^ 1'b0 ;
  assign n20308 = ~x184 & n20307 ;
  assign n20309 = n9600 ^ n4646 ^ 1'b0 ;
  assign n20310 = n13948 & n20309 ;
  assign n20311 = n20041 ^ n18310 ^ 1'b0 ;
  assign n20312 = ~n10236 & n20311 ;
  assign n20313 = n9196 ^ n3127 ^ 1'b0 ;
  assign n20314 = n11920 ^ n9072 ^ n6781 ;
  assign n20315 = ( n13949 & n20313 ) | ( n13949 & n20314 ) | ( n20313 & n20314 ) ;
  assign n20316 = n20315 ^ n17229 ^ n2915 ;
  assign n20317 = n10803 & n20316 ;
  assign n20318 = ( ~n2157 & n3499 ) | ( ~n2157 & n10809 ) | ( n3499 & n10809 ) ;
  assign n20319 = n2549 | n13176 ;
  assign n20320 = n20319 ^ n6593 ^ 1'b0 ;
  assign n20321 = n15491 & ~n20320 ;
  assign n20322 = n20318 & n20321 ;
  assign n20323 = n497 | n13848 ;
  assign n20324 = n20323 ^ n13653 ^ 1'b0 ;
  assign n20325 = n5172 & n15477 ;
  assign n20326 = n20325 ^ n11609 ^ 1'b0 ;
  assign n20327 = n1878 & ~n8219 ;
  assign n20328 = ~n5898 & n20327 ;
  assign n20329 = n1716 & ~n17076 ;
  assign n20330 = n20328 & n20329 ;
  assign n20331 = n18734 | n20330 ;
  assign n20332 = n3279 & ~n20331 ;
  assign n20333 = n10266 & n12244 ;
  assign n20334 = n8182 ^ n2076 ^ 1'b0 ;
  assign n20335 = ~n2600 & n20334 ;
  assign n20336 = ( ~n3293 & n19297 ) | ( ~n3293 & n20335 ) | ( n19297 & n20335 ) ;
  assign n20337 = n18123 ^ n10404 ^ 1'b0 ;
  assign n20338 = n445 & n11167 ;
  assign n20339 = n9246 & n12811 ;
  assign n20340 = n1553 | n15347 ;
  assign n20341 = n838 & n4045 ;
  assign n20342 = n491 & ~n8547 ;
  assign n20345 = n7344 ^ n4400 ^ n420 ;
  assign n20343 = n5803 & n8269 ;
  assign n20344 = ~n13911 & n20343 ;
  assign n20346 = n20345 ^ n20344 ^ 1'b0 ;
  assign n20347 = n1185 & ~n4025 ;
  assign n20348 = n2242 ^ n1674 ^ n1234 ;
  assign n20349 = n20347 & ~n20348 ;
  assign n20350 = n4323 & ~n4639 ;
  assign n20351 = n19344 ^ n14988 ^ n4410 ;
  assign n20352 = n6679 ^ n1081 ^ 1'b0 ;
  assign n20353 = n17899 | n20352 ;
  assign n20354 = n2935 ^ n2627 ^ 1'b0 ;
  assign n20355 = n6906 & n20354 ;
  assign n20356 = n20353 & n20355 ;
  assign n20357 = n15756 ^ n11672 ^ 1'b0 ;
  assign n20358 = n6886 & n20357 ;
  assign n20368 = ( ~n3722 & n10876 ) | ( ~n3722 & n13083 ) | ( n10876 & n13083 ) ;
  assign n20359 = n2322 ^ n1288 ^ 1'b0 ;
  assign n20360 = n5407 & n20359 ;
  assign n20361 = n13452 & n20360 ;
  assign n20362 = n2297 | n2749 ;
  assign n20363 = n8877 ^ n4957 ^ 1'b0 ;
  assign n20364 = n10888 & n20363 ;
  assign n20365 = ( n12573 & n20362 ) | ( n12573 & n20364 ) | ( n20362 & n20364 ) ;
  assign n20366 = n20365 ^ n2518 ^ 1'b0 ;
  assign n20367 = ~n20361 & n20366 ;
  assign n20369 = n20368 ^ n20367 ^ 1'b0 ;
  assign n20370 = n20369 ^ n18800 ^ 1'b0 ;
  assign n20371 = n9094 ^ n5038 ^ 1'b0 ;
  assign n20372 = n8112 & ~n20371 ;
  assign n20373 = n4267 & n13789 ;
  assign n20374 = n9646 & n20373 ;
  assign n20375 = ~n5143 & n14838 ;
  assign n20376 = n1349 | n20375 ;
  assign n20377 = n4914 & ~n14930 ;
  assign n20378 = n6456 ^ n2089 ^ 1'b0 ;
  assign n20379 = n2282 & n19207 ;
  assign n20380 = n9281 | n20379 ;
  assign n20381 = n8210 ^ n3825 ^ 1'b0 ;
  assign n20382 = n13154 ^ n6177 ^ 1'b0 ;
  assign n20383 = ~n12742 & n20382 ;
  assign n20384 = n16098 ^ n11296 ^ n3688 ;
  assign n20385 = ~n14292 & n19522 ;
  assign n20386 = n20385 ^ n12124 ^ 1'b0 ;
  assign n20387 = n17939 | n20386 ;
  assign n20388 = ~n2788 & n4447 ;
  assign n20389 = n14462 ^ n7350 ^ 1'b0 ;
  assign n20390 = n20389 ^ n635 ^ 1'b0 ;
  assign n20391 = ~n5456 & n20390 ;
  assign n20392 = ~n14661 & n20391 ;
  assign n20393 = n6941 | n18082 ;
  assign n20394 = ~n5990 & n20393 ;
  assign n20395 = n17664 ^ x122 ^ 1'b0 ;
  assign n20396 = n3831 ^ n2595 ^ 1'b0 ;
  assign n20398 = n16291 ^ n1999 ^ 1'b0 ;
  assign n20399 = n6057 & n20398 ;
  assign n20397 = ~n1397 & n12442 ;
  assign n20400 = n20399 ^ n20397 ^ 1'b0 ;
  assign n20401 = n1203 | n20400 ;
  assign n20402 = n6321 & ~n20401 ;
  assign n20403 = n17272 ^ n8980 ^ 1'b0 ;
  assign n20404 = ~n20402 & n20403 ;
  assign n20405 = n6306 ^ n5221 ^ 1'b0 ;
  assign n20407 = n9587 & n14222 ;
  assign n20406 = n9336 ^ n911 ^ 1'b0 ;
  assign n20408 = n20407 ^ n20406 ^ n7421 ;
  assign n20410 = n15711 ^ n393 ^ 1'b0 ;
  assign n20409 = n15189 | n15349 ;
  assign n20411 = n20410 ^ n20409 ^ 1'b0 ;
  assign n20412 = n19327 ^ n8714 ^ 1'b0 ;
  assign n20413 = n779 | n20412 ;
  assign n20417 = n2434 & n7378 ;
  assign n20418 = n8736 & n20417 ;
  assign n20419 = n2330 | n20418 ;
  assign n20420 = n20419 ^ n1956 ^ 1'b0 ;
  assign n20414 = ~n7150 & n8633 ;
  assign n20415 = n3038 & n20414 ;
  assign n20416 = n10517 & ~n20415 ;
  assign n20421 = n20420 ^ n20416 ^ n6398 ;
  assign n20422 = n1404 & ~n9302 ;
  assign n20423 = n20422 ^ n11720 ^ 1'b0 ;
  assign n20424 = n1319 & n13613 ;
  assign n20425 = n19375 & n20424 ;
  assign n20426 = n9595 ^ n865 ^ 1'b0 ;
  assign n20427 = ~n20425 & n20426 ;
  assign n20428 = n5216 & ~n7596 ;
  assign n20429 = ~n1980 & n20428 ;
  assign n20430 = n8698 | n20429 ;
  assign n20431 = n20430 ^ n10825 ^ 1'b0 ;
  assign n20433 = ( ~n9016 & n10899 ) | ( ~n9016 & n13124 ) | ( n10899 & n13124 ) ;
  assign n20432 = ~n1956 & n2116 ;
  assign n20434 = n20433 ^ n20432 ^ 1'b0 ;
  assign n20435 = n16010 ^ n1875 ^ 1'b0 ;
  assign n20436 = ~n6040 & n20435 ;
  assign n20437 = n20436 ^ n10914 ^ 1'b0 ;
  assign n20438 = n12104 ^ n10180 ^ 1'b0 ;
  assign n20439 = x177 & n20438 ;
  assign n20440 = n1875 | n11967 ;
  assign n20441 = n1443 | n6525 ;
  assign n20442 = n432 | n5849 ;
  assign n20443 = ( n20168 & ~n20441 ) | ( n20168 & n20442 ) | ( ~n20441 & n20442 ) ;
  assign n20444 = n10801 & ~n12479 ;
  assign n20445 = ~n8941 & n20444 ;
  assign n20446 = n1891 & n20445 ;
  assign n20447 = n5459 ^ n1402 ^ 1'b0 ;
  assign n20448 = n20447 ^ n11770 ^ 1'b0 ;
  assign n20449 = ~n2029 & n4331 ;
  assign n20450 = n10541 | n12007 ;
  assign n20451 = n20450 ^ n20177 ^ 1'b0 ;
  assign n20452 = n1694 & ~n2803 ;
  assign n20453 = ( ~n5197 & n19386 ) | ( ~n5197 & n20452 ) | ( n19386 & n20452 ) ;
  assign n20457 = n18637 ^ n8452 ^ 1'b0 ;
  assign n20458 = n579 | n20457 ;
  assign n20454 = n3672 & ~n17643 ;
  assign n20455 = n20454 ^ n9687 ^ 1'b0 ;
  assign n20456 = ( n825 & n5625 ) | ( n825 & n20455 ) | ( n5625 & n20455 ) ;
  assign n20459 = n20458 ^ n20456 ^ n12736 ;
  assign n20460 = n5180 & n5646 ;
  assign n20461 = n20460 ^ n3806 ^ 1'b0 ;
  assign n20462 = n18028 & n20461 ;
  assign n20463 = n5659 & n9956 ;
  assign n20464 = n5840 & ~n10297 ;
  assign n20465 = ~x194 & n12426 ;
  assign n20466 = n7804 ^ n5602 ^ 1'b0 ;
  assign n20467 = n20109 ^ n8977 ^ 1'b0 ;
  assign n20468 = n12485 & n20467 ;
  assign n20469 = n10569 ^ n9258 ^ 1'b0 ;
  assign n20470 = n3042 & ~n20469 ;
  assign n20474 = x141 & n4085 ;
  assign n20472 = n19990 ^ n6378 ^ 1'b0 ;
  assign n20473 = ~n7558 & n20472 ;
  assign n20475 = n20474 ^ n20473 ^ n5785 ;
  assign n20471 = ~n752 & n4331 ;
  assign n20476 = n20475 ^ n20471 ^ 1'b0 ;
  assign n20477 = ( n4958 & n12698 ) | ( n4958 & n19959 ) | ( n12698 & n19959 ) ;
  assign n20479 = n12400 ^ n579 ^ 1'b0 ;
  assign n20480 = n5531 & ~n20479 ;
  assign n20478 = n558 & n19277 ;
  assign n20481 = n20480 ^ n20478 ^ n20244 ;
  assign n20482 = n10556 | n11072 ;
  assign n20483 = n20481 & ~n20482 ;
  assign n20484 = n15343 ^ n15285 ^ 1'b0 ;
  assign n20485 = n15105 & n20484 ;
  assign n20486 = n3828 | n20485 ;
  assign n20487 = n15235 ^ n3060 ^ n2936 ;
  assign n20488 = n4598 ^ n631 ^ 1'b0 ;
  assign n20489 = n4132 & ~n20488 ;
  assign n20490 = n12085 & n20489 ;
  assign n20491 = n20490 ^ n2863 ^ 1'b0 ;
  assign n20492 = n16008 & n20491 ;
  assign n20494 = x16 & ~n2703 ;
  assign n20493 = ~n294 & n1129 ;
  assign n20495 = n20494 ^ n20493 ^ 1'b0 ;
  assign n20496 = ~n5004 & n17818 ;
  assign n20497 = n11525 & n20496 ;
  assign n20498 = n10991 | n20497 ;
  assign n20499 = n5049 | n20498 ;
  assign n20500 = ~n905 & n20499 ;
  assign n20501 = ~n10966 & n12161 ;
  assign n20502 = n854 & n18310 ;
  assign n20503 = n4267 & ~n11354 ;
  assign n20504 = n20503 ^ n17562 ^ n3462 ;
  assign n20509 = n9878 ^ n8174 ^ 1'b0 ;
  assign n20510 = ~n7811 & n20509 ;
  assign n20505 = n8417 | n12677 ;
  assign n20506 = n20505 ^ n3656 ^ n1391 ;
  assign n20507 = n16801 ^ n2513 ^ 1'b0 ;
  assign n20508 = ~n20506 & n20507 ;
  assign n20511 = n20510 ^ n20508 ^ 1'b0 ;
  assign n20512 = ~n3985 & n19380 ;
  assign n20513 = ~n1204 & n3335 ;
  assign n20514 = ~n3604 & n20513 ;
  assign n20515 = n518 & n15559 ;
  assign n20516 = n12622 & ~n16775 ;
  assign n20517 = n20516 ^ n8200 ^ n3684 ;
  assign n20518 = n20517 ^ n12649 ^ 1'b0 ;
  assign n20519 = n8996 & ~n20518 ;
  assign n20520 = ~n924 & n9002 ;
  assign n20521 = n9273 ^ n5025 ^ 1'b0 ;
  assign n20522 = n20520 | n20521 ;
  assign n20523 = n3678 ^ n2227 ^ 1'b0 ;
  assign n20524 = n13791 & ~n15290 ;
  assign n20525 = x107 | n8983 ;
  assign n20526 = n5646 | n20525 ;
  assign n20527 = ( n3012 & n16624 ) | ( n3012 & ~n20526 ) | ( n16624 & ~n20526 ) ;
  assign n20528 = ~n10043 & n20527 ;
  assign n20529 = ~n20524 & n20528 ;
  assign n20530 = n12627 & n12802 ;
  assign n20531 = n19106 ^ n9696 ^ n9216 ;
  assign n20532 = ~n2367 & n16285 ;
  assign n20533 = n20532 ^ n4424 ^ 1'b0 ;
  assign n20534 = n20533 ^ n9568 ^ 1'b0 ;
  assign n20535 = n5398 & ~n20534 ;
  assign n20536 = n10944 & n20535 ;
  assign n20537 = n17396 | n20536 ;
  assign n20538 = n20531 & ~n20537 ;
  assign n20541 = n1167 & n2204 ;
  assign n20542 = ~n1486 & n20541 ;
  assign n20543 = ~n9680 & n20542 ;
  assign n20539 = ~n3139 & n5788 ;
  assign n20540 = n724 & n20539 ;
  assign n20544 = n20543 ^ n20540 ^ 1'b0 ;
  assign n20545 = ( n3122 & ~n8446 ) | ( n3122 & n16327 ) | ( ~n8446 & n16327 ) ;
  assign n20546 = n8801 & ~n13711 ;
  assign n20547 = n20546 ^ n15503 ^ n4416 ;
  assign n20548 = n20547 ^ n1923 ^ 1'b0 ;
  assign n20549 = ( n845 & ~n5973 ) | ( n845 & n9072 ) | ( ~n5973 & n9072 ) ;
  assign n20550 = n2239 & n20549 ;
  assign n20551 = n20550 ^ n5104 ^ 1'b0 ;
  assign n20552 = n3900 & ~n12574 ;
  assign n20553 = ~n608 & n11879 ;
  assign n20554 = n20553 ^ n786 ^ 1'b0 ;
  assign n20555 = n5806 | n20554 ;
  assign n20556 = n20552 | n20555 ;
  assign n20557 = ~n2378 & n3458 ;
  assign n20558 = ~n2668 & n20557 ;
  assign n20559 = x224 ^ x124 ^ x76 ;
  assign n20560 = n20558 & ~n20559 ;
  assign n20561 = ( ~n5150 & n10477 ) | ( ~n5150 & n19306 ) | ( n10477 & n19306 ) ;
  assign n20562 = ( n378 & ~n7855 ) | ( n378 & n14543 ) | ( ~n7855 & n14543 ) ;
  assign n20563 = n14846 ^ n12721 ^ 1'b0 ;
  assign n20564 = n20562 & ~n20563 ;
  assign n20565 = n8455 | n13101 ;
  assign n20566 = n18404 ^ n5752 ^ 1'b0 ;
  assign n20567 = n20566 ^ n10291 ^ 1'b0 ;
  assign n20568 = n20565 & ~n20567 ;
  assign n20569 = ( n1037 & n2162 ) | ( n1037 & n16940 ) | ( n2162 & n16940 ) ;
  assign n20570 = ( x2 & n1712 ) | ( x2 & ~n12359 ) | ( n1712 & ~n12359 ) ;
  assign n20571 = n5626 ^ n948 ^ 1'b0 ;
  assign n20572 = n6166 ^ n2901 ^ 1'b0 ;
  assign n20573 = n6649 & ~n20572 ;
  assign n20574 = n17129 ^ n13461 ^ 1'b0 ;
  assign n20575 = n20573 & n20574 ;
  assign n20576 = n10766 ^ n7000 ^ 1'b0 ;
  assign n20577 = ~n4997 & n20576 ;
  assign n20578 = x247 & n20577 ;
  assign n20579 = n2039 & n15672 ;
  assign n20580 = n1219 & n4010 ;
  assign n20581 = n6964 | n20580 ;
  assign n20582 = n20581 ^ n3352 ^ 1'b0 ;
  assign n20583 = n20582 ^ n9147 ^ 1'b0 ;
  assign n20584 = n8544 ^ x133 ^ 1'b0 ;
  assign n20585 = ~n2716 & n20584 ;
  assign n20586 = ~n1324 & n20585 ;
  assign n20588 = n5326 | n8695 ;
  assign n20589 = n20588 ^ n17156 ^ 1'b0 ;
  assign n20587 = n19940 & ~n20474 ;
  assign n20590 = n20589 ^ n20587 ^ 1'b0 ;
  assign n20591 = n2045 & n13415 ;
  assign n20592 = n20591 ^ n2378 ^ 1'b0 ;
  assign n20593 = n20592 ^ n737 ^ 1'b0 ;
  assign n20594 = n938 | n20593 ;
  assign n20595 = n19211 ^ n16108 ^ 1'b0 ;
  assign n20596 = n14866 & ~n20595 ;
  assign n20597 = n1733 ^ x185 ^ 1'b0 ;
  assign n20598 = n5560 & ~n20597 ;
  assign n20599 = n8143 ^ n2743 ^ 1'b0 ;
  assign n20600 = n20599 ^ n5713 ^ 1'b0 ;
  assign n20601 = n20598 & ~n20600 ;
  assign n20602 = n4553 | n18786 ;
  assign n20603 = n15962 | n20602 ;
  assign n20604 = n958 & n5103 ;
  assign n20605 = ~n3690 & n20604 ;
  assign n20606 = n9773 ^ n8864 ^ 1'b0 ;
  assign n20607 = x117 & ~n7743 ;
  assign n20608 = n20607 ^ n7271 ^ 1'b0 ;
  assign n20609 = n5208 | n20608 ;
  assign n20610 = n18462 & n20609 ;
  assign n20611 = n5020 & n20610 ;
  assign n20612 = n5556 ^ n5066 ^ 1'b0 ;
  assign n20613 = n17756 | n20612 ;
  assign n20614 = ( n264 & ~n4296 ) | ( n264 & n20613 ) | ( ~n4296 & n20613 ) ;
  assign n20615 = ~n9971 & n10449 ;
  assign n20616 = n20614 & n20615 ;
  assign n20617 = n11186 ^ n8693 ^ 1'b0 ;
  assign n20618 = n1062 | n6088 ;
  assign n20619 = n10176 & ~n20618 ;
  assign n20620 = n18761 | n20619 ;
  assign n20621 = n20620 ^ n18892 ^ 1'b0 ;
  assign n20622 = n20621 ^ n10752 ^ 1'b0 ;
  assign n20623 = n8950 & ~n20622 ;
  assign n20624 = n8772 | n16280 ;
  assign n20625 = n15678 & ~n20624 ;
  assign n20626 = x6 & ~n20625 ;
  assign n20627 = ~n992 & n9951 ;
  assign n20628 = n20627 ^ n9993 ^ 1'b0 ;
  assign n20629 = n7964 ^ n2887 ^ 1'b0 ;
  assign n20630 = ( ~n4890 & n8336 ) | ( ~n4890 & n20629 ) | ( n8336 & n20629 ) ;
  assign n20631 = ( n1829 & n20628 ) | ( n1829 & ~n20630 ) | ( n20628 & ~n20630 ) ;
  assign n20632 = n4254 & ~n15345 ;
  assign n20633 = n16846 & n20632 ;
  assign n20634 = n20631 | n20633 ;
  assign n20635 = n20634 ^ n11994 ^ 1'b0 ;
  assign n20636 = n2506 | n9359 ;
  assign n20637 = n20636 ^ n7397 ^ 1'b0 ;
  assign n20638 = n20637 ^ n6514 ^ 1'b0 ;
  assign n20639 = n20638 ^ n20081 ^ 1'b0 ;
  assign n20640 = n11603 ^ n10606 ^ 1'b0 ;
  assign n20641 = n10441 ^ n7421 ^ 1'b0 ;
  assign n20642 = n20640 & n20641 ;
  assign n20643 = n18664 ^ n3754 ^ 1'b0 ;
  assign n20644 = ~n13695 & n20643 ;
  assign n20645 = n20644 ^ x188 ^ 1'b0 ;
  assign n20646 = n11945 & ~n14769 ;
  assign n20647 = n3589 ^ n3054 ^ n2980 ;
  assign n20648 = n20647 ^ n14533 ^ n6122 ;
  assign n20649 = n20648 ^ n2961 ^ 1'b0 ;
  assign n20650 = n5665 | n10900 ;
  assign n20651 = n3372 | n20650 ;
  assign n20652 = ~n12679 & n20120 ;
  assign n20653 = n10448 ^ n8159 ^ n416 ;
  assign n20654 = n6902 ^ n1208 ^ 1'b0 ;
  assign n20655 = n20653 & n20654 ;
  assign n20656 = ~n8530 & n10168 ;
  assign n20657 = n20656 ^ n20257 ^ 1'b0 ;
  assign n20658 = n4860 | n9276 ;
  assign n20659 = n481 & ~n20658 ;
  assign n20660 = n20659 ^ x248 ^ 1'b0 ;
  assign n20661 = n20657 & n20660 ;
  assign n20662 = n3131 & n9996 ;
  assign n20663 = ~n1133 & n20662 ;
  assign n20664 = n1123 & ~n20663 ;
  assign n20665 = ~n15507 & n20664 ;
  assign n20666 = n20665 ^ n20324 ^ 1'b0 ;
  assign n20667 = n11211 ^ n1741 ^ 1'b0 ;
  assign n20668 = n7511 & ~n7940 ;
  assign n20669 = n20668 ^ n1557 ^ 1'b0 ;
  assign n20670 = n18050 ^ n8594 ^ 1'b0 ;
  assign n20671 = n18190 ^ n17386 ^ n12155 ;
  assign n20672 = n19718 & n20671 ;
  assign n20673 = x45 & n2978 ;
  assign n20674 = n4931 ^ n3653 ^ 1'b0 ;
  assign n20675 = n20673 & ~n20674 ;
  assign n20676 = ~n2993 & n20675 ;
  assign n20677 = ~n20675 & n20676 ;
  assign n20678 = n3696 & ~n20677 ;
  assign n20679 = ~n10360 & n12593 ;
  assign n20680 = n12412 ^ n11353 ^ 1'b0 ;
  assign n20681 = n1590 & ~n19783 ;
  assign n20683 = n11296 & ~n19714 ;
  assign n20682 = n15303 & ~n15952 ;
  assign n20684 = n20683 ^ n20682 ^ 1'b0 ;
  assign n20685 = n5513 & n7219 ;
  assign n20686 = n20685 ^ n3189 ^ 1'b0 ;
  assign n20687 = n8250 | n20686 ;
  assign n20688 = n20687 ^ n3149 ^ 1'b0 ;
  assign n20689 = ~n2870 & n20688 ;
  assign n20690 = n20689 ^ n4852 ^ 1'b0 ;
  assign n20691 = ~n6506 & n11034 ;
  assign n20692 = n4306 ^ x129 ^ 1'b0 ;
  assign n20693 = ( n11615 & n14423 ) | ( n11615 & ~n16967 ) | ( n14423 & ~n16967 ) ;
  assign n20694 = n293 | n20693 ;
  assign n20695 = n20694 ^ n20051 ^ 1'b0 ;
  assign n20696 = ~n2029 & n3011 ;
  assign n20697 = ~n4226 & n8108 ;
  assign n20698 = ~n20696 & n20697 ;
  assign n20699 = n11201 ^ n1077 ^ 1'b0 ;
  assign n20700 = n15650 & n20699 ;
  assign n20701 = ( n11211 & n12428 ) | ( n11211 & ~n12494 ) | ( n12428 & ~n12494 ) ;
  assign n20702 = n8931 ^ n2496 ^ 1'b0 ;
  assign n20703 = n20702 ^ n10006 ^ n9001 ;
  assign n20704 = n7307 & ~n13993 ;
  assign n20705 = n20703 & n20704 ;
  assign n20706 = n20701 | n20705 ;
  assign n20707 = n20706 ^ n451 ^ 1'b0 ;
  assign n20708 = n9009 & ~n10843 ;
  assign n20709 = n20708 ^ n4837 ^ 1'b0 ;
  assign n20710 = n20709 ^ n16573 ^ n12552 ;
  assign n20711 = n9873 | n13953 ;
  assign n20712 = n20711 ^ n12809 ^ 1'b0 ;
  assign n20713 = n7775 ^ n7511 ^ 1'b0 ;
  assign n20714 = n3096 & ~n20713 ;
  assign n20715 = n5540 ^ n2335 ^ 1'b0 ;
  assign n20719 = n8926 & n12754 ;
  assign n20720 = ~n3203 & n20719 ;
  assign n20716 = x1 & ~n486 ;
  assign n20717 = n7513 & n7945 ;
  assign n20718 = n20716 & n20717 ;
  assign n20721 = n20720 ^ n20718 ^ n4393 ;
  assign n20723 = ~n6042 & n16885 ;
  assign n20724 = n20723 ^ n5734 ^ 1'b0 ;
  assign n20725 = n1561 & n20724 ;
  assign n20722 = n9146 & n14794 ;
  assign n20726 = n20725 ^ n20722 ^ 1'b0 ;
  assign n20727 = n6299 ^ n2743 ^ 1'b0 ;
  assign n20728 = n16203 ^ n8792 ^ 1'b0 ;
  assign n20730 = x130 & n7473 ;
  assign n20729 = n3539 | n15596 ;
  assign n20731 = n20730 ^ n20729 ^ 1'b0 ;
  assign n20736 = n6066 ^ n4062 ^ 1'b0 ;
  assign n20737 = ~n5704 & n20736 ;
  assign n20733 = ~n3332 & n7736 ;
  assign n20734 = n2264 & n20733 ;
  assign n20732 = n9096 | n16871 ;
  assign n20735 = n20734 ^ n20732 ^ 1'b0 ;
  assign n20738 = n20737 ^ n20735 ^ n11157 ;
  assign n20739 = n7935 & ~n20738 ;
  assign n20740 = n8731 | n20690 ;
  assign n20741 = n20740 ^ x69 ^ 1'b0 ;
  assign n20743 = n6424 | n8253 ;
  assign n20744 = ( n16221 & n20160 ) | ( n16221 & n20743 ) | ( n20160 & n20743 ) ;
  assign n20742 = n13901 & ~n15733 ;
  assign n20745 = n20744 ^ n20742 ^ n14509 ;
  assign n20746 = n13651 ^ n6238 ^ 1'b0 ;
  assign n20747 = ~n5036 & n20746 ;
  assign n20748 = ( n5594 & n15712 ) | ( n5594 & n20747 ) | ( n15712 & n20747 ) ;
  assign n20749 = n6688 & n7388 ;
  assign n20750 = n20748 & n20749 ;
  assign n20751 = ~n964 & n4124 ;
  assign n20752 = ~n12638 & n20751 ;
  assign n20753 = n8519 & ~n20752 ;
  assign n20754 = n4189 | n5403 ;
  assign n20755 = n20754 ^ n11536 ^ 1'b0 ;
  assign n20756 = n11053 ^ n3012 ^ 1'b0 ;
  assign n20757 = ~n15213 & n20756 ;
  assign n20758 = n6812 ^ n6151 ^ 1'b0 ;
  assign n20759 = n6058 & ~n20758 ;
  assign n20760 = ~n20619 & n20759 ;
  assign n20761 = n20760 ^ n15555 ^ 1'b0 ;
  assign n20762 = ~n792 & n14792 ;
  assign n20763 = n7789 ^ n5385 ^ 1'b0 ;
  assign n20764 = n14972 & ~n20763 ;
  assign n20765 = n20764 ^ n1458 ^ 1'b0 ;
  assign n20766 = x169 | n20765 ;
  assign n20767 = n20766 ^ n19893 ^ 1'b0 ;
  assign n20768 = n3958 & n7602 ;
  assign n20769 = n20768 ^ n3102 ^ 1'b0 ;
  assign n20770 = n20769 ^ n932 ^ 1'b0 ;
  assign n20771 = n4634 & n20770 ;
  assign n20772 = ( n3478 & n3614 ) | ( n3478 & n19465 ) | ( n3614 & n19465 ) ;
  assign n20773 = ( n3231 & ~n7416 ) | ( n3231 & n20772 ) | ( ~n7416 & n20772 ) ;
  assign n20774 = ( n7143 & ~n15852 ) | ( n7143 & n20773 ) | ( ~n15852 & n20773 ) ;
  assign n20775 = n1565 & ~n6811 ;
  assign n20776 = n8415 & n20775 ;
  assign n20777 = n20776 ^ n14302 ^ 1'b0 ;
  assign n20778 = n9627 | n20777 ;
  assign n20779 = n13586 ^ n11981 ^ 1'b0 ;
  assign n20782 = ~n1674 & n3210 ;
  assign n20783 = n1105 & n20782 ;
  assign n20780 = n2343 | n7907 ;
  assign n20781 = ~n624 & n20780 ;
  assign n20784 = n20783 ^ n20781 ^ 1'b0 ;
  assign n20785 = n2142 | n5933 ;
  assign n20786 = n9543 & ~n20785 ;
  assign n20787 = n1440 | n20786 ;
  assign n20788 = n9496 & ~n20787 ;
  assign n20789 = n13706 ^ n5474 ^ 1'b0 ;
  assign n20790 = n18288 ^ n16533 ^ 1'b0 ;
  assign n20791 = n10557 & n20790 ;
  assign n20792 = n20791 ^ n3878 ^ 1'b0 ;
  assign n20793 = n4084 ^ n3942 ^ 1'b0 ;
  assign n20794 = n14466 | n20793 ;
  assign n20795 = n20579 ^ n1137 ^ 1'b0 ;
  assign n20796 = n10041 ^ n5170 ^ 1'b0 ;
  assign n20797 = n13390 & n20796 ;
  assign n20798 = n3930 & ~n14964 ;
  assign n20799 = n16360 & n20798 ;
  assign n20800 = n12708 ^ n1968 ^ 1'b0 ;
  assign n20801 = n20799 | n20800 ;
  assign n20802 = n20801 ^ n8380 ^ 1'b0 ;
  assign n20803 = n8228 ^ n7448 ^ 1'b0 ;
  assign n20804 = n18661 ^ n7458 ^ 1'b0 ;
  assign n20805 = n7547 & ~n20804 ;
  assign n20806 = n8164 & ~n14232 ;
  assign n20807 = n5628 & ~n20759 ;
  assign n20808 = n10294 & n10917 ;
  assign n20809 = n20808 ^ n15733 ^ 1'b0 ;
  assign n20810 = n5825 & ~n20809 ;
  assign n20811 = n12314 | n16271 ;
  assign n20812 = n7520 ^ n518 ^ 1'b0 ;
  assign n20813 = ~n13373 & n20812 ;
  assign n20814 = n20813 ^ n4325 ^ 1'b0 ;
  assign n20815 = ~n13452 & n20814 ;
  assign n20816 = n2812 | n12415 ;
  assign n20817 = ( ~n1705 & n1989 ) | ( ~n1705 & n7706 ) | ( n1989 & n7706 ) ;
  assign n20818 = n20817 ^ x201 ^ 1'b0 ;
  assign n20819 = n3851 | n20818 ;
  assign n20820 = n4447 & ~n5650 ;
  assign n20821 = n20820 ^ n1309 ^ 1'b0 ;
  assign n20822 = n20819 & n20821 ;
  assign n20823 = n3410 | n4649 ;
  assign n20824 = n20823 ^ n15093 ^ 1'b0 ;
  assign n20825 = n17051 ^ n2050 ^ 1'b0 ;
  assign n20826 = n18960 | n20825 ;
  assign n20827 = n4196 & ~n12427 ;
  assign n20828 = n5118 & ~n8699 ;
  assign n20829 = n6879 & n20828 ;
  assign n20830 = x122 | n20829 ;
  assign n20832 = n7069 & ~n14838 ;
  assign n20831 = n11140 & n11677 ;
  assign n20833 = n20832 ^ n20831 ^ 1'b0 ;
  assign n20834 = ( ~n1030 & n20830 ) | ( ~n1030 & n20833 ) | ( n20830 & n20833 ) ;
  assign n20835 = n11511 ^ n1272 ^ 1'b0 ;
  assign n20836 = n20835 ^ n2148 ^ n710 ;
  assign n20837 = n3016 | n5205 ;
  assign n20838 = n931 | n20837 ;
  assign n20839 = n20838 ^ n8990 ^ 1'b0 ;
  assign n20840 = ~n11206 & n20839 ;
  assign n20841 = n8030 & n20442 ;
  assign n20842 = ~n328 & n20841 ;
  assign n20843 = n7884 ^ n483 ^ 1'b0 ;
  assign n20844 = n7689 ^ n4775 ^ 1'b0 ;
  assign n20845 = n14440 & n20844 ;
  assign n20846 = n13738 & ~n20845 ;
  assign n20847 = n12643 ^ n8614 ^ 1'b0 ;
  assign n20848 = n6812 & ~n19538 ;
  assign n20849 = ~n18507 & n20848 ;
  assign n20850 = n842 | n8188 ;
  assign n20851 = n16533 & ~n20850 ;
  assign n20852 = n3586 & ~n20851 ;
  assign n20853 = ~n16923 & n20852 ;
  assign n20854 = n20629 | n20853 ;
  assign n20855 = n20854 ^ n17537 ^ n5195 ;
  assign n20856 = n6058 | n19415 ;
  assign n20857 = n20856 ^ n10475 ^ 1'b0 ;
  assign n20858 = n1632 ^ n722 ^ 1'b0 ;
  assign n20859 = ~n5127 & n18014 ;
  assign n20860 = n13547 & ~n20859 ;
  assign n20861 = ~n5300 & n20860 ;
  assign n20862 = n6979 & n17415 ;
  assign n20863 = ~n1726 & n20862 ;
  assign n20864 = n20647 ^ n12653 ^ 1'b0 ;
  assign n20865 = ~n10101 & n20450 ;
  assign n20866 = n20865 ^ n16778 ^ 1'b0 ;
  assign n20867 = n18306 & n20866 ;
  assign n20868 = n17787 ^ n8210 ^ n3710 ;
  assign n20869 = ~n6311 & n9452 ;
  assign n20870 = n14596 ^ n13912 ^ 1'b0 ;
  assign n20871 = n9012 ^ n1002 ^ n376 ;
  assign n20872 = ~n5924 & n20871 ;
  assign n20873 = n8202 & n10148 ;
  assign n20874 = n18596 & n20873 ;
  assign n20875 = ~n10134 & n12022 ;
  assign n20876 = n20875 ^ n8658 ^ 1'b0 ;
  assign n20877 = n14134 | n20876 ;
  assign n20878 = n5927 ^ n552 ^ 1'b0 ;
  assign n20879 = n3754 | n10451 ;
  assign n20880 = n10451 & ~n20879 ;
  assign n20881 = n2234 | n20880 ;
  assign n20882 = n20880 & ~n20881 ;
  assign n20883 = n5700 | n20882 ;
  assign n20884 = n5700 & ~n20883 ;
  assign n20885 = n6847 & ~n20884 ;
  assign n20886 = ~n20878 & n20885 ;
  assign n20887 = n2705 & ~n3407 ;
  assign n20888 = n20887 ^ n5780 ^ 1'b0 ;
  assign n20889 = n20888 ^ n18268 ^ 1'b0 ;
  assign n20890 = ~n9747 & n20889 ;
  assign n20891 = n20890 ^ n13626 ^ 1'b0 ;
  assign n20892 = n20891 ^ n14669 ^ n7884 ;
  assign n20893 = ~n12445 & n17940 ;
  assign n20894 = n20893 ^ n8907 ^ n8011 ;
  assign n20895 = n19211 ^ n7404 ^ 1'b0 ;
  assign n20896 = n5452 | n20895 ;
  assign n20897 = n12861 & ~n20896 ;
  assign n20898 = n20897 ^ n18773 ^ 1'b0 ;
  assign n20899 = ~n8566 & n17071 ;
  assign n20900 = n11919 & ~n19961 ;
  assign n20901 = n8837 & n19463 ;
  assign n20902 = n20901 ^ n417 ^ 1'b0 ;
  assign n20903 = x162 & n20902 ;
  assign n20904 = n8382 | n13385 ;
  assign n20905 = ~n10847 & n13630 ;
  assign n20906 = n14887 ^ n6731 ^ 1'b0 ;
  assign n20907 = n7912 & n10282 ;
  assign n20908 = n8605 & n20907 ;
  assign n20909 = n7223 ^ n1605 ^ 1'b0 ;
  assign n20910 = n2936 & n20909 ;
  assign n20911 = ~n20908 & n20910 ;
  assign n20912 = n20628 & n20911 ;
  assign n20913 = n13087 ^ n7906 ^ 1'b0 ;
  assign n20914 = ~n5309 & n20913 ;
  assign n20915 = ( n1153 & n7549 ) | ( n1153 & ~n20914 ) | ( n7549 & ~n20914 ) ;
  assign n20916 = ~n6811 & n20915 ;
  assign n20917 = n9938 | n17226 ;
  assign n20918 = n5286 | n20917 ;
  assign n20919 = n759 & n20918 ;
  assign n20920 = n20916 & n20919 ;
  assign n20921 = ~n2406 & n20920 ;
  assign n20922 = n9088 & ~n20921 ;
  assign n20923 = n20922 ^ n12730 ^ 1'b0 ;
  assign n20924 = n13163 ^ n1742 ^ 1'b0 ;
  assign n20926 = ~n3917 & n12969 ;
  assign n20927 = ~n2718 & n20926 ;
  assign n20925 = n2929 & n9218 ;
  assign n20928 = n20927 ^ n20925 ^ 1'b0 ;
  assign n20929 = n1392 | n20928 ;
  assign n20930 = n5169 ^ x244 ^ 1'b0 ;
  assign n20931 = n17029 & ~n20930 ;
  assign n20932 = n1662 & ~n1890 ;
  assign n20933 = n2909 & ~n20932 ;
  assign n20934 = n10048 & ~n20933 ;
  assign n20935 = ~n6572 & n20934 ;
  assign n20936 = n11739 & ~n20935 ;
  assign n20937 = n13643 & n20936 ;
  assign n20938 = n10284 | n20937 ;
  assign n20939 = n9695 | n20938 ;
  assign n20940 = ~n19711 & n20939 ;
  assign n20941 = n6271 ^ n2116 ^ 1'b0 ;
  assign n20942 = ~n11730 & n20941 ;
  assign n20943 = n9897 ^ n361 ^ 1'b0 ;
  assign n20944 = ~n2069 & n2622 ;
  assign n20945 = n12187 ^ x221 ^ 1'b0 ;
  assign n20946 = n20945 ^ n8191 ^ 1'b0 ;
  assign n20947 = ~n20944 & n20946 ;
  assign n20948 = ~n17958 & n20947 ;
  assign n20949 = n20948 ^ n1105 ^ 1'b0 ;
  assign n20952 = ( ~n991 & n6230 ) | ( ~n991 & n6731 ) | ( n6230 & n6731 ) ;
  assign n20950 = x200 & ~n17543 ;
  assign n20951 = n16059 & n20950 ;
  assign n20953 = n20952 ^ n20951 ^ 1'b0 ;
  assign n20954 = n8293 ^ n5142 ^ 1'b0 ;
  assign n20955 = n18502 ^ n16823 ^ 1'b0 ;
  assign n20956 = n294 & ~n7678 ;
  assign n20957 = ~n1664 & n20956 ;
  assign n20958 = n20957 ^ n7243 ^ 1'b0 ;
  assign n20959 = ~x6 & n451 ;
  assign n20960 = ~n862 & n20959 ;
  assign n20961 = n19594 | n20960 ;
  assign n20962 = n10869 ^ n2403 ^ 1'b0 ;
  assign n20963 = n8087 & n20962 ;
  assign n20964 = x70 & ~n6548 ;
  assign n20965 = n20964 ^ n2216 ^ 1'b0 ;
  assign n20966 = n18043 ^ n3012 ^ 1'b0 ;
  assign n20967 = n7174 & n20966 ;
  assign n20968 = n543 & ~n3620 ;
  assign n20969 = ~n10622 & n14029 ;
  assign n20970 = n7994 | n11443 ;
  assign n20971 = n20970 ^ n4210 ^ 1'b0 ;
  assign n20972 = n11044 ^ n6131 ^ 1'b0 ;
  assign n20973 = n9329 ^ n2789 ^ 1'b0 ;
  assign n20974 = n19145 & n20973 ;
  assign n20975 = n13469 & ~n20974 ;
  assign n20976 = ( ~n5497 & n6350 ) | ( ~n5497 & n9977 ) | ( n6350 & n9977 ) ;
  assign n20977 = n20976 ^ n16674 ^ n13673 ;
  assign n20978 = ~n8473 & n9722 ;
  assign n20979 = n20977 & n20978 ;
  assign n20980 = n4018 | n9622 ;
  assign n20981 = n4578 & ~n20980 ;
  assign n20982 = n14445 & ~n20981 ;
  assign n20983 = n16473 & n20982 ;
  assign n20984 = n671 & n10805 ;
  assign n20985 = x247 | n6295 ;
  assign n20986 = n6905 & ~n20985 ;
  assign n20987 = ( n4843 & n5525 ) | ( n4843 & n7501 ) | ( n5525 & n7501 ) ;
  assign n20988 = n20987 ^ x89 ^ 1'b0 ;
  assign n20989 = n18774 ^ n10454 ^ 1'b0 ;
  assign n20990 = ( n1725 & n5294 ) | ( n1725 & ~n7672 ) | ( n5294 & ~n7672 ) ;
  assign n20991 = ~n6603 & n20990 ;
  assign n20992 = n17635 ^ n3899 ^ 1'b0 ;
  assign n20993 = ~n8079 & n13834 ;
  assign n20994 = n20993 ^ n4585 ^ 1'b0 ;
  assign n20995 = n713 & n6340 ;
  assign n20996 = n3023 ^ n1753 ^ 1'b0 ;
  assign n20997 = n11320 ^ n3050 ^ x75 ;
  assign n20998 = n20997 ^ n10418 ^ 1'b0 ;
  assign n20999 = n14913 | n20998 ;
  assign n21000 = n1129 | n20999 ;
  assign n21001 = n15138 ^ n7290 ^ 1'b0 ;
  assign n21002 = n7382 & ~n21001 ;
  assign n21003 = n21002 ^ n5450 ^ 1'b0 ;
  assign n21004 = ( n370 & ~n3806 ) | ( n370 & n12030 ) | ( ~n3806 & n12030 ) ;
  assign n21005 = n3038 & ~n21004 ;
  assign n21006 = n12328 & n21005 ;
  assign n21007 = n16545 | n21006 ;
  assign n21008 = ~n6106 & n21007 ;
  assign n21009 = ~n8632 & n14557 ;
  assign n21010 = n21009 ^ n11547 ^ n9649 ;
  assign n21011 = n20916 ^ n6270 ^ 1'b0 ;
  assign n21012 = n4871 | n20932 ;
  assign n21013 = n4997 & ~n21012 ;
  assign n21014 = n5688 ^ n2890 ^ 1'b0 ;
  assign n21015 = n1851 & n21014 ;
  assign n21016 = n946 & n21015 ;
  assign n21017 = n14227 ^ n1343 ^ 1'b0 ;
  assign n21018 = ~n9986 & n21017 ;
  assign n21019 = n19340 ^ n16214 ^ 1'b0 ;
  assign n21020 = n21018 & ~n21019 ;
  assign n21021 = ~n8571 & n11874 ;
  assign n21022 = n7463 & n21021 ;
  assign n21023 = n19230 & n21022 ;
  assign n21024 = n1496 & n21023 ;
  assign n21025 = ( ~n5118 & n6985 ) | ( ~n5118 & n17153 ) | ( n6985 & n17153 ) ;
  assign n21026 = n9584 & n9992 ;
  assign n21027 = n8002 & n10706 ;
  assign n21028 = n21027 ^ n12956 ^ 1'b0 ;
  assign n21029 = ~n21026 & n21028 ;
  assign n21031 = n18953 ^ n17263 ^ 1'b0 ;
  assign n21030 = n6051 ^ x46 ^ 1'b0 ;
  assign n21032 = n21031 ^ n21030 ^ n9291 ;
  assign n21033 = n21032 ^ n17949 ^ 1'b0 ;
  assign n21034 = n20791 ^ n16087 ^ n11834 ;
  assign n21035 = n2833 & ~n6305 ;
  assign n21036 = n11784 ^ n5342 ^ 1'b0 ;
  assign n21037 = n10048 & ~n21036 ;
  assign n21038 = n13470 ^ n8396 ^ 1'b0 ;
  assign n21039 = n21038 ^ n12700 ^ 1'b0 ;
  assign n21040 = n5188 ^ n880 ^ 1'b0 ;
  assign n21041 = n4255 | n21040 ;
  assign n21042 = n21041 ^ n13845 ^ n12887 ;
  assign n21043 = ~n19465 & n20427 ;
  assign n21044 = ~n21042 & n21043 ;
  assign n21045 = n6849 & ~n19372 ;
  assign n21046 = n21045 ^ n3411 ^ 1'b0 ;
  assign n21049 = ~n1347 & n6616 ;
  assign n21050 = n21049 ^ n6359 ^ 1'b0 ;
  assign n21047 = n1116 | n2697 ;
  assign n21048 = n21047 ^ n6091 ^ 1'b0 ;
  assign n21051 = n21050 ^ n21048 ^ 1'b0 ;
  assign n21056 = n14256 & n14319 ;
  assign n21057 = ~n4608 & n21056 ;
  assign n21055 = ~n3788 & n7482 ;
  assign n21052 = n320 | n10142 ;
  assign n21053 = n6127 & ~n21052 ;
  assign n21054 = n21053 ^ n12190 ^ 1'b0 ;
  assign n21058 = n21057 ^ n21055 ^ n21054 ;
  assign n21059 = n18768 ^ n3508 ^ 1'b0 ;
  assign n21060 = ~n2320 & n19559 ;
  assign n21061 = n7260 & ~n14758 ;
  assign n21062 = n5182 & n21061 ;
  assign n21063 = ~n1554 & n2856 ;
  assign n21064 = n21063 ^ n13812 ^ 1'b0 ;
  assign n21065 = n13151 ^ n3325 ^ 1'b0 ;
  assign n21066 = n8614 | n21065 ;
  assign n21067 = n21066 ^ n10858 ^ 1'b0 ;
  assign n21068 = n21067 ^ n14375 ^ x195 ;
  assign n21069 = n14118 ^ n10489 ^ n2447 ;
  assign n21070 = n21069 ^ n11930 ^ 1'b0 ;
  assign n21071 = n8277 & n21070 ;
  assign n21072 = n19963 ^ n1854 ^ n738 ;
  assign n21073 = n723 & ~n21072 ;
  assign n21074 = ~n20340 & n21073 ;
  assign n21075 = n501 & ~n20703 ;
  assign n21076 = n21075 ^ n7846 ^ 1'b0 ;
  assign n21077 = n18466 ^ n16779 ^ n14083 ;
  assign n21078 = n16615 ^ n3320 ^ 1'b0 ;
  assign n21079 = ~n10961 & n15331 ;
  assign n21080 = n21079 ^ n6412 ^ 1'b0 ;
  assign n21081 = ( x147 & n9808 ) | ( x147 & n14412 ) | ( n9808 & n14412 ) ;
  assign n21082 = ~n2306 & n20186 ;
  assign n21083 = ~n8904 & n21082 ;
  assign n21084 = ( x159 & n882 ) | ( x159 & n8591 ) | ( n882 & n8591 ) ;
  assign n21085 = n14246 & n21084 ;
  assign n21086 = x53 & n15304 ;
  assign n21087 = ~n7065 & n10124 ;
  assign n21088 = n21087 ^ n13116 ^ 1'b0 ;
  assign n21089 = ( ~n11807 & n20146 ) | ( ~n11807 & n21088 ) | ( n20146 & n21088 ) ;
  assign n21090 = ~n1878 & n11149 ;
  assign n21091 = n11112 ^ n9659 ^ 1'b0 ;
  assign n21092 = n310 & n21091 ;
  assign n21093 = ~n21090 & n21092 ;
  assign n21095 = n498 | n5404 ;
  assign n21096 = n6292 | n21095 ;
  assign n21097 = n21096 ^ n17176 ^ n6918 ;
  assign n21094 = n9002 & ~n15948 ;
  assign n21098 = n21097 ^ n21094 ^ 1'b0 ;
  assign n21099 = n2149 | n9088 ;
  assign n21100 = n3895 ^ n1126 ^ 1'b0 ;
  assign n21101 = n21100 ^ n10534 ^ 1'b0 ;
  assign n21102 = x88 & ~n6660 ;
  assign n21103 = n21102 ^ n4230 ^ 1'b0 ;
  assign n21104 = n5540 | n21103 ;
  assign n21105 = n11321 | n20297 ;
  assign n21106 = n21105 ^ n8072 ^ 1'b0 ;
  assign n21107 = n10588 & n16718 ;
  assign n21108 = n21107 ^ n8363 ^ 1'b0 ;
  assign n21109 = n13526 ^ n11415 ^ 1'b0 ;
  assign n21110 = n18813 ^ n16526 ^ 1'b0 ;
  assign n21111 = ~n12384 & n21110 ;
  assign n21112 = n14529 & n21111 ;
  assign n21113 = ~n3775 & n4916 ;
  assign n21114 = n16761 & n21113 ;
  assign n21115 = n21114 ^ n18040 ^ 1'b0 ;
  assign n21116 = ~n12305 & n15669 ;
  assign n21117 = n2857 & ~n21010 ;
  assign n21118 = n8131 & n21117 ;
  assign n21119 = n710 & n2114 ;
  assign n21120 = ~n16946 & n21119 ;
  assign n21121 = n19744 ^ n9218 ^ 1'b0 ;
  assign n21122 = n13870 | n19344 ;
  assign n21123 = n21122 ^ n17168 ^ 1'b0 ;
  assign n21124 = n21121 | n21123 ;
  assign n21125 = ~n6155 & n8677 ;
  assign n21126 = ~n3223 & n21125 ;
  assign n21127 = n9802 ^ n2535 ^ 1'b0 ;
  assign n21128 = n21126 | n21127 ;
  assign n21129 = ~n4342 & n11567 ;
  assign n21130 = ( ~n8336 & n10442 ) | ( ~n8336 & n21129 ) | ( n10442 & n21129 ) ;
  assign n21131 = ~n2970 & n20235 ;
  assign n21132 = n2893 & ~n12538 ;
  assign n21133 = n21132 ^ n7185 ^ 1'b0 ;
  assign n21134 = n16429 & n21133 ;
  assign n21135 = ~n21131 & n21134 ;
  assign n21136 = x48 & n7879 ;
  assign n21137 = ~n9538 & n21136 ;
  assign n21138 = n2369 | n21137 ;
  assign n21139 = n20543 ^ n14935 ^ n7641 ;
  assign n21140 = ~n5160 & n11929 ;
  assign n21141 = ~n9388 & n21140 ;
  assign n21142 = n344 & n6576 ;
  assign n21143 = n21142 ^ n18727 ^ 1'b0 ;
  assign n21144 = n2089 & ~n11627 ;
  assign n21145 = ~n14606 & n21144 ;
  assign n21146 = n21145 ^ n8429 ^ 1'b0 ;
  assign n21147 = n2526 ^ x248 ^ 1'b0 ;
  assign n21148 = n3352 & ~n16735 ;
  assign n21149 = ~n10709 & n21148 ;
  assign n21151 = n4463 ^ n850 ^ 1'b0 ;
  assign n21152 = ~n19200 & n21151 ;
  assign n21150 = n3588 & ~n9263 ;
  assign n21153 = n21152 ^ n21150 ^ 1'b0 ;
  assign n21154 = n15692 ^ n891 ^ 1'b0 ;
  assign n21155 = n12687 & n20726 ;
  assign n21156 = x129 | n5308 ;
  assign n21157 = n21156 ^ n4826 ^ 1'b0 ;
  assign n21158 = n17796 ^ n14752 ^ 1'b0 ;
  assign n21159 = ~n21157 & n21158 ;
  assign n21160 = ( ~n7521 & n10942 ) | ( ~n7521 & n15945 ) | ( n10942 & n15945 ) ;
  assign n21161 = n1621 & n4830 ;
  assign n21162 = n21161 ^ n933 ^ 1'b0 ;
  assign n21163 = n7057 | n21162 ;
  assign n21164 = n5341 | n21163 ;
  assign n21165 = n21164 ^ n7353 ^ 1'b0 ;
  assign n21166 = ~n18098 & n21165 ;
  assign n21167 = n17974 ^ n9551 ^ 1'b0 ;
  assign n21168 = x118 | n11677 ;
  assign n21169 = n3655 & ~n16559 ;
  assign n21170 = n11481 | n21169 ;
  assign n21171 = n21170 ^ n7888 ^ 1'b0 ;
  assign n21172 = n7304 & ~n21171 ;
  assign n21173 = n21172 ^ n6374 ^ n3297 ;
  assign n21174 = ( ~n9630 & n12357 ) | ( ~n9630 & n13154 ) | ( n12357 & n13154 ) ;
  assign n21175 = n19223 ^ n6365 ^ 1'b0 ;
  assign n21176 = n4883 | n21175 ;
  assign n21177 = n15895 ^ n3294 ^ n2868 ;
  assign n21178 = n4673 & n8001 ;
  assign n21179 = n13565 ^ x25 ^ 1'b0 ;
  assign n21180 = n14960 ^ n14012 ^ 1'b0 ;
  assign n21181 = n3400 & n21180 ;
  assign n21182 = n8428 & n21181 ;
  assign n21183 = n21179 & n21182 ;
  assign n21184 = n8733 & ~n8963 ;
  assign n21185 = n516 & n21184 ;
  assign n21186 = n18651 ^ n2296 ^ 1'b0 ;
  assign n21187 = n4993 & ~n21186 ;
  assign n21188 = n21187 ^ n2779 ^ 1'b0 ;
  assign n21189 = n21188 ^ n7818 ^ 1'b0 ;
  assign n21190 = n17395 & ~n21189 ;
  assign n21191 = n4042 | n5851 ;
  assign n21192 = n21190 | n21191 ;
  assign n21193 = n333 | n15999 ;
  assign n21194 = n19768 | n21193 ;
  assign n21195 = n5958 ^ n1729 ^ 1'b0 ;
  assign n21196 = n21194 & n21195 ;
  assign n21197 = n1406 & ~n18200 ;
  assign n21198 = n21197 ^ n7769 ^ 1'b0 ;
  assign n21199 = n21198 ^ n8874 ^ 1'b0 ;
  assign n21200 = n16254 | n21199 ;
  assign n21201 = n14616 & ~n16106 ;
  assign n21202 = n18217 ^ n2948 ^ 1'b0 ;
  assign n21203 = n5450 ^ n3972 ^ 1'b0 ;
  assign n21204 = ~n21202 & n21203 ;
  assign n21205 = n2523 ^ n2319 ^ 1'b0 ;
  assign n21206 = n20533 ^ n2177 ^ 1'b0 ;
  assign n21207 = n21205 & n21206 ;
  assign n21208 = n1875 | n3925 ;
  assign n21209 = n21208 ^ n7707 ^ 1'b0 ;
  assign n21210 = x2 & n10290 ;
  assign n21211 = n14084 & n21210 ;
  assign n21212 = n21211 ^ n12339 ^ 1'b0 ;
  assign n21213 = n7025 | n12070 ;
  assign n21214 = n3030 | n10800 ;
  assign n21215 = x175 | n21214 ;
  assign n21216 = n12998 ^ n6690 ^ 1'b0 ;
  assign n21217 = n2924 & ~n6606 ;
  assign n21218 = n21217 ^ n5203 ^ 1'b0 ;
  assign n21219 = n21218 ^ n18747 ^ 1'b0 ;
  assign n21220 = n2067 & ~n21219 ;
  assign n21221 = n6584 ^ n2013 ^ 1'b0 ;
  assign n21222 = ~n13039 & n21221 ;
  assign n21223 = n1565 & n12603 ;
  assign n21224 = n21223 ^ n10144 ^ 1'b0 ;
  assign n21225 = n15277 & ~n15635 ;
  assign n21226 = n6404 & n10566 ;
  assign n21227 = ~n21225 & n21226 ;
  assign n21228 = n21227 ^ n3574 ^ 1'b0 ;
  assign n21229 = n13311 ^ x6 ^ 1'b0 ;
  assign n21230 = n11013 & n21229 ;
  assign n21231 = n6609 & n8646 ;
  assign n21232 = n12355 ^ n8781 ^ n8667 ;
  assign n21233 = n5559 ^ n3274 ^ 1'b0 ;
  assign n21234 = ( n890 & n10127 ) | ( n890 & n18578 ) | ( n10127 & n18578 ) ;
  assign n21235 = n21234 ^ n16301 ^ n6582 ;
  assign n21236 = n12397 ^ n11316 ^ 1'b0 ;
  assign n21237 = ~n2460 & n21236 ;
  assign n21238 = n21237 ^ n19927 ^ 1'b0 ;
  assign n21239 = n11179 ^ x41 ^ 1'b0 ;
  assign n21240 = n19124 | n21239 ;
  assign n21241 = n7053 & ~n18255 ;
  assign n21242 = n7494 & n21241 ;
  assign n21243 = n19167 | n21242 ;
  assign n21244 = n21243 ^ n2663 ^ 1'b0 ;
  assign n21245 = x24 & ~n8133 ;
  assign n21246 = n21245 ^ n9311 ^ 1'b0 ;
  assign n21247 = n11226 & n21246 ;
  assign n21248 = n3666 & n4799 ;
  assign n21249 = n21247 & n21248 ;
  assign n21250 = n21249 ^ n6563 ^ 1'b0 ;
  assign n21251 = n9958 ^ n6959 ^ 1'b0 ;
  assign n21252 = n932 | n1962 ;
  assign n21253 = n21252 ^ n10999 ^ 1'b0 ;
  assign n21254 = n6195 | n16438 ;
  assign n21255 = x0 & n21254 ;
  assign n21256 = n6333 & n21255 ;
  assign n21257 = ~n7089 & n21256 ;
  assign n21258 = n11375 ^ n4807 ^ n2870 ;
  assign n21259 = n11676 ^ n5023 ^ 1'b0 ;
  assign n21260 = n10082 & n14523 ;
  assign n21261 = n21260 ^ n1550 ^ 1'b0 ;
  assign n21262 = n6991 | n9072 ;
  assign n21263 = n20788 & n21262 ;
  assign n21264 = n8277 & ~n9436 ;
  assign n21265 = n7907 & ~n15122 ;
  assign n21266 = n3739 ^ n2577 ^ n1977 ;
  assign n21267 = n21266 ^ n2789 ^ 1'b0 ;
  assign n21268 = x172 | n21267 ;
  assign n21269 = ~n4541 & n11838 ;
  assign n21270 = n21269 ^ n14288 ^ 1'b0 ;
  assign n21271 = ~n21268 & n21270 ;
  assign n21272 = n2946 & n18326 ;
  assign n21273 = n15212 ^ n5402 ^ n4074 ;
  assign n21274 = ~n5820 & n12725 ;
  assign n21277 = n749 & ~n9762 ;
  assign n21278 = ~n749 & n21277 ;
  assign n21275 = n5853 | n9228 ;
  assign n21276 = n9946 & ~n21275 ;
  assign n21279 = n21278 ^ n21276 ^ 1'b0 ;
  assign n21280 = ~n11883 & n21279 ;
  assign n21281 = n4983 & ~n14998 ;
  assign n21282 = n21281 ^ n4086 ^ 1'b0 ;
  assign n21283 = ~n15123 & n21282 ;
  assign n21284 = n3216 & n14402 ;
  assign n21285 = ~n11019 & n21284 ;
  assign n21286 = ~n8476 & n17650 ;
  assign n21287 = n2771 & n21286 ;
  assign n21288 = n14908 ^ n6317 ^ 1'b0 ;
  assign n21289 = n21266 & ~n21288 ;
  assign n21290 = n21289 ^ n1591 ^ 1'b0 ;
  assign n21291 = n8401 & n21290 ;
  assign n21292 = ( n11061 & ~n12758 ) | ( n11061 & n21291 ) | ( ~n12758 & n21291 ) ;
  assign n21293 = n4610 & ~n9545 ;
  assign n21294 = ~n15932 & n21293 ;
  assign n21295 = n14157 ^ n6759 ^ 1'b0 ;
  assign n21296 = n932 & ~n6964 ;
  assign n21297 = ( ~x117 & n17694 ) | ( ~x117 & n21296 ) | ( n17694 & n21296 ) ;
  assign n21298 = x53 & ~n13810 ;
  assign n21299 = ~n2275 & n21298 ;
  assign n21300 = n8634 & n16080 ;
  assign n21301 = n12201 ^ n2324 ^ 1'b0 ;
  assign n21302 = n21300 & ~n21301 ;
  assign n21303 = n8130 | n19916 ;
  assign n21304 = n11503 ^ n6532 ^ 1'b0 ;
  assign n21305 = n13942 & n21304 ;
  assign n21306 = x51 & n8004 ;
  assign n21307 = n8079 | n21306 ;
  assign n21308 = n14821 ^ n813 ^ n466 ;
  assign n21309 = ~n716 & n11295 ;
  assign n21310 = n17480 & ~n21309 ;
  assign n21311 = n7830 & n12865 ;
  assign n21312 = ~n5385 & n21311 ;
  assign n21313 = ~n3139 & n21312 ;
  assign n21314 = n21313 ^ n1714 ^ 1'b0 ;
  assign n21315 = n3702 & ~n21314 ;
  assign n21316 = n21315 ^ n7087 ^ 1'b0 ;
  assign n21317 = n1132 & ~n21316 ;
  assign n21318 = n10917 & ~n19866 ;
  assign n21319 = n11204 | n21318 ;
  assign n21321 = n4337 & n7420 ;
  assign n21322 = n8276 & n21321 ;
  assign n21320 = n3067 & n11127 ;
  assign n21323 = n21322 ^ n21320 ^ 1'b0 ;
  assign n21324 = n2275 | n9554 ;
  assign n21325 = n21323 & ~n21324 ;
  assign n21326 = ~n3494 & n10949 ;
  assign n21327 = n21326 ^ n9879 ^ 1'b0 ;
  assign n21328 = n9028 | n21327 ;
  assign n21329 = n19148 | n21328 ;
  assign n21331 = n6730 ^ n6317 ^ n2859 ;
  assign n21330 = x46 & ~n765 ;
  assign n21332 = n21331 ^ n21330 ^ 1'b0 ;
  assign n21333 = n5305 & n7506 ;
  assign n21334 = ~n2131 & n11331 ;
  assign n21335 = n1382 & n21334 ;
  assign n21336 = ( n9289 & n14690 ) | ( n9289 & n21335 ) | ( n14690 & n21335 ) ;
  assign n21337 = n5016 & n16758 ;
  assign n21338 = n21337 ^ n16523 ^ 1'b0 ;
  assign n21339 = n12245 ^ n3866 ^ 1'b0 ;
  assign n21340 = ~n11290 & n21339 ;
  assign n21341 = ~n3650 & n13238 ;
  assign n21342 = n21341 ^ n10360 ^ 1'b0 ;
  assign n21343 = n3073 ^ x221 ^ 1'b0 ;
  assign n21344 = ~n3047 & n21343 ;
  assign n21345 = ~n13540 & n21344 ;
  assign n21346 = n21345 ^ n13824 ^ 1'b0 ;
  assign n21347 = n7458 ^ n1633 ^ 1'b0 ;
  assign n21348 = n5579 & ~n21347 ;
  assign n21349 = n6433 ^ n5162 ^ 1'b0 ;
  assign n21350 = n4205 & ~n5894 ;
  assign n21351 = n11439 | n11655 ;
  assign n21352 = n10540 ^ n4343 ^ n4174 ;
  assign n21353 = n3411 & n12138 ;
  assign n21354 = n3319 | n9733 ;
  assign n21355 = n1405 & ~n21354 ;
  assign n21356 = n9632 & ~n21355 ;
  assign n21357 = n21353 | n21356 ;
  assign n21358 = n9366 | n9781 ;
  assign n21359 = n8570 ^ n2400 ^ 1'b0 ;
  assign n21360 = n21358 & ~n21359 ;
  assign n21361 = n920 & n13184 ;
  assign n21362 = n8059 & n21361 ;
  assign n21363 = ~n13829 & n21362 ;
  assign n21364 = n3091 ^ x165 ^ 1'b0 ;
  assign n21365 = n15966 ^ n6964 ^ 1'b0 ;
  assign n21366 = ( n19714 & n21364 ) | ( n19714 & ~n21365 ) | ( n21364 & ~n21365 ) ;
  assign n21367 = ~n21363 & n21366 ;
  assign n21368 = n7298 & n21367 ;
  assign n21369 = n3911 | n10997 ;
  assign n21370 = ( n1854 & n6945 ) | ( n1854 & ~n21369 ) | ( n6945 & ~n21369 ) ;
  assign n21371 = n14669 ^ n5865 ^ 1'b0 ;
  assign n21372 = n3464 & ~n18628 ;
  assign n21373 = n21372 ^ n9572 ^ 1'b0 ;
  assign n21374 = n21171 ^ n8269 ^ 1'b0 ;
  assign n21375 = n9303 | n21374 ;
  assign n21376 = n680 & ~n11891 ;
  assign n21377 = ~n680 & n21376 ;
  assign n21378 = ~n15518 & n21377 ;
  assign n21379 = ~n1667 & n21378 ;
  assign n21380 = n1667 & n21379 ;
  assign n21381 = n11354 ^ n3416 ^ 1'b0 ;
  assign n21382 = x65 & ~n21381 ;
  assign n21383 = ~n21380 & n21382 ;
  assign n21384 = n21383 ^ n12865 ^ 1'b0 ;
  assign n21385 = n16366 & ~n18551 ;
  assign n21386 = n21385 ^ n19626 ^ 1'b0 ;
  assign n21387 = n13360 ^ n10239 ^ 1'b0 ;
  assign n21388 = n10884 & ~n21387 ;
  assign n21391 = n1664 & n5287 ;
  assign n21392 = n3863 ^ n969 ^ 1'b0 ;
  assign n21393 = n21391 | n21392 ;
  assign n21389 = n501 & ~n7135 ;
  assign n21390 = ~n13343 & n21389 ;
  assign n21394 = n21393 ^ n21390 ^ 1'b0 ;
  assign n21395 = n21388 & n21394 ;
  assign n21396 = n10532 & n13077 ;
  assign n21397 = n11863 & ~n18023 ;
  assign n21398 = n21397 ^ n16326 ^ 1'b0 ;
  assign n21399 = n12242 ^ n6053 ^ 1'b0 ;
  assign n21400 = n15880 | n21399 ;
  assign n21401 = n2004 & ~n11264 ;
  assign n21402 = n14302 ^ n9513 ^ 1'b0 ;
  assign n21403 = n20662 ^ n5118 ^ 1'b0 ;
  assign n21404 = ~n4119 & n21403 ;
  assign n21405 = ~n6369 & n21404 ;
  assign n21406 = ~n14754 & n21405 ;
  assign n21407 = n21406 ^ n8147 ^ n1369 ;
  assign n21408 = ~n6623 & n19866 ;
  assign n21409 = ~n21407 & n21408 ;
  assign n21410 = n14451 | n17887 ;
  assign n21411 = n1163 & ~n21410 ;
  assign n21412 = n10208 & ~n21411 ;
  assign n21413 = n21412 ^ n4550 ^ 1'b0 ;
  assign n21414 = n3146 ^ n3142 ^ 1'b0 ;
  assign n21415 = n21414 ^ n13539 ^ 1'b0 ;
  assign n21416 = n21413 & ~n21415 ;
  assign n21417 = n12451 ^ n1682 ^ 1'b0 ;
  assign n21418 = n21417 ^ n8636 ^ n6744 ;
  assign n21419 = n2982 ^ n1813 ^ 1'b0 ;
  assign n21420 = n12269 ^ n3939 ^ 1'b0 ;
  assign n21421 = ~n9654 & n10770 ;
  assign n21422 = n7832 ^ n4638 ^ 1'b0 ;
  assign n21423 = x223 & ~n10840 ;
  assign n21424 = ~n17666 & n21423 ;
  assign n21425 = x8 & n3450 ;
  assign n21426 = n21425 ^ n1833 ^ 1'b0 ;
  assign n21427 = n21426 ^ n10022 ^ 1'b0 ;
  assign n21428 = n5432 | n21427 ;
  assign n21429 = n21428 ^ n7191 ^ 1'b0 ;
  assign n21430 = n7831 | n21429 ;
  assign n21431 = n2356 ^ n2282 ^ 1'b0 ;
  assign n21432 = n289 & ~n21431 ;
  assign n21433 = n1563 & n21432 ;
  assign n21434 = n21433 ^ n13861 ^ 1'b0 ;
  assign n21435 = n14412 | n21434 ;
  assign n21436 = n21435 ^ n10105 ^ 1'b0 ;
  assign n21437 = n7940 ^ n6335 ^ 1'b0 ;
  assign n21438 = n18002 & ~n21437 ;
  assign n21439 = ( ~n14792 & n21436 ) | ( ~n14792 & n21438 ) | ( n21436 & n21438 ) ;
  assign n21442 = n4944 & ~n18551 ;
  assign n21443 = ~n4944 & n21442 ;
  assign n21440 = n17373 ^ n1148 ^ 1'b0 ;
  assign n21441 = n21440 ^ n19128 ^ 1'b0 ;
  assign n21444 = n21443 ^ n21441 ^ 1'b0 ;
  assign n21445 = ~n1855 & n20593 ;
  assign n21446 = n6868 ^ n6526 ^ x115 ;
  assign n21447 = n8801 | n21446 ;
  assign n21448 = n7232 ^ n5851 ^ 1'b0 ;
  assign n21449 = n14341 | n21448 ;
  assign n21450 = n12328 & ~n21449 ;
  assign n21453 = n1600 & ~n2831 ;
  assign n21454 = n21453 ^ n12165 ^ 1'b0 ;
  assign n21451 = n6164 ^ n997 ^ 1'b0 ;
  assign n21452 = n8837 & n21451 ;
  assign n21455 = n21454 ^ n21452 ^ 1'b0 ;
  assign n21456 = n2788 | n15977 ;
  assign n21457 = n17447 | n21456 ;
  assign n21458 = n4315 & ~n17517 ;
  assign n21459 = n15259 & n21458 ;
  assign n21460 = x40 & ~n11134 ;
  assign n21461 = n17728 ^ n14120 ^ n10794 ;
  assign n21462 = n21461 ^ n14053 ^ n8216 ;
  assign n21463 = n13212 ^ n1338 ^ 1'b0 ;
  assign n21464 = ~n2302 & n21463 ;
  assign n21465 = n15760 & ~n21464 ;
  assign n21466 = ~n14177 & n17362 ;
  assign n21467 = ( ~n1272 & n5570 ) | ( ~n1272 & n21466 ) | ( n5570 & n21466 ) ;
  assign n21468 = n19591 & n21467 ;
  assign n21469 = n21465 | n21468 ;
  assign n21470 = n21469 ^ n9061 ^ 1'b0 ;
  assign n21471 = n20914 ^ n7801 ^ 1'b0 ;
  assign n21472 = n17312 & ~n21471 ;
  assign n21473 = n13809 & n21472 ;
  assign n21474 = n1138 & n13031 ;
  assign n21475 = n21474 ^ n12123 ^ n7301 ;
  assign n21476 = ~n15427 & n19309 ;
  assign n21477 = n21476 ^ x4 ^ 1'b0 ;
  assign n21478 = n16967 ^ n3823 ^ 1'b0 ;
  assign n21479 = ~n1971 & n9811 ;
  assign n21480 = n665 & n21479 ;
  assign n21481 = n6954 & n9079 ;
  assign n21482 = ~n1734 & n21481 ;
  assign n21483 = ( n6031 & n14030 ) | ( n6031 & n21482 ) | ( n14030 & n21482 ) ;
  assign n21484 = n21483 ^ n4096 ^ 1'b0 ;
  assign n21485 = n4004 | n9321 ;
  assign n21486 = n21484 & ~n21485 ;
  assign n21487 = n13560 ^ n4795 ^ 1'b0 ;
  assign n21488 = ( n5062 & n16283 ) | ( n5062 & n21487 ) | ( n16283 & n21487 ) ;
  assign n21489 = n3917 | n14448 ;
  assign n21490 = ~n5049 & n8044 ;
  assign n21492 = ~n1551 & n8909 ;
  assign n21491 = n1391 & ~n1855 ;
  assign n21493 = n21492 ^ n21491 ^ n3195 ;
  assign n21494 = ~n11392 & n21493 ;
  assign n21495 = n21490 & n21494 ;
  assign n21496 = n16495 ^ n6701 ^ 1'b0 ;
  assign n21497 = n2262 | n21496 ;
  assign n21498 = n21497 ^ n2446 ^ 1'b0 ;
  assign n21499 = n15889 & ~n21498 ;
  assign n21500 = n1682 & ~n14908 ;
  assign n21501 = n12309 ^ n5237 ^ 1'b0 ;
  assign n21502 = x73 & n19623 ;
  assign n21503 = n21502 ^ n3016 ^ 1'b0 ;
  assign n21504 = n19815 ^ n6603 ^ x55 ;
  assign n21505 = n3776 & ~n7332 ;
  assign n21506 = n21505 ^ n2121 ^ 1'b0 ;
  assign n21507 = ( n943 & n1223 ) | ( n943 & ~n2718 ) | ( n1223 & ~n2718 ) ;
  assign n21508 = ~n2646 & n17426 ;
  assign n21509 = n21508 ^ n9609 ^ 1'b0 ;
  assign n21510 = n6895 | n8408 ;
  assign n21511 = n21509 & ~n21510 ;
  assign n21512 = n8481 & ~n21511 ;
  assign n21513 = ~n21507 & n21512 ;
  assign n21514 = n15187 ^ n812 ^ 1'b0 ;
  assign n21515 = n1328 & ~n21514 ;
  assign n21516 = n2247 | n6304 ;
  assign n21517 = n4666 & ~n21516 ;
  assign n21518 = ~n1032 & n21517 ;
  assign n21519 = ~n2141 & n14202 ;
  assign n21520 = n21518 & n21519 ;
  assign n21521 = ~n4830 & n8112 ;
  assign n21522 = ~n3802 & n13193 ;
  assign n21523 = n10383 & n21522 ;
  assign n21524 = n21521 & ~n21523 ;
  assign n21530 = n6655 ^ n2930 ^ 1'b0 ;
  assign n21531 = n6950 & n21530 ;
  assign n21525 = n12902 ^ n764 ^ 1'b0 ;
  assign n21526 = n2835 & ~n18583 ;
  assign n21527 = n409 & ~n21526 ;
  assign n21528 = ~n21525 & n21527 ;
  assign n21529 = n8342 | n21528 ;
  assign n21532 = n21531 ^ n21529 ^ 1'b0 ;
  assign n21533 = x129 & n10552 ;
  assign n21534 = n1085 & n1249 ;
  assign n21535 = ~n3525 & n21534 ;
  assign n21536 = n11554 | n21535 ;
  assign n21537 = n21536 ^ n9428 ^ 1'b0 ;
  assign n21538 = n21537 ^ n6479 ^ n5614 ;
  assign n21539 = n21538 ^ n19678 ^ 1'b0 ;
  assign n21540 = n12639 | n18535 ;
  assign n21541 = n21540 ^ n10172 ^ 1'b0 ;
  assign n21542 = n4995 & ~n7351 ;
  assign n21543 = n21542 ^ n16853 ^ 1'b0 ;
  assign n21544 = n4970 & ~n21543 ;
  assign n21545 = n21544 ^ n8663 ^ 1'b0 ;
  assign n21546 = n10915 ^ n983 ^ 1'b0 ;
  assign n21547 = ~n5589 & n10432 ;
  assign n21548 = ~n8893 & n21547 ;
  assign n21549 = n15255 & ~n21548 ;
  assign n21550 = n13533 & n21549 ;
  assign n21551 = n21550 ^ n19805 ^ 1'b0 ;
  assign n21552 = n8970 & n18921 ;
  assign n21553 = ~n9996 & n19961 ;
  assign n21554 = n3474 ^ n3106 ^ 1'b0 ;
  assign n21555 = ~n2710 & n21554 ;
  assign n21556 = n21555 ^ n16391 ^ 1'b0 ;
  assign n21557 = ~n1332 & n16906 ;
  assign n21558 = n21556 & n21557 ;
  assign n21559 = ~n4935 & n7683 ;
  assign n21560 = ~n8092 & n21559 ;
  assign n21561 = n20152 ^ n625 ^ 1'b0 ;
  assign n21562 = ~n21560 & n21561 ;
  assign n21563 = n4509 | n6119 ;
  assign n21564 = n1042 & n1484 ;
  assign n21565 = ~n1484 & n21564 ;
  assign n21566 = x58 & ~n21565 ;
  assign n21567 = ~x58 & n21566 ;
  assign n21568 = ~n1067 & n5046 ;
  assign n21569 = n21567 & n21568 ;
  assign n21570 = n21569 ^ n3383 ^ 1'b0 ;
  assign n21571 = n11185 | n21570 ;
  assign n21572 = n4296 & ~n8355 ;
  assign n21573 = ~n6400 & n21572 ;
  assign n21574 = n8141 | n21573 ;
  assign n21575 = n19785 ^ n10710 ^ 1'b0 ;
  assign n21576 = n21575 ^ n10535 ^ 1'b0 ;
  assign n21577 = n6370 ^ n1146 ^ 1'b0 ;
  assign n21578 = n21577 ^ n8016 ^ 1'b0 ;
  assign n21579 = n21578 ^ n7294 ^ 1'b0 ;
  assign n21580 = n21018 ^ n12332 ^ 1'b0 ;
  assign n21581 = ~n15792 & n21580 ;
  assign n21582 = n7358 ^ n2983 ^ n1267 ;
  assign n21583 = ~n6873 & n21582 ;
  assign n21584 = n13079 ^ n9251 ^ 1'b0 ;
  assign n21585 = ~x120 & n21584 ;
  assign n21586 = n1454 & n21585 ;
  assign n21587 = n21586 ^ n5992 ^ 1'b0 ;
  assign n21588 = ~n2647 & n21587 ;
  assign n21589 = n923 & n2485 ;
  assign n21590 = n21589 ^ n10978 ^ 1'b0 ;
  assign n21591 = ~x116 & n21590 ;
  assign n21592 = n17674 | n21591 ;
  assign n21593 = ~n16297 & n19441 ;
  assign n21594 = ( ~x244 & n854 ) | ( ~x244 & n10514 ) | ( n854 & n10514 ) ;
  assign n21595 = n21594 ^ n15998 ^ 1'b0 ;
  assign n21596 = n16968 & ~n21595 ;
  assign n21597 = ~n11042 & n11108 ;
  assign n21598 = n21597 ^ n10610 ^ 1'b0 ;
  assign n21599 = n16668 | n21598 ;
  assign n21603 = n279 & ~n18700 ;
  assign n21604 = n21603 ^ n1336 ^ 1'b0 ;
  assign n21600 = n4175 & n9714 ;
  assign n21601 = n20746 ^ n16513 ^ n5025 ;
  assign n21602 = ( n7269 & n21600 ) | ( n7269 & ~n21601 ) | ( n21600 & ~n21601 ) ;
  assign n21605 = n21604 ^ n21602 ^ 1'b0 ;
  assign n21606 = n11755 & n21605 ;
  assign n21607 = n2672 & n21606 ;
  assign n21608 = ~x82 & n21607 ;
  assign n21609 = n17643 ^ n15275 ^ 1'b0 ;
  assign n21610 = n21609 ^ n12659 ^ 1'b0 ;
  assign n21611 = ( n7273 & n9062 ) | ( n7273 & n18205 ) | ( n9062 & n18205 ) ;
  assign n21612 = n10872 ^ n2988 ^ 1'b0 ;
  assign n21613 = n6526 & ~n21612 ;
  assign n21614 = n5771 | n13357 ;
  assign n21615 = n4031 & ~n21614 ;
  assign n21616 = n21615 ^ n5983 ^ n4249 ;
  assign n21617 = ( n5078 & n9755 ) | ( n5078 & n16915 ) | ( n9755 & n16915 ) ;
  assign n21618 = ~n9220 & n9264 ;
  assign n21619 = n19525 ^ n9664 ^ 1'b0 ;
  assign n21620 = n15071 | n21619 ;
  assign n21621 = n11892 ^ n9990 ^ 1'b0 ;
  assign n21622 = ~n15668 & n21621 ;
  assign n21623 = n21622 ^ n16377 ^ n318 ;
  assign n21624 = ~n13214 & n13641 ;
  assign n21625 = n21624 ^ n15055 ^ 1'b0 ;
  assign n21626 = ~n593 & n8301 ;
  assign n21627 = n5421 & ~n6897 ;
  assign n21628 = n21626 & n21627 ;
  assign n21629 = n14285 ^ n6797 ^ 1'b0 ;
  assign n21630 = n21629 ^ n10124 ^ 1'b0 ;
  assign n21631 = n4992 | n21630 ;
  assign n21632 = n738 & n17127 ;
  assign n21633 = ~n6049 & n21632 ;
  assign n21634 = n21633 ^ n462 ^ x36 ;
  assign n21635 = n14846 & n17411 ;
  assign n21636 = n4432 & n9113 ;
  assign n21637 = n21636 ^ n10551 ^ 1'b0 ;
  assign n21638 = n15737 | n21066 ;
  assign n21639 = n21637 | n21638 ;
  assign n21640 = n6270 ^ n2167 ^ 1'b0 ;
  assign n21641 = n15612 & n21640 ;
  assign n21643 = n3106 & ~n17374 ;
  assign n21642 = x205 & ~n9808 ;
  assign n21644 = n21643 ^ n21642 ^ 1'b0 ;
  assign n21645 = n21644 ^ n19422 ^ 1'b0 ;
  assign n21646 = n11659 ^ n7685 ^ 1'b0 ;
  assign n21647 = n267 | n14341 ;
  assign n21648 = n7330 ^ n5315 ^ 1'b0 ;
  assign n21649 = n4932 & ~n21648 ;
  assign n21650 = ( n17517 & n21647 ) | ( n17517 & n21649 ) | ( n21647 & n21649 ) ;
  assign n21651 = n3913 & ~n21650 ;
  assign n21652 = n17562 ^ n5231 ^ 1'b0 ;
  assign n21653 = ~n11699 & n21652 ;
  assign n21654 = n7128 & ~n8198 ;
  assign n21655 = n9526 | n21654 ;
  assign n21656 = n1659 & n15514 ;
  assign n21657 = n5700 & n21656 ;
  assign n21658 = ( n8071 & n12361 ) | ( n8071 & n19310 ) | ( n12361 & n19310 ) ;
  assign n21659 = n4691 | n7828 ;
  assign n21660 = n21659 ^ n2062 ^ 1'b0 ;
  assign n21661 = ( ~n9377 & n19237 ) | ( ~n9377 & n21660 ) | ( n19237 & n21660 ) ;
  assign n21662 = n7329 & n18296 ;
  assign n21663 = n2122 & n21662 ;
  assign n21668 = n11813 & ~n17918 ;
  assign n21669 = n16491 & n21668 ;
  assign n21670 = n21669 ^ n18838 ^ 1'b0 ;
  assign n21664 = n638 | n4648 ;
  assign n21665 = n18171 | n21664 ;
  assign n21666 = n21665 ^ n9154 ^ 1'b0 ;
  assign n21667 = n6476 & ~n21666 ;
  assign n21671 = n21670 ^ n21667 ^ 1'b0 ;
  assign n21672 = n5713 & n10385 ;
  assign n21673 = n17040 & n21672 ;
  assign n21674 = ( ~n1085 & n8426 ) | ( ~n1085 & n20144 ) | ( n8426 & n20144 ) ;
  assign n21675 = n21674 ^ n14283 ^ n2951 ;
  assign n21676 = n4025 | n7482 ;
  assign n21677 = n2535 & n9724 ;
  assign n21678 = n3124 & n21677 ;
  assign n21679 = n15372 | n21678 ;
  assign n21680 = n17926 | n21679 ;
  assign n21681 = ~n14518 & n21680 ;
  assign n21682 = n407 & n21681 ;
  assign n21683 = n4245 | n7902 ;
  assign n21684 = ~n2016 & n3014 ;
  assign n21686 = n8834 | n13813 ;
  assign n21685 = n4902 & ~n5305 ;
  assign n21687 = n21686 ^ n21685 ^ n8104 ;
  assign n21688 = n3838 & ~n21687 ;
  assign n21689 = ( n8424 & n10622 ) | ( n8424 & n21688 ) | ( n10622 & n21688 ) ;
  assign n21690 = n4172 & ~n6701 ;
  assign n21691 = n21690 ^ n3238 ^ 1'b0 ;
  assign n21692 = n21691 ^ n4067 ^ n961 ;
  assign n21693 = n21692 ^ n11986 ^ 1'b0 ;
  assign n21694 = n2484 & n21693 ;
  assign n21695 = n5118 | n6957 ;
  assign n21696 = ~n3243 & n18343 ;
  assign n21697 = n19557 & ~n21696 ;
  assign n21698 = n21695 & n21697 ;
  assign n21699 = n16215 ^ n11374 ^ 1'b0 ;
  assign n21700 = ~n1756 & n10059 ;
  assign n21701 = ~n8244 & n21700 ;
  assign n21702 = n3169 & n21701 ;
  assign n21703 = ~n21347 & n21702 ;
  assign n21704 = n10646 & ~n11191 ;
  assign n21705 = n21704 ^ n12737 ^ 1'b0 ;
  assign n21706 = n11366 | n21016 ;
  assign n21707 = n8873 | n21706 ;
  assign n21708 = n3875 | n10414 ;
  assign n21709 = n18546 ^ n4397 ^ 1'b0 ;
  assign n21710 = n21708 & n21709 ;
  assign n21711 = n8667 ^ n1598 ^ 1'b0 ;
  assign n21712 = n6015 & n21711 ;
  assign n21713 = n8814 & ~n21712 ;
  assign n21714 = n18142 & n21713 ;
  assign n21715 = n6797 & n17488 ;
  assign n21716 = n21714 & n21715 ;
  assign n21717 = n10915 | n19191 ;
  assign n21718 = n21717 ^ n5847 ^ 1'b0 ;
  assign n21719 = n4051 & n6190 ;
  assign n21720 = n13861 ^ n2940 ^ 1'b0 ;
  assign n21721 = ~n17349 & n21720 ;
  assign n21722 = n5517 & n12446 ;
  assign n21723 = n21722 ^ n8305 ^ 1'b0 ;
  assign n21724 = n21723 ^ n991 ^ 1'b0 ;
  assign n21725 = n4132 & ~n4821 ;
  assign n21726 = n21725 ^ n6331 ^ 1'b0 ;
  assign n21727 = n14571 & n21726 ;
  assign n21728 = n13022 & ~n21727 ;
  assign n21729 = n3425 & ~n13357 ;
  assign n21730 = n10988 & n21729 ;
  assign n21731 = n20536 | n21730 ;
  assign n21732 = n5813 & ~n21731 ;
  assign n21733 = n6470 & ~n9973 ;
  assign n21734 = n21733 ^ n8770 ^ 1'b0 ;
  assign n21735 = n21734 ^ n11678 ^ 1'b0 ;
  assign n21736 = n19619 & ~n21735 ;
  assign n21737 = n618 & n3695 ;
  assign n21738 = n21737 ^ n5895 ^ 1'b0 ;
  assign n21739 = n389 | n21738 ;
  assign n21740 = n21739 ^ n256 ^ 1'b0 ;
  assign n21741 = n6342 & n7798 ;
  assign n21742 = n12932 ^ n6298 ^ 1'b0 ;
  assign n21743 = n12713 & n21742 ;
  assign n21744 = n21743 ^ n11849 ^ n1945 ;
  assign n21750 = n10480 & n18180 ;
  assign n21745 = n19624 ^ n1405 ^ n809 ;
  assign n21746 = n5402 ^ n4443 ^ 1'b0 ;
  assign n21747 = x100 & n21746 ;
  assign n21748 = n655 & n21747 ;
  assign n21749 = n21745 & n21748 ;
  assign n21751 = n21750 ^ n21749 ^ 1'b0 ;
  assign n21752 = n389 & n9792 ;
  assign n21753 = n3349 & ~n21752 ;
  assign n21754 = n14912 ^ n9892 ^ 1'b0 ;
  assign n21755 = n3876 & ~n18011 ;
  assign n21756 = n6853 | n11414 ;
  assign n21757 = n21756 ^ n8666 ^ 1'b0 ;
  assign n21758 = n20410 & n21757 ;
  assign n21759 = n17224 ^ n12766 ^ 1'b0 ;
  assign n21760 = n15547 & n21759 ;
  assign n21761 = n21397 | n21760 ;
  assign n21762 = ~n7447 & n20582 ;
  assign n21763 = ~n11994 & n21762 ;
  assign n21764 = n11155 ^ n8302 ^ 1'b0 ;
  assign n21765 = n1010 | n5168 ;
  assign n21766 = n21765 ^ n6060 ^ 1'b0 ;
  assign n21767 = x114 & ~n21766 ;
  assign n21768 = ~n9175 & n21767 ;
  assign n21769 = n13487 & ~n21768 ;
  assign n21770 = n21769 ^ n10627 ^ 1'b0 ;
  assign n21771 = n3266 ^ n1028 ^ 1'b0 ;
  assign n21772 = n20913 ^ n14666 ^ 1'b0 ;
  assign n21773 = x110 & n2250 ;
  assign n21774 = ~n2250 & n21773 ;
  assign n21775 = n886 & n1626 ;
  assign n21776 = ~n886 & n21775 ;
  assign n21777 = ~n5241 & n21776 ;
  assign n21778 = n21774 | n21777 ;
  assign n21779 = n21778 ^ n10460 ^ 1'b0 ;
  assign n21780 = n15802 ^ n2089 ^ 1'b0 ;
  assign n21781 = n16095 ^ n15234 ^ 1'b0 ;
  assign n21782 = ( ~n8666 & n21780 ) | ( ~n8666 & n21781 ) | ( n21780 & n21781 ) ;
  assign n21783 = x149 & ~n21291 ;
  assign n21784 = n10310 ^ n5195 ^ 1'b0 ;
  assign n21785 = ~n17001 & n21784 ;
  assign n21786 = n7510 | n21785 ;
  assign n21787 = n3853 & ~n6807 ;
  assign n21788 = ~n19497 & n21787 ;
  assign n21789 = n6611 & ~n21788 ;
  assign n21790 = n21789 ^ n13731 ^ 1'b0 ;
  assign n21791 = n5318 ^ n2362 ^ 1'b0 ;
  assign n21792 = n11656 | n21791 ;
  assign n21793 = n20614 ^ n4739 ^ 1'b0 ;
  assign n21794 = ~n1583 & n21793 ;
  assign n21795 = n21616 | n21794 ;
  assign n21796 = ~n6957 & n14788 ;
  assign n21797 = n13452 ^ n11142 ^ n1867 ;
  assign n21798 = n10336 ^ n2812 ^ 1'b0 ;
  assign n21799 = n9933 ^ n6886 ^ 1'b0 ;
  assign n21800 = n3576 & ~n21799 ;
  assign n21801 = n1092 & ~n21800 ;
  assign n21802 = ( n16390 & n19656 ) | ( n16390 & n21801 ) | ( n19656 & n21801 ) ;
  assign n21803 = n15316 & n21802 ;
  assign n21804 = ~n15299 & n21803 ;
  assign n21805 = n7345 ^ n2061 ^ 1'b0 ;
  assign n21806 = n1328 ^ x230 ^ 1'b0 ;
  assign n21807 = n4698 ^ n3685 ^ n2903 ;
  assign n21808 = ~n4896 & n21807 ;
  assign n21809 = n13116 | n14263 ;
  assign n21810 = n21808 | n21809 ;
  assign n21811 = n5216 & n5385 ;
  assign n21812 = ~n15275 & n21811 ;
  assign n21813 = n10738 | n21483 ;
  assign n21814 = n5602 ^ n3493 ^ n1997 ;
  assign n21815 = n21814 ^ n12411 ^ 1'b0 ;
  assign n21816 = ~n12288 & n21815 ;
  assign n21817 = ~n13856 & n21816 ;
  assign n21818 = n2235 | n5977 ;
  assign n21819 = n21818 ^ n6278 ^ 1'b0 ;
  assign n21820 = n7066 & ~n21819 ;
  assign n21821 = n21820 ^ n19198 ^ 1'b0 ;
  assign n21822 = ( n3564 & ~n21817 ) | ( n3564 & n21821 ) | ( ~n21817 & n21821 ) ;
  assign n21823 = n8186 ^ n7752 ^ 1'b0 ;
  assign n21824 = n21823 ^ n15850 ^ n2655 ;
  assign n21825 = n7241 | n21824 ;
  assign n21826 = n21825 ^ n9397 ^ x82 ;
  assign n21827 = ~n5566 & n6920 ;
  assign n21828 = n1409 & n21827 ;
  assign n21829 = n7906 & ~n21828 ;
  assign n21830 = n21829 ^ n4527 ^ 1'b0 ;
  assign n21831 = n12792 & n21830 ;
  assign n21832 = n3199 & ~n11369 ;
  assign n21833 = n11369 & n21832 ;
  assign n21834 = n2687 & n7190 ;
  assign n21835 = n4875 | n5323 ;
  assign n21836 = n21835 ^ n15008 ^ 1'b0 ;
  assign n21837 = n21834 & n21836 ;
  assign n21838 = ~n15533 & n19971 ;
  assign n21839 = n11772 ^ n8330 ^ 1'b0 ;
  assign n21841 = n16877 ^ n11381 ^ 1'b0 ;
  assign n21842 = n1992 ^ n1590 ^ 1'b0 ;
  assign n21843 = ~n21841 & n21842 ;
  assign n21840 = n7418 & ~n9844 ;
  assign n21844 = n21843 ^ n21840 ^ 1'b0 ;
  assign n21845 = n2383 | n19349 ;
  assign n21846 = n4325 & n16246 ;
  assign n21847 = ~n1023 & n21846 ;
  assign n21848 = ~n14430 & n14484 ;
  assign n21849 = ~x103 & n7476 ;
  assign n21850 = n6504 & n21643 ;
  assign n21851 = n21849 & n21850 ;
  assign n21852 = n6429 & ~n20332 ;
  assign n21853 = n4447 & ~n7036 ;
  assign n21854 = n21853 ^ n20817 ^ 1'b0 ;
  assign n21855 = n3626 | n13049 ;
  assign n21856 = n21854 & ~n21855 ;
  assign n21857 = n2167 & n15692 ;
  assign n21858 = ~n7304 & n21857 ;
  assign n21859 = ~n5416 & n21858 ;
  assign n21860 = n21859 ^ n16088 ^ 1'b0 ;
  assign n21861 = n14152 ^ n7737 ^ 1'b0 ;
  assign n21862 = n7148 & n8902 ;
  assign n21863 = n5531 ^ n618 ^ 1'b0 ;
  assign n21864 = n21863 ^ n5479 ^ 1'b0 ;
  assign n21865 = n4883 | n11290 ;
  assign n21866 = n21864 & ~n21865 ;
  assign n21867 = n21862 & ~n21866 ;
  assign n21868 = ~n14703 & n21867 ;
  assign n21869 = n699 & ~n13476 ;
  assign n21870 = ~n1454 & n10615 ;
  assign n21872 = n3629 & ~n12534 ;
  assign n21873 = n13981 & n21872 ;
  assign n21874 = n21873 ^ n13060 ^ 1'b0 ;
  assign n21871 = n4301 & ~n5895 ;
  assign n21875 = n21874 ^ n21871 ^ 1'b0 ;
  assign n21876 = n15898 | n16728 ;
  assign n21877 = n4177 & ~n11282 ;
  assign n21878 = n5734 | n17922 ;
  assign n21879 = x159 & n1039 ;
  assign n21880 = n15863 & n21879 ;
  assign n21881 = n3866 & n7197 ;
  assign n21882 = n21881 ^ n11331 ^ 1'b0 ;
  assign n21883 = ( n819 & n14568 ) | ( n819 & ~n21882 ) | ( n14568 & ~n21882 ) ;
  assign n21884 = n10424 & ~n13026 ;
  assign n21886 = n2857 ^ n1491 ^ 1'b0 ;
  assign n21887 = n3481 | n21886 ;
  assign n21885 = ~n6508 & n8545 ;
  assign n21888 = n21887 ^ n21885 ^ 1'b0 ;
  assign n21889 = n12517 & n16307 ;
  assign n21890 = n21889 ^ n4105 ^ 1'b0 ;
  assign n21891 = n6813 & n21890 ;
  assign n21892 = n3235 & ~n9375 ;
  assign n21893 = n21892 ^ n5941 ^ 1'b0 ;
  assign n21894 = n3932 | n21893 ;
  assign n21895 = n21891 | n21894 ;
  assign n21896 = ~n4612 & n21895 ;
  assign n21897 = n2400 & n21896 ;
  assign n21898 = n21748 ^ n2076 ^ x195 ;
  assign n21899 = ( x187 & n7948 ) | ( x187 & ~n14109 ) | ( n7948 & ~n14109 ) ;
  assign n21900 = n6735 & ~n10331 ;
  assign n21901 = n21900 ^ n357 ^ 1'b0 ;
  assign n21902 = n13693 & ~n21901 ;
  assign n21903 = n21902 ^ n13608 ^ 1'b0 ;
  assign n21904 = n7128 & ~n13303 ;
  assign n21905 = n21904 ^ x1 ^ 1'b0 ;
  assign n21906 = n4130 | n9336 ;
  assign n21907 = n11983 | n21906 ;
  assign n21908 = n11337 ^ n8333 ^ 1'b0 ;
  assign n21909 = n8056 & ~n20435 ;
  assign n21910 = n21908 & ~n21909 ;
  assign n21911 = ~n12321 & n12857 ;
  assign n21912 = n12321 & n21911 ;
  assign n21913 = n16493 ^ n9225 ^ 1'b0 ;
  assign n21914 = ~n1086 & n14902 ;
  assign n21915 = n8277 & ~n20348 ;
  assign n21916 = n21915 ^ n404 ^ 1'b0 ;
  assign n21917 = n11055 | n21916 ;
  assign n21918 = n7263 & ~n12409 ;
  assign n21919 = n21917 | n21918 ;
  assign n21920 = n3582 | n8440 ;
  assign n21921 = n21919 & ~n21920 ;
  assign n21922 = ~n1398 & n5754 ;
  assign n21923 = n11186 & n17518 ;
  assign n21924 = n6818 & n21923 ;
  assign n21930 = ~n3076 & n9549 ;
  assign n21931 = n21930 ^ n338 ^ 1'b0 ;
  assign n21932 = ~n922 & n21931 ;
  assign n21933 = ~n21931 & n21932 ;
  assign n21925 = n5216 & n14499 ;
  assign n21926 = n5980 & n21925 ;
  assign n21927 = x100 & ~n886 ;
  assign n21928 = n4842 & n21927 ;
  assign n21929 = ( n9006 & ~n21926 ) | ( n9006 & n21928 ) | ( ~n21926 & n21928 ) ;
  assign n21934 = n21933 ^ n21929 ^ 1'b0 ;
  assign n21935 = n16829 | n21934 ;
  assign n21936 = n9329 ^ n7867 ^ 1'b0 ;
  assign n21937 = ( n4540 & n11701 ) | ( n4540 & n21936 ) | ( n11701 & n21936 ) ;
  assign n21938 = n4649 | n13271 ;
  assign n21939 = n4036 ^ n2716 ^ 1'b0 ;
  assign n21940 = n9067 ^ n3016 ^ 1'b0 ;
  assign n21941 = n2716 ^ n1647 ^ 1'b0 ;
  assign n21942 = n1770 & n21941 ;
  assign n21943 = n21942 ^ n9134 ^ 1'b0 ;
  assign n21944 = n19692 ^ n10636 ^ 1'b0 ;
  assign n21945 = n11185 | n17930 ;
  assign n21946 = n21944 | n21945 ;
  assign n21947 = n3453 & n21946 ;
  assign n21948 = n21943 & n21947 ;
  assign n21949 = ~n2281 & n6613 ;
  assign n21950 = ( n4562 & ~n6954 ) | ( n4562 & n14455 ) | ( ~n6954 & n14455 ) ;
  assign n21955 = n10995 ^ n1426 ^ 1'b0 ;
  assign n21956 = n3547 & ~n21955 ;
  assign n21957 = n20656 & n21956 ;
  assign n21958 = ~n20656 & n21957 ;
  assign n21954 = n6522 & ~n7942 ;
  assign n21959 = n21958 ^ n21954 ^ 1'b0 ;
  assign n21951 = n663 & n7472 ;
  assign n21952 = n21951 ^ n15906 ^ 1'b0 ;
  assign n21953 = n7220 & ~n21952 ;
  assign n21960 = n21959 ^ n21953 ^ 1'b0 ;
  assign n21961 = n2024 | n5301 ;
  assign n21962 = n21961 ^ n16250 ^ 1'b0 ;
  assign n21963 = ~n5462 & n9225 ;
  assign n21964 = n888 | n14887 ;
  assign n21965 = n21963 & ~n21964 ;
  assign n21966 = n21650 ^ n5806 ^ 1'b0 ;
  assign n21967 = n1856 | n4678 ;
  assign n21968 = ~n2809 & n21967 ;
  assign n21969 = n21968 ^ n19575 ^ 1'b0 ;
  assign n21970 = n9081 ^ n3614 ^ 1'b0 ;
  assign n21971 = n17478 ^ n4009 ^ 1'b0 ;
  assign n21972 = n5402 & ~n10713 ;
  assign n21973 = n21972 ^ n3161 ^ 1'b0 ;
  assign n21974 = ( ~n11624 & n15258 ) | ( ~n11624 & n21973 ) | ( n15258 & n21973 ) ;
  assign n21975 = n2900 & n15464 ;
  assign n21976 = n5732 & n21975 ;
  assign n21977 = n21976 ^ n3121 ^ 1'b0 ;
  assign n21978 = n18697 | n19273 ;
  assign n21979 = n11760 ^ n5796 ^ 1'b0 ;
  assign n21980 = n10015 | n21979 ;
  assign n21981 = n14862 & n20177 ;
  assign n21984 = n4985 ^ n4610 ^ n2520 ;
  assign n21982 = n6416 ^ n2358 ^ 1'b0 ;
  assign n21983 = n5859 & ~n21982 ;
  assign n21985 = n21984 ^ n21983 ^ 1'b0 ;
  assign n21986 = n16956 & ~n20866 ;
  assign n21987 = ~n840 & n21891 ;
  assign n21988 = n21987 ^ n20146 ^ 1'b0 ;
  assign n21989 = ~n3346 & n3395 ;
  assign n21990 = n2948 ^ n466 ^ 1'b0 ;
  assign n21991 = n21990 ^ n8333 ^ n742 ;
  assign n21992 = n2262 & ~n7147 ;
  assign n21993 = n21992 ^ n7261 ^ 1'b0 ;
  assign n21994 = n12569 ^ n8818 ^ n6311 ;
  assign n21995 = n21993 & ~n21994 ;
  assign n21996 = n15196 & ~n21995 ;
  assign n21997 = ~n3509 & n21996 ;
  assign n21998 = n4367 | n5229 ;
  assign n21999 = n21998 ^ n1204 ^ 1'b0 ;
  assign n22000 = n10149 & ~n21999 ;
  assign n22001 = n12714 & n22000 ;
  assign n22002 = n12446 ^ n3256 ^ 1'b0 ;
  assign n22003 = n22001 | n22002 ;
  assign n22004 = n10180 | n11683 ;
  assign n22005 = n7732 & n12002 ;
  assign n22006 = n1330 | n6410 ;
  assign n22007 = n4584 ^ n3215 ^ 1'b0 ;
  assign n22008 = n22006 & n22007 ;
  assign n22009 = ~n12605 & n13828 ;
  assign n22010 = n12050 | n12730 ;
  assign n22011 = n5033 ^ n3615 ^ 1'b0 ;
  assign n22012 = n1577 | n22011 ;
  assign n22013 = n4874 | n6746 ;
  assign n22014 = n22013 ^ n5277 ^ 1'b0 ;
  assign n22015 = n12555 ^ n637 ^ 1'b0 ;
  assign n22016 = n22015 ^ x102 ^ 1'b0 ;
  assign n22017 = n3329 ^ n1871 ^ 1'b0 ;
  assign n22018 = ~n22016 & n22017 ;
  assign n22019 = ~n2968 & n4248 ;
  assign n22020 = n20267 & n22019 ;
  assign n22021 = n22020 ^ n4642 ^ 1'b0 ;
  assign n22022 = n22021 ^ n2411 ^ 1'b0 ;
  assign n22023 = n5252 | n22022 ;
  assign n22024 = n13720 ^ n10604 ^ n638 ;
  assign n22025 = n1660 & ~n5481 ;
  assign n22026 = n22025 ^ n9438 ^ 1'b0 ;
  assign n22027 = n22026 ^ n4933 ^ 1'b0 ;
  assign n22028 = n1186 & ~n6750 ;
  assign n22029 = n11262 ^ x176 ^ 1'b0 ;
  assign n22030 = ~n14089 & n17919 ;
  assign n22031 = n6465 & ~n14565 ;
  assign n22032 = n4266 & ~n10974 ;
  assign n22033 = n22032 ^ n420 ^ 1'b0 ;
  assign n22034 = ~n13437 & n22033 ;
  assign n22035 = n14605 & n22034 ;
  assign n22036 = n9816 ^ n2411 ^ 1'b0 ;
  assign n22037 = n22035 | n22036 ;
  assign n22038 = n14379 & ~n19767 ;
  assign n22039 = n22038 ^ n9971 ^ 1'b0 ;
  assign n22040 = n13773 ^ n10484 ^ 1'b0 ;
  assign n22041 = n12380 & n22040 ;
  assign n22042 = ~n10834 & n22041 ;
  assign n22043 = ~n8018 & n22042 ;
  assign n22044 = ~n18278 & n20613 ;
  assign n22045 = ~n963 & n15515 ;
  assign n22046 = n22045 ^ n8863 ^ 1'b0 ;
  assign n22047 = n22044 & ~n22046 ;
  assign n22048 = ( n2349 & n8143 ) | ( n2349 & ~n16153 ) | ( n8143 & ~n16153 ) ;
  assign n22049 = n16346 | n22048 ;
  assign n22050 = n10039 ^ n9357 ^ 1'b0 ;
  assign n22051 = n395 & n2255 ;
  assign n22052 = n22051 ^ n3202 ^ 1'b0 ;
  assign n22053 = ~n11976 & n22052 ;
  assign n22054 = x134 & ~n22053 ;
  assign n22055 = n14486 | n22054 ;
  assign n22056 = n14282 & n22055 ;
  assign n22057 = n22056 ^ x181 ^ 1'b0 ;
  assign n22058 = n7405 | n19430 ;
  assign n22059 = x195 & ~n22058 ;
  assign n22060 = n6844 & ~n22059 ;
  assign n22061 = n1723 & ~n3016 ;
  assign n22062 = ~n1723 & n22061 ;
  assign n22063 = n15055 | n22062 ;
  assign n22064 = n466 & n7174 ;
  assign n22065 = n22064 ^ n5498 ^ 1'b0 ;
  assign n22066 = n6770 & ~n22065 ;
  assign n22067 = ~n16695 & n22066 ;
  assign n22068 = n22063 & n22067 ;
  assign n22069 = n4038 & ~n7581 ;
  assign n22070 = n3234 | n20933 ;
  assign n22071 = n22070 ^ n20392 ^ 1'b0 ;
  assign n22072 = n4460 & n14529 ;
  assign n22073 = n6138 & ~n13423 ;
  assign n22074 = ( n1021 & n4677 ) | ( n1021 & ~n13568 ) | ( n4677 & ~n13568 ) ;
  assign n22075 = n8850 | n22074 ;
  assign n22076 = n574 & ~n7577 ;
  assign n22077 = n571 & ~n22076 ;
  assign n22078 = ~n1738 & n10960 ;
  assign n22079 = n14788 & n22078 ;
  assign n22081 = n6842 ^ n6604 ^ 1'b0 ;
  assign n22082 = n709 | n22081 ;
  assign n22080 = ~n5034 & n7513 ;
  assign n22083 = n22082 ^ n22080 ^ 1'b0 ;
  assign n22084 = n8495 & ~n8895 ;
  assign n22085 = n13245 ^ n7778 ^ 1'b0 ;
  assign n22086 = n22085 ^ n9043 ^ 1'b0 ;
  assign n22087 = n22084 & n22086 ;
  assign n22088 = n17887 | n22087 ;
  assign n22089 = n9224 ^ n6242 ^ 1'b0 ;
  assign n22090 = ~n4430 & n22089 ;
  assign n22091 = n3643 | n12634 ;
  assign n22092 = n22091 ^ n6920 ^ 1'b0 ;
  assign n22093 = n18651 ^ n16521 ^ 1'b0 ;
  assign n22094 = n11801 & ~n22093 ;
  assign n22095 = n15878 ^ n5797 ^ 1'b0 ;
  assign n22096 = n3571 & n7275 ;
  assign n22097 = ~n298 & n22096 ;
  assign n22098 = n20819 ^ n10291 ^ 1'b0 ;
  assign n22099 = ~n14494 & n22098 ;
  assign n22100 = n5333 ^ n1389 ^ 1'b0 ;
  assign n22101 = n1261 | n22100 ;
  assign n22102 = n22101 ^ n20747 ^ 1'b0 ;
  assign n22103 = n22099 & n22102 ;
  assign n22104 = ~n5182 & n22103 ;
  assign n22105 = n7170 ^ n3581 ^ 1'b0 ;
  assign n22106 = n6534 & n22105 ;
  assign n22107 = n17690 ^ x176 ^ 1'b0 ;
  assign n22108 = n7295 & ~n22107 ;
  assign n22109 = n22106 & n22108 ;
  assign n22110 = n14852 & ~n17728 ;
  assign n22111 = n22110 ^ n5437 ^ 1'b0 ;
  assign n22112 = n6731 | n7813 ;
  assign n22113 = n22112 ^ n2715 ^ 1'b0 ;
  assign n22114 = n4665 & n22113 ;
  assign n22115 = n10805 ^ x229 ^ 1'b0 ;
  assign n22116 = n21700 | n22115 ;
  assign n22117 = n22116 ^ n10059 ^ n2572 ;
  assign n22118 = n14729 & ~n22117 ;
  assign n22119 = n22118 ^ n3067 ^ 1'b0 ;
  assign n22120 = ~n6343 & n14347 ;
  assign n22121 = n22120 ^ n14865 ^ 1'b0 ;
  assign n22122 = n13125 & n20241 ;
  assign n22123 = n6555 ^ n6518 ^ 1'b0 ;
  assign n22124 = n5507 & n22123 ;
  assign n22125 = ~n18794 & n19712 ;
  assign n22126 = n22125 ^ n16969 ^ 1'b0 ;
  assign n22127 = n10702 & ~n10724 ;
  assign n22128 = n22127 ^ n20914 ^ 1'b0 ;
  assign n22129 = ~n2165 & n7597 ;
  assign n22130 = n12989 & n17912 ;
  assign n22131 = n22129 & n22130 ;
  assign n22132 = n4762 | n16135 ;
  assign n22133 = n22132 ^ n9365 ^ 1'b0 ;
  assign n22134 = n6417 ^ n4807 ^ 1'b0 ;
  assign n22135 = n10150 & n22134 ;
  assign n22136 = n22135 ^ n10209 ^ 1'b0 ;
  assign n22137 = n13861 & ~n22136 ;
  assign n22138 = n14666 ^ n10532 ^ n4571 ;
  assign n22139 = n9429 ^ n3032 ^ 1'b0 ;
  assign n22140 = n1997 | n22139 ;
  assign n22141 = n19347 ^ n17441 ^ 1'b0 ;
  assign n22142 = n3606 | n13176 ;
  assign n22143 = n9444 ^ n4470 ^ 1'b0 ;
  assign n22144 = n7349 & n22143 ;
  assign n22145 = n6965 | n22144 ;
  assign n22146 = n22145 ^ n1170 ^ 1'b0 ;
  assign n22147 = n2034 | n2821 ;
  assign n22148 = ~n11563 & n22147 ;
  assign n22149 = n8984 & n22148 ;
  assign n22150 = ~n22146 & n22149 ;
  assign n22151 = n5763 & ~n7902 ;
  assign n22152 = n20835 ^ n15059 ^ 1'b0 ;
  assign n22153 = n8519 ^ n5163 ^ 1'b0 ;
  assign n22156 = n5140 & n10865 ;
  assign n22157 = n22156 ^ n21647 ^ 1'b0 ;
  assign n22158 = n3557 & ~n22157 ;
  assign n22159 = n20527 & ~n22158 ;
  assign n22154 = n14514 ^ n4553 ^ 1'b0 ;
  assign n22155 = ~n5034 & n22154 ;
  assign n22160 = n22159 ^ n22155 ^ 1'b0 ;
  assign n22161 = n22153 & ~n22160 ;
  assign n22162 = n7873 ^ x218 ^ 1'b0 ;
  assign n22163 = n17643 | n22162 ;
  assign n22164 = n4443 & n9852 ;
  assign n22165 = n22163 & n22164 ;
  assign n22166 = ~n3771 & n19763 ;
  assign n22167 = ~n860 & n22166 ;
  assign n22168 = n1525 & ~n15278 ;
  assign n22170 = n15227 ^ n9225 ^ 1'b0 ;
  assign n22169 = ~n9589 & n12115 ;
  assign n22171 = n22170 ^ n22169 ^ 1'b0 ;
  assign n22172 = n3626 & ~n17815 ;
  assign n22173 = ( ~n1674 & n2383 ) | ( ~n1674 & n8584 ) | ( n2383 & n8584 ) ;
  assign n22174 = n22173 ^ n2464 ^ 1'b0 ;
  assign n22176 = n9664 ^ n4038 ^ 1'b0 ;
  assign n22177 = n11297 & ~n13620 ;
  assign n22178 = n5248 & n22177 ;
  assign n22179 = ~n22176 & n22178 ;
  assign n22175 = n5978 & ~n7674 ;
  assign n22180 = n22179 ^ n22175 ^ 1'b0 ;
  assign n22181 = n17872 ^ n16606 ^ n1103 ;
  assign n22184 = x247 & n14617 ;
  assign n22185 = n8662 & n22184 ;
  assign n22182 = ~x31 & n13303 ;
  assign n22183 = n16543 & ~n22182 ;
  assign n22186 = n22185 ^ n22183 ^ 1'b0 ;
  assign n22187 = n6514 ^ n3431 ^ 1'b0 ;
  assign n22188 = ( n8945 & n20878 ) | ( n8945 & n22187 ) | ( n20878 & n22187 ) ;
  assign n22190 = n5316 ^ x84 ^ 1'b0 ;
  assign n22189 = n8838 & n12517 ;
  assign n22191 = n22190 ^ n22189 ^ 1'b0 ;
  assign n22192 = n16920 ^ n15473 ^ 1'b0 ;
  assign n22193 = n4325 & n11170 ;
  assign n22194 = ( n16614 & n22192 ) | ( n16614 & n22193 ) | ( n22192 & n22193 ) ;
  assign n22195 = n4871 | n9149 ;
  assign n22196 = x124 | n22195 ;
  assign n22197 = n5690 & n10731 ;
  assign n22198 = n2528 & n22197 ;
  assign n22199 = n8557 ^ n6155 ^ 1'b0 ;
  assign n22200 = n14206 | n15733 ;
  assign n22201 = n7089 | n22200 ;
  assign n22202 = ~n22199 & n22201 ;
  assign n22203 = n22202 ^ n14398 ^ n2075 ;
  assign n22204 = ( ~x45 & n6789 ) | ( ~x45 & n12610 ) | ( n6789 & n12610 ) ;
  assign n22205 = n22204 ^ n14578 ^ 1'b0 ;
  assign n22206 = n22205 ^ n3207 ^ 1'b0 ;
  assign n22207 = n4629 ^ n2406 ^ 1'b0 ;
  assign n22208 = ( n3639 & n9302 ) | ( n3639 & n22207 ) | ( n9302 & n22207 ) ;
  assign n22209 = n16943 | n20898 ;
  assign n22210 = n9792 | n22209 ;
  assign n22211 = n16170 ^ n7873 ^ 1'b0 ;
  assign n22212 = n5650 | n12935 ;
  assign n22213 = n22212 ^ n5769 ^ 1'b0 ;
  assign n22214 = n12342 & ~n22213 ;
  assign n22215 = ~n17562 & n22214 ;
  assign n22216 = n20516 | n20896 ;
  assign n22217 = n22216 ^ n3680 ^ 1'b0 ;
  assign n22218 = n17483 ^ n10731 ^ 1'b0 ;
  assign n22219 = n22217 | n22218 ;
  assign n22220 = n22069 & ~n22219 ;
  assign n22221 = x55 & n6083 ;
  assign n22222 = n5898 & ~n21949 ;
  assign n22223 = n22222 ^ n4247 ^ 1'b0 ;
  assign n22225 = n19963 ^ n7092 ^ 1'b0 ;
  assign n22224 = n5513 & ~n17643 ;
  assign n22226 = n22225 ^ n22224 ^ 1'b0 ;
  assign n22227 = n7109 & ~n8963 ;
  assign n22228 = n22227 ^ n6654 ^ 1'b0 ;
  assign n22229 = ~n6027 & n22228 ;
  assign n22230 = n1279 & n22229 ;
  assign n22231 = n5729 & ~n6678 ;
  assign n22232 = n22231 ^ n11041 ^ 1'b0 ;
  assign n22233 = n22232 ^ n14398 ^ 1'b0 ;
  assign n22234 = n1021 | n1284 ;
  assign n22235 = n5557 | n22234 ;
  assign n22236 = n2901 | n22235 ;
  assign n22237 = n21738 & ~n22236 ;
  assign n22238 = ( n3868 & ~n14463 ) | ( n3868 & n22237 ) | ( ~n14463 & n22237 ) ;
  assign n22239 = n20481 ^ n10534 ^ n8785 ;
  assign n22240 = n11118 ^ n585 ^ 1'b0 ;
  assign n22241 = ~n19709 & n22240 ;
  assign n22242 = n22241 ^ n8634 ^ 1'b0 ;
  assign n22250 = n12058 & ~n12870 ;
  assign n22243 = n14516 ^ n5328 ^ 1'b0 ;
  assign n22244 = n3915 ^ x61 ^ 1'b0 ;
  assign n22245 = ~n4352 & n22244 ;
  assign n22246 = n4036 & n22245 ;
  assign n22247 = n22246 ^ n15544 ^ 1'b0 ;
  assign n22248 = n22247 ^ n11909 ^ 1'b0 ;
  assign n22249 = n22243 & ~n22248 ;
  assign n22251 = n22250 ^ n22249 ^ 1'b0 ;
  assign n22252 = n11734 ^ n7674 ^ 1'b0 ;
  assign n22253 = n11379 | n22252 ;
  assign n22254 = ( n10309 & n13524 ) | ( n10309 & n22253 ) | ( n13524 & n22253 ) ;
  assign n22255 = n2112 ^ x43 ^ 1'b0 ;
  assign n22256 = x61 & ~n22255 ;
  assign n22257 = n2613 | n5119 ;
  assign n22258 = n22256 | n22257 ;
  assign n22259 = n15469 ^ n9207 ^ 1'b0 ;
  assign n22260 = n20930 | n22259 ;
  assign n22261 = n2180 & ~n4624 ;
  assign n22262 = n22261 ^ n5900 ^ 1'b0 ;
  assign n22263 = n8011 ^ n4450 ^ 1'b0 ;
  assign n22264 = n6391 & ~n22263 ;
  assign n22265 = n22264 ^ n9507 ^ n4559 ;
  assign n22266 = n9336 ^ n9001 ^ n8974 ;
  assign n22267 = ( n22262 & ~n22265 ) | ( n22262 & n22266 ) | ( ~n22265 & n22266 ) ;
  assign n22268 = n781 & n4345 ;
  assign n22269 = ~n1471 & n19813 ;
  assign n22270 = n22269 ^ n6391 ^ 1'b0 ;
  assign n22271 = n2879 & ~n16424 ;
  assign n22272 = n22271 ^ n1182 ^ 1'b0 ;
  assign n22273 = n2215 & ~n22272 ;
  assign n22274 = n22273 ^ n13144 ^ n10169 ;
  assign n22275 = n11076 ^ n6994 ^ 1'b0 ;
  assign n22276 = n22275 ^ n17438 ^ n12029 ;
  assign n22277 = n22276 ^ n19319 ^ 1'b0 ;
  assign n22278 = x56 & ~n15240 ;
  assign n22279 = n22277 & ~n22278 ;
  assign n22280 = n7664 & n10606 ;
  assign n22281 = n22280 ^ n7652 ^ 1'b0 ;
  assign n22282 = n22281 ^ n3855 ^ 1'b0 ;
  assign n22283 = n18915 ^ n7168 ^ 1'b0 ;
  assign n22284 = n19330 ^ n6737 ^ 1'b0 ;
  assign n22285 = n6679 & ~n22284 ;
  assign n22286 = n4367 ^ n2618 ^ 1'b0 ;
  assign n22287 = n8581 & n22286 ;
  assign n22288 = n8638 & ~n22287 ;
  assign n22289 = x91 & ~n21515 ;
  assign n22290 = n22289 ^ x204 ^ 1'b0 ;
  assign n22292 = n13725 ^ n12124 ^ 1'b0 ;
  assign n22293 = n9928 | n22292 ;
  assign n22291 = ~n7359 & n19028 ;
  assign n22294 = n22293 ^ n22291 ^ 1'b0 ;
  assign n22295 = n498 | n4413 ;
  assign n22296 = n10001 & n22295 ;
  assign n22297 = n10719 & n22296 ;
  assign n22298 = n14392 & n22297 ;
  assign n22299 = n20406 ^ n17043 ^ n12554 ;
  assign n22300 = n11749 & n22299 ;
  assign n22301 = n3337 & n22300 ;
  assign n22302 = n20073 & n21507 ;
  assign n22303 = n22302 ^ n20766 ^ 1'b0 ;
  assign n22304 = n10552 ^ x180 ^ 1'b0 ;
  assign n22305 = n4878 | n22304 ;
  assign n22307 = n19966 ^ n6421 ^ 1'b0 ;
  assign n22306 = n16408 ^ n13293 ^ 1'b0 ;
  assign n22308 = n22307 ^ n22306 ^ 1'b0 ;
  assign n22309 = n18518 ^ n3817 ^ 1'b0 ;
  assign n22310 = n8252 & ~n13738 ;
  assign n22311 = ~n376 & n22310 ;
  assign n22312 = ~n7476 & n22311 ;
  assign n22313 = n22312 ^ n15999 ^ 1'b0 ;
  assign n22314 = ~n12592 & n22313 ;
  assign n22315 = ~n5560 & n11262 ;
  assign n22316 = n22315 ^ n2447 ^ 1'b0 ;
  assign n22317 = ~n15839 & n22316 ;
  assign n22318 = n5055 & n5497 ;
  assign n22319 = n3674 & n22318 ;
  assign n22320 = ~n22317 & n22319 ;
  assign n22321 = n11056 ^ n4677 ^ n2992 ;
  assign n22322 = n22321 ^ n9527 ^ 1'b0 ;
  assign n22323 = n21682 | n22322 ;
  assign n22324 = n1353 & n3142 ;
  assign n22325 = n22324 ^ n20361 ^ 1'b0 ;
  assign n22326 = ~n17710 & n22325 ;
  assign n22327 = n4647 & ~n10229 ;
  assign n22328 = ( n2950 & n11114 ) | ( n2950 & n19972 ) | ( n11114 & n19972 ) ;
  assign n22329 = n2482 & n20659 ;
  assign n22330 = ~n12736 & n18453 ;
  assign n22331 = ~n1065 & n22330 ;
  assign n22332 = ( n1103 & n7557 ) | ( n1103 & n7742 ) | ( n7557 & n7742 ) ;
  assign n22333 = n5243 & n22332 ;
  assign n22334 = n7266 ^ n5317 ^ 1'b0 ;
  assign n22335 = n22334 ^ n1397 ^ 1'b0 ;
  assign n22337 = n11450 & n18741 ;
  assign n22338 = ~n20956 & n22337 ;
  assign n22339 = n8254 | n22338 ;
  assign n22336 = n12632 ^ n11024 ^ 1'b0 ;
  assign n22340 = n22339 ^ n22336 ^ 1'b0 ;
  assign n22341 = ~n2696 & n22340 ;
  assign n22342 = n9706 ^ n8244 ^ 1'b0 ;
  assign n22343 = ~n5353 & n22342 ;
  assign n22344 = ~n6414 & n22343 ;
  assign n22345 = n15414 | n22344 ;
  assign n22346 = n22345 ^ n1841 ^ 1'b0 ;
  assign n22347 = n2188 | n10273 ;
  assign n22348 = n22347 ^ n14739 ^ 1'b0 ;
  assign n22349 = n15838 & ~n22348 ;
  assign n22350 = ~n9064 & n22349 ;
  assign n22351 = n3771 & n22350 ;
  assign n22352 = n14842 ^ n1723 ^ 1'b0 ;
  assign n22353 = n4347 & n22352 ;
  assign n22354 = n12924 | n22353 ;
  assign n22355 = n20701 ^ n17543 ^ n5474 ;
  assign n22356 = n5413 & ~n10135 ;
  assign n22357 = n22356 ^ n10937 ^ 1'b0 ;
  assign n22358 = n3797 & ~n22357 ;
  assign n22359 = n22358 ^ n14256 ^ 1'b0 ;
  assign n22360 = n7903 & n14160 ;
  assign n22361 = n12288 & ~n16237 ;
  assign n22362 = n22361 ^ n15150 ^ 1'b0 ;
  assign n22363 = n2687 & ~n19532 ;
  assign n22364 = n5967 | n9614 ;
  assign n22365 = n2556 | n22364 ;
  assign n22366 = n7880 & n22365 ;
  assign n22367 = n9611 & n22366 ;
  assign n22368 = n14752 ^ n375 ^ 1'b0 ;
  assign n22369 = ~n12922 & n22368 ;
  assign n22370 = n6187 & ~n9958 ;
  assign n22371 = n22370 ^ n711 ^ 1'b0 ;
  assign n22372 = x101 & ~n15279 ;
  assign n22373 = n2701 | n12218 ;
  assign n22374 = n16663 & ~n22373 ;
  assign n22375 = n12414 ^ n1680 ^ 1'b0 ;
  assign n22376 = n21360 ^ n20389 ^ 1'b0 ;
  assign n22377 = ~n992 & n6453 ;
  assign n22378 = n22377 ^ n12359 ^ 1'b0 ;
  assign n22379 = n22378 ^ n18812 ^ 1'b0 ;
  assign n22380 = n20330 ^ n10407 ^ 1'b0 ;
  assign n22381 = n2035 & ~n22380 ;
  assign n22382 = n8039 & n22381 ;
  assign n22383 = n22382 ^ n8725 ^ 1'b0 ;
  assign n22384 = n4839 & n14645 ;
  assign n22385 = n16421 & n22384 ;
  assign n22386 = n5349 & n8125 ;
  assign n22387 = n22386 ^ n20595 ^ 1'b0 ;
  assign n22388 = n20845 ^ n11105 ^ 1'b0 ;
  assign n22389 = ~x196 & n19765 ;
  assign n22390 = n22389 ^ n7609 ^ 1'b0 ;
  assign n22391 = n18364 ^ n15689 ^ 1'b0 ;
  assign n22392 = ~n3908 & n22391 ;
  assign n22393 = n22392 ^ n7619 ^ 1'b0 ;
  assign n22394 = ~n3186 & n11440 ;
  assign n22395 = n4070 & ~n18856 ;
  assign n22396 = n22395 ^ n17985 ^ 1'b0 ;
  assign n22397 = x178 | n5912 ;
  assign n22398 = n22397 ^ n7223 ^ 1'b0 ;
  assign n22399 = n22398 ^ n11901 ^ n6257 ;
  assign n22400 = n7603 & n22399 ;
  assign n22401 = n22396 & n22400 ;
  assign n22402 = n11170 ^ n7328 ^ 1'b0 ;
  assign n22403 = x172 & n22402 ;
  assign n22404 = n22403 ^ n11007 ^ 1'b0 ;
  assign n22405 = n21523 ^ n8766 ^ 1'b0 ;
  assign n22406 = n14895 ^ n8841 ^ n5188 ;
  assign n22407 = n842 | n22406 ;
  assign n22408 = n22407 ^ n12262 ^ 1'b0 ;
  assign n22409 = n1547 & ~n10929 ;
  assign n22410 = n18551 ^ n5908 ^ 1'b0 ;
  assign n22411 = n22410 ^ n16203 ^ 1'b0 ;
  assign n22412 = n22411 ^ n8007 ^ n535 ;
  assign n22413 = n11957 ^ n8321 ^ 1'b0 ;
  assign n22414 = n22412 & n22413 ;
  assign n22415 = n7340 | n22233 ;
  assign n22416 = n4267 & ~n22415 ;
  assign n22417 = n12325 ^ n3982 ^ n1077 ;
  assign n22418 = n5723 & n10242 ;
  assign n22419 = n2657 & n22418 ;
  assign n22420 = n22417 | n22419 ;
  assign n22421 = n22420 ^ n7271 ^ 1'b0 ;
  assign n22422 = ~n8251 & n18011 ;
  assign n22424 = ~n10726 & n11381 ;
  assign n22425 = ~n1634 & n22424 ;
  assign n22423 = n9359 & n14765 ;
  assign n22426 = n22425 ^ n22423 ^ 1'b0 ;
  assign n22427 = n22422 & n22426 ;
  assign n22428 = n11462 & n13239 ;
  assign n22429 = n16300 ^ n2231 ^ 1'b0 ;
  assign n22430 = n10062 & ~n22429 ;
  assign n22431 = n15777 ^ n11331 ^ 1'b0 ;
  assign n22432 = n2939 | n22431 ;
  assign n22434 = n11295 ^ n3837 ^ 1'b0 ;
  assign n22435 = n4562 & n22434 ;
  assign n22433 = n784 & n11127 ;
  assign n22436 = n22435 ^ n22433 ^ 1'b0 ;
  assign n22437 = n22432 | n22436 ;
  assign n22438 = n22437 ^ n16657 ^ 1'b0 ;
  assign n22439 = ~n2646 & n9054 ;
  assign n22440 = n22439 ^ n8446 ^ 1'b0 ;
  assign n22441 = n3255 | n22440 ;
  assign n22442 = ~n274 & n619 ;
  assign n22443 = n22442 ^ n21701 ^ n4703 ;
  assign n22444 = n5748 ^ x45 ^ 1'b0 ;
  assign n22445 = n6526 & n22444 ;
  assign n22446 = n22445 ^ n9659 ^ 1'b0 ;
  assign n22447 = n1500 & n22446 ;
  assign n22448 = x40 & ~n13476 ;
  assign n22449 = n22448 ^ n7968 ^ 1'b0 ;
  assign n22450 = n5452 ^ n831 ^ 1'b0 ;
  assign n22451 = n21882 & ~n22450 ;
  assign n22453 = x96 & n817 ;
  assign n22454 = ~x96 & n22453 ;
  assign n22455 = n1554 | n22454 ;
  assign n22456 = n1554 & ~n22455 ;
  assign n22457 = n705 & ~n22456 ;
  assign n22458 = n22457 ^ n1730 ^ 1'b0 ;
  assign n22452 = n4740 & n8289 ;
  assign n22459 = n22458 ^ n22452 ^ 1'b0 ;
  assign n22460 = x13 & ~n22459 ;
  assign n22461 = n2609 & ~n22460 ;
  assign n22462 = n4040 & ~n4708 ;
  assign n22463 = n8503 & n18948 ;
  assign n22464 = n10162 & n18410 ;
  assign n22465 = n1474 | n9255 ;
  assign n22466 = n10097 | n22465 ;
  assign n22467 = n14546 ^ n9401 ^ n3729 ;
  assign n22468 = ~n608 & n22467 ;
  assign n22469 = n15326 ^ n10146 ^ 1'b0 ;
  assign n22470 = n5223 | n22469 ;
  assign n22471 = n12022 | n22470 ;
  assign n22473 = n4827 & ~n21487 ;
  assign n22474 = n22473 ^ n11703 ^ 1'b0 ;
  assign n22475 = n22474 ^ n17091 ^ 1'b0 ;
  assign n22476 = ~n14359 & n22475 ;
  assign n22472 = n638 | n14009 ;
  assign n22477 = n22476 ^ n22472 ^ 1'b0 ;
  assign n22478 = n10014 ^ n9698 ^ 1'b0 ;
  assign n22479 = n4742 & n22478 ;
  assign n22480 = n5016 & n22479 ;
  assign n22481 = n22480 ^ n15405 ^ 1'b0 ;
  assign n22482 = n22477 & n22481 ;
  assign n22484 = n8584 | n12218 ;
  assign n22485 = n8919 | n22484 ;
  assign n22483 = n3868 | n16794 ;
  assign n22486 = n22485 ^ n22483 ^ n20625 ;
  assign n22487 = n4657 | n18088 ;
  assign n22488 = n22487 ^ n11316 ^ 1'b0 ;
  assign n22489 = ~n7999 & n22488 ;
  assign n22490 = n11459 & n20927 ;
  assign n22491 = ( n5413 & ~n8863 ) | ( n5413 & n22490 ) | ( ~n8863 & n22490 ) ;
  assign n22492 = n920 | n8980 ;
  assign n22493 = n5839 ^ n4502 ^ 1'b0 ;
  assign n22494 = n22493 ^ n16017 ^ 1'b0 ;
  assign n22495 = ~x46 & n3197 ;
  assign n22496 = n871 & ~n20249 ;
  assign n22497 = ~n7934 & n8322 ;
  assign n22498 = n5429 | n15783 ;
  assign n22499 = n10215 | n15387 ;
  assign n22500 = n16682 & ~n22499 ;
  assign n22501 = n22500 ^ n9580 ^ 1'b0 ;
  assign n22502 = n6711 ^ n2903 ^ 1'b0 ;
  assign n22503 = n836 & n22502 ;
  assign n22504 = n6483 & n22503 ;
  assign n22505 = n8378 & ~n14555 ;
  assign n22506 = n6331 & ~n22505 ;
  assign n22507 = n21468 ^ n9783 ^ 1'b0 ;
  assign n22508 = n16703 | n21048 ;
  assign n22509 = n11981 & ~n22508 ;
  assign n22510 = ~n11981 & n22509 ;
  assign n22513 = x43 & n1230 ;
  assign n22514 = ~n1230 & n22513 ;
  assign n22515 = n4840 | n22514 ;
  assign n22511 = n3506 & n21361 ;
  assign n22512 = n22511 ^ n1608 ^ 1'b0 ;
  assign n22516 = n22515 ^ n22512 ^ 1'b0 ;
  assign n22517 = ~n22510 & n22516 ;
  assign n22518 = n7586 ^ n6483 ^ 1'b0 ;
  assign n22519 = n22518 ^ n5138 ^ n4215 ;
  assign n22521 = n5497 & n20743 ;
  assign n22520 = ~n497 & n13896 ;
  assign n22522 = n22521 ^ n22520 ^ 1'b0 ;
  assign n22523 = n17526 ^ n14448 ^ n871 ;
  assign n22524 = n22523 ^ n12487 ^ 1'b0 ;
  assign n22525 = n5576 & n22524 ;
  assign n22526 = n8103 ^ n2184 ^ 1'b0 ;
  assign n22527 = n22418 ^ x12 ^ 1'b0 ;
  assign n22528 = n3509 | n22527 ;
  assign n22529 = n14760 ^ n12515 ^ 1'b0 ;
  assign n22530 = ~n3780 & n4757 ;
  assign n22531 = ~n11602 & n19975 ;
  assign n22532 = ~n11769 & n22531 ;
  assign n22533 = n9803 | n22532 ;
  assign n22534 = n22530 & ~n22533 ;
  assign n22535 = n2697 & n20764 ;
  assign n22536 = ( ~n6655 & n22534 ) | ( ~n6655 & n22535 ) | ( n22534 & n22535 ) ;
  assign n22544 = n10247 & ~n19416 ;
  assign n22537 = n1300 ^ n1100 ^ 1'b0 ;
  assign n22538 = n22537 ^ n1966 ^ 1'b0 ;
  assign n22539 = ( n617 & ~n11730 ) | ( n617 & n22538 ) | ( ~n11730 & n22538 ) ;
  assign n22540 = n5091 ^ n3074 ^ 1'b0 ;
  assign n22541 = x40 | n22540 ;
  assign n22542 = n10040 & n22541 ;
  assign n22543 = n22539 & ~n22542 ;
  assign n22545 = n22544 ^ n22543 ^ 1'b0 ;
  assign n22547 = n22442 ^ n14267 ^ n11049 ;
  assign n22548 = n20896 | n22547 ;
  assign n22546 = ~n12643 & n17029 ;
  assign n22549 = n22548 ^ n22546 ^ 1'b0 ;
  assign n22551 = n5856 ^ x86 ^ 1'b0 ;
  assign n22550 = ~n2248 & n17566 ;
  assign n22552 = n22551 ^ n22550 ^ 1'b0 ;
  assign n22553 = ~n7065 & n18482 ;
  assign n22554 = n22553 ^ x155 ^ 1'b0 ;
  assign n22557 = ~n606 & n2620 ;
  assign n22555 = n4107 & n14681 ;
  assign n22556 = n22555 ^ n11683 ^ 1'b0 ;
  assign n22558 = n22557 ^ n22556 ^ 1'b0 ;
  assign n22559 = n22558 ^ n21714 ^ n4222 ;
  assign n22560 = n15416 & ~n17633 ;
  assign n22561 = n3416 & n13502 ;
  assign n22562 = n22561 ^ n1696 ^ 1'b0 ;
  assign n22563 = ( n11436 & n15739 ) | ( n11436 & n21008 ) | ( n15739 & n21008 ) ;
  assign n22564 = ~n13714 & n22563 ;
  assign n22565 = n8927 & n11974 ;
  assign n22566 = n2622 | n5625 ;
  assign n22567 = n11337 | n22566 ;
  assign n22568 = n20888 & n21834 ;
  assign n22569 = n9412 & n22568 ;
  assign n22570 = n645 | n22569 ;
  assign n22571 = n22570 ^ n6415 ^ 1'b0 ;
  assign n22572 = n8236 ^ n2986 ^ 1'b0 ;
  assign n22573 = n17730 & n22572 ;
  assign n22574 = n7552 & n22573 ;
  assign n22575 = x135 & ~n6301 ;
  assign n22576 = n22575 ^ n17091 ^ 1'b0 ;
  assign n22577 = ~n583 & n11041 ;
  assign n22578 = ~n13452 & n22577 ;
  assign n22581 = ( ~n8690 & n9715 ) | ( ~n8690 & n12864 ) | ( n9715 & n12864 ) ;
  assign n22579 = n4865 ^ n2338 ^ x213 ;
  assign n22580 = n3421 & n22579 ;
  assign n22582 = n22581 ^ n22580 ^ 1'b0 ;
  assign n22583 = n8559 & n22582 ;
  assign n22584 = ~n1324 & n22583 ;
  assign n22585 = n11696 ^ n8042 ^ 1'b0 ;
  assign n22586 = n21258 & n22585 ;
  assign n22587 = ( n2702 & n8155 ) | ( n2702 & ~n11901 ) | ( n8155 & ~n11901 ) ;
  assign n22588 = n5754 ^ n4989 ^ 1'b0 ;
  assign n22589 = n22587 & ~n22588 ;
  assign n22590 = n5851 | n11863 ;
  assign n22591 = n22590 ^ n1589 ^ 1'b0 ;
  assign n22592 = n7428 ^ n6534 ^ 1'b0 ;
  assign n22593 = ~n3946 & n22592 ;
  assign n22594 = n22593 ^ n13515 ^ 1'b0 ;
  assign n22595 = n2743 ^ n451 ^ 1'b0 ;
  assign n22596 = n7813 | n22595 ;
  assign n22597 = n22596 ^ n10402 ^ 1'b0 ;
  assign n22598 = n1726 & n20160 ;
  assign n22599 = n1227 & ~n10317 ;
  assign n22600 = n2887 & ~n8248 ;
  assign n22601 = ~n7347 & n22600 ;
  assign n22602 = n9157 & ~n13433 ;
  assign n22603 = n2687 & n22602 ;
  assign n22604 = n14843 ^ n7263 ^ 1'b0 ;
  assign n22605 = n22604 ^ n12784 ^ 1'b0 ;
  assign n22606 = n19704 & ~n20830 ;
  assign n22607 = n5675 & n22606 ;
  assign n22608 = n2104 & ~n17455 ;
  assign n22609 = n2376 & n22608 ;
  assign n22610 = n6177 & ~n18381 ;
  assign n22611 = n22610 ^ n5890 ^ 1'b0 ;
  assign n22612 = n22609 | n22611 ;
  assign n22613 = n6990 & ~n11608 ;
  assign n22614 = n6604 & n22613 ;
  assign n22615 = n22614 ^ n21177 ^ n15602 ;
  assign n22616 = ~x154 & n19297 ;
  assign n22617 = n9523 & n12575 ;
  assign n22618 = n22617 ^ n1815 ^ 1'b0 ;
  assign n22619 = n15289 ^ n3203 ^ 1'b0 ;
  assign n22620 = n8452 | n16353 ;
  assign n22621 = n22620 ^ n3923 ^ 1'b0 ;
  assign n22622 = n22621 ^ n4222 ^ 1'b0 ;
  assign n22623 = n22619 | n22622 ;
  assign n22624 = n22623 ^ n14017 ^ 1'b0 ;
  assign n22625 = n15622 ^ n9804 ^ 1'b0 ;
  assign n22626 = n2950 & n8717 ;
  assign n22627 = n3137 & n22626 ;
  assign n22628 = n22627 ^ n11049 ^ n9919 ;
  assign n22629 = n6439 ^ n3598 ^ 1'b0 ;
  assign n22630 = n1575 & ~n22629 ;
  assign n22631 = ~x9 & n22630 ;
  assign n22632 = ( n11000 & ~n19575 ) | ( n11000 & n22631 ) | ( ~n19575 & n22631 ) ;
  assign n22633 = n12721 ^ n2623 ^ 1'b0 ;
  assign n22634 = n2128 & n22633 ;
  assign n22635 = n8632 ^ n3736 ^ 1'b0 ;
  assign n22636 = n22634 & n22635 ;
  assign n22637 = n2328 ^ n1956 ^ 1'b0 ;
  assign n22638 = n22636 & n22637 ;
  assign n22639 = n22638 ^ n5607 ^ 1'b0 ;
  assign n22640 = ~x89 & n4229 ;
  assign n22641 = n22640 ^ n17486 ^ 1'b0 ;
  assign n22642 = ~n13657 & n22641 ;
  assign n22643 = n9678 ^ n2338 ^ 1'b0 ;
  assign n22644 = n3421 & n22643 ;
  assign n22645 = ~n13557 & n22644 ;
  assign n22646 = ~n7180 & n22645 ;
  assign n22647 = n22646 ^ n8462 ^ 1'b0 ;
  assign n22648 = n12892 ^ n5350 ^ 1'b0 ;
  assign n22649 = ~n16521 & n22648 ;
  assign n22650 = n547 | n13805 ;
  assign n22651 = n12355 & ~n13256 ;
  assign n22652 = n22651 ^ n15348 ^ 1'b0 ;
  assign n22653 = n5654 ^ n4343 ^ 1'b0 ;
  assign n22654 = ~n17842 & n22653 ;
  assign n22655 = n22654 ^ n20195 ^ 1'b0 ;
  assign n22657 = n1522 & n2878 ;
  assign n22656 = ~n4430 & n6252 ;
  assign n22658 = n22657 ^ n22656 ^ n2219 ;
  assign n22659 = n9562 | n22658 ;
  assign n22660 = n20611 ^ n5357 ^ 1'b0 ;
  assign n22661 = ~n5243 & n9333 ;
  assign n22662 = n5621 | n5895 ;
  assign n22663 = ( n2975 & ~n14215 ) | ( n2975 & n18847 ) | ( ~n14215 & n18847 ) ;
  assign n22664 = ~n1402 & n8816 ;
  assign n22665 = n3066 & n22664 ;
  assign n22666 = n18315 & n22665 ;
  assign n22667 = ~n5225 & n20487 ;
  assign n22668 = n1982 & n6709 ;
  assign n22669 = n22668 ^ n2117 ^ 1'b0 ;
  assign n22670 = n22669 ^ n1937 ^ 1'b0 ;
  assign n22671 = n22667 | n22670 ;
  assign n22672 = n817 & ~n15807 ;
  assign n22673 = n22672 ^ n9691 ^ 1'b0 ;
  assign n22674 = n6425 | n22673 ;
  assign n22675 = n12515 ^ n1225 ^ 1'b0 ;
  assign n22676 = n937 & n13679 ;
  assign n22677 = n22675 & n22676 ;
  assign n22678 = ( x180 & n19754 ) | ( x180 & n22677 ) | ( n19754 & n22677 ) ;
  assign n22679 = n6750 | n8785 ;
  assign n22680 = n13490 | n22679 ;
  assign n22681 = n22680 ^ n19983 ^ 1'b0 ;
  assign n22682 = n1512 & ~n22681 ;
  assign n22685 = n19530 ^ n18640 ^ 1'b0 ;
  assign n22683 = n12366 ^ n9844 ^ 1'b0 ;
  assign n22684 = ( n3954 & n15656 ) | ( n3954 & n22683 ) | ( n15656 & n22683 ) ;
  assign n22686 = n22685 ^ n22684 ^ 1'b0 ;
  assign n22687 = n10744 & ~n14944 ;
  assign n22688 = n7640 & ~n22687 ;
  assign n22689 = ~n6618 & n18382 ;
  assign n22690 = n1338 & ~n2746 ;
  assign n22691 = n18325 ^ n16682 ^ 1'b0 ;
  assign n22692 = ~n10944 & n22691 ;
  assign n22693 = ~n6335 & n15337 ;
  assign n22694 = ~n984 & n22693 ;
  assign n22695 = n22694 ^ n15056 ^ 1'b0 ;
  assign n22696 = n2544 & ~n3750 ;
  assign n22697 = n17537 | n17877 ;
  assign n22699 = ( ~x88 & n2772 ) | ( ~x88 & n5323 ) | ( n2772 & n5323 ) ;
  assign n22698 = ~n21145 & n22587 ;
  assign n22700 = n22699 ^ n22698 ^ 1'b0 ;
  assign n22701 = n2073 & n10808 ;
  assign n22702 = n22701 ^ n4716 ^ 1'b0 ;
  assign n22703 = n22702 ^ n8633 ^ 1'b0 ;
  assign n22704 = n8284 | n11911 ;
  assign n22706 = n6301 ^ n3305 ^ 1'b0 ;
  assign n22707 = n6812 & ~n22706 ;
  assign n22708 = ~n14736 & n22707 ;
  assign n22709 = n22708 ^ n15779 ^ 1'b0 ;
  assign n22710 = n10275 ^ n6733 ^ 1'b0 ;
  assign n22711 = ~n22709 & n22710 ;
  assign n22705 = n4145 | n4218 ;
  assign n22712 = n22711 ^ n22705 ^ 1'b0 ;
  assign n22713 = n977 & ~n20893 ;
  assign n22714 = n15428 ^ n5846 ^ n5622 ;
  assign n22715 = n22714 ^ n8733 ^ n5212 ;
  assign n22716 = n3702 & ~n5359 ;
  assign n22717 = n8945 | n9938 ;
  assign n22718 = n1738 & n11168 ;
  assign n22719 = n22718 ^ n6693 ^ 1'b0 ;
  assign n22720 = n4669 & n11178 ;
  assign n22721 = n22720 ^ n1345 ^ 1'b0 ;
  assign n22722 = n9475 ^ n276 ^ 1'b0 ;
  assign n22723 = ~n2450 & n22722 ;
  assign n22724 = n3223 & n8647 ;
  assign n22725 = ~n1376 & n1983 ;
  assign n22726 = n13144 & n22725 ;
  assign n22727 = n4637 ^ n2264 ^ 1'b0 ;
  assign n22728 = n22726 | n22727 ;
  assign n22729 = ~n5475 & n21050 ;
  assign n22730 = ~n3843 & n22729 ;
  assign n22731 = n1125 ^ n682 ^ 1'b0 ;
  assign n22732 = n510 & ~n22731 ;
  assign n22733 = n22732 ^ n14126 ^ 1'b0 ;
  assign n22734 = x209 & n22700 ;
  assign n22735 = n22734 ^ n597 ^ 1'b0 ;
  assign n22736 = ~n1271 & n9168 ;
  assign n22737 = ~n5576 & n22736 ;
  assign n22738 = ~n4114 & n5686 ;
  assign n22739 = ~n11051 & n22738 ;
  assign n22740 = n6916 & ~n22739 ;
  assign n22741 = n22737 | n22740 ;
  assign n22742 = n3642 | n9733 ;
  assign n22743 = ( n7093 & ~n7890 ) | ( n7093 & n14856 ) | ( ~n7890 & n14856 ) ;
  assign n22744 = n22743 ^ n17107 ^ n15543 ;
  assign n22745 = n12305 | n22744 ;
  assign n22746 = n11834 & ~n22313 ;
  assign n22747 = n16792 & n22746 ;
  assign n22748 = ~n3828 & n8885 ;
  assign n22749 = n22748 ^ n13433 ^ 1'b0 ;
  assign n22750 = ~n2848 & n5114 ;
  assign n22751 = n22750 ^ n6370 ^ 1'b0 ;
  assign n22752 = n22751 ^ n2089 ^ 1'b0 ;
  assign n22753 = n7456 ^ n6536 ^ 1'b0 ;
  assign n22754 = n16988 & ~n22753 ;
  assign n22755 = ~n13363 & n22754 ;
  assign n22756 = n22755 ^ n8730 ^ 1'b0 ;
  assign n22757 = n7421 & ~n16622 ;
  assign n22758 = n6885 & ~n12962 ;
  assign n22759 = n22757 & ~n22758 ;
  assign n22760 = x214 & n22759 ;
  assign n22761 = n22756 & n22760 ;
  assign n22762 = x28 & ~n10246 ;
  assign n22763 = n14421 ^ n6116 ^ 1'b0 ;
  assign n22764 = n14705 & ~n22763 ;
  assign n22765 = n11726 & ~n21250 ;
  assign n22766 = ~n22764 & n22765 ;
  assign n22767 = ~n10410 & n12085 ;
  assign n22768 = ~n5540 & n22767 ;
  assign n22769 = ( n6398 & n6731 ) | ( n6398 & n17056 ) | ( n6731 & n17056 ) ;
  assign n22770 = n22082 | n22769 ;
  assign n22771 = n22770 ^ n13895 ^ 1'b0 ;
  assign n22772 = n8850 ^ n4868 ^ n2140 ;
  assign n22773 = n2995 & ~n9397 ;
  assign n22774 = n22773 ^ n2264 ^ 1'b0 ;
  assign n22775 = ~n378 & n2580 ;
  assign n22776 = n22775 ^ n6160 ^ 1'b0 ;
  assign n22777 = n7121 | n22776 ;
  assign n22778 = n22777 ^ n3258 ^ 1'b0 ;
  assign n22779 = n813 ^ x10 ^ 1'b0 ;
  assign n22780 = n4985 & ~n22779 ;
  assign n22781 = ~x2 & n466 ;
  assign n22782 = ~n4919 & n13074 ;
  assign n22783 = n13949 ^ n10582 ^ 1'b0 ;
  assign n22784 = n6485 | n22783 ;
  assign n22785 = n1859 | n22784 ;
  assign n22786 = n606 & ~n22785 ;
  assign n22787 = ~n4150 & n22786 ;
  assign n22788 = ~n2225 & n22787 ;
  assign n22789 = n11760 & n22788 ;
  assign n22790 = n1651 & n8016 ;
  assign n22791 = n274 & ~n3491 ;
  assign n22792 = n11460 ^ n9173 ^ 1'b0 ;
  assign n22793 = n6090 & ~n8738 ;
  assign n22794 = n22792 | n22793 ;
  assign n22795 = n11114 ^ n4568 ^ 1'b0 ;
  assign n22796 = n17395 & n22795 ;
  assign n22797 = n281 | n5756 ;
  assign n22798 = n22797 ^ n7467 ^ 1'b0 ;
  assign n22799 = n22798 ^ n10475 ^ 1'b0 ;
  assign n22800 = ( n1664 & ~n3970 ) | ( n1664 & n15500 ) | ( ~n3970 & n15500 ) ;
  assign n22801 = n22800 ^ n5265 ^ 1'b0 ;
  assign n22802 = n17201 | n22801 ;
  assign n22803 = n13882 & ~n22802 ;
  assign n22804 = ~n9612 & n15288 ;
  assign n22805 = n22804 ^ n7455 ^ 1'b0 ;
  assign n22806 = ~n15954 & n22805 ;
  assign n22807 = n20387 ^ n20065 ^ 1'b0 ;
  assign n22808 = ~n2263 & n22807 ;
  assign n22809 = n3158 ^ x192 ^ 1'b0 ;
  assign n22810 = ~n12298 & n22809 ;
  assign n22811 = ( n7067 & n19922 ) | ( n7067 & n22810 ) | ( n19922 & n22810 ) ;
  assign n22812 = n20665 ^ n14086 ^ n11660 ;
  assign n22813 = n16145 ^ n2846 ^ 1'b0 ;
  assign n22814 = n19469 | n22813 ;
  assign n22815 = n22812 | n22814 ;
  assign n22821 = n2450 ^ n1014 ^ 1'b0 ;
  assign n22816 = n4914 ^ n723 ^ 1'b0 ;
  assign n22817 = n1170 & n22816 ;
  assign n22818 = n5380 | n7183 ;
  assign n22819 = n7154 | n22818 ;
  assign n22820 = n22817 & n22819 ;
  assign n22822 = n22821 ^ n22820 ^ 1'b0 ;
  assign n22823 = ~n3003 & n5187 ;
  assign n22824 = n20916 & n22823 ;
  assign n22825 = ( ~n677 & n12080 ) | ( ~n677 & n22824 ) | ( n12080 & n22824 ) ;
  assign n22826 = n4842 & n15078 ;
  assign n22827 = n10184 | n22826 ;
  assign n22828 = ~n432 & n16796 ;
  assign n22829 = ~n9193 & n22828 ;
  assign n22831 = n5300 & ~n8268 ;
  assign n22832 = n22831 ^ n19592 ^ 1'b0 ;
  assign n22830 = n1982 & n19695 ;
  assign n22833 = n22832 ^ n22830 ^ 1'b0 ;
  assign n22834 = n22829 & ~n22833 ;
  assign n22835 = n22834 ^ n16256 ^ 1'b0 ;
  assign n22836 = n18953 ^ n9965 ^ 1'b0 ;
  assign n22837 = n11581 ^ n10807 ^ n10559 ;
  assign n22838 = n8545 ^ n2968 ^ 1'b0 ;
  assign n22839 = ~n22837 & n22838 ;
  assign n22840 = n5418 & ~n10407 ;
  assign n22841 = ( n7210 & ~n19213 ) | ( n7210 & n22840 ) | ( ~n19213 & n22840 ) ;
  assign n22842 = n6149 & ~n8546 ;
  assign n22843 = n22842 ^ n9347 ^ 1'b0 ;
  assign n22844 = n16871 ^ n7463 ^ 1'b0 ;
  assign n22845 = ~n19454 & n22844 ;
  assign n22846 = n14052 | n22845 ;
  assign n22847 = n3685 | n17349 ;
  assign n22848 = n5333 ^ n2007 ^ 1'b0 ;
  assign n22849 = n22847 & ~n22848 ;
  assign n22850 = ~n3996 & n17666 ;
  assign n22851 = n3034 | n11576 ;
  assign n22852 = n1059 & ~n22851 ;
  assign n22853 = n10594 & n11994 ;
  assign n22854 = n22853 ^ n17852 ^ 1'b0 ;
  assign n22855 = n11601 & n22854 ;
  assign n22856 = n503 & ~n3645 ;
  assign n22857 = n7319 | n20010 ;
  assign n22858 = ~n22856 & n22857 ;
  assign n22859 = ~n17285 & n22858 ;
  assign n22860 = n530 & ~n16872 ;
  assign n22861 = n619 | n8103 ;
  assign n22862 = n575 & n3915 ;
  assign n22863 = n22862 ^ n1899 ^ 1'b0 ;
  assign n22864 = n22863 ^ n14445 ^ 1'b0 ;
  assign n22865 = n3941 | n11516 ;
  assign n22866 = n8513 & ~n11000 ;
  assign n22867 = ~n801 & n4936 ;
  assign n22868 = n22867 ^ n12075 ^ 1'b0 ;
  assign n22869 = n9306 | n17082 ;
  assign n22870 = n18730 ^ n5835 ^ 1'b0 ;
  assign n22871 = n18145 & n22870 ;
  assign n22872 = n19337 ^ n5004 ^ 1'b0 ;
  assign n22873 = n10854 ^ n7710 ^ 1'b0 ;
  assign n22874 = n3670 | n22873 ;
  assign n22875 = n4520 & ~n22874 ;
  assign n22876 = ~n13238 & n22875 ;
  assign n22877 = n1759 ^ n1730 ^ 1'b0 ;
  assign n22883 = n2617 ^ x190 ^ 1'b0 ;
  assign n22884 = n2594 | n22883 ;
  assign n22878 = n420 | n3039 ;
  assign n22879 = n4830 | n22878 ;
  assign n22880 = n2589 & ~n22879 ;
  assign n22881 = ~n3257 & n22880 ;
  assign n22882 = n14021 & ~n22881 ;
  assign n22885 = n22884 ^ n22882 ^ 1'b0 ;
  assign n22886 = n998 | n6204 ;
  assign n22887 = n22886 ^ n1231 ^ 1'b0 ;
  assign n22888 = n4639 | n22887 ;
  assign n22889 = n1997 & n6609 ;
  assign n22890 = n527 & n22889 ;
  assign n22891 = n22890 ^ n13954 ^ n5371 ;
  assign n22892 = n22888 | n22891 ;
  assign n22893 = n5163 & n9935 ;
  assign n22894 = n22893 ^ n11472 ^ 1'b0 ;
  assign n22895 = n9200 & n10495 ;
  assign n22896 = n17911 ^ n3235 ^ 1'b0 ;
  assign n22897 = n3686 ^ n3670 ^ 1'b0 ;
  assign n22898 = n7701 | n11564 ;
  assign n22899 = n6659 & n11492 ;
  assign n22900 = n1232 & n22899 ;
  assign n22902 = n21516 ^ n3264 ^ 1'b0 ;
  assign n22901 = n2011 | n8072 ;
  assign n22903 = n22902 ^ n22901 ^ n13277 ;
  assign n22904 = ~n14361 & n15264 ;
  assign n22909 = n1138 | n9159 ;
  assign n22905 = n8322 ^ n6119 ^ 1'b0 ;
  assign n22906 = n13540 ^ n13164 ^ 1'b0 ;
  assign n22907 = n22905 | n22906 ;
  assign n22908 = n344 | n22907 ;
  assign n22910 = n22909 ^ n22908 ^ n1170 ;
  assign n22911 = n11116 ^ n6914 ^ 1'b0 ;
  assign n22912 = n22910 & n22911 ;
  assign n22913 = ~n4515 & n14433 ;
  assign n22914 = n19064 & ~n22913 ;
  assign n22915 = n22914 ^ n20408 ^ 1'b0 ;
  assign n22916 = ~n2783 & n12246 ;
  assign n22917 = n21730 & n22916 ;
  assign n22918 = n3688 ^ n3090 ^ 1'b0 ;
  assign n22919 = ~n2192 & n21918 ;
  assign n22921 = n1848 & ~n16508 ;
  assign n22922 = x17 & ~n22921 ;
  assign n22920 = ~x48 & n17359 ;
  assign n22923 = n22922 ^ n22920 ^ 1'b0 ;
  assign n22924 = n10510 & ~n22702 ;
  assign n22925 = ~n20629 & n22924 ;
  assign n22926 = n21366 ^ n8110 ^ n6208 ;
  assign n22927 = n22926 ^ n19751 ^ 1'b0 ;
  assign n22928 = n18952 & ~n22927 ;
  assign n22929 = n18653 ^ n10428 ^ n9958 ;
  assign n22936 = n296 | n10820 ;
  assign n22937 = n22936 ^ n5367 ^ 1'b0 ;
  assign n22934 = n909 | n4029 ;
  assign n22930 = x133 & ~n21072 ;
  assign n22931 = ~n6796 & n22930 ;
  assign n22932 = n372 | n10168 ;
  assign n22933 = n22931 & ~n22932 ;
  assign n22935 = n22934 ^ n22933 ^ 1'b0 ;
  assign n22938 = n22937 ^ n22935 ^ 1'b0 ;
  assign n22939 = ~n22929 & n22938 ;
  assign n22940 = n22939 ^ n3114 ^ 1'b0 ;
  assign n22942 = n3855 | n6895 ;
  assign n22943 = n2387 | n4239 ;
  assign n22944 = n22943 ^ n5896 ^ 1'b0 ;
  assign n22945 = n22944 ^ n11453 ^ 1'b0 ;
  assign n22946 = n6433 & n22945 ;
  assign n22947 = n22942 & n22946 ;
  assign n22941 = n4293 & n9872 ;
  assign n22948 = n22947 ^ n22941 ^ 1'b0 ;
  assign n22949 = ~n7173 & n22948 ;
  assign n22950 = ~n11270 & n18526 ;
  assign n22951 = ~n22949 & n22950 ;
  assign n22952 = n21510 ^ n7401 ^ 1'b0 ;
  assign n22953 = n12854 ^ n351 ^ 1'b0 ;
  assign n22954 = n8592 & ~n13427 ;
  assign n22955 = ~n4152 & n22954 ;
  assign n22956 = n10513 & ~n22955 ;
  assign n22957 = n21718 & n22956 ;
  assign n22958 = ~n13095 & n19417 ;
  assign n22959 = n22958 ^ n13657 ^ 1'b0 ;
  assign n22960 = ~n4046 & n20067 ;
  assign n22961 = n3815 ^ n3251 ^ 1'b0 ;
  assign n22962 = ~n18543 & n20585 ;
  assign n22963 = n22962 ^ n3417 ^ 1'b0 ;
  assign n22964 = n22963 ^ n3845 ^ 1'b0 ;
  assign n22965 = n22964 ^ n16329 ^ 1'b0 ;
  assign n22966 = n22961 & n22965 ;
  assign n22967 = ( ~n21942 & n22960 ) | ( ~n21942 & n22966 ) | ( n22960 & n22966 ) ;
  assign n22968 = n21347 ^ n1439 ^ 1'b0 ;
  assign n22969 = n6834 ^ n1960 ^ 1'b0 ;
  assign n22970 = n11342 & ~n22969 ;
  assign n22971 = n7987 & ~n22970 ;
  assign n22972 = ~n11957 & n22971 ;
  assign n22973 = n3588 & ~n4069 ;
  assign n22974 = n4981 & n22973 ;
  assign n22975 = n19952 & n22974 ;
  assign n22976 = n7638 | n22975 ;
  assign n22977 = n22976 ^ n9074 ^ 1'b0 ;
  assign n22978 = n5678 & n13071 ;
  assign n22979 = n22977 & n22978 ;
  assign n22980 = n13521 & ~n21688 ;
  assign n22981 = n19377 ^ n9412 ^ 1'b0 ;
  assign n22982 = n4109 & ~n21396 ;
  assign n22983 = n13031 & ~n22982 ;
  assign n22984 = n8816 | n9093 ;
  assign n22985 = n22840 ^ n3223 ^ 1'b0 ;
  assign n22986 = n2629 & ~n8594 ;
  assign n22987 = ( n4813 & n22615 ) | ( n4813 & ~n22986 ) | ( n22615 & ~n22986 ) ;
  assign n22988 = n649 & n794 ;
  assign n22989 = ~n21780 & n22988 ;
  assign n22990 = x159 | n2939 ;
  assign n22991 = n6018 & ~n22990 ;
  assign n22992 = x17 | n1762 ;
  assign n22993 = n3642 ^ n3639 ^ 1'b0 ;
  assign n22994 = n577 | n22993 ;
  assign n22995 = n22994 ^ n14561 ^ 1'b0 ;
  assign n22996 = n22995 ^ n15088 ^ n2487 ;
  assign n22997 = n1211 | n7714 ;
  assign n22998 = n22570 & ~n22997 ;
  assign n22999 = n22998 ^ n15097 ^ n815 ;
  assign n23000 = n9632 & ~n19927 ;
  assign n23001 = n23000 ^ n3425 ^ 1'b0 ;
  assign n23002 = n19924 ^ n10152 ^ 1'b0 ;
  assign n23003 = ( ~n14865 & n14974 ) | ( ~n14865 & n18455 ) | ( n14974 & n18455 ) ;
  assign n23004 = n23003 ^ n957 ^ 1'b0 ;
  assign n23005 = n842 | n23004 ;
  assign n23006 = ~n23002 & n23005 ;
  assign n23007 = ~n363 & n23006 ;
  assign n23008 = ~n20684 & n23007 ;
  assign n23009 = ~n6386 & n14955 ;
  assign n23010 = n23009 ^ n14206 ^ 1'b0 ;
  assign n23011 = n23010 ^ n9792 ^ 1'b0 ;
  assign n23012 = ~n7979 & n23011 ;
  assign n23013 = n23012 ^ n10244 ^ 1'b0 ;
  assign n23014 = n3265 & ~n6424 ;
  assign n23015 = n23014 ^ n5709 ^ 1'b0 ;
  assign n23016 = n3458 & n4047 ;
  assign n23017 = n23016 ^ n3693 ^ 1'b0 ;
  assign n23018 = x202 & n23017 ;
  assign n23019 = n890 & n23018 ;
  assign n23020 = x163 | n23019 ;
  assign n23021 = n12515 & ~n15214 ;
  assign n23022 = n9056 & ~n14690 ;
  assign n23023 = n14094 & ~n17161 ;
  assign n23024 = n8371 ^ n4005 ^ 1'b0 ;
  assign n23025 = n23024 ^ n11810 ^ n8431 ;
  assign n23026 = n3001 & ~n23025 ;
  assign n23027 = n23026 ^ x198 ^ 1'b0 ;
  assign n23028 = n12962 | n16627 ;
  assign n23029 = n12632 | n23028 ;
  assign n23030 = n1738 & n4754 ;
  assign n23031 = n9586 & n23030 ;
  assign n23032 = n23031 ^ n22490 ^ n9967 ;
  assign n23033 = ~n3823 & n7677 ;
  assign n23034 = n7882 ^ n6430 ^ 1'b0 ;
  assign n23035 = n8676 & ~n23034 ;
  assign n23036 = n23035 ^ n4733 ^ n2920 ;
  assign n23037 = ~n3177 & n23036 ;
  assign n23038 = n8844 | n14647 ;
  assign n23039 = n17401 ^ n16142 ^ 1'b0 ;
  assign n23040 = ~n10196 & n23039 ;
  assign n23041 = n23038 & n23040 ;
  assign n23042 = n3475 & ~n12447 ;
  assign n23043 = n7432 & n23042 ;
  assign n23044 = n18141 & n23043 ;
  assign n23045 = n5163 ^ n1027 ^ 1'b0 ;
  assign n23046 = n455 | n23045 ;
  assign n23048 = n4705 & ~n5855 ;
  assign n23049 = n23048 ^ n19166 ^ 1'b0 ;
  assign n23050 = n14141 & n23049 ;
  assign n23051 = n23050 ^ n1170 ^ 1'b0 ;
  assign n23047 = ~n8015 & n14739 ;
  assign n23052 = n23051 ^ n23047 ^ 1'b0 ;
  assign n23053 = n1866 & ~n20540 ;
  assign n23054 = n4100 & n23053 ;
  assign n23055 = n3044 & ~n23054 ;
  assign n23056 = ~n9065 & n13047 ;
  assign n23057 = n17705 & ~n22376 ;
  assign n23060 = n10341 ^ n8100 ^ 1'b0 ;
  assign n23061 = n2928 & n23060 ;
  assign n23058 = n8011 & ~n19328 ;
  assign n23059 = n10682 & n23058 ;
  assign n23062 = n23061 ^ n23059 ^ n11702 ;
  assign n23063 = ~n12703 & n16739 ;
  assign n23065 = n7581 & ~n9470 ;
  assign n23064 = x152 & ~n3686 ;
  assign n23066 = n23065 ^ n23064 ^ 1'b0 ;
  assign n23069 = n13063 & n15269 ;
  assign n23067 = n1737 | n17238 ;
  assign n23068 = n7717 & ~n23067 ;
  assign n23070 = n23069 ^ n23068 ^ 1'b0 ;
  assign n23071 = n16106 & n19947 ;
  assign n23072 = ~n6725 & n23071 ;
  assign n23073 = n6907 & ~n8136 ;
  assign n23074 = n7602 & n23073 ;
  assign n23075 = ~n19656 & n23074 ;
  assign n23076 = n13125 & n17378 ;
  assign n23077 = n6202 & ~n14844 ;
  assign n23078 = ( ~n786 & n6725 ) | ( ~n786 & n23077 ) | ( n6725 & n23077 ) ;
  assign n23079 = ~x129 & n23078 ;
  assign n23080 = n23079 ^ n5953 ^ 1'b0 ;
  assign n23081 = n11181 ^ n1199 ^ 1'b0 ;
  assign n23082 = ( ~n11063 & n17932 ) | ( ~n11063 & n23081 ) | ( n17932 & n23081 ) ;
  assign n23083 = n1885 & n3315 ;
  assign n23084 = n14865 | n23083 ;
  assign n23085 = x205 | n23084 ;
  assign n23086 = n2928 & ~n22483 ;
  assign n23087 = ~n23085 & n23086 ;
  assign n23088 = n13894 ^ n5093 ^ 1'b0 ;
  assign n23089 = n5201 | n23088 ;
  assign n23090 = ~n8138 & n12914 ;
  assign n23091 = n15738 ^ n10746 ^ n4432 ;
  assign n23092 = ( n3850 & ~n7110 ) | ( n3850 & n23091 ) | ( ~n7110 & n23091 ) ;
  assign n23093 = n16481 & n17012 ;
  assign n23094 = n16805 & n19178 ;
  assign n23095 = n9100 ^ n5630 ^ 1'b0 ;
  assign n23096 = n16037 ^ n11732 ^ n938 ;
  assign n23097 = ~x130 & n19695 ;
  assign n23098 = ~n20236 & n23097 ;
  assign n23099 = n23098 ^ n1381 ^ 1'b0 ;
  assign n23100 = n22277 & ~n23099 ;
  assign n23102 = n2035 ^ n1237 ^ 1'b0 ;
  assign n23101 = n8388 | n13917 ;
  assign n23103 = n23102 ^ n23101 ^ 1'b0 ;
  assign n23104 = n14699 | n16329 ;
  assign n23105 = n23104 ^ n1749 ^ 1'b0 ;
  assign n23106 = n3820 | n23105 ;
  assign n23107 = n23106 ^ n458 ^ 1'b0 ;
  assign n23108 = n3568 & n5515 ;
  assign n23109 = n5391 & ~n18235 ;
  assign n23110 = n23109 ^ n12548 ^ 1'b0 ;
  assign n23111 = n23108 | n23110 ;
  assign n23112 = n4576 & n8513 ;
  assign n23113 = ( x242 & n23111 ) | ( x242 & n23112 ) | ( n23111 & n23112 ) ;
  assign n23114 = n5356 ^ n2051 ^ 1'b0 ;
  assign n23115 = n10509 & n21954 ;
  assign n23116 = n14166 & ~n16238 ;
  assign n23117 = n7443 & ~n22942 ;
  assign n23118 = ~n10947 & n23117 ;
  assign n23119 = ~n11997 & n17157 ;
  assign n23120 = n10137 & n23119 ;
  assign n23121 = n21471 ^ n12295 ^ n8233 ;
  assign n23122 = n21426 ^ n11454 ^ 1'b0 ;
  assign n23126 = n583 & ~n15948 ;
  assign n23127 = n2633 | n23126 ;
  assign n23128 = n5652 | n23127 ;
  assign n23123 = n10066 & ~n18617 ;
  assign n23124 = n9824 ^ n4218 ^ 1'b0 ;
  assign n23125 = n23123 & ~n23124 ;
  assign n23129 = n23128 ^ n23125 ^ 1'b0 ;
  assign n23130 = n14972 | n16288 ;
  assign n23131 = ( ~n15260 & n22942 ) | ( ~n15260 & n23130 ) | ( n22942 & n23130 ) ;
  assign n23132 = n23131 ^ n9123 ^ 1'b0 ;
  assign n23133 = n6812 & n23132 ;
  assign n23134 = ~n17586 & n23133 ;
  assign n23135 = ~n18796 & n23134 ;
  assign n23136 = n23135 ^ n9887 ^ 1'b0 ;
  assign n23139 = n7856 ^ n6813 ^ 1'b0 ;
  assign n23140 = n6120 & n23139 ;
  assign n23137 = n1080 & n18286 ;
  assign n23138 = n23137 ^ n14982 ^ 1'b0 ;
  assign n23141 = n23140 ^ n23138 ^ n22840 ;
  assign n23142 = ~n19684 & n22556 ;
  assign n23143 = n16935 ^ n16566 ^ 1'b0 ;
  assign n23144 = n5535 ^ n2228 ^ 1'b0 ;
  assign n23145 = n4202 | n23144 ;
  assign n23146 = n983 | n23145 ;
  assign n23147 = n23146 ^ n3790 ^ 1'b0 ;
  assign n23148 = n2679 ^ n509 ^ 1'b0 ;
  assign n23149 = n23148 ^ n6115 ^ 1'b0 ;
  assign n23150 = ~n23147 & n23149 ;
  assign n23151 = x172 | n9104 ;
  assign n23152 = n8307 | n23151 ;
  assign n23153 = n16768 ^ n3266 ^ n725 ;
  assign n23154 = n17764 ^ n2883 ^ 1'b0 ;
  assign n23155 = n4957 | n20904 ;
  assign n23156 = ( n3549 & n8566 ) | ( n3549 & ~n10099 ) | ( n8566 & ~n10099 ) ;
  assign n23157 = n23156 ^ n7051 ^ 1'b0 ;
  assign n23158 = n6483 | n9700 ;
  assign n23159 = n21780 | n23158 ;
  assign n23160 = n19591 ^ n6856 ^ 1'b0 ;
  assign n23161 = ~n691 & n23160 ;
  assign n23162 = n14433 & n23161 ;
  assign n23163 = n2771 & ~n23162 ;
  assign n23164 = n2975 ^ n725 ^ 1'b0 ;
  assign n23165 = n19952 ^ n3850 ^ 1'b0 ;
  assign n23166 = ~n2928 & n13549 ;
  assign n23167 = n8921 & n13538 ;
  assign n23171 = n12736 ^ n4403 ^ 1'b0 ;
  assign n23168 = n3446 ^ n2314 ^ 1'b0 ;
  assign n23169 = n3070 & n23168 ;
  assign n23170 = n22628 & n23169 ;
  assign n23172 = n23171 ^ n23170 ^ 1'b0 ;
  assign n23173 = n17471 ^ n537 ^ 1'b0 ;
  assign n23174 = n11883 | n23173 ;
  assign n23175 = ( n2769 & ~n14034 ) | ( n2769 & n23174 ) | ( ~n14034 & n23174 ) ;
  assign n23176 = n23175 ^ n4453 ^ 1'b0 ;
  assign n23177 = n11097 | n23176 ;
  assign n23178 = n13650 & ~n23177 ;
  assign n23179 = ~n3967 & n4357 ;
  assign n23180 = ~n9215 & n23179 ;
  assign n23181 = n14206 | n23180 ;
  assign n23182 = ~n5437 & n12557 ;
  assign n23183 = n1727 | n21516 ;
  assign n23184 = n12242 | n23183 ;
  assign n23185 = ~n8815 & n23184 ;
  assign n23186 = n23185 ^ n9264 ^ 1'b0 ;
  assign n23187 = n23186 ^ n18408 ^ 1'b0 ;
  assign n23188 = n3648 & n23187 ;
  assign n23189 = n15671 ^ n8163 ^ 1'b0 ;
  assign n23190 = n6510 | n18142 ;
  assign n23191 = n7665 & n22375 ;
  assign n23192 = ~x253 & n23191 ;
  assign n23193 = n21690 ^ n16385 ^ n9623 ;
  assign n23194 = n23193 ^ n15027 ^ 1'b0 ;
  assign n23195 = n2929 ^ n1935 ^ 1'b0 ;
  assign n23196 = n13849 & n23195 ;
  assign n23197 = x254 & ~n23196 ;
  assign n23198 = n13107 ^ n4128 ^ 1'b0 ;
  assign n23199 = ~n9898 & n23198 ;
  assign n23200 = n2901 & n23199 ;
  assign n23201 = n5453 & n10254 ;
  assign n23202 = n23201 ^ n10443 ^ 1'b0 ;
  assign n23203 = n23202 ^ n4459 ^ 1'b0 ;
  assign n23204 = n1592 | n23203 ;
  assign n23205 = n12884 ^ n1220 ^ 1'b0 ;
  assign n23206 = n21705 & n23205 ;
  assign n23209 = n831 & n17449 ;
  assign n23207 = n21110 ^ n11988 ^ 1'b0 ;
  assign n23208 = n11091 & ~n23207 ;
  assign n23210 = n23209 ^ n23208 ^ n5891 ;
  assign n23211 = ~x204 & n13787 ;
  assign n23212 = n23211 ^ n20592 ^ 1'b0 ;
  assign n23213 = n10246 ^ n2271 ^ 1'b0 ;
  assign n23214 = n8452 | n23213 ;
  assign n23215 = n23214 ^ n3158 ^ 1'b0 ;
  assign n23216 = n23215 ^ n17750 ^ 1'b0 ;
  assign n23217 = n9030 ^ n4178 ^ 1'b0 ;
  assign n23220 = n1328 & ~n9933 ;
  assign n23221 = n23220 ^ n8177 ^ 1'b0 ;
  assign n23218 = n3810 & ~n10959 ;
  assign n23219 = n23218 ^ n1571 ^ 1'b0 ;
  assign n23222 = n23221 ^ n23219 ^ 1'b0 ;
  assign n23223 = n11945 & n23222 ;
  assign n23224 = n15410 & ~n16270 ;
  assign n23225 = ~n15537 & n23224 ;
  assign n23226 = n15051 & ~n23225 ;
  assign n23227 = n5800 & n8447 ;
  assign n23228 = ~n14227 & n23227 ;
  assign n23233 = n15080 ^ n3419 ^ 1'b0 ;
  assign n23234 = n11534 & n23233 ;
  assign n23235 = ~n1262 & n23234 ;
  assign n23229 = n16419 ^ n4185 ^ 1'b0 ;
  assign n23230 = n23229 ^ n13521 ^ 1'b0 ;
  assign n23231 = n20987 & n23230 ;
  assign n23232 = ~n14699 & n23231 ;
  assign n23236 = n23235 ^ n23232 ^ 1'b0 ;
  assign n23237 = x155 & n3978 ;
  assign n23238 = n23237 ^ n7977 ^ 1'b0 ;
  assign n23239 = n23238 ^ n17633 ^ 1'b0 ;
  assign n23240 = n17401 ^ n7600 ^ 1'b0 ;
  assign n23241 = n9595 ^ n4215 ^ 1'b0 ;
  assign n23242 = n15912 ^ n1503 ^ 1'b0 ;
  assign n23243 = n18115 | n23242 ;
  assign n23244 = n5132 ^ n421 ^ 1'b0 ;
  assign n23245 = n23244 ^ n9290 ^ 1'b0 ;
  assign n23246 = n7294 | n11717 ;
  assign n23247 = n23246 ^ n8197 ^ 1'b0 ;
  assign n23248 = n23247 ^ n2746 ^ 1'b0 ;
  assign n23249 = n872 | n4721 ;
  assign n23250 = n23249 ^ n7724 ^ 1'b0 ;
  assign n23251 = n3581 & n10606 ;
  assign n23252 = n23251 ^ n1938 ^ 1'b0 ;
  assign n23253 = n1093 & ~n3348 ;
  assign n23254 = ( ~n1591 & n9955 ) | ( ~n1591 & n13131 ) | ( n9955 & n13131 ) ;
  assign n23255 = n913 | n23254 ;
  assign n23256 = n10794 & n18630 ;
  assign n23257 = ~n23255 & n23256 ;
  assign n23258 = n23253 & ~n23257 ;
  assign n23259 = n16940 & n23258 ;
  assign n23260 = n11470 ^ n4779 ^ 1'b0 ;
  assign n23261 = n5189 | n23260 ;
  assign n23262 = n8977 ^ n8025 ^ 1'b0 ;
  assign n23263 = n4830 & n23262 ;
  assign n23264 = n23263 ^ n6437 ^ 1'b0 ;
  assign n23265 = n4703 & ~n14389 ;
  assign n23266 = n7295 ^ n1250 ^ 1'b0 ;
  assign n23267 = n5607 & ~n23266 ;
  assign n23268 = n6532 & ~n21826 ;
  assign n23270 = ~n1336 & n9271 ;
  assign n23269 = n15669 & n16427 ;
  assign n23271 = n23270 ^ n23269 ^ 1'b0 ;
  assign n23272 = n18773 | n23271 ;
  assign n23273 = n5493 & ~n22881 ;
  assign n23274 = n14282 ^ n4836 ^ 1'b0 ;
  assign n23275 = n7516 & ~n23274 ;
  assign n23276 = n6212 | n6436 ;
  assign n23277 = n434 | n23276 ;
  assign n23278 = n5316 ^ n2203 ^ 1'b0 ;
  assign n23279 = n9532 & n23278 ;
  assign n23280 = ( ~n1575 & n7705 ) | ( ~n1575 & n9155 ) | ( n7705 & n9155 ) ;
  assign n23281 = n23280 ^ n3372 ^ n1853 ;
  assign n23282 = n7936 & n10149 ;
  assign n23283 = n10978 & n23282 ;
  assign n23284 = n16431 ^ n12792 ^ 1'b0 ;
  assign n23285 = n23284 ^ n3977 ^ 1'b0 ;
  assign n23286 = n19682 | n23285 ;
  assign n23287 = n23286 ^ n464 ^ 1'b0 ;
  assign n23288 = n18580 ^ n17388 ^ 1'b0 ;
  assign n23289 = ~n17116 & n23288 ;
  assign n23290 = n23289 ^ n6864 ^ n5039 ;
  assign n23292 = ~n5262 & n15598 ;
  assign n23291 = n18763 & ~n20927 ;
  assign n23293 = n23292 ^ n23291 ^ 1'b0 ;
  assign n23294 = n8180 ^ n1344 ^ 1'b0 ;
  assign n23295 = n7813 | n23294 ;
  assign n23296 = n18092 ^ n6235 ^ 1'b0 ;
  assign n23297 = n23295 | n23296 ;
  assign n23298 = n5678 | n23297 ;
  assign n23299 = n23293 | n23298 ;
  assign n23300 = n1125 & ~n9538 ;
  assign n23301 = n267 & n23300 ;
  assign n23302 = n2240 | n19973 ;
  assign n23303 = n1738 & ~n23011 ;
  assign n23304 = n725 ^ x225 ^ 1'b0 ;
  assign n23305 = ~n564 & n23304 ;
  assign n23306 = n2370 | n17972 ;
  assign n23307 = n8454 ^ n6868 ^ 1'b0 ;
  assign n23308 = n9773 ^ n7506 ^ 1'b0 ;
  assign n23309 = n16283 & ~n23308 ;
  assign n23310 = n15230 ^ n7464 ^ 1'b0 ;
  assign n23311 = n3944 & ~n23310 ;
  assign n23312 = n8483 & n9275 ;
  assign n23313 = ( n7094 & n7123 ) | ( n7094 & ~n14663 ) | ( n7123 & ~n14663 ) ;
  assign n23314 = n23313 ^ n21500 ^ 1'b0 ;
  assign n23315 = ~n7716 & n21574 ;
  assign n23316 = n23315 ^ n11569 ^ 1'b0 ;
  assign n23317 = ~n4001 & n5016 ;
  assign n23318 = n23317 ^ n18314 ^ 1'b0 ;
  assign n23319 = n23318 ^ n12963 ^ n6180 ;
  assign n23320 = n6857 & n7109 ;
  assign n23321 = n23320 ^ n3407 ^ 1'b0 ;
  assign n23322 = n23321 ^ n6357 ^ 1'b0 ;
  assign n23323 = n13119 ^ n2733 ^ 1'b0 ;
  assign n23324 = n4718 & ~n23323 ;
  assign n23325 = ~n5589 & n19866 ;
  assign n23326 = ~n1039 & n23325 ;
  assign n23327 = n9210 | n23326 ;
  assign n23328 = n14522 | n23327 ;
  assign n23329 = n9584 & n23328 ;
  assign n23330 = n14423 & n23329 ;
  assign n23331 = n19576 ^ n1867 ^ 1'b0 ;
  assign n23332 = ( n8282 & n11853 ) | ( n8282 & ~n21666 ) | ( n11853 & ~n21666 ) ;
  assign n23334 = n12961 ^ n9836 ^ n8353 ;
  assign n23333 = ( ~n7998 & n11283 ) | ( ~n7998 & n19388 ) | ( n11283 & n19388 ) ;
  assign n23335 = n23334 ^ n23333 ^ 1'b0 ;
  assign n23336 = n1919 & ~n23335 ;
  assign n23337 = n23336 ^ n21004 ^ 1'b0 ;
  assign n23338 = n9946 | n22970 ;
  assign n23339 = n21353 | n21363 ;
  assign n23340 = n6970 & n21546 ;
  assign n23341 = ~n1261 & n18184 ;
  assign n23342 = ~n1073 & n1569 ;
  assign n23344 = n9028 | n20400 ;
  assign n23345 = n23344 ^ n14762 ^ 1'b0 ;
  assign n23346 = n23345 ^ n7957 ^ n6049 ;
  assign n23347 = n10120 & n11804 ;
  assign n23348 = n23346 & n23347 ;
  assign n23343 = n11719 ^ n10414 ^ 1'b0 ;
  assign n23349 = n23348 ^ n23343 ^ 1'b0 ;
  assign n23350 = ~n23342 & n23349 ;
  assign n23351 = n2716 | n13030 ;
  assign n23352 = ~n860 & n23351 ;
  assign n23353 = n23352 ^ n11677 ^ 1'b0 ;
  assign n23354 = n1197 | n7874 ;
  assign n23355 = x46 | n23354 ;
  assign n23356 = n23355 ^ n2827 ^ 1'b0 ;
  assign n23357 = n10151 ^ n9753 ^ 1'b0 ;
  assign n23358 = n23357 ^ n6889 ^ 1'b0 ;
  assign n23359 = n18326 & ~n23358 ;
  assign n23360 = n17805 ^ n12371 ^ 1'b0 ;
  assign n23361 = ~n11747 & n23360 ;
  assign n23362 = n22669 ^ n1804 ^ 1'b0 ;
  assign n23363 = n19218 | n23362 ;
  assign n23364 = n12766 | n23363 ;
  assign n23365 = n19994 ^ n14071 ^ 1'b0 ;
  assign n23366 = ( n17499 & ~n20340 ) | ( n17499 & n20392 ) | ( ~n20340 & n20392 ) ;
  assign n23367 = n14744 & ~n22921 ;
  assign n23368 = n2335 ^ n1413 ^ 1'b0 ;
  assign n23369 = ~n20944 & n23368 ;
  assign n23370 = n23369 ^ n22634 ^ 1'b0 ;
  assign n23371 = x166 & n1563 ;
  assign n23372 = n8583 & n23371 ;
  assign n23373 = n8975 & n11841 ;
  assign n23374 = n23372 & n23373 ;
  assign n23375 = n22677 ^ n2067 ^ 1'b0 ;
  assign n23376 = n18601 & ~n23375 ;
  assign n23377 = n23376 ^ n18598 ^ n6202 ;
  assign n23378 = n10451 | n13682 ;
  assign n23379 = n13726 ^ n9998 ^ 1'b0 ;
  assign n23380 = n10303 & n23379 ;
  assign n23381 = n16066 | n20148 ;
  assign n23382 = n18385 ^ n9192 ^ 1'b0 ;
  assign n23383 = x40 & ~n23382 ;
  assign n23384 = n18340 ^ n16203 ^ 1'b0 ;
  assign n23385 = n927 | n10356 ;
  assign n23386 = n23385 ^ n12828 ^ 1'b0 ;
  assign n23387 = n7736 & n23386 ;
  assign n23388 = n8490 & ~n23387 ;
  assign n23389 = n710 & n6381 ;
  assign n23390 = n318 & n23389 ;
  assign n23391 = n23390 ^ n7825 ^ 1'b0 ;
  assign n23392 = n5208 & n23391 ;
  assign n23393 = ~n19815 & n22599 ;
  assign n23394 = n17077 ^ n8613 ^ 1'b0 ;
  assign n23395 = n16986 | n23394 ;
  assign n23396 = n19435 ^ n3934 ^ n3114 ;
  assign n23397 = n10066 & n23396 ;
  assign n23398 = n1556 & n23397 ;
  assign n23403 = n2481 & n7552 ;
  assign n23399 = n2761 & ~n6908 ;
  assign n23400 = ~n14165 & n23399 ;
  assign n23401 = n15574 & ~n23400 ;
  assign n23402 = n1912 & n23401 ;
  assign n23404 = n23403 ^ n23402 ^ n6257 ;
  assign n23405 = n10846 ^ n5218 ^ n675 ;
  assign n23406 = n13716 | n23405 ;
  assign n23407 = ~n6555 & n23406 ;
  assign n23408 = n23407 ^ n16252 ^ 1'b0 ;
  assign n23409 = n2064 & n16108 ;
  assign n23410 = n23409 ^ n15097 ^ 1'b0 ;
  assign n23411 = n23410 ^ n4562 ^ 1'b0 ;
  assign n23412 = n2054 & n8745 ;
  assign n23413 = n9754 | n23412 ;
  assign n23415 = n11146 & n21613 ;
  assign n23414 = x100 & ~n21999 ;
  assign n23416 = n23415 ^ n23414 ^ 1'b0 ;
  assign n23417 = n4473 | n20474 ;
  assign n23418 = n1556 & ~n23417 ;
  assign n23419 = n21946 ^ n19888 ^ 1'b0 ;
  assign n23420 = n21573 ^ n14259 ^ 1'b0 ;
  assign n23421 = ~n22709 & n23420 ;
  assign n23422 = n3761 ^ n1523 ^ 1'b0 ;
  assign n23423 = ~n333 & n23422 ;
  assign n23424 = ~x222 & n8544 ;
  assign n23425 = ~n7419 & n23424 ;
  assign n23426 = n3565 & n9450 ;
  assign n23427 = n13398 | n13964 ;
  assign n23428 = n5225 | n23427 ;
  assign n23429 = n9456 ^ x185 ^ 1'b0 ;
  assign n23430 = n11830 & n23429 ;
  assign n23431 = n19617 & n23430 ;
  assign n23432 = n20730 & n23431 ;
  assign n23433 = ~n5316 & n5806 ;
  assign n23434 = n23433 ^ n2293 ^ 1'b0 ;
  assign n23435 = n15251 | n23434 ;
  assign n23436 = n13629 ^ n455 ^ 1'b0 ;
  assign n23437 = ~n15689 & n23436 ;
  assign n23438 = ~n21231 & n23437 ;
  assign n23439 = x59 & ~n699 ;
  assign n23440 = n23439 ^ n5703 ^ 1'b0 ;
  assign n23441 = n23440 ^ n21269 ^ n20058 ;
  assign n23442 = n18397 ^ n8673 ^ 1'b0 ;
  assign n23443 = n3858 | n4088 ;
  assign n23444 = n15264 | n23443 ;
  assign n23445 = n1379 & n8127 ;
  assign n23446 = n569 & n7863 ;
  assign n23447 = n23445 & n23446 ;
  assign n23448 = n14010 | n23447 ;
  assign n23449 = n13830 & ~n23448 ;
  assign n23450 = n10529 ^ n6322 ^ 1'b0 ;
  assign n23451 = n23450 ^ n19422 ^ n5219 ;
  assign n23452 = ( ~n3134 & n7246 ) | ( ~n3134 & n11739 ) | ( n7246 & n11739 ) ;
  assign n23454 = n14873 ^ n6235 ^ 1'b0 ;
  assign n23455 = ~n5683 & n23454 ;
  assign n23453 = n5604 | n20039 ;
  assign n23456 = n23455 ^ n23453 ^ 1'b0 ;
  assign n23457 = n6475 ^ n2114 ^ 1'b0 ;
  assign n23458 = n15923 | n23457 ;
  assign n23459 = ~n14109 & n23458 ;
  assign n23460 = ~n3039 & n13668 ;
  assign n23461 = n11976 & n23460 ;
  assign n23462 = n4716 & n5409 ;
  assign n23463 = n11043 & n23462 ;
  assign n23464 = n10809 | n12326 ;
  assign n23465 = n23463 & ~n23464 ;
  assign n23466 = n7241 | n15359 ;
  assign n23467 = n10139 & n19952 ;
  assign n23468 = n7846 & ~n8258 ;
  assign n23469 = n23468 ^ n3695 ^ 1'b0 ;
  assign n23470 = n23469 ^ n6347 ^ 1'b0 ;
  assign n23471 = n16598 & n18902 ;
  assign n23472 = n12922 & ~n23141 ;
  assign n23474 = n6473 ^ n5723 ^ 1'b0 ;
  assign n23475 = ~n3853 & n23474 ;
  assign n23473 = n8449 | n20516 ;
  assign n23476 = n23475 ^ n23473 ^ n12587 ;
  assign n23477 = n19227 ^ n10292 ^ 1'b0 ;
  assign n23480 = n11919 ^ n10264 ^ 1'b0 ;
  assign n23481 = n4532 & ~n23480 ;
  assign n23482 = n23481 ^ n2276 ^ 1'b0 ;
  assign n23483 = n8564 & ~n23482 ;
  assign n23484 = n23483 ^ n7643 ^ 1'b0 ;
  assign n23478 = n8001 ^ x46 ^ 1'b0 ;
  assign n23479 = n2569 & ~n23478 ;
  assign n23485 = n23484 ^ n23479 ^ 1'b0 ;
  assign n23486 = n23485 ^ n10225 ^ 1'b0 ;
  assign n23487 = n14462 & n23486 ;
  assign n23488 = n3601 | n18126 ;
  assign n23489 = n13602 ^ n12971 ^ n8127 ;
  assign n23490 = n23489 ^ n8391 ^ 1'b0 ;
  assign n23491 = n20630 & ~n23490 ;
  assign n23492 = n22504 ^ n874 ^ 1'b0 ;
  assign n23493 = n4308 & n23492 ;
  assign n23494 = ~n6744 & n17650 ;
  assign n23495 = n23494 ^ n20918 ^ 1'b0 ;
  assign n23496 = n4714 | n14649 ;
  assign n23497 = x52 & ~n3745 ;
  assign n23498 = ~n7384 & n23497 ;
  assign n23499 = n17027 ^ n3672 ^ n1788 ;
  assign n23500 = ~n1086 & n23499 ;
  assign n23501 = ~n18613 & n23500 ;
  assign n23502 = n23501 ^ n11671 ^ 1'b0 ;
  assign n23503 = n8997 ^ n6597 ^ 1'b0 ;
  assign n23504 = n2691 & n23503 ;
  assign n23505 = n7123 & ~n11195 ;
  assign n23506 = ~n23504 & n23505 ;
  assign n23507 = n23506 ^ n19546 ^ 1'b0 ;
  assign n23508 = n18859 ^ n2272 ^ 1'b0 ;
  assign n23510 = n2993 ^ n580 ^ 1'b0 ;
  assign n23509 = n3705 | n12846 ;
  assign n23511 = n23510 ^ n23509 ^ 1'b0 ;
  assign n23513 = n22726 ^ n17808 ^ 1'b0 ;
  assign n23512 = n22163 ^ n15169 ^ 1'b0 ;
  assign n23514 = n23513 ^ n23512 ^ 1'b0 ;
  assign n23515 = n23511 & ~n23514 ;
  assign n23516 = ( n5364 & ~n6701 ) | ( n5364 & n14865 ) | ( ~n6701 & n14865 ) ;
  assign n23517 = n2317 & ~n23516 ;
  assign n23518 = n13085 & n23517 ;
  assign n23519 = ~n1606 & n23518 ;
  assign n23520 = n18040 & n18796 ;
  assign n23521 = n22758 ^ n7166 ^ 1'b0 ;
  assign n23525 = ~n8454 & n11663 ;
  assign n23526 = n6655 & n23525 ;
  assign n23522 = n2531 | n3266 ;
  assign n23523 = n23522 ^ n3806 ^ 1'b0 ;
  assign n23524 = ~n20292 & n23523 ;
  assign n23527 = n23526 ^ n23524 ^ 1'b0 ;
  assign n23528 = n1059 | n23527 ;
  assign n23529 = n16023 | n23068 ;
  assign n23530 = ( n2001 & n8331 ) | ( n2001 & ~n21347 ) | ( n8331 & ~n21347 ) ;
  assign n23531 = ~n6282 & n23530 ;
  assign n23532 = n22341 ^ n7020 ^ 1'b0 ;
  assign n23533 = n6352 & ~n12123 ;
  assign n23534 = n23533 ^ n6781 ^ 1'b0 ;
  assign n23535 = n425 & n2755 ;
  assign n23536 = ~n21874 & n23535 ;
  assign n23537 = n12746 ^ n7137 ^ 1'b0 ;
  assign n23538 = n23537 ^ n9416 ^ n4169 ;
  assign n23539 = n21794 ^ n13708 ^ n10352 ;
  assign n23540 = n23538 & n23539 ;
  assign n23541 = n8424 ^ n351 ^ 1'b0 ;
  assign n23542 = n23541 ^ n20956 ^ 1'b0 ;
  assign n23543 = n13370 & n23542 ;
  assign n23544 = ~n3210 & n21107 ;
  assign n23545 = n23544 ^ n19109 ^ 1'b0 ;
  assign n23546 = n2178 | n8028 ;
  assign n23547 = ~n728 & n16244 ;
  assign n23548 = n1995 & n8600 ;
  assign n23549 = ~n2355 & n23548 ;
  assign n23550 = n3491 & ~n4319 ;
  assign n23551 = n2995 & ~n23550 ;
  assign n23552 = ~n4611 & n19515 ;
  assign n23553 = n23552 ^ n23097 ^ 1'b0 ;
  assign n23554 = n22235 ^ n10416 ^ n8766 ;
  assign n23555 = n23554 ^ n16440 ^ 1'b0 ;
  assign n23556 = n12975 | n23555 ;
  assign n23559 = n12955 | n14398 ;
  assign n23560 = n19718 | n23559 ;
  assign n23557 = n2489 & n3235 ;
  assign n23558 = ~n2712 & n23557 ;
  assign n23561 = n23560 ^ n23558 ^ 1'b0 ;
  assign n23564 = n7519 & ~n8026 ;
  assign n23565 = n23564 ^ n682 ^ 1'b0 ;
  assign n23566 = ~n5519 & n23565 ;
  assign n23567 = n11349 & n23566 ;
  assign n23562 = n764 & ~n15647 ;
  assign n23563 = n23562 ^ n23186 ^ 1'b0 ;
  assign n23568 = n23567 ^ n23563 ^ 1'b0 ;
  assign n23569 = n16822 | n23568 ;
  assign n23570 = n11965 ^ n5181 ^ 1'b0 ;
  assign n23571 = n6931 | n23570 ;
  assign n23573 = ~n7786 & n10730 ;
  assign n23574 = ~n9905 & n23573 ;
  assign n23575 = n8493 ^ n3518 ^ 1'b0 ;
  assign n23576 = ( n3542 & ~n23574 ) | ( n3542 & n23575 ) | ( ~n23574 & n23575 ) ;
  assign n23572 = n4239 | n9115 ;
  assign n23577 = n23576 ^ n23572 ^ 1'b0 ;
  assign n23578 = n5553 & n12677 ;
  assign n23579 = n2787 & n23578 ;
  assign n23580 = n23579 ^ n10870 ^ 1'b0 ;
  assign n23581 = n7992 & n23580 ;
  assign n23582 = n1027 & ~n6514 ;
  assign n23583 = n23582 ^ n13574 ^ 1'b0 ;
  assign n23584 = n2011 | n8930 ;
  assign n23585 = n1628 & ~n23584 ;
  assign n23586 = n8838 ^ n8505 ^ 1'b0 ;
  assign n23587 = ~n23585 & n23586 ;
  assign n23588 = n1142 & n2055 ;
  assign n23589 = n4597 ^ n384 ^ 1'b0 ;
  assign n23590 = n4568 & n9705 ;
  assign n23591 = n14542 ^ n10407 ^ 1'b0 ;
  assign n23592 = ~n23590 & n23591 ;
  assign n23593 = n20279 ^ n4407 ^ 1'b0 ;
  assign n23594 = n12622 & ~n23593 ;
  assign n23595 = ~n4699 & n6340 ;
  assign n23596 = n3600 & n23595 ;
  assign n23597 = x107 & ~n23596 ;
  assign n23598 = n23597 ^ n9307 ^ 1'b0 ;
  assign n23599 = ( n2672 & ~n11181 ) | ( n2672 & n13997 ) | ( ~n11181 & n13997 ) ;
  assign n23600 = ~n11321 & n23599 ;
  assign n23601 = n23600 ^ n8336 ^ 1'b0 ;
  assign n23602 = n2576 & n10781 ;
  assign n23603 = ~n425 & n4824 ;
  assign n23604 = ( n19966 & ~n22975 ) | ( n19966 & n23603 ) | ( ~n22975 & n23603 ) ;
  assign n23605 = n21302 ^ n1738 ^ 1'b0 ;
  assign n23607 = n13037 ^ n4205 ^ 1'b0 ;
  assign n23606 = n3975 | n8690 ;
  assign n23608 = n23607 ^ n23606 ^ 1'b0 ;
  assign n23609 = n23608 ^ n5426 ^ 1'b0 ;
  assign n23610 = n2615 & ~n5070 ;
  assign n23611 = n10761 ^ n3413 ^ n1532 ;
  assign n23612 = n21393 & ~n23611 ;
  assign n23613 = n23612 ^ n15141 ^ 1'b0 ;
  assign n23615 = ~n8381 & n15429 ;
  assign n23616 = ~n8781 & n23615 ;
  assign n23614 = n10518 | n17334 ;
  assign n23617 = n23616 ^ n23614 ^ 1'b0 ;
  assign n23618 = n10499 ^ x169 ^ 1'b0 ;
  assign n23619 = ~n270 & n12222 ;
  assign n23620 = n23618 & n23619 ;
  assign n23621 = n23620 ^ n4844 ^ 1'b0 ;
  assign n23622 = n16970 | n21345 ;
  assign n23623 = n23622 ^ n1324 ^ 1'b0 ;
  assign n23624 = n8892 ^ n5010 ^ 1'b0 ;
  assign n23625 = n6148 & n23624 ;
  assign n23626 = ( ~n2439 & n13633 ) | ( ~n2439 & n22113 ) | ( n13633 & n22113 ) ;
  assign n23632 = n10034 ^ n2728 ^ 1'b0 ;
  assign n23627 = n8336 ^ n4327 ^ 1'b0 ;
  assign n23628 = ~n872 & n23627 ;
  assign n23629 = n19641 ^ n6102 ^ 1'b0 ;
  assign n23630 = n23629 ^ n11730 ^ n2988 ;
  assign n23631 = n23628 & n23630 ;
  assign n23633 = n23632 ^ n23631 ^ 1'b0 ;
  assign n23634 = n23626 & ~n23633 ;
  assign n23635 = ~n23625 & n23634 ;
  assign n23638 = n11087 & n12173 ;
  assign n23639 = n23638 ^ n16401 ^ 1'b0 ;
  assign n23636 = n11511 | n13354 ;
  assign n23637 = n2001 | n23636 ;
  assign n23640 = n23639 ^ n23637 ^ 1'b0 ;
  assign n23641 = n5421 ^ n1557 ^ 1'b0 ;
  assign n23642 = n19200 ^ n6574 ^ 1'b0 ;
  assign n23643 = n3019 & n23642 ;
  assign n23644 = n4134 ^ n2934 ^ 1'b0 ;
  assign n23645 = n11511 | n23644 ;
  assign n23646 = n23645 ^ n7663 ^ n2785 ;
  assign n23647 = n23643 & n23646 ;
  assign n23648 = ~x6 & n2110 ;
  assign n23649 = n23648 ^ n18050 ^ 1'b0 ;
  assign n23650 = n483 | n1301 ;
  assign n23651 = n23650 ^ n6900 ^ 1'b0 ;
  assign n23652 = n11992 ^ n6001 ^ 1'b0 ;
  assign n23653 = n14350 ^ n2056 ^ 1'b0 ;
  assign n23654 = n22236 ^ n14756 ^ n2409 ;
  assign n23655 = n23653 & ~n23654 ;
  assign n23656 = ~n369 & n954 ;
  assign n23657 = n23656 ^ n13280 ^ 1'b0 ;
  assign n23658 = n12998 ^ n11517 ^ 1'b0 ;
  assign n23659 = n11274 ^ n432 ^ 1'b0 ;
  assign n23660 = n23659 ^ n3825 ^ 1'b0 ;
  assign n23662 = ~n3945 & n4230 ;
  assign n23661 = n3462 | n8517 ;
  assign n23663 = n23662 ^ n23661 ^ 1'b0 ;
  assign n23664 = ( n9973 & ~n10383 ) | ( n9973 & n14641 ) | ( ~n10383 & n14641 ) ;
  assign n23665 = ( n14902 & ~n15078 ) | ( n14902 & n19940 ) | ( ~n15078 & n19940 ) ;
  assign n23666 = ~n599 & n4646 ;
  assign n23667 = ~n3150 & n23666 ;
  assign n23668 = n3297 ^ x164 ^ 1'b0 ;
  assign n23669 = n3184 | n23668 ;
  assign n23670 = n19937 | n23669 ;
  assign n23671 = n23667 & ~n23670 ;
  assign n23672 = n1523 | n2988 ;
  assign n23673 = n22123 & ~n23672 ;
  assign n23674 = ~n3453 & n7381 ;
  assign n23677 = n4421 & n11191 ;
  assign n23678 = n23677 ^ n7015 ^ 1'b0 ;
  assign n23675 = n1813 & ~n7933 ;
  assign n23676 = ~n11125 & n23675 ;
  assign n23679 = n23678 ^ n23676 ^ 1'b0 ;
  assign n23680 = n4635 & ~n11961 ;
  assign n23681 = n23680 ^ n4597 ^ 1'b0 ;
  assign n23682 = n23219 | n23681 ;
  assign n23683 = n5416 | n23682 ;
  assign n23684 = n1333 & n11786 ;
  assign n23685 = n1519 & n2801 ;
  assign n23686 = n23685 ^ n6413 ^ 1'b0 ;
  assign n23688 = ~n865 & n9400 ;
  assign n23687 = ~n11522 & n17664 ;
  assign n23689 = n23688 ^ n23687 ^ 1'b0 ;
  assign n23690 = n23686 & n23689 ;
  assign n23692 = n22053 ^ n15970 ^ 1'b0 ;
  assign n23693 = n10698 & n23692 ;
  assign n23691 = x248 & ~n15370 ;
  assign n23694 = n23693 ^ n23691 ^ 1'b0 ;
  assign n23695 = ~x76 & n12146 ;
  assign n23696 = ~n567 & n16334 ;
  assign n23697 = n23696 ^ n8943 ^ 1'b0 ;
  assign n23698 = n539 & ~n23697 ;
  assign n23700 = n20996 ^ n12162 ^ 1'b0 ;
  assign n23699 = n19319 | n23590 ;
  assign n23701 = n23700 ^ n23699 ^ 1'b0 ;
  assign n23702 = n16254 & ~n23701 ;
  assign n23703 = ( n3209 & n4934 ) | ( n3209 & n9072 ) | ( n4934 & n9072 ) ;
  assign n23704 = n23703 ^ n404 ^ 1'b0 ;
  assign n23705 = n1442 & ~n23704 ;
  assign n23706 = n23705 ^ n17981 ^ 1'b0 ;
  assign n23707 = n6551 & n7703 ;
  assign n23708 = ~n18237 & n23707 ;
  assign n23709 = n23708 ^ n20140 ^ 1'b0 ;
  assign n23710 = n18131 | n20542 ;
  assign n23711 = n2085 & ~n23710 ;
  assign n23712 = n298 ^ x47 ^ 1'b0 ;
  assign n23713 = n23711 | n23712 ;
  assign n23714 = n11069 ^ n8415 ^ 1'b0 ;
  assign n23715 = n4428 & n23714 ;
  assign n23716 = n6951 | n11231 ;
  assign n23717 = ~n7040 & n10730 ;
  assign n23718 = n23717 ^ n11662 ^ 1'b0 ;
  assign n23719 = ~n4868 & n10655 ;
  assign n23720 = n10532 & n23719 ;
  assign n23721 = n23720 ^ n9876 ^ 1'b0 ;
  assign n23722 = n23718 | n23721 ;
  assign n23723 = n4433 | n21188 ;
  assign n23724 = n15486 & ~n23723 ;
  assign n23725 = n23724 ^ n4082 ^ 1'b0 ;
  assign n23728 = n10145 ^ n8454 ^ 1'b0 ;
  assign n23726 = n4701 ^ n611 ^ 1'b0 ;
  assign n23727 = n281 | n23726 ;
  assign n23729 = n23728 ^ n23727 ^ 1'b0 ;
  assign n23730 = n13940 ^ n8438 ^ 1'b0 ;
  assign n23731 = n5735 & n23730 ;
  assign n23732 = n3985 | n17801 ;
  assign n23734 = n7629 ^ n7370 ^ 1'b0 ;
  assign n23735 = n8957 | n23734 ;
  assign n23736 = n16481 & ~n23735 ;
  assign n23737 = n23736 ^ n2689 ^ 1'b0 ;
  assign n23733 = n2819 & ~n10827 ;
  assign n23738 = n23737 ^ n23733 ^ n17267 ;
  assign n23739 = n23738 ^ n258 ^ 1'b0 ;
  assign n23740 = ~n3319 & n22821 ;
  assign n23741 = ~n18953 & n23740 ;
  assign n23742 = n21609 ^ n9531 ^ 1'b0 ;
  assign n23743 = ( n3850 & n9347 ) | ( n3850 & n12522 ) | ( n9347 & n12522 ) ;
  assign n23744 = n4520 & n5282 ;
  assign n23745 = n23744 ^ n5802 ^ 1'b0 ;
  assign n23746 = n14380 | n15761 ;
  assign n23747 = n14992 & n16885 ;
  assign n23748 = n12133 ^ n8414 ^ 1'b0 ;
  assign n23749 = x116 & n14840 ;
  assign n23750 = n11877 ^ n9461 ^ 1'b0 ;
  assign n23751 = ( n3536 & n5667 ) | ( n3536 & n7455 ) | ( n5667 & n7455 ) ;
  assign n23752 = n23751 ^ n11685 ^ 1'b0 ;
  assign n23753 = n16708 ^ n14905 ^ n12655 ;
  assign n23754 = n3098 & ~n3155 ;
  assign n23755 = ~n4460 & n23754 ;
  assign n23756 = n997 | n20033 ;
  assign n23757 = n10297 | n23756 ;
  assign n23758 = ~n22925 & n23757 ;
  assign n23759 = n23758 ^ n7199 ^ 1'b0 ;
  assign n23760 = n4684 & ~n22557 ;
  assign n23761 = ~n6759 & n23760 ;
  assign n23762 = n23761 ^ n731 ^ 1'b0 ;
  assign n23763 = n13918 & n23762 ;
  assign n23764 = n23763 ^ n10907 ^ 1'b0 ;
  assign n23765 = n23737 | n23764 ;
  assign n23766 = ~n3009 & n16128 ;
  assign n23767 = n23765 & n23766 ;
  assign n23768 = ( n2710 & n13236 ) | ( n2710 & ~n23767 ) | ( n13236 & ~n23767 ) ;
  assign n23771 = n7276 | n17707 ;
  assign n23769 = n6359 & n16308 ;
  assign n23770 = n23769 ^ n6627 ^ 1'b0 ;
  assign n23772 = n23771 ^ n23770 ^ 1'b0 ;
  assign n23773 = n15276 & n22604 ;
  assign n23774 = n4931 & ~n9989 ;
  assign n23775 = n9138 & n23774 ;
  assign n23776 = n2531 | n10043 ;
  assign n23777 = n23776 ^ n17033 ^ 1'b0 ;
  assign n23779 = ~n3140 & n5122 ;
  assign n23778 = n1416 | n17825 ;
  assign n23780 = n23779 ^ n23778 ^ 1'b0 ;
  assign n23781 = n12262 | n23780 ;
  assign n23782 = n23781 ^ n920 ^ 1'b0 ;
  assign n23783 = n23782 ^ n13603 ^ 1'b0 ;
  assign n23784 = n9767 & n23783 ;
  assign n23785 = n16524 ^ n9889 ^ 1'b0 ;
  assign n23786 = n9293 | n23785 ;
  assign n23787 = n8873 | n23786 ;
  assign n23792 = ~n1086 & n18985 ;
  assign n23788 = n949 & ~n5054 ;
  assign n23789 = ~n949 & n23788 ;
  assign n23790 = n23789 ^ n16314 ^ 1'b0 ;
  assign n23791 = n754 | n23790 ;
  assign n23793 = n23792 ^ n23791 ^ 1'b0 ;
  assign n23794 = n9903 ^ n4083 ^ 1'b0 ;
  assign n23795 = n4294 ^ n1398 ^ 1'b0 ;
  assign n23796 = n1599 & n23795 ;
  assign n23797 = ~n10485 & n13451 ;
  assign n23798 = n23797 ^ n13607 ^ 1'b0 ;
  assign n23799 = ~n11643 & n14375 ;
  assign n23800 = n16204 & n23799 ;
  assign n23801 = n1245 & ~n2325 ;
  assign n23802 = n3081 & n23801 ;
  assign n23803 = ~n1749 & n23802 ;
  assign n23805 = n1125 & n16967 ;
  assign n23806 = n11230 & n23805 ;
  assign n23804 = n16829 ^ n5705 ^ 1'b0 ;
  assign n23807 = n23806 ^ n23804 ^ 1'b0 ;
  assign n23808 = ~n13494 & n13539 ;
  assign n23809 = n13198 & ~n16463 ;
  assign n23810 = n13858 & n23809 ;
  assign n23811 = n17607 ^ n5339 ^ 1'b0 ;
  assign n23812 = n767 & ~n23811 ;
  assign n23813 = n18852 & n23812 ;
  assign n23814 = n3806 | n5333 ;
  assign n23815 = n3124 & ~n23814 ;
  assign n23816 = ( ~n5084 & n16267 ) | ( ~n5084 & n23815 ) | ( n16267 & n23815 ) ;
  assign n23822 = ~n3367 & n4340 ;
  assign n23823 = ~n4340 & n23822 ;
  assign n23824 = n3864 & ~n23823 ;
  assign n23825 = n23823 & n23824 ;
  assign n23826 = n17872 | n23825 ;
  assign n23817 = n4011 ^ n874 ^ 1'b0 ;
  assign n23818 = n556 & n23817 ;
  assign n23819 = n9342 & n11369 ;
  assign n23820 = ~n23818 & n23819 ;
  assign n23821 = n19538 | n23820 ;
  assign n23827 = n23826 ^ n23821 ^ 1'b0 ;
  assign n23828 = n14324 ^ n9679 ^ 1'b0 ;
  assign n23829 = n15094 ^ n1599 ^ 1'b0 ;
  assign n23830 = ( ~n2856 & n3081 ) | ( ~n2856 & n23829 ) | ( n3081 & n23829 ) ;
  assign n23831 = n1799 & ~n23830 ;
  assign n23832 = n23831 ^ n4277 ^ 1'b0 ;
  assign n23833 = n7796 ^ n2646 ^ 1'b0 ;
  assign n23834 = n23833 ^ x230 ^ 1'b0 ;
  assign n23835 = n3355 & n23834 ;
  assign n23836 = n6649 & n17264 ;
  assign n23837 = n23836 ^ n1509 ^ 1'b0 ;
  assign n23838 = n16463 ^ n14065 ^ 1'b0 ;
  assign n23839 = n3588 & n23838 ;
  assign n23840 = n4739 ^ n2086 ^ x74 ;
  assign n23841 = ~n4925 & n23840 ;
  assign n23842 = n1086 & n23841 ;
  assign n23843 = n1121 & ~n7000 ;
  assign n23844 = n23843 ^ x206 ^ 1'b0 ;
  assign n23845 = n3073 & ~n5705 ;
  assign n23846 = ~n3607 & n23845 ;
  assign n23847 = n23846 ^ n14846 ^ 1'b0 ;
  assign n23848 = ~n23844 & n23847 ;
  assign n23849 = n671 & ~n19800 ;
  assign n23850 = ( n10628 & n19306 ) | ( n10628 & n21577 ) | ( n19306 & n21577 ) ;
  assign n23851 = ~n2598 & n15282 ;
  assign n23852 = n23851 ^ n651 ^ 1'b0 ;
  assign n23853 = n10756 ^ n2743 ^ 1'b0 ;
  assign n23854 = n23852 & ~n23853 ;
  assign n23855 = n545 & ~n2013 ;
  assign n23856 = n23855 ^ n7119 ^ 1'b0 ;
  assign n23857 = n22445 & n23856 ;
  assign n23858 = n21615 & n23857 ;
  assign n23859 = n3498 | n3725 ;
  assign n23860 = n23859 ^ n9676 ^ 1'b0 ;
  assign n23861 = ~n3984 & n23860 ;
  assign n23862 = n23861 ^ n11952 ^ 1'b0 ;
  assign n23863 = n6707 ^ n4788 ^ 1'b0 ;
  assign n23869 = n3956 | n4022 ;
  assign n23864 = n14569 ^ n8904 ^ 1'b0 ;
  assign n23865 = n4656 | n10084 ;
  assign n23866 = n23081 | n23865 ;
  assign n23867 = n23069 & ~n23866 ;
  assign n23868 = ~n23864 & n23867 ;
  assign n23870 = n23869 ^ n23868 ^ 1'b0 ;
  assign n23871 = n23863 | n23870 ;
  assign n23877 = ~n624 & n756 ;
  assign n23878 = n624 & n23877 ;
  assign n23872 = n11954 ^ n11348 ^ n8974 ;
  assign n23873 = n1633 | n23872 ;
  assign n23874 = n23872 & ~n23873 ;
  assign n23875 = n5812 & ~n8806 ;
  assign n23876 = ~n23874 & n23875 ;
  assign n23879 = n23878 ^ n23876 ^ 1'b0 ;
  assign n23880 = ~n13074 & n19952 ;
  assign n23881 = ~n6219 & n10742 ;
  assign n23883 = ~n2390 & n2624 ;
  assign n23884 = ~n13689 & n23883 ;
  assign n23885 = n4489 & n23884 ;
  assign n23882 = ~n8649 & n19064 ;
  assign n23886 = n23885 ^ n23882 ^ 1'b0 ;
  assign n23887 = n4436 | n5443 ;
  assign n23888 = n23887 ^ n14510 ^ 1'b0 ;
  assign n23889 = n13737 & n16372 ;
  assign n23890 = n872 | n6421 ;
  assign n23891 = n420 & n23662 ;
  assign n23892 = n1091 & n23891 ;
  assign n23893 = n23892 ^ n23701 ^ 1'b0 ;
  assign n23894 = n21361 ^ n17639 ^ 1'b0 ;
  assign n23895 = n9714 & ~n23894 ;
  assign n23896 = n13629 & ~n19200 ;
  assign n23901 = n359 & ~n1034 ;
  assign n23902 = n23901 ^ n9385 ^ 1'b0 ;
  assign n23903 = n8113 & n21225 ;
  assign n23904 = ~n23902 & n23903 ;
  assign n23897 = n1309 | n6826 ;
  assign n23898 = n23897 ^ n4394 ^ 1'b0 ;
  assign n23899 = n1388 & n20630 ;
  assign n23900 = ~n23898 & n23899 ;
  assign n23905 = n23904 ^ n23900 ^ n946 ;
  assign n23906 = n4393 | n7084 ;
  assign n23907 = n11841 | n23906 ;
  assign n23908 = n23907 ^ n18087 ^ 1'b0 ;
  assign n23909 = n17315 & n23908 ;
  assign n23910 = n7597 ^ n4144 ^ 1'b0 ;
  assign n23911 = n23910 ^ n10429 ^ 1'b0 ;
  assign n23925 = n1682 & ~n5235 ;
  assign n23926 = ~n1682 & n23925 ;
  assign n23927 = n716 | n23926 ;
  assign n23928 = n13210 & ~n23927 ;
  assign n23929 = n1671 & ~n5316 ;
  assign n23930 = ~n1671 & n23929 ;
  assign n23931 = n23930 ^ n8950 ^ 1'b0 ;
  assign n23932 = n23928 | n23931 ;
  assign n23923 = n10325 | n18786 ;
  assign n23924 = n23923 ^ n9017 ^ 1'b0 ;
  assign n23912 = ~n3494 & n4417 ;
  assign n23913 = ~n4417 & n23912 ;
  assign n23914 = n2693 | n23913 ;
  assign n23915 = n2693 & ~n23914 ;
  assign n23916 = n11714 | n15616 ;
  assign n23917 = n23915 & ~n23916 ;
  assign n23918 = x100 & ~n3359 ;
  assign n23919 = ~x100 & n23918 ;
  assign n23920 = n23919 ^ n2055 ^ 1'b0 ;
  assign n23921 = ~n6510 & n23920 ;
  assign n23922 = n23917 & n23921 ;
  assign n23933 = n23932 ^ n23924 ^ n23922 ;
  assign n23934 = n7449 & ~n11628 ;
  assign n23935 = n8829 | n18781 ;
  assign n23936 = n15177 | n23935 ;
  assign n23937 = ~n2783 & n20351 ;
  assign n23938 = n14235 ^ n875 ^ 1'b0 ;
  assign n23939 = n18459 ^ n7643 ^ n671 ;
  assign n23940 = n5296 & ~n13622 ;
  assign n23941 = n11196 ^ n8252 ^ 1'b0 ;
  assign n23942 = n7141 & n23941 ;
  assign n23943 = ~n4747 & n6633 ;
  assign n23944 = ~n9693 & n23943 ;
  assign n23945 = n23944 ^ n14777 ^ 1'b0 ;
  assign n23946 = n6171 & n23945 ;
  assign n23947 = n11186 ^ n983 ^ 1'b0 ;
  assign n23948 = n6921 | n7573 ;
  assign n23949 = n23948 ^ n11965 ^ 1'b0 ;
  assign n23956 = n16871 ^ n4424 ^ 1'b0 ;
  assign n23957 = n3592 | n23956 ;
  assign n23950 = n5438 & n19957 ;
  assign n23951 = n23950 ^ n15564 ^ 1'b0 ;
  assign n23952 = ~n1809 & n2048 ;
  assign n23953 = n12956 & n23952 ;
  assign n23954 = n23951 & ~n23953 ;
  assign n23955 = ~n14890 & n23954 ;
  assign n23958 = n23957 ^ n23955 ^ 1'b0 ;
  assign n23959 = n16903 & n23958 ;
  assign n23960 = ~n4949 & n12597 ;
  assign n23961 = n13110 & n23960 ;
  assign n23962 = n3946 | n18733 ;
  assign n23963 = ( n879 & n1859 ) | ( n879 & ~n7128 ) | ( n1859 & ~n7128 ) ;
  assign n23964 = n23963 ^ n3184 ^ 1'b0 ;
  assign n23965 = ( n3298 & ~n11446 ) | ( n3298 & n23964 ) | ( ~n11446 & n23964 ) ;
  assign n23966 = n20927 ^ n10172 ^ 1'b0 ;
  assign n23967 = n344 & n23966 ;
  assign n23968 = n22737 & n23967 ;
  assign n23969 = n1034 | n10435 ;
  assign n23970 = n23969 ^ n12569 ^ 1'b0 ;
  assign n23971 = n21296 ^ n4321 ^ 1'b0 ;
  assign n23972 = n4519 & n23971 ;
  assign n23973 = n14222 & ~n17693 ;
  assign n23974 = n23973 ^ n5933 ^ 1'b0 ;
  assign n23975 = x8 & ~n16943 ;
  assign n23976 = ~n4519 & n23975 ;
  assign n23977 = n23976 ^ n7045 ^ 1'b0 ;
  assign n23978 = n4496 ^ n3594 ^ 1'b0 ;
  assign n23979 = ~n7298 & n20648 ;
  assign n23980 = ( x254 & ~n6701 ) | ( x254 & n20637 ) | ( ~n6701 & n20637 ) ;
  assign n23981 = ~n2050 & n19866 ;
  assign n23982 = n23981 ^ n6819 ^ n3419 ;
  assign n23983 = n3432 ^ n2434 ^ x26 ;
  assign n23984 = n5831 & ~n8097 ;
  assign n23985 = ~n23983 & n23984 ;
  assign n23986 = n13842 ^ x18 ^ 1'b0 ;
  assign n23987 = n7201 | n23986 ;
  assign n23988 = n8850 | n10095 ;
  assign n23989 = n23988 ^ n17984 ^ 1'b0 ;
  assign n23990 = n6131 & n7069 ;
  assign n23991 = ~n7069 & n23990 ;
  assign n23992 = n23991 ^ n17491 ^ 1'b0 ;
  assign n23993 = n2214 & n10218 ;
  assign n23994 = n23993 ^ n3724 ^ 1'b0 ;
  assign n23995 = n23994 ^ n17728 ^ n9054 ;
  assign n23996 = n4405 | n13079 ;
  assign n23997 = ~n2070 & n23996 ;
  assign n23998 = n615 | n13442 ;
  assign n23999 = n23998 ^ n10547 ^ 1'b0 ;
  assign n24000 = n3142 ^ n1789 ^ 1'b0 ;
  assign n24001 = n2331 & n24000 ;
  assign n24002 = n23999 & n24001 ;
  assign n24003 = n6531 & ~n19564 ;
  assign n24004 = n24003 ^ n3978 ^ 1'b0 ;
  assign n24005 = n4150 ^ x50 ^ 1'b0 ;
  assign n24006 = n21956 ^ n19162 ^ 1'b0 ;
  assign n24007 = n4668 | n24006 ;
  assign n24008 = n14757 & n16329 ;
  assign n24009 = n24008 ^ n4750 ^ 1'b0 ;
  assign n24011 = n5033 ^ n4793 ^ 1'b0 ;
  assign n24012 = n12839 ^ n8422 ^ 1'b0 ;
  assign n24013 = n24011 | n24012 ;
  assign n24014 = n24013 ^ x241 ^ 1'b0 ;
  assign n24010 = x235 & ~n19430 ;
  assign n24015 = n24014 ^ n24010 ^ 1'b0 ;
  assign n24016 = n3709 | n6653 ;
  assign n24017 = n3709 & ~n24016 ;
  assign n24018 = n14267 ^ n9993 ^ n2098 ;
  assign n24019 = n1342 | n7627 ;
  assign n24020 = n7627 & ~n24019 ;
  assign n24021 = n23219 | n24020 ;
  assign n24022 = n24021 ^ n5573 ^ 1'b0 ;
  assign n24023 = ~n3740 & n23839 ;
  assign n24024 = n13600 & n24023 ;
  assign n24025 = n20876 ^ n11105 ^ 1'b0 ;
  assign n24026 = n710 & n18800 ;
  assign n24027 = n18357 ^ n5987 ^ 1'b0 ;
  assign n24028 = n15125 ^ n3805 ^ 1'b0 ;
  assign n24029 = n8030 & ~n12133 ;
  assign n24030 = n23538 ^ n15275 ^ 1'b0 ;
  assign n24031 = n24029 & ~n24030 ;
  assign n24032 = n12802 & n24031 ;
  assign n24033 = n8005 ^ n4899 ^ 1'b0 ;
  assign n24034 = n24032 | n24033 ;
  assign n24035 = n15937 & n16388 ;
  assign n24036 = n11660 & n24035 ;
  assign n24037 = n5704 & n20688 ;
  assign n24038 = ~n6387 & n24037 ;
  assign n24039 = ( n9199 & ~n16069 ) | ( n9199 & n24038 ) | ( ~n16069 & n24038 ) ;
  assign n24040 = n9856 ^ n1846 ^ 1'b0 ;
  assign n24043 = n9739 ^ n520 ^ x92 ;
  assign n24041 = ~n3590 & n17311 ;
  assign n24042 = n6273 & n24041 ;
  assign n24044 = n24043 ^ n24042 ^ 1'b0 ;
  assign n24045 = n6278 | n24044 ;
  assign n24046 = n24045 ^ n5175 ^ 1'b0 ;
  assign n24047 = n10657 & n24046 ;
  assign n24048 = ~n3150 & n3419 ;
  assign n24049 = n18828 ^ x154 ^ 1'b0 ;
  assign n24050 = n2540 & n24049 ;
  assign n24051 = ( ~n3150 & n10578 ) | ( ~n3150 & n20308 ) | ( n10578 & n20308 ) ;
  assign n24052 = n5680 ^ x230 ^ 1'b0 ;
  assign n24053 = n5994 & ~n24052 ;
  assign n24054 = n19765 & n24053 ;
  assign n24055 = n23765 & n24054 ;
  assign n24056 = n7243 ^ n6921 ^ 1'b0 ;
  assign n24057 = n19385 & n24056 ;
  assign n24058 = ~n20067 & n24057 ;
  assign n24059 = n10702 ^ n10495 ^ 1'b0 ;
  assign n24060 = ~n3042 & n12714 ;
  assign n24061 = n10837 & n24060 ;
  assign n24062 = n24061 ^ n688 ^ 1'b0 ;
  assign n24063 = n4999 ^ n1129 ^ n348 ;
  assign n24064 = n1759 & ~n2098 ;
  assign n24065 = ~n21665 & n24064 ;
  assign n24066 = x81 & ~n11151 ;
  assign n24067 = n24066 ^ n9496 ^ 1'b0 ;
  assign n24068 = n4579 ^ n3094 ^ n3070 ;
  assign n24069 = n24068 ^ n19038 ^ n8616 ;
  assign n24070 = n15392 ^ n1148 ^ 1'b0 ;
  assign n24071 = n24070 ^ n18177 ^ 1'b0 ;
  assign n24072 = ~n16521 & n24071 ;
  assign n24073 = n5474 ^ n3139 ^ 1'b0 ;
  assign n24074 = n24073 ^ n14752 ^ 1'b0 ;
  assign n24075 = n3721 | n14002 ;
  assign n24076 = n24075 ^ n17075 ^ 1'b0 ;
  assign n24077 = n3383 & n4622 ;
  assign n24078 = ~n10180 & n24077 ;
  assign n24079 = n1125 & ~n24078 ;
  assign n24080 = n8679 ^ n3121 ^ n2924 ;
  assign n24081 = n9754 | n24080 ;
  assign n24082 = n24079 & ~n24081 ;
  assign n24083 = n1391 & ~n6748 ;
  assign n24085 = ~n3477 & n5432 ;
  assign n24084 = n8139 & n10691 ;
  assign n24086 = n24085 ^ n24084 ^ 1'b0 ;
  assign n24087 = n11566 ^ n5003 ^ 1'b0 ;
  assign n24088 = n13251 | n17887 ;
  assign n24089 = n6309 & ~n24088 ;
  assign n24091 = n9608 | n17981 ;
  assign n24092 = n466 | n24091 ;
  assign n24090 = x73 & n13657 ;
  assign n24093 = n24092 ^ n24090 ^ 1'b0 ;
  assign n24094 = ( n3234 & n12865 ) | ( n3234 & n17649 ) | ( n12865 & n17649 ) ;
  assign n24095 = n8001 ^ n7109 ^ 1'b0 ;
  assign n24100 = n15275 ^ n2055 ^ 1'b0 ;
  assign n24096 = ~n4380 & n4447 ;
  assign n24097 = n7791 & ~n24096 ;
  assign n24098 = n24097 ^ n8865 ^ 1'b0 ;
  assign n24099 = n9433 & ~n24098 ;
  assign n24101 = n24100 ^ n24099 ^ 1'b0 ;
  assign n24102 = n12673 & ~n21169 ;
  assign n24103 = n20554 ^ n20519 ^ n6135 ;
  assign n24104 = n260 | n9605 ;
  assign n24105 = n24104 ^ n8702 ^ 1'b0 ;
  assign n24106 = ~n3814 & n14253 ;
  assign n24107 = ~n1123 & n24106 ;
  assign n24114 = n333 | n522 ;
  assign n24115 = n333 & ~n24114 ;
  assign n24116 = n676 & ~n813 ;
  assign n24117 = n24115 & n24116 ;
  assign n24118 = n12765 | n24117 ;
  assign n24119 = n24117 & ~n24118 ;
  assign n24120 = n11868 | n24119 ;
  assign n24108 = ~n1805 & n3395 ;
  assign n24109 = ~n3395 & n24108 ;
  assign n24110 = n2211 | n3156 ;
  assign n24111 = n24109 & ~n24110 ;
  assign n24112 = n2189 & n24111 ;
  assign n24113 = ~n13191 & n24112 ;
  assign n24121 = n24120 ^ n24113 ^ 1'b0 ;
  assign n24122 = n1219 | n4510 ;
  assign n24123 = n2326 | n20834 ;
  assign n24124 = n24122 & ~n24123 ;
  assign n24125 = n14014 ^ n4688 ^ 1'b0 ;
  assign n24126 = n7731 ^ n567 ^ 1'b0 ;
  assign n24127 = ~n2783 & n8496 ;
  assign n24128 = n24127 ^ n7298 ^ 1'b0 ;
  assign n24129 = n24128 ^ n10431 ^ 1'b0 ;
  assign n24130 = n1025 & ~n3850 ;
  assign n24132 = n3555 ^ n359 ^ 1'b0 ;
  assign n24131 = n2102 ^ n1112 ^ 1'b0 ;
  assign n24133 = n24132 ^ n24131 ^ 1'b0 ;
  assign n24134 = n4268 | n14468 ;
  assign n24135 = n9576 & ~n24134 ;
  assign n24137 = ~n471 & n6093 ;
  assign n24136 = ~n1591 & n7478 ;
  assign n24138 = n24137 ^ n24136 ^ 1'b0 ;
  assign n24140 = n7179 ^ n671 ^ 1'b0 ;
  assign n24141 = n1129 & n24140 ;
  assign n24139 = n11147 ^ n3034 ^ 1'b0 ;
  assign n24142 = n24141 ^ n24139 ^ 1'b0 ;
  assign n24143 = n15153 & n16490 ;
  assign n24144 = ( n3761 & n5849 ) | ( n3761 & ~n11942 ) | ( n5849 & ~n11942 ) ;
  assign n24145 = n2725 & ~n24144 ;
  assign n24146 = ~n1195 & n7686 ;
  assign n24147 = ~n1306 & n13727 ;
  assign n24148 = ~n24146 & n24147 ;
  assign n24149 = n6490 & ~n10733 ;
  assign n24150 = ~n5582 & n24149 ;
  assign n24151 = n844 & ~n3457 ;
  assign n24152 = n4511 & n24151 ;
  assign n24157 = ~n4663 & n5067 ;
  assign n24153 = n12140 ^ n7734 ^ 1'b0 ;
  assign n24154 = n3106 & n24153 ;
  assign n24155 = ~n21448 & n24154 ;
  assign n24156 = ~n19888 & n24155 ;
  assign n24158 = n24157 ^ n24156 ^ 1'b0 ;
  assign n24160 = ~n724 & n735 ;
  assign n24159 = n10268 ^ n3699 ^ 1'b0 ;
  assign n24161 = n24160 ^ n24159 ^ n11747 ;
  assign n24162 = n21446 ^ n3804 ^ 1'b0 ;
  assign n24163 = ~n10096 & n21694 ;
  assign n24164 = n24162 & n24163 ;
  assign n24165 = n4263 ^ n2140 ^ 1'b0 ;
  assign n24166 = n10809 ^ n6155 ^ 1'b0 ;
  assign n24169 = n7723 ^ n1739 ^ 1'b0 ;
  assign n24170 = n8954 ^ n2211 ^ 1'b0 ;
  assign n24171 = n24169 & n24170 ;
  assign n24168 = n608 | n1788 ;
  assign n24167 = n16686 ^ n13678 ^ 1'b0 ;
  assign n24172 = n24171 ^ n24168 ^ n24167 ;
  assign n24173 = n4128 & n24172 ;
  assign n24174 = n1204 | n10096 ;
  assign n24175 = n24174 ^ n9529 ^ 1'b0 ;
  assign n24176 = x159 | n1242 ;
  assign n24177 = n9230 & ~n24176 ;
  assign n24178 = n24177 ^ n19444 ^ 1'b0 ;
  assign n24179 = n7788 & ~n15194 ;
  assign n24180 = n24179 ^ x164 ^ 1'b0 ;
  assign n24181 = n4633 ^ n3620 ^ 1'b0 ;
  assign n24182 = n24181 ^ n21014 ^ 1'b0 ;
  assign n24183 = ~n7020 & n24182 ;
  assign n24184 = n3619 & ~n24183 ;
  assign n24185 = n3410 | n17089 ;
  assign n24186 = n3410 & ~n24185 ;
  assign n24187 = ~n3915 & n15875 ;
  assign n24188 = n7504 & n13981 ;
  assign n24189 = n8216 & n24188 ;
  assign n24190 = ( n7608 & n20575 ) | ( n7608 & ~n24189 ) | ( n20575 & ~n24189 ) ;
  assign n24191 = n17056 | n18492 ;
  assign n24193 = n9456 ^ n9215 ^ 1'b0 ;
  assign n24192 = n8265 & n14573 ;
  assign n24194 = n24193 ^ n24192 ^ n13759 ;
  assign n24195 = ~n13054 & n24194 ;
  assign n24196 = ~n6206 & n24195 ;
  assign n24197 = n5253 ^ n3313 ^ 1'b0 ;
  assign n24198 = n2433 & n24197 ;
  assign n24199 = ( ~n328 & n10034 ) | ( ~n328 & n24198 ) | ( n10034 & n24198 ) ;
  assign n24200 = n24199 ^ n19055 ^ 1'b0 ;
  assign n24201 = ~n7497 & n24200 ;
  assign n24202 = n6385 | n16532 ;
  assign n24203 = n4094 & ~n24202 ;
  assign n24204 = ( n3975 & n22114 ) | ( n3975 & ~n24203 ) | ( n22114 & ~n24203 ) ;
  assign n24205 = n4903 & ~n17197 ;
  assign n24206 = n24205 ^ n4042 ^ 1'b0 ;
  assign n24207 = n8508 ^ n8477 ^ 1'b0 ;
  assign n24208 = n6690 & n24207 ;
  assign n24209 = n24208 ^ n14227 ^ 1'b0 ;
  assign n24210 = n5984 ^ n3888 ^ 1'b0 ;
  assign n24211 = n14462 & n24210 ;
  assign n24212 = n10963 | n21048 ;
  assign n24213 = x215 & ~n1471 ;
  assign n24214 = ~n7005 & n24213 ;
  assign n24215 = n8224 | n9110 ;
  assign n24216 = n24215 ^ n10489 ^ 1'b0 ;
  assign n24217 = ( n2424 & n24214 ) | ( n2424 & n24216 ) | ( n24214 & n24216 ) ;
  assign n24218 = n5802 ^ n2625 ^ 1'b0 ;
  assign n24219 = n2064 & ~n24218 ;
  assign n24220 = n24219 ^ n15540 ^ 1'b0 ;
  assign n24221 = n9465 & n10303 ;
  assign n24222 = n24221 ^ n2246 ^ 1'b0 ;
  assign n24223 = n16332 & n24222 ;
  assign n24224 = n24223 ^ n23295 ^ 1'b0 ;
  assign n24225 = n8506 | n11880 ;
  assign n24226 = n14125 & ~n24225 ;
  assign n24228 = n23852 ^ n3011 ^ 1'b0 ;
  assign n24227 = n532 & n4037 ;
  assign n24229 = n24228 ^ n24227 ^ n8228 ;
  assign n24230 = n16622 ^ n15318 ^ 1'b0 ;
  assign n24231 = n3509 | n22732 ;
  assign n24232 = n24231 ^ n2043 ^ 1'b0 ;
  assign n24233 = n24230 & n24232 ;
  assign n24234 = n24233 ^ n13204 ^ 1'b0 ;
  assign n24235 = n24229 & n24234 ;
  assign n24237 = ~n804 & n7423 ;
  assign n24238 = n24237 ^ n3294 ^ 1'b0 ;
  assign n24236 = ~n14105 & n19549 ;
  assign n24239 = n24238 ^ n24236 ^ 1'b0 ;
  assign n24240 = n4425 & n6506 ;
  assign n24241 = n15693 & n24240 ;
  assign n24242 = n14371 | n24241 ;
  assign n24243 = n19458 | n24242 ;
  assign n24244 = n12928 | n23947 ;
  assign n24245 = n20314 ^ n296 ^ 1'b0 ;
  assign n24246 = ~n8963 & n17543 ;
  assign n24247 = n1848 & ~n24246 ;
  assign n24248 = n2798 & ~n10395 ;
  assign n24249 = ~n24247 & n24248 ;
  assign n24250 = n1620 | n2950 ;
  assign n24251 = n2881 & ~n24250 ;
  assign n24252 = n8440 & ~n24251 ;
  assign n24253 = n2466 ^ n1238 ^ 1'b0 ;
  assign n24254 = n17003 & n24253 ;
  assign n24255 = n18096 ^ n15765 ^ 1'b0 ;
  assign n24256 = n24254 & n24255 ;
  assign n24257 = ~n5500 & n11979 ;
  assign n24258 = ( ~n7130 & n13508 ) | ( ~n7130 & n24257 ) | ( n13508 & n24257 ) ;
  assign n24259 = n12754 & n24258 ;
  assign n24260 = n14234 ^ n4433 ^ 1'b0 ;
  assign n24262 = n9028 | n11316 ;
  assign n24263 = n6428 | n24262 ;
  assign n24261 = n13420 & ~n14064 ;
  assign n24264 = n24263 ^ n24261 ^ 1'b0 ;
  assign n24265 = n11607 ^ n9813 ^ 1'b0 ;
  assign n24266 = n3925 | n11000 ;
  assign n24267 = n17027 ^ n7906 ^ n3230 ;
  assign n24268 = n24267 ^ n5857 ^ 1'b0 ;
  assign n24269 = n24266 | n24268 ;
  assign n24270 = n6826 ^ n4970 ^ 1'b0 ;
  assign n24271 = n2098 & n24270 ;
  assign n24272 = n3397 & ~n16644 ;
  assign n24273 = n24272 ^ n15918 ^ 1'b0 ;
  assign n24274 = n4173 & n5269 ;
  assign n24275 = ( n5422 & n7825 ) | ( n5422 & ~n24274 ) | ( n7825 & ~n24274 ) ;
  assign n24276 = n24275 ^ n9998 ^ x187 ;
  assign n24277 = n24276 ^ n20908 ^ 1'b0 ;
  assign n24278 = n8613 ^ n2097 ^ 1'b0 ;
  assign n24280 = n14982 ^ n10822 ^ 1'b0 ;
  assign n24281 = n9873 | n24280 ;
  assign n24279 = n6791 | n16246 ;
  assign n24282 = n24281 ^ n24279 ^ 1'b0 ;
  assign n24283 = n20096 & n24282 ;
  assign n24284 = ~n2560 & n14296 ;
  assign n24285 = n9642 & ~n21814 ;
  assign n24286 = ~n8940 & n24285 ;
  assign n24287 = ~n24284 & n24286 ;
  assign n24288 = ( n9321 & n11465 ) | ( n9321 & ~n21909 ) | ( n11465 & ~n21909 ) ;
  assign n24289 = n8816 & ~n22363 ;
  assign n24290 = n22035 ^ n16801 ^ 1'b0 ;
  assign n24291 = n17543 & n24290 ;
  assign n24292 = n8216 | n10560 ;
  assign n24293 = n24292 ^ n13363 ^ n10663 ;
  assign n24294 = n16522 | n24293 ;
  assign n24295 = n17175 ^ n8140 ^ 1'b0 ;
  assign n24297 = n10275 & n11059 ;
  assign n24296 = n14312 & ~n24127 ;
  assign n24298 = n24297 ^ n24296 ^ n6421 ;
  assign n24299 = n22928 & n24298 ;
  assign n24300 = n13672 ^ n2466 ^ n2062 ;
  assign n24301 = n5245 ^ n4635 ^ 1'b0 ;
  assign n24302 = n842 | n24301 ;
  assign n24303 = n7266 ^ n2226 ^ 1'b0 ;
  assign n24304 = n739 & n12513 ;
  assign n24305 = n24304 ^ n6571 ^ 1'b0 ;
  assign n24306 = n914 | n15319 ;
  assign n24307 = n24306 ^ n6023 ^ 1'b0 ;
  assign n24308 = ~n14313 & n24307 ;
  assign n24309 = n24308 ^ n4370 ^ 1'b0 ;
  assign n24310 = ( n13275 & n15368 ) | ( n13275 & n22940 ) | ( n15368 & n22940 ) ;
  assign n24311 = n15977 & n22235 ;
  assign n24312 = n10007 ^ x10 ^ 1'b0 ;
  assign n24313 = n19066 ^ n6886 ^ 1'b0 ;
  assign n24314 = n24312 & n24313 ;
  assign n24315 = ( n21365 & ~n24311 ) | ( n21365 & n24314 ) | ( ~n24311 & n24314 ) ;
  assign n24316 = n9958 & ~n13217 ;
  assign n24317 = ~n4260 & n24316 ;
  assign n24318 = n24317 ^ n8582 ^ 1'b0 ;
  assign n24319 = n8921 & ~n24318 ;
  assign n24320 = n958 & ~n14525 ;
  assign n24321 = n19225 ^ n9967 ^ 1'b0 ;
  assign n24322 = n11256 & n18557 ;
  assign n24323 = n24322 ^ n5398 ^ 1'b0 ;
  assign n24324 = n24323 ^ n9691 ^ 1'b0 ;
  assign n24325 = n24324 ^ n13000 ^ n5847 ;
  assign n24326 = n1512 | n24325 ;
  assign n24327 = n13547 & n14957 ;
  assign n24328 = n24327 ^ n23806 ^ 1'b0 ;
  assign n24329 = n16479 ^ n5248 ^ 1'b0 ;
  assign n24330 = x140 & ~n300 ;
  assign n24331 = ~n9076 & n24330 ;
  assign n24332 = n24331 ^ n9623 ^ n3795 ;
  assign n24333 = n17894 ^ n5780 ^ n4031 ;
  assign n24334 = n24332 & ~n24333 ;
  assign n24335 = n1067 & n24334 ;
  assign n24336 = x233 & n1569 ;
  assign n24337 = ( ~n270 & n17035 ) | ( ~n270 & n24336 ) | ( n17035 & n24336 ) ;
  assign n24338 = n14994 ^ n13871 ^ 1'b0 ;
  assign n24339 = n18326 & n19440 ;
  assign n24340 = n24339 ^ n19169 ^ 1'b0 ;
  assign n24341 = ~n11863 & n13863 ;
  assign n24342 = n6155 & n24341 ;
  assign n24343 = n23856 ^ x194 ^ 1'b0 ;
  assign n24344 = n2400 | n6495 ;
  assign n24345 = n24344 ^ n19042 ^ 1'b0 ;
  assign n24346 = n24343 & ~n24345 ;
  assign n24347 = n22332 ^ n18221 ^ 1'b0 ;
  assign n24348 = n19386 & n24347 ;
  assign n24349 = n14350 ^ n5509 ^ 1'b0 ;
  assign n24350 = ~n16958 & n24349 ;
  assign n24351 = n24348 & n24350 ;
  assign n24352 = n14488 ^ n3288 ^ 1'b0 ;
  assign n24353 = n11002 | n24352 ;
  assign n24354 = n24353 ^ n4568 ^ n1121 ;
  assign n24355 = n7501 & ~n22523 ;
  assign n24356 = n12204 & n24355 ;
  assign n24357 = ~n7912 & n24356 ;
  assign n24358 = n5437 | n22879 ;
  assign n24359 = n5587 & n9496 ;
  assign n24360 = n17061 & n24359 ;
  assign n24361 = n6404 & ~n22675 ;
  assign n24362 = ~n6527 & n24361 ;
  assign n24363 = n16451 & n24362 ;
  assign n24364 = n2995 & n17638 ;
  assign n24365 = n4484 & n24364 ;
  assign n24366 = n24365 ^ n3817 ^ 1'b0 ;
  assign n24367 = ~n1500 & n9067 ;
  assign n24368 = n24367 ^ n5130 ^ n2452 ;
  assign n24369 = n20744 ^ n1561 ^ 1'b0 ;
  assign n24370 = ~n6220 & n24355 ;
  assign n24371 = n11558 | n17537 ;
  assign n24372 = n24030 ^ n16031 ^ 1'b0 ;
  assign n24373 = n3509 | n9902 ;
  assign n24374 = ~n6802 & n8766 ;
  assign n24375 = n9475 & n24374 ;
  assign n24376 = n24375 ^ n20249 ^ n6413 ;
  assign n24377 = ( n2794 & n5101 ) | ( n2794 & ~n19819 ) | ( n5101 & ~n19819 ) ;
  assign n24378 = n20444 ^ n15143 ^ n13533 ;
  assign n24379 = ~n3704 & n24378 ;
  assign n24380 = n12148 ^ n8011 ^ 1'b0 ;
  assign n24381 = ~n589 & n5339 ;
  assign n24382 = n9981 ^ n8772 ^ 1'b0 ;
  assign n24383 = ( n9256 & n11722 ) | ( n9256 & n24382 ) | ( n11722 & n24382 ) ;
  assign n24384 = n7872 & n14711 ;
  assign n24385 = n15637 ^ n13552 ^ 1'b0 ;
  assign n24386 = n15730 ^ n3198 ^ n2790 ;
  assign n24387 = n12539 ^ n3425 ^ 1'b0 ;
  assign n24388 = n24386 & ~n24387 ;
  assign n24389 = n10849 ^ n8428 ^ 1'b0 ;
  assign n24390 = n16614 ^ n13221 ^ n11206 ;
  assign n24391 = n19741 ^ n19640 ^ 1'b0 ;
  assign n24392 = n11660 ^ n7002 ^ 1'b0 ;
  assign n24393 = n4315 & n6252 ;
  assign n24394 = n10840 & n24393 ;
  assign n24395 = n24394 ^ n12471 ^ 1'b0 ;
  assign n24396 = n7605 & ~n19583 ;
  assign n24397 = ~n309 & n24396 ;
  assign n24398 = n7561 ^ n6376 ^ 1'b0 ;
  assign n24399 = n751 | n24398 ;
  assign n24400 = n4220 & n24399 ;
  assign n24403 = n4031 | n6350 ;
  assign n24404 = ( n6060 & n12198 ) | ( n6060 & n24403 ) | ( n12198 & n24403 ) ;
  assign n24401 = n5607 & n19535 ;
  assign n24402 = n23832 & n24401 ;
  assign n24405 = n24404 ^ n24402 ^ 1'b0 ;
  assign n24406 = n18630 ^ n3915 ^ 1'b0 ;
  assign n24407 = ~n1680 & n24406 ;
  assign n24408 = n8048 | n18267 ;
  assign n24409 = ~n4282 & n13317 ;
  assign n24410 = ~n4424 & n24409 ;
  assign n24411 = n24410 ^ n12111 ^ 1'b0 ;
  assign n24412 = x29 & ~n2254 ;
  assign n24413 = n24412 ^ n3444 ^ 1'b0 ;
  assign n24414 = n24413 ^ n8839 ^ 1'b0 ;
  assign n24415 = n19897 ^ n10247 ^ 1'b0 ;
  assign n24416 = n1833 & n24415 ;
  assign n24417 = n21538 & n24416 ;
  assign n24418 = n24417 ^ n21351 ^ 1'b0 ;
  assign n24419 = ~n18136 & n24418 ;
  assign n24420 = n24414 & n24419 ;
  assign n24421 = n14312 | n24420 ;
  assign n24422 = n24421 ^ n1589 ^ 1'b0 ;
  assign n24423 = n5596 & n9623 ;
  assign n24424 = ~n3274 & n24423 ;
  assign n24425 = n6093 | n8352 ;
  assign n24426 = n24424 & ~n24425 ;
  assign n24427 = n7582 ^ n5690 ^ n1267 ;
  assign n24428 = n2580 & n24427 ;
  assign n24429 = n23396 & n24428 ;
  assign n24430 = n16536 ^ x112 ^ 1'b0 ;
  assign n24431 = ~n24286 & n24430 ;
  assign n24432 = ~n24429 & n24431 ;
  assign n24433 = n2872 ^ n2149 ^ n928 ;
  assign n24434 = ( ~x130 & n18492 ) | ( ~x130 & n24433 ) | ( n18492 & n24433 ) ;
  assign n24435 = n13981 ^ n10244 ^ 1'b0 ;
  assign n24436 = n8363 | n11810 ;
  assign n24437 = n1846 & ~n24436 ;
  assign n24438 = n19394 & ~n24437 ;
  assign n24439 = n12413 & n21580 ;
  assign n24440 = n24439 ^ n14852 ^ 1'b0 ;
  assign n24441 = n24440 ^ n8729 ^ 1'b0 ;
  assign n24442 = n24438 & n24441 ;
  assign n24443 = n1680 | n7596 ;
  assign n24444 = n24443 ^ n12922 ^ 1'b0 ;
  assign n24445 = n20915 | n24444 ;
  assign n24446 = n3416 | n14504 ;
  assign n24447 = n2041 & n23955 ;
  assign n24448 = n2959 & ~n11868 ;
  assign n24449 = ~n1964 & n9701 ;
  assign n24450 = n1664 & ~n24449 ;
  assign n24453 = n20014 ^ n7871 ^ n6286 ;
  assign n24451 = n5511 ^ n5018 ^ 1'b0 ;
  assign n24452 = n3769 & n24451 ;
  assign n24454 = n24453 ^ n24452 ^ n20249 ;
  assign n24455 = n11519 ^ n7939 ^ n6707 ;
  assign n24456 = n1634 & ~n24455 ;
  assign n24457 = n24456 ^ n5610 ^ 1'b0 ;
  assign n24458 = n24457 ^ n12210 ^ 1'b0 ;
  assign n24459 = n23255 & ~n24458 ;
  assign n24460 = n4875 ^ n1749 ^ 1'b0 ;
  assign n24461 = n22520 & ~n24460 ;
  assign n24462 = n13006 & ~n24461 ;
  assign n24463 = n24462 ^ n2330 ^ 1'b0 ;
  assign n24464 = n17305 & n20118 ;
  assign n24465 = n24464 ^ n5659 ^ 1'b0 ;
  assign n24466 = n24465 ^ n14789 ^ 1'b0 ;
  assign n24467 = n7219 & n11260 ;
  assign n24468 = ~n4340 & n24467 ;
  assign n24469 = n2362 & ~n24468 ;
  assign n24470 = n24469 ^ n17033 ^ 1'b0 ;
  assign n24471 = n17968 ^ n5811 ^ 1'b0 ;
  assign n24472 = n12170 ^ n10840 ^ 1'b0 ;
  assign n24473 = n19641 & ~n24472 ;
  assign n24474 = n10377 ^ n4811 ^ n703 ;
  assign n24475 = n18732 ^ n3081 ^ 1'b0 ;
  assign n24476 = ~n24474 & n24475 ;
  assign n24477 = n24476 ^ n18444 ^ 1'b0 ;
  assign n24478 = n3589 | n24477 ;
  assign n24479 = n24473 | n24478 ;
  assign n24480 = n11059 | n12541 ;
  assign n24481 = n24480 ^ n11285 ^ 1'b0 ;
  assign n24483 = n6991 ^ n6043 ^ n2502 ;
  assign n24484 = n5307 | n24483 ;
  assign n24482 = ~n11382 & n19837 ;
  assign n24485 = n24484 ^ n24482 ^ 1'b0 ;
  assign n24486 = ( n4871 & ~n5423 ) | ( n4871 & n5717 ) | ( ~n5423 & n5717 ) ;
  assign n24487 = n4386 & ~n19603 ;
  assign n24488 = ~n24486 & n24487 ;
  assign n24489 = n1138 & n17288 ;
  assign n24490 = n4285 & ~n9276 ;
  assign n24491 = n24490 ^ n430 ^ 1'b0 ;
  assign n24492 = n24491 ^ n7117 ^ 1'b0 ;
  assign n24493 = n12053 & ~n24063 ;
  assign n24494 = n24493 ^ n17369 ^ 1'b0 ;
  assign n24495 = n19501 ^ n1440 ^ 1'b0 ;
  assign n24496 = n23728 | n24495 ;
  assign n24497 = x40 | n24331 ;
  assign n24498 = n19528 ^ n1729 ^ 1'b0 ;
  assign n24499 = n11371 | n24498 ;
  assign n24500 = ( n3546 & ~n8167 ) | ( n3546 & n15857 ) | ( ~n8167 & n15857 ) ;
  assign n24501 = ~n1633 & n12562 ;
  assign n24502 = n8300 | n24501 ;
  assign n24503 = n24502 ^ n15300 ^ 1'b0 ;
  assign n24504 = n15088 & n24503 ;
  assign n24505 = ~n11905 & n24504 ;
  assign n24506 = n24505 ^ n655 ^ 1'b0 ;
  assign n24507 = n21145 & n24506 ;
  assign n24508 = n20211 ^ n3172 ^ 1'b0 ;
  assign n24509 = n12775 ^ n11130 ^ 1'b0 ;
  assign n24510 = n11609 & n24509 ;
  assign n24511 = n22951 ^ n1101 ^ 1'b0 ;
  assign n24512 = x196 & n23036 ;
  assign n24513 = n1405 & n24512 ;
  assign n24514 = n24513 ^ n15240 ^ 1'b0 ;
  assign n24515 = n15332 ^ n2815 ^ 1'b0 ;
  assign n24516 = ~n24514 & n24515 ;
  assign n24517 = n973 | n19504 ;
  assign n24518 = n24516 | n24517 ;
  assign n24519 = n6868 ^ n5847 ^ 1'b0 ;
  assign n24520 = ~x181 & n24519 ;
  assign n24521 = n8473 | n10194 ;
  assign n24522 = n21592 | n24521 ;
  assign n24524 = n1112 | n3801 ;
  assign n24525 = n812 | n24524 ;
  assign n24523 = n3989 & n9076 ;
  assign n24526 = n24525 ^ n24523 ^ 1'b0 ;
  assign n24527 = n10114 & n11068 ;
  assign n24528 = n3696 & n24527 ;
  assign n24529 = ( n716 & n24526 ) | ( n716 & n24528 ) | ( n24526 & n24528 ) ;
  assign n24530 = n11091 | n12004 ;
  assign n24531 = n7387 ^ n5261 ^ n1135 ;
  assign n24532 = n13796 & ~n24531 ;
  assign n24533 = ( n2807 & n6432 ) | ( n2807 & ~n22122 ) | ( n6432 & ~n22122 ) ;
  assign n24534 = n877 & ~n7550 ;
  assign n24535 = n20071 & n24534 ;
  assign n24536 = n4149 & n13317 ;
  assign n24537 = ~n12798 & n24536 ;
  assign n24538 = n8664 & ~n24537 ;
  assign n24539 = n24538 ^ n16020 ^ 1'b0 ;
  assign n24540 = n20898 ^ n14705 ^ n2409 ;
  assign n24541 = n13942 & n24540 ;
  assign n24542 = n2949 & ~n16575 ;
  assign n24543 = ~n19064 & n24542 ;
  assign n24544 = n7407 & n10556 ;
  assign n24545 = n24544 ^ n15088 ^ n5665 ;
  assign n24546 = n8730 ^ n4420 ^ n749 ;
  assign n24547 = ~n1874 & n24546 ;
  assign n24548 = n24545 & n24547 ;
  assign n24549 = n8959 ^ n825 ^ 1'b0 ;
  assign n24550 = ~n7405 & n9180 ;
  assign n24551 = n24549 & n24550 ;
  assign n24552 = n6064 & ~n6415 ;
  assign n24553 = n8974 | n24552 ;
  assign n24554 = n7704 ^ n2120 ^ n527 ;
  assign n24555 = ~n3631 & n8356 ;
  assign n24557 = ( n1553 & n11755 ) | ( n1553 & n11935 ) | ( n11755 & n11935 ) ;
  assign n24556 = n6271 & ~n18894 ;
  assign n24558 = n24557 ^ n24556 ^ 1'b0 ;
  assign n24559 = ~n3213 & n11605 ;
  assign n24560 = n24558 & n24559 ;
  assign n24561 = ~n5829 & n8976 ;
  assign n24562 = n24561 ^ n14589 ^ 1'b0 ;
  assign n24563 = n15003 | n16379 ;
  assign n24564 = n24563 ^ n2622 ^ 1'b0 ;
  assign n24565 = n5927 & n19005 ;
  assign n24566 = n19885 ^ n378 ^ 1'b0 ;
  assign n24567 = n2978 & n8891 ;
  assign n24568 = ~n6581 & n24567 ;
  assign n24569 = n24568 ^ n21750 ^ 1'b0 ;
  assign n24570 = n6826 | n12308 ;
  assign n24571 = n1206 | n1365 ;
  assign n24572 = n8595 | n24571 ;
  assign n24573 = x119 & ~n3007 ;
  assign n24574 = n24573 ^ n8275 ^ 1'b0 ;
  assign n24575 = n24572 & ~n24574 ;
  assign n24576 = x159 & ~n6226 ;
  assign n24577 = x143 & n24576 ;
  assign n24578 = n13258 & ~n24577 ;
  assign n24579 = n16593 & n24578 ;
  assign n24581 = ~n1797 & n2208 ;
  assign n24580 = n10397 & n19535 ;
  assign n24582 = n24581 ^ n24580 ^ 1'b0 ;
  assign n24583 = n10934 & n15294 ;
  assign n24584 = n24583 ^ n2768 ^ 1'b0 ;
  assign n24585 = n1935 ^ n366 ^ 1'b0 ;
  assign n24586 = n24584 & ~n24585 ;
  assign n24587 = ~n10215 & n13077 ;
  assign n24588 = n996 & n24587 ;
  assign n24589 = n12308 & n16923 ;
  assign n24590 = ~n13309 & n18350 ;
  assign n24591 = ~n21373 & n24590 ;
  assign n24592 = n12680 ^ n11743 ^ 1'b0 ;
  assign n24593 = n24592 ^ n15979 ^ 1'b0 ;
  assign n24594 = ~n12148 & n24593 ;
  assign n24595 = n22618 ^ n19344 ^ 1'b0 ;
  assign n24596 = n19901 ^ n2067 ^ 1'b0 ;
  assign n24597 = n24595 & n24596 ;
  assign n24598 = n23070 ^ n13230 ^ 1'b0 ;
  assign n24599 = n8172 | n24598 ;
  assign n24601 = n1671 ^ x73 ^ 1'b0 ;
  assign n24602 = n2041 & n24601 ;
  assign n24600 = ( ~n1749 & n10526 ) | ( ~n1749 & n12576 ) | ( n10526 & n12576 ) ;
  assign n24603 = n24602 ^ n24600 ^ 1'b0 ;
  assign n24604 = n12123 | n19673 ;
  assign n24605 = n24603 & ~n24604 ;
  assign n24606 = n7940 & n7996 ;
  assign n24607 = ~n4047 & n24606 ;
  assign n24609 = ~n5195 & n21188 ;
  assign n24610 = ~n4799 & n24609 ;
  assign n24611 = n24610 ^ n4498 ^ 1'b0 ;
  assign n24612 = n2920 | n24611 ;
  assign n24608 = n1312 & n19035 ;
  assign n24613 = n24612 ^ n24608 ^ 1'b0 ;
  assign n24614 = n3106 | n20753 ;
  assign n24615 = n24614 ^ n15192 ^ 1'b0 ;
  assign n24616 = n3454 & ~n7638 ;
  assign n24617 = ~n24615 & n24616 ;
  assign n24618 = n24617 ^ n23871 ^ 1'b0 ;
  assign n24619 = n1931 ^ n1286 ^ 1'b0 ;
  assign n24620 = n3944 & n20010 ;
  assign n24621 = ~n10834 & n24620 ;
  assign n24622 = n24621 ^ n4139 ^ 1'b0 ;
  assign n24623 = n17555 ^ n5556 ^ 1'b0 ;
  assign n24625 = n10871 ^ n3532 ^ 1'b0 ;
  assign n24624 = n1803 ^ n1369 ^ 1'b0 ;
  assign n24626 = n24625 ^ n24624 ^ 1'b0 ;
  assign n24627 = n24626 ^ n9189 ^ 1'b0 ;
  assign n24628 = n18653 & ~n24627 ;
  assign n24629 = ~n15711 & n18219 ;
  assign n24630 = ~n24628 & n24629 ;
  assign n24631 = n729 | n8587 ;
  assign n24632 = n24631 ^ n8663 ^ 1'b0 ;
  assign n24633 = n10805 ^ n1008 ^ 1'b0 ;
  assign n24634 = n8291 & ~n11730 ;
  assign n24635 = ~n24633 & n24634 ;
  assign n24636 = n19443 ^ n7939 ^ 1'b0 ;
  assign n24637 = n24635 | n24636 ;
  assign n24638 = n1899 & ~n12703 ;
  assign n24639 = n2469 & ~n5537 ;
  assign n24640 = n9024 & ~n13411 ;
  assign n24641 = n4677 & ~n19980 ;
  assign n24642 = n24641 ^ n10042 ^ 1'b0 ;
  assign n24643 = n6088 ^ n4417 ^ 1'b0 ;
  assign n24644 = n1534 & ~n24643 ;
  assign n24645 = n9461 & ~n18502 ;
  assign n24646 = ~n4553 & n24645 ;
  assign n24647 = n24646 ^ n1219 ^ 1'b0 ;
  assign n24648 = n4222 & ~n24647 ;
  assign n24649 = n6853 & n24648 ;
  assign n24650 = ( n19075 & ~n24644 ) | ( n19075 & n24649 ) | ( ~n24644 & n24649 ) ;
  assign n24651 = n2681 | n7751 ;
  assign n24652 = n6527 & ~n16663 ;
  assign n24653 = n9965 & n19145 ;
  assign n24654 = n2338 | n18590 ;
  assign n24655 = n24654 ^ n6201 ^ 1'b0 ;
  assign n24658 = n20818 ^ n13845 ^ 1'b0 ;
  assign n24656 = n12074 & ~n13070 ;
  assign n24657 = n2972 & n24656 ;
  assign n24659 = n24658 ^ n24657 ^ n4612 ;
  assign n24660 = n1137 ^ n1083 ^ x31 ;
  assign n24661 = n24660 ^ n13373 ^ 1'b0 ;
  assign n24663 = ~n3791 & n6470 ;
  assign n24664 = n3791 & n24663 ;
  assign n24665 = n1328 | n24664 ;
  assign n24666 = n1328 & ~n24665 ;
  assign n24667 = n24666 ^ n18813 ^ 1'b0 ;
  assign n24662 = n1701 | n22218 ;
  assign n24668 = n24667 ^ n24662 ^ 1'b0 ;
  assign n24669 = n13892 ^ n10520 ^ 1'b0 ;
  assign n24670 = n13991 ^ n7212 ^ 1'b0 ;
  assign n24671 = n20292 | n24670 ;
  assign n24672 = ( ~n13144 & n24669 ) | ( ~n13144 & n24671 ) | ( n24669 & n24671 ) ;
  assign n24673 = n9605 & n23073 ;
  assign n24674 = n13976 & ~n24136 ;
  assign n24675 = n14514 | n19839 ;
  assign n24676 = n24675 ^ n2525 ^ 1'b0 ;
  assign n24677 = n13776 ^ n4621 ^ 1'b0 ;
  assign n24681 = ~n9931 & n18259 ;
  assign n24682 = ~n7632 & n24681 ;
  assign n24678 = n24053 ^ n8004 ^ 1'b0 ;
  assign n24679 = ~n14756 & n21810 ;
  assign n24680 = n24678 & n24679 ;
  assign n24683 = n24682 ^ n24680 ^ 1'b0 ;
  assign n24684 = n11511 & ~n19208 ;
  assign n24685 = n7328 ^ n4092 ^ n564 ;
  assign n24686 = n1535 | n22824 ;
  assign n24687 = n829 | n6572 ;
  assign n24688 = n13664 & n24687 ;
  assign n24689 = n10024 ^ n5585 ^ 1'b0 ;
  assign n24690 = n5462 & ~n24689 ;
  assign n24691 = n10414 & n12266 ;
  assign n24692 = n6794 & ~n17977 ;
  assign n24693 = ~n20219 & n24692 ;
  assign n24694 = n24623 & ~n24693 ;
  assign n24695 = n24691 & n24694 ;
  assign n24696 = n15240 ^ n8970 ^ 1'b0 ;
  assign n24697 = n3420 & n9064 ;
  assign n24698 = n1600 ^ n309 ^ 1'b0 ;
  assign n24699 = n5097 | n24698 ;
  assign n24700 = n11366 ^ n4326 ^ 1'b0 ;
  assign n24701 = ~n13104 & n16177 ;
  assign n24702 = n4554 & ~n5401 ;
  assign n24703 = ~n16030 & n24702 ;
  assign n24704 = n11810 & ~n16187 ;
  assign n24705 = ( n940 & n5626 ) | ( n940 & ~n14259 ) | ( n5626 & ~n14259 ) ;
  assign n24706 = ~n7745 & n24705 ;
  assign n24707 = n16439 & n24706 ;
  assign n24708 = ~n679 & n9264 ;
  assign n24709 = ~n8005 & n9290 ;
  assign n24710 = n14428 ^ n7355 ^ n3680 ;
  assign n24711 = n9636 & ~n10809 ;
  assign n24712 = n24711 ^ n21686 ^ 1'b0 ;
  assign n24713 = n3038 ^ n2951 ^ x94 ;
  assign n24714 = n625 & n24713 ;
  assign n24715 = n24714 ^ n3694 ^ 1'b0 ;
  assign n24716 = n14062 & ~n24715 ;
  assign n24717 = n24716 ^ n1882 ^ 1'b0 ;
  assign n24718 = n16944 & n23856 ;
  assign n24719 = n4627 & n23051 ;
  assign n24720 = n24719 ^ n2615 ^ 1'b0 ;
  assign n24721 = n5104 & ~n11531 ;
  assign n24722 = n24721 ^ n19110 ^ n3761 ;
  assign n24723 = n1968 & n1993 ;
  assign n24724 = n6745 & n17789 ;
  assign n24725 = ~n4117 & n5216 ;
  assign n24726 = n24725 ^ n2903 ^ 1'b0 ;
  assign n24727 = n24726 ^ n11935 ^ 1'b0 ;
  assign n24728 = ~n24724 & n24727 ;
  assign n24729 = n2532 & ~n16225 ;
  assign n24730 = n10864 ^ n8969 ^ 1'b0 ;
  assign n24731 = n22599 ^ n1170 ^ 1'b0 ;
  assign n24732 = n24183 | n24731 ;
  assign n24733 = n11649 ^ n6121 ^ 1'b0 ;
  assign n24734 = n642 | n3039 ;
  assign n24735 = n24702 & ~n24734 ;
  assign n24736 = n24735 ^ x40 ^ 1'b0 ;
  assign n24737 = ~n3592 & n24736 ;
  assign n24738 = n24737 ^ n3685 ^ 1'b0 ;
  assign n24739 = n15308 & n24738 ;
  assign n24740 = ( ~n15348 & n24733 ) | ( ~n15348 & n24739 ) | ( n24733 & n24739 ) ;
  assign n24741 = ~n4488 & n6376 ;
  assign n24742 = n24741 ^ n7212 ^ 1'b0 ;
  assign n24743 = n5927 | n24742 ;
  assign n24744 = n2898 & ~n18256 ;
  assign n24745 = ~n14183 & n24744 ;
  assign n24746 = n16300 & ~n24745 ;
  assign n24747 = n3861 & ~n14830 ;
  assign n24748 = n21104 ^ n5704 ^ 1'b0 ;
  assign n24749 = n4197 | n6405 ;
  assign n24750 = n1586 | n3908 ;
  assign n24751 = n1728 & ~n24750 ;
  assign n24752 = n24751 ^ n6423 ^ 1'b0 ;
  assign n24753 = n11839 & n24752 ;
  assign n24754 = n15979 ^ n14055 ^ 1'b0 ;
  assign n24755 = n22800 & n24754 ;
  assign n24756 = ( n17183 & ~n21600 ) | ( n17183 & n24755 ) | ( ~n21600 & n24755 ) ;
  assign n24757 = n15886 | n24756 ;
  assign n24758 = n24757 ^ n9651 ^ 1'b0 ;
  assign n24759 = n16439 ^ n2958 ^ 1'b0 ;
  assign n24760 = n3196 & n24759 ;
  assign n24761 = n7107 & ~n15228 ;
  assign n24762 = ~n3860 & n24761 ;
  assign n24763 = n6826 ^ n4875 ^ 1'b0 ;
  assign n24764 = n24763 ^ n5528 ^ 1'b0 ;
  assign n24765 = n24764 ^ n17274 ^ 1'b0 ;
  assign n24766 = ~n10331 & n24765 ;
  assign n24767 = n24766 ^ n18857 ^ 1'b0 ;
  assign n24768 = ~n8820 & n24767 ;
  assign n24769 = ~n17943 & n24768 ;
  assign n24770 = n5833 & n15245 ;
  assign n24771 = n6278 ^ n372 ^ 1'b0 ;
  assign n24772 = n24770 & n24771 ;
  assign n24773 = n2022 ^ n854 ^ 1'b0 ;
  assign n24774 = n17262 & n24773 ;
  assign n24775 = ~n9679 & n24774 ;
  assign n24776 = n8297 & ~n11862 ;
  assign n24777 = n24776 ^ n2657 ^ 1'b0 ;
  assign n24778 = n24775 | n24777 ;
  assign n24779 = n14464 ^ n858 ^ 1'b0 ;
  assign n24780 = n24735 ^ n11860 ^ n8474 ;
  assign n24781 = n3380 ^ n3081 ^ 1'b0 ;
  assign n24782 = n4712 | n17925 ;
  assign n24783 = ~n3770 & n16196 ;
  assign n24784 = n20241 ^ n12696 ^ n12536 ;
  assign n24788 = n283 & n880 ;
  assign n24789 = ~n880 & n24788 ;
  assign n24790 = n1748 & n1813 ;
  assign n24791 = n24789 & n24790 ;
  assign n24785 = n885 | n2395 ;
  assign n24786 = n2395 & ~n24785 ;
  assign n24787 = n2988 | n24786 ;
  assign n24792 = n24791 ^ n24787 ^ 1'b0 ;
  assign n24793 = n1161 & ~n9679 ;
  assign n24794 = n9679 & n24793 ;
  assign n24795 = n4420 & ~n24794 ;
  assign n24796 = n24792 & n24795 ;
  assign n24797 = n10374 ^ n6431 ^ 1'b0 ;
  assign n24798 = n20769 & ~n24797 ;
  assign n24799 = n7358 & ~n14522 ;
  assign n24800 = n12078 & n19832 ;
  assign n24801 = n6557 & ~n15826 ;
  assign n24802 = n24801 ^ n8258 ^ 1'b0 ;
  assign n24803 = n13300 & ~n24545 ;
  assign n24804 = n20295 ^ n2330 ^ 1'b0 ;
  assign n24805 = n24759 ^ n11487 ^ n2529 ;
  assign n24806 = n2959 & ~n24805 ;
  assign n24807 = n24806 ^ n21919 ^ 1'b0 ;
  assign n24808 = n3704 ^ n792 ^ 1'b0 ;
  assign n24809 = x247 | n24808 ;
  assign n24810 = n24809 ^ n14795 ^ n3760 ;
  assign n24811 = n8632 & ~n16674 ;
  assign n24812 = ~n3327 & n6230 ;
  assign n24813 = ~n1454 & n24812 ;
  assign n24814 = n9510 & ~n24813 ;
  assign n24816 = n18679 ^ n14964 ^ 1'b0 ;
  assign n24817 = n10639 & n24816 ;
  assign n24815 = n14612 | n22632 ;
  assign n24818 = n24817 ^ n24815 ^ 1'b0 ;
  assign n24819 = n8256 & ~n13849 ;
  assign n24820 = n5994 & ~n20245 ;
  assign n24821 = n2248 & n24820 ;
  assign n24822 = ~n1062 & n11459 ;
  assign n24823 = n24822 ^ n13962 ^ 1'b0 ;
  assign n24824 = n3649 & n24823 ;
  assign n24825 = n16882 & n24824 ;
  assign n24826 = n24825 ^ n24011 ^ 1'b0 ;
  assign n24827 = n899 & n11839 ;
  assign n24828 = n8843 | n17343 ;
  assign n24829 = n24827 | n24828 ;
  assign n24830 = n7863 & ~n15789 ;
  assign n24831 = ~n11416 & n24830 ;
  assign n24832 = n2657 | n24831 ;
  assign n24833 = n20832 | n24832 ;
  assign n24834 = x61 & ~n9847 ;
  assign n24835 = n1588 ^ n1352 ^ 1'b0 ;
  assign n24836 = n5625 & n24835 ;
  assign n24837 = ~n21705 & n24836 ;
  assign n24843 = n15282 & n18562 ;
  assign n24844 = ~n6912 & n24843 ;
  assign n24838 = ( ~n1351 & n3180 ) | ( ~n1351 & n22122 ) | ( n3180 & n22122 ) ;
  assign n24839 = n24838 ^ n10554 ^ 1'b0 ;
  assign n24840 = n21674 ^ n18856 ^ 1'b0 ;
  assign n24841 = n24839 & ~n24840 ;
  assign n24842 = ~n15074 & n24841 ;
  assign n24845 = n24844 ^ n24842 ^ 1'b0 ;
  assign n24846 = n4220 & n6499 ;
  assign n24847 = n1956 | n12765 ;
  assign n24848 = n1189 & ~n24847 ;
  assign n24849 = ~n20233 & n24848 ;
  assign n24850 = n5971 ^ n361 ^ 1'b0 ;
  assign n24851 = n11026 & ~n24850 ;
  assign n24852 = n24851 ^ x198 ^ 1'b0 ;
  assign n24853 = ~n16753 & n20715 ;
  assign n24854 = n3795 ^ n3435 ^ 1'b0 ;
  assign n24855 = n20075 ^ n14016 ^ 1'b0 ;
  assign n24856 = n20236 ^ n10882 ^ 1'b0 ;
  assign n24857 = n12300 & n13011 ;
  assign n24858 = ~n14930 & n24857 ;
  assign n24859 = n24858 ^ n3329 ^ 1'b0 ;
  assign n24860 = n8489 ^ n4074 ^ 1'b0 ;
  assign n24861 = n4686 & n12994 ;
  assign n24862 = n8375 & n24861 ;
  assign n24863 = n24862 ^ n10250 ^ 1'b0 ;
  assign n24864 = n5117 & ~n24863 ;
  assign n24865 = n10932 & ~n14511 ;
  assign n24866 = ~n6951 & n13231 ;
  assign n24867 = n24866 ^ n1748 ^ 1'b0 ;
  assign n24868 = n24867 ^ n16801 ^ 1'b0 ;
  assign n24869 = n24865 | n24868 ;
  assign n24870 = ~n3288 & n10809 ;
  assign n24871 = n3922 & n24870 ;
  assign n24872 = n6186 & n6718 ;
  assign n24873 = ~n24871 & n24872 ;
  assign n24874 = n9916 ^ n6522 ^ 1'b0 ;
  assign n24875 = n6644 ^ n5050 ^ n1290 ;
  assign n24876 = n24875 ^ n1982 ^ 1'b0 ;
  assign n24877 = n754 | n24876 ;
  assign n24880 = ~n3427 & n4964 ;
  assign n24881 = ~n6064 & n24880 ;
  assign n24878 = n2946 & ~n13476 ;
  assign n24879 = n24878 ^ n11685 ^ 1'b0 ;
  assign n24882 = n24881 ^ n24879 ^ 1'b0 ;
  assign n24883 = ~n24877 & n24882 ;
  assign n24884 = n3970 | n5165 ;
  assign n24885 = n731 & ~n24884 ;
  assign n24886 = n6289 ^ n1495 ^ 1'b0 ;
  assign n24887 = n4303 & ~n24886 ;
  assign n24888 = ~n24885 & n24887 ;
  assign n24889 = n24888 ^ n858 ^ 1'b0 ;
  assign n24890 = n853 ^ n842 ^ 1'b0 ;
  assign n24891 = n10775 & ~n24890 ;
  assign n24892 = n24891 ^ n12140 ^ 1'b0 ;
  assign n24893 = n3440 & n24892 ;
  assign n24894 = n9829 & n16318 ;
  assign n24895 = ~n11542 & n24894 ;
  assign n24896 = n14471 & n22719 ;
  assign n24897 = n24896 ^ n18168 ^ 1'b0 ;
  assign n24898 = n7866 & ~n21800 ;
  assign n24899 = n11078 ^ n545 ^ 1'b0 ;
  assign n24900 = n12128 | n24899 ;
  assign n24901 = n2576 | n4632 ;
  assign n24902 = n8629 & n14829 ;
  assign n24903 = n10201 & n24902 ;
  assign n24904 = n3565 & ~n24903 ;
  assign n24905 = ~n24901 & n24904 ;
  assign n24906 = n9872 ^ n4621 ^ 1'b0 ;
  assign n24907 = n7022 | n15479 ;
  assign n24908 = n7450 & n24907 ;
  assign n24909 = n12590 & n24908 ;
  assign n24910 = n24909 ^ n24372 ^ 1'b0 ;
  assign n24911 = n12142 ^ n2446 ^ 1'b0 ;
  assign n24912 = n9281 | n24911 ;
  assign n24913 = ~x162 & n7329 ;
  assign n24914 = x80 & ~n3496 ;
  assign n24915 = ( ~n6773 & n8311 ) | ( ~n6773 & n9959 ) | ( n8311 & n9959 ) ;
  assign n24916 = n4022 & ~n24915 ;
  assign n24917 = n24916 ^ n291 ^ 1'b0 ;
  assign n24918 = n17791 ^ n10839 ^ 1'b0 ;
  assign n24919 = n24917 & n24918 ;
  assign n24920 = ( ~n7145 & n7562 ) | ( ~n7145 & n14456 ) | ( n7562 & n14456 ) ;
  assign n24921 = n24920 ^ n10010 ^ 1'b0 ;
  assign n24922 = ~n9777 & n24921 ;
  assign n24923 = n7662 & ~n15003 ;
  assign n24924 = n24923 ^ n21319 ^ 1'b0 ;
  assign n24925 = n6059 & n24924 ;
  assign n24926 = ~n12627 & n17283 ;
  assign n24927 = n15027 ^ n14642 ^ n7916 ;
  assign n24928 = ~n7594 & n7911 ;
  assign n24932 = ~n16968 & n18476 ;
  assign n24929 = n7196 | n9700 ;
  assign n24930 = ( n4721 & ~n15840 ) | ( n4721 & n21179 ) | ( ~n15840 & n21179 ) ;
  assign n24931 = n24929 | n24930 ;
  assign n24933 = n24932 ^ n24931 ^ 1'b0 ;
  assign n24934 = n1754 | n1778 ;
  assign n24935 = n264 ^ x125 ^ 1'b0 ;
  assign n24936 = n7846 & ~n24935 ;
  assign n24937 = ~n12369 & n24936 ;
  assign n24938 = n24934 & n24937 ;
  assign n24939 = n5909 ^ n3294 ^ 1'b0 ;
  assign n24940 = n10529 & n13615 ;
  assign n24941 = n24940 ^ n16214 ^ 1'b0 ;
  assign n24942 = n24941 ^ n16370 ^ 1'b0 ;
  assign n24943 = n11719 & n21282 ;
  assign n24944 = n24943 ^ n18034 ^ 1'b0 ;
  assign n24945 = n20141 ^ n14935 ^ 1'b0 ;
  assign n24946 = n18367 ^ n11473 ^ 1'b0 ;
  assign n24947 = n24678 | n24946 ;
  assign n24948 = n24947 ^ n915 ^ 1'b0 ;
  assign n24949 = n1890 | n9783 ;
  assign n24950 = n24949 ^ n3825 ^ 1'b0 ;
  assign n24951 = n21045 & n24950 ;
  assign n24952 = n7792 & n24951 ;
  assign n24953 = n16025 ^ n13375 ^ 1'b0 ;
  assign n24954 = n8842 & n24953 ;
  assign n24955 = n10277 & ~n24954 ;
  assign n24956 = n11563 ^ n3647 ^ n1051 ;
  assign n24957 = n24554 & n24956 ;
  assign n24958 = n24957 ^ n20043 ^ 1'b0 ;
  assign n24959 = n11177 ^ n1133 ^ 1'b0 ;
  assign n24960 = n4260 & ~n24959 ;
  assign n24961 = ~n4111 & n24960 ;
  assign n24962 = ~n16037 & n24961 ;
  assign n24965 = n7181 ^ n1854 ^ 1'b0 ;
  assign n24966 = n24965 ^ n5205 ^ 1'b0 ;
  assign n24967 = n4493 | n24966 ;
  assign n24968 = n14141 & ~n24967 ;
  assign n24969 = n6905 & n24968 ;
  assign n24970 = n24969 ^ n9628 ^ n5884 ;
  assign n24963 = n16572 | n20256 ;
  assign n24964 = n3467 & n24963 ;
  assign n24971 = n24970 ^ n24964 ^ 1'b0 ;
  assign n24972 = n7332 & n24971 ;
  assign n24973 = ~n1921 & n4033 ;
  assign n24974 = n14717 & n24973 ;
  assign n24976 = ~n7771 & n8559 ;
  assign n24977 = n24976 ^ n17420 ^ 1'b0 ;
  assign n24975 = ~n13065 & n16122 ;
  assign n24978 = n24977 ^ n24975 ^ 1'b0 ;
  assign n24979 = n1544 | n4083 ;
  assign n24980 = n24979 ^ n14147 ^ 1'b0 ;
  assign n24981 = n11362 ^ n3388 ^ 1'b0 ;
  assign n24982 = n24981 ^ n1945 ^ 1'b0 ;
  assign n24983 = ~n22551 & n24982 ;
  assign n24984 = n8024 ^ n2170 ^ 1'b0 ;
  assign n24985 = n11881 & n24984 ;
  assign n24986 = n2900 & n20219 ;
  assign n24987 = n12652 & n24986 ;
  assign n24988 = n24987 ^ n1182 ^ 1'b0 ;
  assign n24989 = n24985 & ~n24988 ;
  assign n24990 = ( n11632 & n12850 ) | ( n11632 & ~n21647 ) | ( n12850 & ~n21647 ) ;
  assign n24991 = n24990 ^ n19639 ^ n3568 ;
  assign n24992 = n6788 & ~n9696 ;
  assign n24993 = n5948 | n24992 ;
  assign n24994 = n11029 ^ n10142 ^ 1'b0 ;
  assign n24995 = ~n1671 & n24994 ;
  assign n24996 = n3666 ^ n1186 ^ 1'b0 ;
  assign n24997 = n1059 | n2304 ;
  assign n24998 = n2584 & ~n24997 ;
  assign n24999 = n24996 | n24998 ;
  assign n25000 = ~n22669 & n24999 ;
  assign n25001 = n25000 ^ n22567 ^ n13370 ;
  assign n25002 = n15022 ^ n8820 ^ n7912 ;
  assign n25003 = n3646 & ~n25002 ;
  assign n25004 = n25003 ^ n10532 ^ 1'b0 ;
  assign n25005 = n9970 | n19699 ;
  assign n25006 = n2644 & ~n25005 ;
  assign n25007 = n1815 ^ n1307 ^ 1'b0 ;
  assign n25008 = n14573 | n25007 ;
  assign n25009 = ( n5241 & n6204 ) | ( n5241 & n11651 ) | ( n6204 & n11651 ) ;
  assign n25010 = ~n5143 & n25009 ;
  assign n25011 = ~n11030 & n14752 ;
  assign n25012 = n25011 ^ n9806 ^ 1'b0 ;
  assign n25013 = n9630 & ~n25012 ;
  assign n25014 = n8966 & n25013 ;
  assign n25015 = ( ~n2514 & n2584 ) | ( ~n2514 & n25014 ) | ( n2584 & n25014 ) ;
  assign n25016 = n22403 ^ n11053 ^ 1'b0 ;
  assign n25017 = n22551 | n25016 ;
  assign n25018 = n25017 ^ n22064 ^ 1'b0 ;
  assign n25019 = ( n25010 & n25015 ) | ( n25010 & n25018 ) | ( n25015 & n25018 ) ;
  assign n25020 = n12657 & ~n23418 ;
  assign n25021 = ~n13697 & n25020 ;
  assign n25022 = n1738 ^ x32 ^ 1'b0 ;
  assign n25023 = n3184 & n24891 ;
  assign n25024 = ~n7520 & n25023 ;
  assign n25025 = ~n16515 & n25024 ;
  assign n25026 = ~x100 & n25025 ;
  assign n25027 = n24715 ^ n7601 ^ 1'b0 ;
  assign n25028 = ~n5650 & n11411 ;
  assign n25029 = ~n12132 & n25028 ;
  assign n25030 = n7260 & n24532 ;
  assign n25031 = n25029 & n25030 ;
  assign n25032 = ~n4341 & n7363 ;
  assign n25033 = n25032 ^ n5876 ^ 1'b0 ;
  assign n25034 = n7143 ^ x2 ^ 1'b0 ;
  assign n25035 = ~n9028 & n16818 ;
  assign n25036 = n25035 ^ n8807 ^ 1'b0 ;
  assign n25037 = n9767 ^ n1367 ^ 1'b0 ;
  assign n25038 = ( n25034 & n25036 ) | ( n25034 & ~n25037 ) | ( n25036 & ~n25037 ) ;
  assign n25039 = ~n3819 & n10381 ;
  assign n25040 = n25039 ^ n15759 ^ 1'b0 ;
  assign n25041 = n25040 ^ n445 ^ 1'b0 ;
  assign n25042 = ~n2844 & n4603 ;
  assign n25043 = n25042 ^ n3088 ^ 1'b0 ;
  assign n25044 = n13628 | n17233 ;
  assign n25045 = n10803 | n14679 ;
  assign n25046 = n25045 ^ n25018 ^ 1'b0 ;
  assign n25047 = ~n6284 & n18288 ;
  assign n25048 = n25047 ^ n6838 ^ 1'b0 ;
  assign n25049 = n17811 & n25048 ;
  assign n25052 = ~n5683 & n18758 ;
  assign n25053 = ~n16218 & n25052 ;
  assign n25054 = n1010 | n25053 ;
  assign n25055 = n25054 ^ n7810 ^ 1'b0 ;
  assign n25056 = n22966 & ~n25055 ;
  assign n25057 = n25056 ^ n2559 ^ 1'b0 ;
  assign n25050 = n16934 ^ n270 ^ 1'b0 ;
  assign n25051 = n25050 ^ n7976 ^ n2154 ;
  assign n25058 = n25057 ^ n25051 ^ 1'b0 ;
  assign n25059 = n980 | n25058 ;
  assign n25060 = n8499 & n16430 ;
  assign n25061 = n25060 ^ n5425 ^ 1'b0 ;
  assign n25062 = n5038 & n23405 ;
  assign n25063 = n16296 ^ n6414 ^ 1'b0 ;
  assign n25064 = ~n4698 & n17732 ;
  assign n25065 = n22825 ^ n11859 ^ 1'b0 ;
  assign n25066 = n6146 & n25065 ;
  assign n25067 = ~n6908 & n17881 ;
  assign n25068 = ~n18541 & n25067 ;
  assign n25069 = n17078 ^ n2622 ^ 1'b0 ;
  assign n25070 = n13303 & n25069 ;
  assign n25074 = ~n5650 & n13317 ;
  assign n25075 = n25074 ^ n1523 ^ 1'b0 ;
  assign n25076 = n10877 | n25075 ;
  assign n25077 = n25076 ^ n12668 ^ 1'b0 ;
  assign n25071 = n8707 & ~n18569 ;
  assign n25072 = ~n18865 & n25071 ;
  assign n25073 = n6587 & ~n25072 ;
  assign n25078 = n25077 ^ n25073 ^ 1'b0 ;
  assign n25079 = n6925 & n25078 ;
  assign n25080 = ~n25070 & n25079 ;
  assign n25081 = n7899 & n24127 ;
  assign n25082 = ~n9027 & n25081 ;
  assign n25083 = n20571 ^ n10268 ^ 1'b0 ;
  assign n25084 = ~n19767 & n25083 ;
  assign n25085 = n3028 & n3465 ;
  assign n25086 = n25085 ^ n14821 ^ 1'b0 ;
  assign n25087 = x160 & ~n1183 ;
  assign n25088 = n25087 ^ n3137 ^ 1'b0 ;
  assign n25089 = n2301 & n25088 ;
  assign n25090 = ~n8713 & n25089 ;
  assign n25091 = n16250 & n25090 ;
  assign n25092 = n906 & n9199 ;
  assign n25093 = n10108 | n22894 ;
  assign n25094 = n15332 ^ x13 ^ 1'b0 ;
  assign n25095 = n25094 ^ n8136 ^ 1'b0 ;
  assign n25096 = n4178 & n25095 ;
  assign n25097 = n8723 & n12036 ;
  assign n25098 = n18150 & n25097 ;
  assign n25099 = n3159 | n9977 ;
  assign n25100 = n20699 & ~n25099 ;
  assign n25104 = n6707 & ~n18277 ;
  assign n25101 = n2366 & ~n4168 ;
  assign n25102 = n5084 & n25101 ;
  assign n25103 = n25102 ^ n6805 ^ 1'b0 ;
  assign n25105 = n25104 ^ n25103 ^ n15995 ;
  assign n25106 = ~n4714 & n4936 ;
  assign n25107 = n25106 ^ n7445 ^ 1'b0 ;
  assign n25108 = n25107 ^ n3577 ^ 1'b0 ;
  assign n25109 = n2317 & n25108 ;
  assign n25110 = n17736 & ~n25109 ;
  assign n25111 = ~n797 & n25110 ;
  assign n25112 = ~n19227 & n25111 ;
  assign n25113 = n9623 | n16882 ;
  assign n25114 = n3809 ^ n1589 ^ 1'b0 ;
  assign n25115 = n9465 ^ n3594 ^ 1'b0 ;
  assign n25116 = n25114 & ~n25115 ;
  assign n25117 = n12522 ^ n5800 ^ 1'b0 ;
  assign n25118 = n18070 & ~n25117 ;
  assign n25119 = n25118 ^ n22592 ^ n10884 ;
  assign n25120 = n15526 & ~n23087 ;
  assign n25121 = n25120 ^ n13673 ^ 1'b0 ;
  assign n25122 = n12638 ^ n11181 ^ n10676 ;
  assign n25123 = n2726 | n11668 ;
  assign n25124 = n25122 | n25123 ;
  assign n25125 = n14749 | n25124 ;
  assign n25126 = n25125 ^ n638 ^ 1'b0 ;
  assign n25127 = n17505 & ~n19686 ;
  assign n25128 = n25127 ^ n20093 ^ 1'b0 ;
  assign n25129 = n6022 & n7702 ;
  assign n25130 = ~n5966 & n25129 ;
  assign n25131 = n25130 ^ n10907 ^ 1'b0 ;
  assign n25132 = n10113 & n25131 ;
  assign n25133 = ~n1152 & n25132 ;
  assign n25134 = n25133 ^ n2243 ^ 1'b0 ;
  assign n25135 = ( ~n4968 & n8436 ) | ( ~n4968 & n10890 ) | ( n8436 & n10890 ) ;
  assign n25136 = n25134 | n25135 ;
  assign n25137 = n10333 & ~n16794 ;
  assign n25138 = n580 & ~n5236 ;
  assign n25139 = n2611 & n25138 ;
  assign n25140 = n492 | n25139 ;
  assign n25141 = n25140 ^ n25062 ^ 1'b0 ;
  assign n25142 = ~n25137 & n25141 ;
  assign n25143 = n11187 | n17352 ;
  assign n25144 = ~n4301 & n5798 ;
  assign n25145 = n10376 & n18420 ;
  assign n25146 = n25145 ^ n1844 ^ 1'b0 ;
  assign n25147 = ~n23366 & n25146 ;
  assign n25148 = n3886 & n24484 ;
  assign n25149 = ~n8007 & n25148 ;
  assign n25150 = n2542 & ~n8438 ;
  assign n25151 = ( n4551 & n19344 ) | ( n4551 & n25150 ) | ( n19344 & n25150 ) ;
  assign n25152 = n23012 & n25151 ;
  assign n25153 = n7934 ^ n2125 ^ 1'b0 ;
  assign n25154 = n15991 ^ n922 ^ 1'b0 ;
  assign n25155 = ~n3300 & n25154 ;
  assign n25156 = n25153 | n25155 ;
  assign n25157 = n12607 ^ n4309 ^ 1'b0 ;
  assign n25158 = n20910 ^ n7222 ^ 1'b0 ;
  assign n25159 = n1866 & n25158 ;
  assign n25160 = ( n2099 & n4406 ) | ( n2099 & n11061 ) | ( n4406 & n11061 ) ;
  assign n25161 = n13157 | n14398 ;
  assign n25162 = n25161 ^ n7115 ^ 1'b0 ;
  assign n25163 = n6079 ^ n4750 ^ 1'b0 ;
  assign n25164 = n21396 ^ n10575 ^ 1'b0 ;
  assign n25165 = n1586 ^ n1538 ^ 1'b0 ;
  assign n25166 = ~n2714 & n25165 ;
  assign n25167 = n4607 ^ n535 ^ 1'b0 ;
  assign n25168 = ~n9468 & n25167 ;
  assign n25169 = n7373 & ~n13394 ;
  assign n25170 = ~n25168 & n25169 ;
  assign n25171 = n8532 & ~n13734 ;
  assign n25172 = n876 & n25171 ;
  assign n25173 = ( n1682 & ~n6177 ) | ( n1682 & n16739 ) | ( ~n6177 & n16739 ) ;
  assign n25174 = n5387 & n25009 ;
  assign n25175 = n6327 & ~n25174 ;
  assign n25176 = n11301 & n13445 ;
  assign n25177 = ~n5786 & n25176 ;
  assign n25178 = n446 | n25177 ;
  assign n25179 = n25175 & n25178 ;
  assign n25180 = n1705 | n18365 ;
  assign n25181 = n25180 ^ n5373 ^ 1'b0 ;
  assign n25182 = n8456 & n24871 ;
  assign n25183 = n24290 ^ n2604 ^ 1'b0 ;
  assign n25184 = n25183 ^ n15278 ^ 1'b0 ;
  assign n25185 = n4712 & ~n25184 ;
  assign n25186 = n5838 ^ n4931 ^ 1'b0 ;
  assign n25187 = x252 & n25186 ;
  assign n25188 = n3105 & ~n15050 ;
  assign n25189 = n25188 ^ n4612 ^ 1'b0 ;
  assign n25190 = n25187 & ~n25189 ;
  assign n25191 = n3604 & n25190 ;
  assign n25192 = n9531 & n25191 ;
  assign n25193 = n22945 & ~n25192 ;
  assign n25194 = n6119 & ~n10805 ;
  assign n25195 = ~n3123 & n25194 ;
  assign n25196 = n14462 | n25195 ;
  assign n25197 = n7071 & n8754 ;
  assign n25198 = n25197 ^ n22991 ^ 1'b0 ;
  assign n25199 = ~n8778 & n16763 ;
  assign n25200 = n25199 ^ n8937 ^ 1'b0 ;
  assign n25201 = ~n11665 & n25200 ;
  assign n25202 = n16037 & n25201 ;
  assign n25203 = n3054 ^ n2400 ^ 1'b0 ;
  assign n25204 = n21471 | n25203 ;
  assign n25205 = x74 & ~n1591 ;
  assign n25206 = n18886 | n25205 ;
  assign n25207 = n2623 ^ n464 ^ 1'b0 ;
  assign n25208 = ~n3772 & n14311 ;
  assign n25209 = n2807 | n25208 ;
  assign n25210 = ( ~n2928 & n3757 ) | ( ~n2928 & n11796 ) | ( n3757 & n11796 ) ;
  assign n25211 = n12571 ^ n9612 ^ n8159 ;
  assign n25212 = n25211 ^ n11650 ^ 1'b0 ;
  assign n25213 = n4449 ^ n3335 ^ x13 ;
  assign n25214 = n14036 | n25213 ;
  assign n25215 = n10648 & n13662 ;
  assign n25216 = ~n9754 & n10055 ;
  assign n25217 = n25216 ^ n15609 ^ 1'b0 ;
  assign n25218 = n7145 ^ x228 ^ 1'b0 ;
  assign n25219 = n5896 | n25218 ;
  assign n25220 = n20609 | n25219 ;
  assign n25221 = n7050 & ~n17892 ;
  assign n25222 = n25221 ^ n20211 ^ 1'b0 ;
  assign n25223 = n20830 | n25222 ;
  assign n25224 = n659 ^ n613 ^ 1'b0 ;
  assign n25225 = n7996 & ~n25224 ;
  assign n25226 = n6146 & ~n20328 ;
  assign n25227 = n25226 ^ n2926 ^ 1'b0 ;
  assign n25228 = n25227 ^ n16039 ^ 1'b0 ;
  assign n25229 = n924 & n2322 ;
  assign n25230 = n23562 & n25229 ;
  assign n25231 = n5269 ^ n2867 ^ 1'b0 ;
  assign n25232 = n2294 & n4665 ;
  assign n25233 = n25231 | n25232 ;
  assign n25234 = n15718 | n25233 ;
  assign n25235 = n7702 | n25234 ;
  assign n25236 = n2041 & n25235 ;
  assign n25237 = x152 & ~n25236 ;
  assign n25238 = n22102 ^ n4165 ^ 1'b0 ;
  assign n25239 = ~n4721 & n14703 ;
  assign n25240 = n25239 ^ n3589 ^ 1'b0 ;
  assign n25241 = n25240 ^ n12473 ^ 1'b0 ;
  assign n25242 = n25241 ^ n18974 ^ 1'b0 ;
  assign n25243 = ~n11636 & n25242 ;
  assign n25244 = n5051 & ~n15003 ;
  assign n25245 = n17033 & n25244 ;
  assign n25246 = ( n17056 & n22537 ) | ( n17056 & ~n25245 ) | ( n22537 & ~n25245 ) ;
  assign n25247 = n15801 ^ n13083 ^ n9606 ;
  assign n25248 = n6434 | n15247 ;
  assign n25249 = n19589 | n25248 ;
  assign n25250 = n4027 ^ n825 ^ 1'b0 ;
  assign n25251 = n5504 & n10313 ;
  assign n25252 = ~n25250 & n25251 ;
  assign n25253 = n12095 ^ n8185 ^ n6746 ;
  assign n25254 = n10770 & ~n25253 ;
  assign n25255 = n3011 | n6609 ;
  assign n25256 = ~n8105 & n10288 ;
  assign n25257 = ( n22686 & n25255 ) | ( n22686 & n25256 ) | ( n25255 & n25256 ) ;
  assign n25258 = ~n12880 & n25257 ;
  assign n25259 = x180 | n266 ;
  assign n25260 = n9012 | n25259 ;
  assign n25261 = n5746 | n25260 ;
  assign n25262 = ( n9094 & ~n15162 ) | ( n9094 & n20799 ) | ( ~n15162 & n20799 ) ;
  assign n25263 = n15066 & n25262 ;
  assign n25264 = n9199 & ~n11769 ;
  assign n25265 = n4716 ^ x211 ^ 1'b0 ;
  assign n25266 = ~n14456 & n25265 ;
  assign n25267 = n1211 & n3174 ;
  assign n25268 = n4951 & ~n12887 ;
  assign n25269 = n25267 & n25268 ;
  assign n25270 = n17801 & ~n25269 ;
  assign n25271 = n4691 ^ n4069 ^ 1'b0 ;
  assign n25277 = n15518 ^ n7079 ^ 1'b0 ;
  assign n25272 = n15775 ^ n1922 ^ 1'b0 ;
  assign n25273 = ~n3092 & n25272 ;
  assign n25274 = n15311 & ~n25273 ;
  assign n25275 = ~n7418 & n25274 ;
  assign n25276 = n1909 & ~n25275 ;
  assign n25278 = n25277 ^ n25276 ^ 1'b0 ;
  assign n25279 = n4056 & ~n25278 ;
  assign n25280 = ~n2966 & n14096 ;
  assign n25281 = n25280 ^ n17674 ^ 1'b0 ;
  assign n25282 = n24892 & ~n25281 ;
  assign n25283 = n6339 & n6655 ;
  assign n25284 = ~n8452 & n14663 ;
  assign n25285 = ~n862 & n25284 ;
  assign n25286 = n2699 & n8490 ;
  assign n25287 = n7199 | n7719 ;
  assign n25288 = ~n16969 & n25287 ;
  assign n25289 = n3460 & n17609 ;
  assign n25290 = n19888 ^ n428 ^ 1'b0 ;
  assign n25291 = n25290 ^ n13920 ^ 1'b0 ;
  assign n25292 = n12725 | n25291 ;
  assign n25293 = n15826 | n25292 ;
  assign n25294 = n1671 & ~n25293 ;
  assign n25295 = n6187 & n16801 ;
  assign n25296 = ~n15760 & n25295 ;
  assign n25297 = n24484 ^ n13611 ^ 1'b0 ;
  assign n25298 = ~n25296 & n25297 ;
  assign n25299 = n25294 & n25298 ;
  assign n25300 = n2263 & ~n22095 ;
  assign n25301 = n25300 ^ n9076 ^ n2949 ;
  assign n25302 = n13102 & n18092 ;
  assign n25303 = n25302 ^ n10399 ^ 1'b0 ;
  assign n25304 = n8365 & n25303 ;
  assign n25305 = n24956 ^ n14965 ^ 1'b0 ;
  assign n25306 = n5537 | n12633 ;
  assign n25307 = n11585 | n25306 ;
  assign n25308 = n23473 ^ n10178 ^ 1'b0 ;
  assign n25309 = n847 & ~n5980 ;
  assign n25310 = n25309 ^ n8117 ^ 1'b0 ;
  assign n25311 = n1324 & n9601 ;
  assign n25312 = n25311 ^ n1309 ^ 1'b0 ;
  assign n25313 = n25312 ^ n10960 ^ 1'b0 ;
  assign n25314 = n25310 & ~n25313 ;
  assign n25315 = n25314 ^ n12794 ^ 1'b0 ;
  assign n25316 = ~n4379 & n10937 ;
  assign n25317 = n8301 & ~n17075 ;
  assign n25318 = n13088 | n25317 ;
  assign n25319 = n25318 ^ n18461 ^ 1'b0 ;
  assign n25320 = n25319 ^ n9867 ^ 1'b0 ;
  assign n25321 = n25316 & n25320 ;
  assign n25322 = n2691 & n9717 ;
  assign n25323 = n4639 & n25322 ;
  assign n25324 = n25323 ^ n11333 ^ 1'b0 ;
  assign n25325 = ~n23102 & n25324 ;
  assign n25326 = ( ~n3127 & n17462 ) | ( ~n3127 & n19792 ) | ( n17462 & n19792 ) ;
  assign n25327 = n3645 ^ n2895 ^ 1'b0 ;
  assign n25328 = ~n12356 & n25327 ;
  assign n25329 = n3873 & ~n25328 ;
  assign n25330 = n1630 | n5725 ;
  assign n25331 = n25330 ^ n11784 ^ 1'b0 ;
  assign n25332 = n4433 & n6540 ;
  assign n25333 = n25331 & n25332 ;
  assign n25334 = n12840 | n19536 ;
  assign n25335 = n11571 ^ n940 ^ 1'b0 ;
  assign n25336 = n2080 & ~n6895 ;
  assign n25337 = ~n22908 & n25336 ;
  assign n25345 = ~n7452 & n17021 ;
  assign n25346 = ~n9200 & n25345 ;
  assign n25341 = n6311 | n9903 ;
  assign n25342 = n12251 ^ n5016 ^ 1'b0 ;
  assign n25343 = ~n25341 & n25342 ;
  assign n25338 = n4086 ^ x250 ^ 1'b0 ;
  assign n25339 = n25338 ^ n13330 ^ n10451 ;
  assign n25340 = n17100 & n25339 ;
  assign n25344 = n25343 ^ n25340 ^ 1'b0 ;
  assign n25347 = n25346 ^ n25344 ^ 1'b0 ;
  assign n25348 = n16989 ^ n4145 ^ n944 ;
  assign n25349 = n14376 | n25348 ;
  assign n25351 = n572 & ~n8752 ;
  assign n25352 = n25351 ^ n3785 ^ 1'b0 ;
  assign n25350 = n10345 ^ n2885 ^ 1'b0 ;
  assign n25353 = n25352 ^ n25350 ^ n20851 ;
  assign n25354 = n19552 & n20212 ;
  assign n25355 = ~n15623 & n25354 ;
  assign n25356 = n2096 | n10537 ;
  assign n25357 = n25356 ^ n16805 ^ 1'b0 ;
  assign n25358 = ~n15743 & n25357 ;
  assign n25359 = n1114 & n25358 ;
  assign n25360 = n14306 ^ n11146 ^ n4426 ;
  assign n25361 = ( n3424 & n4031 ) | ( n3424 & ~n25360 ) | ( n4031 & ~n25360 ) ;
  assign n25362 = n4135 & ~n25361 ;
  assign n25363 = ~n17633 & n25362 ;
  assign n25364 = n17053 ^ n8155 ^ 1'b0 ;
  assign n25365 = n7329 & n25364 ;
  assign n25366 = ~n1914 & n17858 ;
  assign n25367 = n25366 ^ n5911 ^ 1'b0 ;
  assign n25368 = n25365 & n25367 ;
  assign n25370 = ~n1267 & n7941 ;
  assign n25371 = n25370 ^ n7746 ^ 1'b0 ;
  assign n25369 = n4633 & ~n8957 ;
  assign n25372 = n25371 ^ n25369 ^ 1'b0 ;
  assign n25373 = n25372 ^ x240 ^ 1'b0 ;
  assign n25374 = n8783 ^ n928 ^ 1'b0 ;
  assign n25375 = ~n2093 & n25374 ;
  assign n25376 = n5080 & n25375 ;
  assign n25377 = ~n4701 & n18708 ;
  assign n25378 = n20373 & n25377 ;
  assign n25379 = n923 & ~n7355 ;
  assign n25380 = n1354 ^ n1353 ^ 1'b0 ;
  assign n25381 = n23036 & n25380 ;
  assign n25382 = n22940 | n23404 ;
  assign n25383 = n23408 ^ n11551 ^ 1'b0 ;
  assign n25384 = ~n8085 & n11055 ;
  assign n25385 = n25384 ^ n11199 ^ 1'b0 ;
  assign n25386 = ( n8418 & n19075 ) | ( n8418 & n25385 ) | ( n19075 & n25385 ) ;
  assign n25387 = n10510 & n25386 ;
  assign n25388 = n14413 ^ n11155 ^ 1'b0 ;
  assign n25390 = n21475 & ~n22245 ;
  assign n25389 = n22334 ^ n12656 ^ 1'b0 ;
  assign n25391 = n25390 ^ n25389 ^ 1'b0 ;
  assign n25394 = n7738 ^ n3629 ^ 1'b0 ;
  assign n25392 = n13155 ^ n1936 ^ 1'b0 ;
  assign n25393 = n11747 | n25392 ;
  assign n25395 = n25394 ^ n25393 ^ 1'b0 ;
  assign n25396 = ~n1754 & n6088 ;
  assign n25397 = n10682 | n25396 ;
  assign n25398 = n15968 & ~n25397 ;
  assign n25399 = x175 & n935 ;
  assign n25400 = n25399 ^ n16238 ^ 1'b0 ;
  assign n25401 = n3281 & n25400 ;
  assign n25402 = n25401 ^ n16227 ^ 1'b0 ;
  assign n25403 = n3439 ^ n1680 ^ 1'b0 ;
  assign n25404 = ~n25402 & n25403 ;
  assign n25405 = n20748 ^ n3666 ^ x153 ;
  assign n25406 = n25405 ^ n4979 ^ 1'b0 ;
  assign n25407 = n19474 | n22307 ;
  assign n25408 = n25407 ^ n9083 ^ 1'b0 ;
  assign n25409 = n10556 ^ n8676 ^ 1'b0 ;
  assign n25410 = n756 & ~n12719 ;
  assign n25411 = ~n22365 & n25410 ;
  assign n25412 = n4845 & n25411 ;
  assign n25413 = n9076 & n11389 ;
  assign n25414 = n12445 | n25413 ;
  assign n25415 = ~n17962 & n24437 ;
  assign n25416 = n3850 & n11843 ;
  assign n25417 = ~n14840 & n25416 ;
  assign n25418 = n4184 | n23726 ;
  assign n25419 = n25418 ^ n24063 ^ 1'b0 ;
  assign n25420 = ~n2633 & n4733 ;
  assign n25421 = n17247 ^ n6483 ^ 1'b0 ;
  assign n25422 = n25420 & ~n25421 ;
  assign n25423 = n25422 ^ n5608 ^ 1'b0 ;
  assign n25424 = n7722 & n25423 ;
  assign n25425 = n17259 ^ n8287 ^ 1'b0 ;
  assign n25426 = ~n11129 & n23924 ;
  assign n25427 = ( ~n335 & n25425 ) | ( ~n335 & n25426 ) | ( n25425 & n25426 ) ;
  assign n25428 = n5746 & n25427 ;
  assign n25429 = x35 & ~n9185 ;
  assign n25430 = n10150 & n25429 ;
  assign n25431 = ~n25429 & n25430 ;
  assign n25432 = n5061 & n25431 ;
  assign n25435 = x62 & n1132 ;
  assign n25436 = ~x62 & n25435 ;
  assign n25433 = n17285 & n23751 ;
  assign n25434 = ~n23751 & n25433 ;
  assign n25437 = n25436 ^ n25434 ^ 1'b0 ;
  assign n25438 = ~n25432 & n25437 ;
  assign n25439 = n509 & ~n1731 ;
  assign n25440 = n25439 ^ n8488 ^ 1'b0 ;
  assign n25441 = n14620 & ~n25440 ;
  assign n25442 = n25441 ^ n15904 ^ 1'b0 ;
  assign n25443 = n25442 ^ n24038 ^ 1'b0 ;
  assign n25444 = ~n4871 & n6963 ;
  assign n25445 = ~n1660 & n25444 ;
  assign n25446 = n25445 ^ n1530 ^ 1'b0 ;
  assign n25447 = n4014 & n9299 ;
  assign n25448 = n25447 ^ n4493 ^ 1'b0 ;
  assign n25449 = n25448 ^ n1882 ^ 1'b0 ;
  assign n25450 = n19427 ^ n5812 ^ 1'b0 ;
  assign n25451 = ~n18653 & n25450 ;
  assign n25453 = ~n1023 & n4014 ;
  assign n25454 = n475 & n25453 ;
  assign n25455 = n22884 | n25454 ;
  assign n25456 = n21747 | n25455 ;
  assign n25452 = ~n11764 & n18791 ;
  assign n25457 = n25456 ^ n25452 ^ 1'b0 ;
  assign n25458 = n3828 | n22699 ;
  assign n25459 = n11775 | n25458 ;
  assign n25460 = n25459 ^ n20453 ^ n18391 ;
  assign n25461 = n7179 ^ n2372 ^ 1'b0 ;
  assign n25462 = n12083 ^ n8217 ^ 1'b0 ;
  assign n25463 = n10781 & ~n25462 ;
  assign n25464 = n6177 & ~n9085 ;
  assign n25465 = n17187 ^ n6621 ^ 1'b0 ;
  assign n25466 = ~n24470 & n25465 ;
  assign n25469 = n10264 & n19399 ;
  assign n25470 = n25469 ^ n5318 ^ 1'b0 ;
  assign n25467 = n14729 ^ n8050 ^ 1'b0 ;
  assign n25468 = n25467 ^ n17541 ^ n4602 ;
  assign n25471 = n25470 ^ n25468 ^ 1'b0 ;
  assign n25474 = n671 & ~n6881 ;
  assign n25475 = n12280 | n25474 ;
  assign n25476 = n3915 | n25475 ;
  assign n25472 = ( n15303 & ~n18207 ) | ( n15303 & n23346 ) | ( ~n18207 & n23346 ) ;
  assign n25473 = n10211 | n25472 ;
  assign n25477 = n25476 ^ n25473 ^ 1'b0 ;
  assign n25478 = n16990 & n20384 ;
  assign n25479 = ~n6114 & n25478 ;
  assign n25480 = n7586 | n20818 ;
  assign n25481 = ~n9719 & n9727 ;
  assign n25482 = ~n4193 & n8182 ;
  assign n25483 = ~n25481 & n25482 ;
  assign n25484 = n11702 | n25483 ;
  assign n25485 = n24331 ^ n23659 ^ 1'b0 ;
  assign n25486 = n18146 ^ n4330 ^ 1'b0 ;
  assign n25487 = n19409 & n25486 ;
  assign n25488 = n25487 ^ n23608 ^ 1'b0 ;
  assign n25489 = n8235 ^ n4802 ^ n2927 ;
  assign n25495 = ~n4069 & n11834 ;
  assign n25490 = n17801 ^ n7608 ^ 1'b0 ;
  assign n25491 = n1639 ^ x242 ^ 1'b0 ;
  assign n25492 = n6311 | n25491 ;
  assign n25493 = n25490 & ~n25492 ;
  assign n25494 = ~n14117 & n25493 ;
  assign n25496 = n25495 ^ n25494 ^ n11255 ;
  assign n25497 = n20489 ^ n4845 ^ n1513 ;
  assign n25498 = n25497 ^ n2821 ^ 1'b0 ;
  assign n25499 = ~n486 & n19894 ;
  assign n25500 = n17394 & ~n25499 ;
  assign n25501 = ~n5104 & n25500 ;
  assign n25502 = n11913 ^ n6099 ^ 1'b0 ;
  assign n25503 = n25502 ^ n14145 ^ n2378 ;
  assign n25504 = n21333 ^ n4011 ^ 1'b0 ;
  assign n25505 = n4840 & ~n25504 ;
  assign n25506 = n4972 & ~n11360 ;
  assign n25507 = ~n7672 & n12409 ;
  assign n25508 = ~n8592 & n25507 ;
  assign n25509 = n9207 ^ n983 ^ 1'b0 ;
  assign n25510 = n25509 ^ n12491 ^ n9560 ;
  assign n25511 = n25510 ^ n18057 ^ 1'b0 ;
  assign n25512 = n1635 & ~n15056 ;
  assign n25513 = n14929 & ~n25512 ;
  assign n25514 = ~n25511 & n25513 ;
  assign n25516 = n15665 ^ n6739 ^ 1'b0 ;
  assign n25517 = n11342 & ~n25516 ;
  assign n25515 = n15495 ^ n2167 ^ 1'b0 ;
  assign n25518 = n25517 ^ n25515 ^ 1'b0 ;
  assign n25519 = n2708 & n11897 ;
  assign n25520 = n25519 ^ n7508 ^ 1'b0 ;
  assign n25521 = n25520 ^ n22548 ^ 1'b0 ;
  assign n25522 = n9801 & ~n25521 ;
  assign n25523 = n10024 ^ n1393 ^ 1'b0 ;
  assign n25524 = ~n1871 & n25523 ;
  assign n25525 = n13498 ^ n3090 ^ 1'b0 ;
  assign n25526 = n25524 & n25525 ;
  assign n25527 = n25526 ^ n14424 ^ 1'b0 ;
  assign n25528 = n2458 ^ x230 ^ 1'b0 ;
  assign n25529 = n25527 | n25528 ;
  assign n25530 = n21429 ^ n8349 ^ 1'b0 ;
  assign n25531 = n25530 ^ n15793 ^ 1'b0 ;
  assign n25532 = x126 & n25531 ;
  assign n25534 = n6398 & ~n25130 ;
  assign n25535 = ~n14823 & n25534 ;
  assign n25536 = n8868 & n13887 ;
  assign n25537 = n25535 & n25536 ;
  assign n25533 = n13671 | n23259 ;
  assign n25538 = n25537 ^ n25533 ^ 1'b0 ;
  assign n25539 = n23169 ^ n4445 ^ n2053 ;
  assign n25540 = ~n7613 & n25539 ;
  assign n25541 = n25538 & n25540 ;
  assign n25542 = n8713 ^ n5606 ^ 1'b0 ;
  assign n25543 = n25542 ^ n10674 ^ n6203 ;
  assign n25544 = ( x99 & n932 ) | ( x99 & ~n11450 ) | ( n932 & ~n11450 ) ;
  assign n25545 = n25544 ^ n7058 ^ n4402 ;
  assign n25546 = n25545 ^ n8237 ^ 1'b0 ;
  assign n25547 = n25546 ^ n17054 ^ 1'b0 ;
  assign n25548 = n2317 & ~n23289 ;
  assign n25549 = n25548 ^ n6453 ^ 1'b0 ;
  assign n25550 = n984 & ~n8046 ;
  assign n25551 = n25550 ^ n12132 ^ 1'b0 ;
  assign n25552 = n2403 | n11357 ;
  assign n25553 = n25551 & ~n25552 ;
  assign n25554 = n8791 & ~n11747 ;
  assign n25555 = n24799 | n25554 ;
  assign n25556 = n16730 & ~n25555 ;
  assign n25557 = n1866 & n3506 ;
  assign n25558 = n25557 ^ n13267 ^ 1'b0 ;
  assign n25559 = ~n23259 & n24256 ;
  assign n25560 = n12749 ^ n9775 ^ 1'b0 ;
  assign n25561 = ~n19536 & n25560 ;
  assign n25562 = n25561 ^ n12161 ^ 1'b0 ;
  assign n25563 = n2509 & ~n25562 ;
  assign n25564 = n7141 & ~n13098 ;
  assign n25565 = ~n12878 & n25564 ;
  assign n25568 = x78 & ~n21854 ;
  assign n25569 = n1048 & n25568 ;
  assign n25566 = n24293 ^ n3036 ^ 1'b0 ;
  assign n25567 = n10721 & n25566 ;
  assign n25570 = n25569 ^ n25567 ^ 1'b0 ;
  assign n25571 = ~n25565 & n25570 ;
  assign n25572 = ~n25563 & n25571 ;
  assign n25573 = n13509 & n14428 ;
  assign n25574 = n25573 ^ n5294 ^ 1'b0 ;
  assign n25575 = ( n4210 & n6646 ) | ( n4210 & n16753 ) | ( n6646 & n16753 ) ;
  assign n25576 = n10973 ^ n3160 ^ 1'b0 ;
  assign n25577 = ~n25575 & n25576 ;
  assign n25578 = ~n5749 & n25577 ;
  assign n25579 = ~n17134 & n25578 ;
  assign n25580 = ( n10299 & ~n25174 ) | ( n10299 & n25579 ) | ( ~n25174 & n25579 ) ;
  assign n25581 = n25580 ^ n19192 ^ 1'b0 ;
  assign n25582 = n3424 | n4803 ;
  assign n25583 = n445 | n25582 ;
  assign n25584 = n372 | n25583 ;
  assign n25585 = x180 | n6585 ;
  assign n25586 = n25257 & ~n25585 ;
  assign n25587 = n25586 ^ n13762 ^ 1'b0 ;
  assign n25588 = x241 | n13586 ;
  assign n25589 = n25588 ^ n1689 ^ 1'b0 ;
  assign n25590 = n21227 & ~n21965 ;
  assign n25592 = n9634 ^ n1497 ^ 1'b0 ;
  assign n25593 = n2890 | n25592 ;
  assign n25591 = n5984 & ~n6333 ;
  assign n25594 = n25593 ^ n25591 ^ 1'b0 ;
  assign n25595 = n3342 & ~n25594 ;
  assign n25600 = n13803 ^ n7668 ^ 1'b0 ;
  assign n25596 = ~n3297 & n17398 ;
  assign n25597 = n19269 ^ n2247 ^ 1'b0 ;
  assign n25598 = n25596 & n25597 ;
  assign n25599 = n19393 & n25598 ;
  assign n25601 = n25600 ^ n25599 ^ 1'b0 ;
  assign n25602 = n15387 ^ n6881 ^ 1'b0 ;
  assign n25603 = n18707 ^ n14695 ^ 1'b0 ;
  assign n25604 = n14727 & ~n25603 ;
  assign n25605 = n10713 | n25604 ;
  assign n25606 = n25605 ^ n5129 ^ 1'b0 ;
  assign n25607 = n2188 | n14578 ;
  assign n25608 = n25607 ^ n5949 ^ 1'b0 ;
  assign n25609 = n13003 & ~n25608 ;
  assign n25610 = n5704 & ~n14845 ;
  assign n25611 = n25610 ^ n9347 ^ 1'b0 ;
  assign n25612 = n21441 ^ n2332 ^ n2092 ;
  assign n25613 = n914 & n25612 ;
  assign n25614 = n25613 ^ n7819 ^ 1'b0 ;
  assign n25615 = n6825 ^ n4766 ^ 1'b0 ;
  assign n25616 = n19489 | n25615 ;
  assign n25617 = n11903 | n13953 ;
  assign n25618 = n13049 & ~n25617 ;
  assign n25619 = ( ~n1869 & n2192 ) | ( ~n1869 & n25618 ) | ( n2192 & n25618 ) ;
  assign n25620 = n25616 & ~n25619 ;
  assign n25621 = n25620 ^ n1521 ^ 1'b0 ;
  assign n25622 = n6286 & ~n11201 ;
  assign n25623 = n11260 & ~n25622 ;
  assign n25624 = n25623 ^ n4496 ^ 1'b0 ;
  assign n25625 = ~n13293 & n21344 ;
  assign n25626 = n1342 | n4269 ;
  assign n25627 = n25626 ^ n1398 ^ 1'b0 ;
  assign n25628 = x218 & ~n13562 ;
  assign n25629 = ( ~n11353 & n21429 ) | ( ~n11353 & n21606 ) | ( n21429 & n21606 ) ;
  assign n25630 = n2082 ^ n1132 ^ 1'b0 ;
  assign n25631 = n25630 ^ n5353 ^ 1'b0 ;
  assign n25632 = ~n8100 & n25631 ;
  assign n25633 = n11578 & ~n15037 ;
  assign n25634 = ~n3686 & n25633 ;
  assign n25635 = n5206 & n25634 ;
  assign n25636 = n8917 & n24484 ;
  assign n25637 = n25636 ^ n16114 ^ 1'b0 ;
  assign n25638 = n9905 & ~n25637 ;
  assign n25639 = ~n25635 & n25638 ;
  assign n25640 = ~n25632 & n25639 ;
  assign n25641 = n522 & n6998 ;
  assign n25642 = n13857 ^ n7454 ^ n1475 ;
  assign n25645 = ~n2798 & n3782 ;
  assign n25643 = n2606 & n2757 ;
  assign n25644 = ~n20480 & n25643 ;
  assign n25646 = n25645 ^ n25644 ^ n23955 ;
  assign n25652 = n13399 ^ n2646 ^ 1'b0 ;
  assign n25647 = n3535 | n5089 ;
  assign n25648 = n25647 ^ n13602 ^ 1'b0 ;
  assign n25649 = n24041 & ~n25648 ;
  assign n25650 = n22990 ^ n15260 ^ n9852 ;
  assign n25651 = n25649 & ~n25650 ;
  assign n25653 = n25652 ^ n25651 ^ 1'b0 ;
  assign n25654 = n23724 ^ n22800 ^ 1'b0 ;
  assign n25655 = n25653 | n25654 ;
  assign n25656 = n1470 & ~n5284 ;
  assign n25657 = n25656 ^ n4432 ^ 1'b0 ;
  assign n25658 = n19795 ^ n708 ^ 1'b0 ;
  assign n25659 = n2743 | n25658 ;
  assign n25660 = n16579 ^ n5767 ^ 1'b0 ;
  assign n25661 = n25659 & n25660 ;
  assign n25662 = n25657 & n25661 ;
  assign n25663 = n7419 & ~n8028 ;
  assign n25664 = ~n3385 & n15690 ;
  assign n25665 = ~n21218 & n25664 ;
  assign n25666 = n361 | n17546 ;
  assign n25667 = n15824 | n25666 ;
  assign n25668 = n5515 | n17398 ;
  assign n25669 = n18447 & n25668 ;
  assign n25670 = n6786 ^ n2334 ^ 1'b0 ;
  assign n25671 = n17127 & n25670 ;
  assign n25672 = n25671 ^ n8421 ^ 1'b0 ;
  assign n25673 = n1856 & n25672 ;
  assign n25674 = n10770 & ~n25673 ;
  assign n25675 = n4046 & n9936 ;
  assign n25676 = n25675 ^ n12373 ^ 1'b0 ;
  assign n25677 = n25676 ^ n632 ^ 1'b0 ;
  assign n25678 = n25677 ^ n11617 ^ 1'b0 ;
  assign n25679 = n492 & n25678 ;
  assign n25680 = ~n3432 & n4293 ;
  assign n25683 = n7641 & ~n9510 ;
  assign n25684 = n25683 ^ n4489 ^ 1'b0 ;
  assign n25681 = n2798 ^ x231 ^ 1'b0 ;
  assign n25682 = ~n1365 & n25681 ;
  assign n25685 = n25684 ^ n25682 ^ n1585 ;
  assign n25686 = n25685 ^ n23697 ^ n5621 ;
  assign n25687 = n14846 ^ n14250 ^ 1'b0 ;
  assign n25688 = ~n12519 & n13051 ;
  assign n25689 = n12355 & ~n25122 ;
  assign n25690 = ~n25688 & n25689 ;
  assign n25691 = n9881 | n19788 ;
  assign n25692 = n12936 & ~n25691 ;
  assign n25693 = n25692 ^ n7117 ^ 1'b0 ;
  assign n25694 = n20856 | n25693 ;
  assign n25695 = n6612 ^ n5820 ^ 1'b0 ;
  assign n25696 = ~n5835 & n25695 ;
  assign n25697 = n25696 ^ n3313 ^ 1'b0 ;
  assign n25698 = n15607 ^ n14009 ^ n13003 ;
  assign n25699 = n22905 ^ x24 ^ 1'b0 ;
  assign n25700 = ( n16764 & n19185 ) | ( n16764 & ~n25699 ) | ( n19185 & ~n25699 ) ;
  assign n25701 = n2399 | n25700 ;
  assign n25702 = n2244 & ~n5679 ;
  assign n25703 = n25702 ^ n825 ^ 1'b0 ;
  assign n25704 = ~n1146 & n25703 ;
  assign n25705 = n6310 & ~n23461 ;
  assign n25706 = ~n10249 & n25705 ;
  assign n25707 = n22934 ^ n17728 ^ 1'b0 ;
  assign n25708 = x92 & ~n25707 ;
  assign n25709 = n22520 ^ n16750 ^ 1'b0 ;
  assign n25710 = n25708 & n25709 ;
  assign n25711 = x164 & ~n10111 ;
  assign n25712 = ~n25710 & n25711 ;
  assign n25713 = ~n9914 & n19017 ;
  assign n25714 = n24215 & n25713 ;
  assign n25715 = n25714 ^ n16237 ^ 1'b0 ;
  assign n25716 = n25715 ^ n13402 ^ 1'b0 ;
  assign n25717 = n19218 | n25716 ;
  assign n25718 = n8508 ^ n4497 ^ n1344 ;
  assign n25719 = n6607 | n25718 ;
  assign n25720 = n14998 & ~n25719 ;
  assign n25721 = n25720 ^ n12704 ^ 1'b0 ;
  assign n25722 = ( ~x219 & n9905 ) | ( ~x219 & n25721 ) | ( n9905 & n25721 ) ;
  assign n25724 = n2703 & n7179 ;
  assign n25725 = n25724 ^ n14582 ^ 1'b0 ;
  assign n25723 = n6844 & ~n14716 ;
  assign n25726 = n25725 ^ n25723 ^ 1'b0 ;
  assign n25727 = n21757 & ~n25610 ;
  assign n25729 = n15995 ^ n1055 ^ 1'b0 ;
  assign n25728 = ~n287 & n15857 ;
  assign n25730 = n25729 ^ n25728 ^ 1'b0 ;
  assign n25731 = n4271 & ~n17711 ;
  assign n25732 = n25731 ^ n18059 ^ 1'b0 ;
  assign n25733 = ~n6748 & n25732 ;
  assign n25734 = ~n7150 & n25733 ;
  assign n25735 = n8079 & n25734 ;
  assign n25736 = n4859 & ~n17710 ;
  assign n25737 = n25736 ^ n24611 ^ 1'b0 ;
  assign n25738 = n10928 & n15156 ;
  assign n25739 = n16598 & n25738 ;
  assign n25740 = n4657 | n25739 ;
  assign n25741 = n3320 | n25740 ;
  assign n25742 = n10941 | n15718 ;
  assign n25743 = n4132 ^ n3959 ^ n1034 ;
  assign n25744 = n15638 ^ n10498 ^ 1'b0 ;
  assign n25745 = n25744 ^ n11737 ^ 1'b0 ;
  assign n25746 = n3890 & ~n23802 ;
  assign n25749 = n1639 & ~n8758 ;
  assign n25747 = n993 & ~n15752 ;
  assign n25748 = n5936 | n25747 ;
  assign n25750 = n25749 ^ n25748 ^ 1'b0 ;
  assign n25751 = ~n1680 & n10732 ;
  assign n25752 = n25751 ^ n9930 ^ 1'b0 ;
  assign n25753 = ( ~n8444 & n25750 ) | ( ~n8444 & n25752 ) | ( n25750 & n25752 ) ;
  assign n25754 = n25753 ^ n7945 ^ 1'b0 ;
  assign n25755 = n24763 | n25754 ;
  assign n25756 = n13093 | n25755 ;
  assign n25757 = n25746 & ~n25756 ;
  assign n25758 = n12235 & ~n12476 ;
  assign n25759 = n5513 ^ n3860 ^ 1'b0 ;
  assign n25760 = n869 & n16863 ;
  assign n25761 = n22085 ^ n14417 ^ 1'b0 ;
  assign n25762 = n25760 & n25761 ;
  assign n25763 = n5517 ^ n518 ^ 1'b0 ;
  assign n25764 = ~n12578 & n19988 ;
  assign n25765 = n19069 ^ n9180 ^ 1'b0 ;
  assign n25766 = n7134 | n25765 ;
  assign n25767 = n19684 ^ n9377 ^ 1'b0 ;
  assign n25768 = ~n3888 & n5788 ;
  assign n25769 = ( n5195 & n9270 ) | ( n5195 & n13562 ) | ( n9270 & n13562 ) ;
  assign n25770 = n3496 & n8666 ;
  assign n25771 = ~n25769 & n25770 ;
  assign n25772 = n25771 ^ n15161 ^ 1'b0 ;
  assign n25773 = n25768 & ~n25772 ;
  assign n25774 = n2263 | n21990 ;
  assign n25775 = n25774 ^ n3357 ^ 1'b0 ;
  assign n25776 = n3007 & n7051 ;
  assign n25777 = n5497 | n22035 ;
  assign n25778 = n25776 | n25777 ;
  assign n25779 = n17936 ^ n6387 ^ 1'b0 ;
  assign n25780 = n17302 & n25779 ;
  assign n25781 = n5937 ^ n5246 ^ 1'b0 ;
  assign n25782 = n8831 ^ n2837 ^ 1'b0 ;
  assign n25783 = ~n7219 & n11765 ;
  assign n25784 = n4905 ^ n2646 ^ 1'b0 ;
  assign n25785 = n21305 ^ n15069 ^ 1'b0 ;
  assign n25786 = n2872 & n7041 ;
  assign n25787 = n25786 ^ n11649 ^ 1'b0 ;
  assign n25788 = n25787 ^ n3049 ^ 1'b0 ;
  assign n25789 = n14059 ^ n6118 ^ 1'b0 ;
  assign n25790 = n25789 ^ n13521 ^ 1'b0 ;
  assign n25791 = n11035 ^ n8842 ^ 1'b0 ;
  assign n25792 = n25791 ^ n21485 ^ 1'b0 ;
  assign n25793 = n4631 & ~n25792 ;
  assign n25794 = n19681 ^ n19480 ^ 1'b0 ;
  assign n25795 = n11561 & ~n25794 ;
  assign n25796 = n25795 ^ n17041 ^ 1'b0 ;
  assign n25797 = n18732 | n25796 ;
  assign n25798 = n11902 & n17898 ;
  assign n25799 = n2301 & ~n5160 ;
  assign n25800 = n6070 & n25799 ;
  assign n25801 = n11992 ^ n5664 ^ 1'b0 ;
  assign n25802 = n5021 & ~n25801 ;
  assign n25803 = n1369 | n23610 ;
  assign n25804 = n25802 | n25803 ;
  assign n25805 = x206 & n7204 ;
  assign n25806 = n2055 & ~n7419 ;
  assign n25807 = ~n2462 & n25806 ;
  assign n25808 = n3429 & ~n17949 ;
  assign n25809 = n20418 & n25808 ;
  assign n25810 = n4745 & n17226 ;
  assign n25811 = n25810 ^ n16213 ^ 1'b0 ;
  assign n25812 = n6789 & n25811 ;
  assign n25813 = ~n25809 & n25812 ;
  assign n25814 = n448 & n25813 ;
  assign n25815 = n3508 & n17588 ;
  assign n25816 = n1589 & ~n17778 ;
  assign n25817 = ~n12448 & n12737 ;
  assign n25818 = n25817 ^ n10490 ^ 1'b0 ;
  assign n25819 = n20108 ^ n12163 ^ 1'b0 ;
  assign n25820 = n8499 ^ n2500 ^ 1'b0 ;
  assign n25821 = n25819 & ~n25820 ;
  assign n25822 = n16340 ^ n11280 ^ 1'b0 ;
  assign n25823 = n1635 | n25822 ;
  assign n25824 = n11825 & ~n14723 ;
  assign n25825 = n1671 & ~n3284 ;
  assign n25829 = ( x63 & n1632 ) | ( x63 & ~n3744 ) | ( n1632 & ~n3744 ) ;
  assign n25826 = n535 & ~n1367 ;
  assign n25827 = n25826 ^ n6618 ^ 1'b0 ;
  assign n25828 = ~n22739 & n25827 ;
  assign n25830 = n25829 ^ n25828 ^ 1'b0 ;
  assign n25831 = ~n613 & n3146 ;
  assign n25832 = n10670 & n25831 ;
  assign n25833 = ~n10111 & n25832 ;
  assign n25836 = x246 & ~n725 ;
  assign n25837 = ~x246 & n25836 ;
  assign n25838 = n25837 ^ n1311 ^ 1'b0 ;
  assign n25839 = n574 | n1664 ;
  assign n25840 = n574 & ~n25839 ;
  assign n25841 = n2050 & n25840 ;
  assign n25842 = n25838 & ~n25841 ;
  assign n25843 = ~n25838 & n25842 ;
  assign n25844 = ~n15204 & n25843 ;
  assign n25834 = ~n5925 & n11216 ;
  assign n25835 = n8391 & ~n25834 ;
  assign n25845 = n25844 ^ n25835 ^ 1'b0 ;
  assign n25846 = n25845 ^ n18387 ^ 1'b0 ;
  assign n25847 = n5413 & ~n13779 ;
  assign n25848 = n13368 & n25847 ;
  assign n25849 = ~n25847 & n25848 ;
  assign n25850 = n7496 & ~n25849 ;
  assign n25851 = n25846 & n25850 ;
  assign n25852 = n2114 | n6116 ;
  assign n25856 = n2590 & ~n16915 ;
  assign n25857 = n25856 ^ n5193 ^ 1'b0 ;
  assign n25853 = ~n7952 & n19464 ;
  assign n25854 = ~n2879 & n25853 ;
  assign n25855 = n11852 & ~n25854 ;
  assign n25858 = n25857 ^ n25855 ^ 1'b0 ;
  assign n25859 = n12165 ^ n5582 ^ 1'b0 ;
  assign n25860 = n18146 & ~n25859 ;
  assign n25861 = ~n17616 & n25860 ;
  assign n25862 = n774 | n9316 ;
  assign n25863 = n25862 ^ n15079 ^ 1'b0 ;
  assign n25864 = n21573 ^ n7197 ^ 1'b0 ;
  assign n25865 = n25863 | n25864 ;
  assign n25866 = n8555 ^ x218 ^ 1'b0 ;
  assign n25867 = n13892 ^ n3942 ^ 1'b0 ;
  assign n25868 = n25866 & n25867 ;
  assign n25869 = n10066 & ~n13666 ;
  assign n25870 = ( n3159 & ~n8819 ) | ( n3159 & n25869 ) | ( ~n8819 & n25869 ) ;
  assign n25871 = x204 & n7581 ;
  assign n25872 = ~n15880 & n25871 ;
  assign n25873 = n713 & ~n4003 ;
  assign n25874 = n25873 ^ n24428 ^ 1'b0 ;
  assign n25878 = n5711 ^ n271 ^ 1'b0 ;
  assign n25879 = ~n7022 & n25878 ;
  assign n25876 = n11094 & ~n13576 ;
  assign n25877 = ~n13927 & n25876 ;
  assign n25880 = n25879 ^ n25877 ^ n24705 ;
  assign n25875 = n16863 & ~n19998 ;
  assign n25881 = n25880 ^ n25875 ^ 1'b0 ;
  assign n25882 = ~n11270 & n18314 ;
  assign n25883 = ~n4594 & n25882 ;
  assign n25884 = n10142 | n14209 ;
  assign n25885 = n17806 ^ n16374 ^ 1'b0 ;
  assign n25886 = n13861 ^ n13018 ^ 1'b0 ;
  assign n25887 = ~n25885 & n25886 ;
  assign n25888 = n3717 & n11702 ;
  assign n25889 = n19470 ^ n5392 ^ 1'b0 ;
  assign n25890 = n25889 ^ n13912 ^ n886 ;
  assign n25891 = n15015 ^ n6600 ^ 1'b0 ;
  assign n25892 = n23527 ^ n11703 ^ 1'b0 ;
  assign n25896 = n5349 ^ x38 ^ 1'b0 ;
  assign n25897 = ~n4880 & n25896 ;
  assign n25893 = n3460 | n10973 ;
  assign n25894 = n25893 ^ n13382 ^ 1'b0 ;
  assign n25895 = n15137 | n25894 ;
  assign n25898 = n25897 ^ n25895 ^ n24923 ;
  assign n25899 = ~n6219 & n8975 ;
  assign n25900 = n25899 ^ n10182 ^ 1'b0 ;
  assign n25901 = n9113 & n25900 ;
  assign n25902 = n12068 & n25901 ;
  assign n25903 = n16037 & n25902 ;
  assign n25904 = n483 | n1254 ;
  assign n25905 = n9013 ^ n2317 ^ 1'b0 ;
  assign n25906 = ~n2029 & n25905 ;
  assign n25907 = n25906 ^ n17421 ^ 1'b0 ;
  assign n25908 = n6284 & ~n7204 ;
  assign n25909 = n24987 | n25908 ;
  assign n25910 = n8771 | n25909 ;
  assign n25911 = n25910 ^ n20202 ^ 1'b0 ;
  assign n25912 = n17283 & ~n25911 ;
  assign n25913 = n3704 & n17753 ;
  assign n25914 = n25913 ^ n9889 ^ 1'b0 ;
  assign n25915 = n11551 | n25914 ;
  assign n25916 = n4762 | n7619 ;
  assign n25917 = n25916 ^ n17340 ^ n1557 ;
  assign n25918 = n2736 & n22581 ;
  assign n25919 = n2109 & n25918 ;
  assign n25920 = ~n814 & n4025 ;
  assign n25921 = n25920 ^ n15699 ^ 1'b0 ;
  assign n25922 = n25241 & n25921 ;
  assign n25923 = n25922 ^ n17524 ^ 1'b0 ;
  assign n25924 = n3382 | n12605 ;
  assign n25925 = n1415 & ~n4430 ;
  assign n25926 = ~n8847 & n25925 ;
  assign n25927 = n25170 ^ n8042 ^ 1'b0 ;
  assign n25928 = n12876 ^ n12164 ^ n6525 ;
  assign n25929 = n25927 & n25928 ;
  assign n25930 = n5210 | n25055 ;
  assign n25931 = n9085 & ~n17588 ;
  assign n25932 = n5272 & ~n17548 ;
  assign n25933 = n25932 ^ n21515 ^ 1'b0 ;
  assign n25934 = n20205 ^ n7875 ^ n6075 ;
  assign n25935 = n25934 ^ n19235 ^ 1'b0 ;
  assign n25936 = n15481 | n25935 ;
  assign n25937 = n1598 ^ n1238 ^ x2 ;
  assign n25938 = n7328 ^ n3795 ^ 1'b0 ;
  assign n25939 = n10445 & n20505 ;
  assign n25940 = ~n8354 & n25939 ;
  assign n25941 = ( ~n25937 & n25938 ) | ( ~n25937 & n25940 ) | ( n25938 & n25940 ) ;
  assign n25942 = x213 & n1245 ;
  assign n25943 = n25942 ^ n18100 ^ 1'b0 ;
  assign n25944 = n25943 ^ n3104 ^ 1'b0 ;
  assign n25945 = n11570 ^ n9256 ^ n7148 ;
  assign n25946 = n25945 ^ n1694 ^ 1'b0 ;
  assign n25947 = ~n13121 & n15570 ;
  assign n25948 = n5539 & ~n19545 ;
  assign n25949 = ( n774 & n6224 ) | ( n774 & n23720 ) | ( n6224 & n23720 ) ;
  assign n25950 = n659 & ~n8728 ;
  assign n25951 = n12756 & n25365 ;
  assign n25952 = n25236 ^ n6974 ^ n1118 ;
  assign n25953 = ~n2787 & n9456 ;
  assign n25954 = n4503 & n5908 ;
  assign n25955 = n679 & n25954 ;
  assign n25956 = n3115 ^ n1345 ^ 1'b0 ;
  assign n25957 = n4265 | n25956 ;
  assign n25958 = n25957 ^ n12160 ^ 1'b0 ;
  assign n25959 = n25958 ^ n14854 ^ 1'b0 ;
  assign n25960 = n7163 ^ n6510 ^ 1'b0 ;
  assign n25961 = ( ~n6394 & n21644 ) | ( ~n6394 & n25960 ) | ( n21644 & n25960 ) ;
  assign n25962 = n1741 & n8904 ;
  assign n25963 = ( n3294 & n4481 ) | ( n3294 & ~n25962 ) | ( n4481 & ~n25962 ) ;
  assign n25964 = n4046 | n5635 ;
  assign n25965 = n25964 ^ n17166 ^ 1'b0 ;
  assign n25966 = ~n25963 & n25965 ;
  assign n25967 = n25130 ^ n23808 ^ 1'b0 ;
  assign n25968 = n13887 ^ n9781 ^ 1'b0 ;
  assign n25969 = n16140 ^ n12421 ^ 1'b0 ;
  assign n25970 = n25968 & n25969 ;
  assign n25971 = n7648 & n14842 ;
  assign n25972 = n7942 ^ n7252 ^ 1'b0 ;
  assign n25973 = n12627 & n25972 ;
  assign n25974 = ~n12846 & n25973 ;
  assign n25975 = n10320 & n25974 ;
  assign n25976 = n16216 | n25975 ;
  assign n25977 = n25976 ^ n16885 ^ 1'b0 ;
  assign n25978 = n9577 & ~n25977 ;
  assign n25979 = n2674 & ~n25978 ;
  assign n25980 = ~n25971 & n25979 ;
  assign n25981 = n9098 ^ n2116 ^ n830 ;
  assign n25982 = ( n566 & n16058 ) | ( n566 & n25981 ) | ( n16058 & n25981 ) ;
  assign n25983 = n271 & ~n4506 ;
  assign n25986 = n9002 & ~n21038 ;
  assign n25987 = n17054 & n25986 ;
  assign n25984 = ( n6508 & n8220 ) | ( n6508 & n12861 ) | ( n8220 & n12861 ) ;
  assign n25985 = ~n10317 & n25984 ;
  assign n25988 = n25987 ^ n25985 ^ 1'b0 ;
  assign n25989 = n5771 | n13472 ;
  assign n25990 = n25989 ^ n11318 ^ 1'b0 ;
  assign n25991 = n25990 ^ n18506 ^ 1'b0 ;
  assign n25992 = n6259 & ~n13779 ;
  assign n25993 = n22941 & n25992 ;
  assign n25994 = n3626 | n6305 ;
  assign n25995 = n25994 ^ n8778 ^ 1'b0 ;
  assign n25996 = n8754 | n25995 ;
  assign n25997 = n4546 ^ n296 ^ 1'b0 ;
  assign n25998 = n17946 & n25997 ;
  assign n25999 = n17287 ^ n3739 ^ 1'b0 ;
  assign n26000 = n25998 & ~n25999 ;
  assign n26001 = n2095 | n15631 ;
  assign n26002 = n16735 & ~n26001 ;
  assign n26003 = n22957 & ~n26002 ;
  assign n26004 = n1997 | n9404 ;
  assign n26005 = n10314 & ~n26004 ;
  assign n26006 = n26005 ^ n7562 ^ 1'b0 ;
  assign n26007 = n20905 | n26006 ;
  assign n26008 = n274 | n26007 ;
  assign n26009 = ( n4972 & n7700 ) | ( n4972 & n21649 ) | ( n7700 & n21649 ) ;
  assign n26010 = n26009 ^ n18273 ^ 1'b0 ;
  assign n26011 = n4714 & n5818 ;
  assign n26012 = n5103 & ~n26011 ;
  assign n26013 = ~n11195 & n26012 ;
  assign n26014 = n26013 ^ n13953 ^ 1'b0 ;
  assign n26015 = ~n1075 & n14898 ;
  assign n26016 = n26015 ^ n22258 ^ 1'b0 ;
  assign n26017 = n12948 ^ n12857 ^ 1'b0 ;
  assign n26018 = n26017 ^ n5452 ^ n4868 ;
  assign n26019 = n7245 & n15648 ;
  assign n26020 = ~n4468 & n9996 ;
  assign n26021 = ~n3160 & n26020 ;
  assign n26022 = n26021 ^ n3788 ^ 1'b0 ;
  assign n26023 = ~n26019 & n26022 ;
  assign n26024 = n5392 & ~n11587 ;
  assign n26025 = n13372 & ~n26024 ;
  assign n26026 = n26023 & n26025 ;
  assign n26027 = n428 | n7658 ;
  assign n26028 = n3520 & n26027 ;
  assign n26029 = n23226 ^ n19757 ^ n1748 ;
  assign n26030 = n22451 ^ n6408 ^ 1'b0 ;
  assign n26031 = n13692 & n23055 ;
  assign n26032 = n8476 & n26031 ;
  assign n26033 = n23872 ^ n3082 ^ 1'b0 ;
  assign n26034 = n15069 ^ n9258 ^ 1'b0 ;
  assign n26035 = n1140 & n10480 ;
  assign n26036 = n15648 ^ n3573 ^ 1'b0 ;
  assign n26037 = ~n13773 & n26036 ;
  assign n26038 = ~n6017 & n26037 ;
  assign n26039 = n26038 ^ n3594 ^ 1'b0 ;
  assign n26040 = n1097 & ~n19809 ;
  assign n26041 = n5383 ^ n5031 ^ 1'b0 ;
  assign n26042 = n445 & n26041 ;
  assign n26043 = ~n1772 & n26042 ;
  assign n26044 = ~n5660 & n26043 ;
  assign n26045 = n4520 & ~n5990 ;
  assign n26046 = n7316 & n26045 ;
  assign n26047 = n26046 ^ n7541 ^ n2688 ;
  assign n26048 = n25535 ^ n3461 ^ 1'b0 ;
  assign n26049 = n1028 & ~n2606 ;
  assign n26050 = n26049 ^ n12773 ^ 1'b0 ;
  assign n26056 = n865 & ~n13073 ;
  assign n26057 = ~n19825 & n26056 ;
  assign n26058 = ~n26056 & n26057 ;
  assign n26059 = x46 & ~n1527 ;
  assign n26060 = ~x46 & n26059 ;
  assign n26061 = n2426 & n26060 ;
  assign n26062 = ~n14937 & n26061 ;
  assign n26063 = n14937 & n26062 ;
  assign n26064 = ( n15327 & n26058 ) | ( n15327 & ~n26063 ) | ( n26058 & ~n26063 ) ;
  assign n26051 = ~n1347 & n6650 ;
  assign n26052 = ~n19589 & n26051 ;
  assign n26053 = n26052 ^ n14448 ^ n2466 ;
  assign n26054 = n26053 ^ n19377 ^ n6363 ;
  assign n26055 = n10378 & ~n26054 ;
  assign n26065 = n26064 ^ n26055 ^ 1'b0 ;
  assign n26066 = n8475 ^ n2215 ^ 1'b0 ;
  assign n26067 = n19159 ^ n18390 ^ n1952 ;
  assign n26069 = n8250 ^ n7275 ^ 1'b0 ;
  assign n26068 = n2382 | n9998 ;
  assign n26070 = n26069 ^ n26068 ^ 1'b0 ;
  assign n26071 = ~n2828 & n15131 ;
  assign n26072 = n26071 ^ n16837 ^ 1'b0 ;
  assign n26073 = n16944 ^ n3882 ^ 1'b0 ;
  assign n26075 = n1845 | n2848 ;
  assign n26074 = ~n2726 & n8994 ;
  assign n26076 = n26075 ^ n26074 ^ 1'b0 ;
  assign n26077 = ( n9475 & ~n13661 ) | ( n9475 & n25506 ) | ( ~n13661 & n25506 ) ;
  assign n26080 = n4003 ^ n1648 ^ 1'b0 ;
  assign n26081 = n17765 | n26080 ;
  assign n26078 = n1387 & ~n9967 ;
  assign n26079 = ~n23738 & n26078 ;
  assign n26082 = n26081 ^ n26079 ^ 1'b0 ;
  assign n26083 = n8937 ^ x163 ^ 1'b0 ;
  assign n26084 = n5692 & ~n12576 ;
  assign n26085 = n26084 ^ n4347 ^ 1'b0 ;
  assign n26086 = n7015 & n10690 ;
  assign n26087 = n26085 & n26086 ;
  assign n26089 = ~n7145 & n7442 ;
  assign n26088 = n3755 & ~n20715 ;
  assign n26090 = n26089 ^ n26088 ^ 1'b0 ;
  assign n26091 = n21541 ^ n7707 ^ 1'b0 ;
  assign n26094 = n6680 & n17682 ;
  assign n26093 = ( n1328 & n6920 ) | ( n1328 & n15248 ) | ( n6920 & n15248 ) ;
  assign n26095 = n26094 ^ n26093 ^ 1'b0 ;
  assign n26092 = ~n12301 & n18394 ;
  assign n26096 = n26095 ^ n26092 ^ 1'b0 ;
  assign n26097 = ~n20190 & n24214 ;
  assign n26098 = n9990 & n17580 ;
  assign n26099 = n26098 ^ n8765 ^ 1'b0 ;
  assign n26100 = ~n15003 & n20629 ;
  assign n26101 = n3490 & n26100 ;
  assign n26102 = ( n18300 & n26099 ) | ( n18300 & n26101 ) | ( n26099 & n26101 ) ;
  assign n26104 = n4410 ^ n3413 ^ 1'b0 ;
  assign n26105 = n7312 & ~n26104 ;
  assign n26106 = n20435 ^ x39 ^ 1'b0 ;
  assign n26107 = ( n9751 & n26105 ) | ( n9751 & n26106 ) | ( n26105 & n26106 ) ;
  assign n26103 = n2077 | n23963 ;
  assign n26108 = n26107 ^ n26103 ^ 1'b0 ;
  assign n26109 = n7105 & n23065 ;
  assign n26110 = ~n8087 & n26109 ;
  assign n26111 = n2463 & n11371 ;
  assign n26112 = n21682 & n26111 ;
  assign n26113 = n26112 ^ n13068 ^ 1'b0 ;
  assign n26114 = n8815 | n26113 ;
  assign n26115 = n11769 ^ n1017 ^ 1'b0 ;
  assign n26116 = n21007 & ~n26115 ;
  assign n26117 = ~n2532 & n4249 ;
  assign n26118 = n8182 ^ n6524 ^ 1'b0 ;
  assign n26119 = n9115 | n13505 ;
  assign n26120 = n26118 | n26119 ;
  assign n26121 = n7576 ^ n1413 ^ 1'b0 ;
  assign n26122 = n6772 & n26121 ;
  assign n26123 = n13666 & n26122 ;
  assign n26124 = ~n26120 & n26123 ;
  assign n26127 = n7557 | n8351 ;
  assign n26125 = n5794 & ~n7001 ;
  assign n26126 = n21077 & ~n26125 ;
  assign n26128 = n26127 ^ n26126 ^ 1'b0 ;
  assign n26129 = n5958 ^ n4642 ^ 1'b0 ;
  assign n26130 = n2325 & n26129 ;
  assign n26131 = ~n5195 & n6880 ;
  assign n26132 = n26131 ^ n4585 ^ 1'b0 ;
  assign n26133 = n17711 ^ n9022 ^ 1'b0 ;
  assign n26134 = n1623 | n26133 ;
  assign n26135 = n26132 | n26134 ;
  assign n26136 = n2651 ^ n1295 ^ 1'b0 ;
  assign n26137 = n4840 ^ n3296 ^ 1'b0 ;
  assign n26138 = ~n17646 & n18308 ;
  assign n26139 = n26138 ^ n24733 ^ 1'b0 ;
  assign n26140 = n5602 | n22182 ;
  assign n26141 = n11400 & ~n26140 ;
  assign n26142 = n829 | n9036 ;
  assign n26143 = n18258 ^ n596 ^ 1'b0 ;
  assign n26144 = n26143 ^ n1623 ^ 1'b0 ;
  assign n26145 = n7123 | n11371 ;
  assign n26146 = n26145 ^ n12945 ^ 1'b0 ;
  assign n26147 = n19957 & ~n26146 ;
  assign n26148 = n8632 ^ n7026 ^ 1'b0 ;
  assign n26149 = ~n3763 & n26148 ;
  assign n26150 = x168 & n16923 ;
  assign n26151 = ~n26149 & n26150 ;
  assign n26152 = x139 & n3757 ;
  assign n26153 = ~n7819 & n26152 ;
  assign n26154 = x153 & n26153 ;
  assign n26155 = n23761 ^ n2936 ^ 1'b0 ;
  assign n26156 = n4441 ^ n4387 ^ 1'b0 ;
  assign n26157 = n26155 & n26156 ;
  assign n26158 = n7051 & n10795 ;
  assign n26159 = ~n26157 & n26158 ;
  assign n26160 = ~n9507 & n16198 ;
  assign n26161 = n13789 ^ n503 ^ 1'b0 ;
  assign n26162 = n26161 ^ n18194 ^ 1'b0 ;
  assign n26163 = n7319 ^ n1741 ^ 1'b0 ;
  assign n26164 = n16092 | n26163 ;
  assign n26165 = n1006 & n17179 ;
  assign n26166 = n2929 ^ n839 ^ 1'b0 ;
  assign n26167 = n18392 | n26166 ;
  assign n26168 = n26167 ^ n7353 ^ n7086 ;
  assign n26169 = n26168 ^ n6629 ^ 1'b0 ;
  assign n26172 = ( ~n492 & n1839 ) | ( ~n492 & n9194 ) | ( n1839 & n9194 ) ;
  assign n26170 = n2992 & ~n4267 ;
  assign n26171 = n3699 & n26170 ;
  assign n26173 = n26172 ^ n26171 ^ 1'b0 ;
  assign n26174 = n7147 | n25361 ;
  assign n26175 = n26174 ^ n17907 ^ 1'b0 ;
  assign n26176 = n12694 & ~n13382 ;
  assign n26177 = n13331 & n26176 ;
  assign n26178 = n14429 | n26177 ;
  assign n26179 = ( n1051 & n2043 ) | ( n1051 & n6400 ) | ( n2043 & n6400 ) ;
  assign n26180 = n13283 ^ n10372 ^ 1'b0 ;
  assign n26181 = n5420 & ~n13845 ;
  assign n26182 = n18774 & n26181 ;
  assign n26183 = n11084 & ~n26182 ;
  assign n26184 = n9911 | n26183 ;
  assign n26185 = n4117 & ~n22173 ;
  assign n26186 = n26185 ^ n18655 ^ 1'b0 ;
  assign n26187 = n2463 & n26186 ;
  assign n26188 = n16415 ^ n16059 ^ n14716 ;
  assign n26190 = n7353 ^ n2247 ^ 1'b0 ;
  assign n26189 = n16885 & ~n18110 ;
  assign n26191 = n26190 ^ n26189 ^ 1'b0 ;
  assign n26192 = n4462 & n5525 ;
  assign n26193 = ( ~n6340 & n19546 ) | ( ~n6340 & n26192 ) | ( n19546 & n26192 ) ;
  assign n26194 = n11116 & ~n13061 ;
  assign n26195 = n26194 ^ x131 ^ 1'b0 ;
  assign n26196 = n26195 ^ n8380 ^ 1'b0 ;
  assign n26197 = n5176 & ~n26196 ;
  assign n26198 = n4594 & ~n9348 ;
  assign n26199 = n26198 ^ n4509 ^ n4330 ;
  assign n26200 = ~n11778 & n11941 ;
  assign n26201 = n21441 | n26200 ;
  assign n26202 = n26201 ^ n6921 ^ 1'b0 ;
  assign n26203 = n3622 | n15674 ;
  assign n26204 = n26203 ^ n9661 ^ 1'b0 ;
  assign n26205 = ( n5934 & ~n7804 ) | ( n5934 & n26204 ) | ( ~n7804 & n26204 ) ;
  assign n26206 = n5325 ^ n4964 ^ 1'b0 ;
  assign n26207 = n24781 ^ n11820 ^ 1'b0 ;
  assign n26208 = ( n3161 & n12607 ) | ( n3161 & ~n26207 ) | ( n12607 & ~n26207 ) ;
  assign n26211 = n2106 & n10634 ;
  assign n26209 = n4078 & n4403 ;
  assign n26210 = n3253 & n26209 ;
  assign n26212 = n26211 ^ n26210 ^ 1'b0 ;
  assign n26213 = ~n19166 & n22819 ;
  assign n26214 = n26213 ^ n9605 ^ 1'b0 ;
  assign n26215 = n22375 | n25940 ;
  assign n26216 = n26215 ^ n6830 ^ n5525 ;
  assign n26217 = n17065 ^ n12188 ^ n1521 ;
  assign n26218 = n26217 ^ n14501 ^ 1'b0 ;
  assign n26219 = n3966 & ~n26218 ;
  assign n26220 = n3841 ^ n2411 ^ 1'b0 ;
  assign n26221 = n8087 & ~n26220 ;
  assign n26222 = ~n1474 & n4520 ;
  assign n26223 = n4319 | n26222 ;
  assign n26224 = n26223 ^ n13607 ^ 1'b0 ;
  assign n26225 = n26221 & n26224 ;
  assign n26226 = n7430 | n18580 ;
  assign n26227 = n24781 & ~n26226 ;
  assign n26228 = n26227 ^ n21781 ^ n10368 ;
  assign n26229 = ~n1720 & n18336 ;
  assign n26230 = ~n11087 & n26229 ;
  assign n26231 = n20935 ^ n18384 ^ 1'b0 ;
  assign n26232 = ~n26230 & n26231 ;
  assign n26233 = x113 & n21583 ;
  assign n26234 = ~n4193 & n6359 ;
  assign n26235 = n26234 ^ n7932 ^ 1'b0 ;
  assign n26236 = ~n18828 & n26235 ;
  assign n26237 = n18286 ^ n9355 ^ 1'b0 ;
  assign n26238 = n20653 & n26237 ;
  assign n26239 = n2946 | n24150 ;
  assign n26240 = n26238 | n26239 ;
  assign n26241 = n4840 & ~n13661 ;
  assign n26242 = n26241 ^ n12643 ^ 1'b0 ;
  assign n26243 = n451 | n22032 ;
  assign n26244 = n9440 ^ n1817 ^ 1'b0 ;
  assign n26245 = ( n1940 & ~n2257 ) | ( n1940 & n26244 ) | ( ~n2257 & n26244 ) ;
  assign n26249 = n1065 & ~n4638 ;
  assign n26250 = n9359 & n26249 ;
  assign n26246 = ~n4400 & n6638 ;
  assign n26247 = ~n23608 & n26246 ;
  assign n26248 = n9580 & n26247 ;
  assign n26251 = n26250 ^ n26248 ^ 1'b0 ;
  assign n26252 = ~n2433 & n8907 ;
  assign n26253 = n23782 ^ n10176 ^ 1'b0 ;
  assign n26254 = n26253 ^ n889 ^ x169 ;
  assign n26255 = n5773 ^ n917 ^ 1'b0 ;
  assign n26256 = n21802 & n26255 ;
  assign n26257 = ( n1876 & n13445 ) | ( n1876 & n14416 ) | ( n13445 & n14416 ) ;
  assign n26258 = n26257 ^ n13432 ^ 1'b0 ;
  assign n26259 = n18917 & ~n26005 ;
  assign n26260 = ~n3848 & n26259 ;
  assign n26261 = n13658 & n16487 ;
  assign n26262 = n14220 & n26261 ;
  assign n26263 = ( n19411 & n26260 ) | ( n19411 & ~n26262 ) | ( n26260 & ~n26262 ) ;
  assign n26264 = n11855 ^ n1778 ^ 1'b0 ;
  assign n26265 = n20360 ^ n6020 ^ n5509 ;
  assign n26266 = n26265 ^ n6049 ^ 1'b0 ;
  assign n26267 = n22847 & n26266 ;
  assign n26268 = ~n8425 & n9243 ;
  assign n26269 = ~n15360 & n26268 ;
  assign n26270 = n26269 ^ n2559 ^ 1'b0 ;
  assign n26271 = n17501 ^ n3590 ^ 1'b0 ;
  assign n26272 = n26270 | n26271 ;
  assign n26273 = ~n3234 & n3922 ;
  assign n26274 = n26273 ^ n25928 ^ 1'b0 ;
  assign n26275 = x0 | n3032 ;
  assign n26276 = n3651 & n26275 ;
  assign n26277 = n26276 ^ n16355 ^ 1'b0 ;
  assign n26278 = n5936 | n21718 ;
  assign n26279 = n26277 | n26278 ;
  assign n26280 = n3716 ^ n3328 ^ 1'b0 ;
  assign n26281 = ( n11981 & n24581 ) | ( n11981 & n26280 ) | ( n24581 & n26280 ) ;
  assign n26282 = n26281 ^ n17676 ^ n17544 ;
  assign n26283 = n3206 ^ n1589 ^ 1'b0 ;
  assign n26284 = n26283 ^ n15080 ^ n5392 ;
  assign n26285 = n15213 | n21754 ;
  assign n26286 = n6492 ^ n3451 ^ x3 ;
  assign n26287 = ~n26285 & n26286 ;
  assign n26288 = n10145 & n26287 ;
  assign n26289 = n6319 & n22198 ;
  assign n26290 = n13585 ^ n11253 ^ 1'b0 ;
  assign n26291 = ~n2574 & n26290 ;
  assign n26292 = n4871 & ~n15135 ;
  assign n26293 = n26292 ^ n21976 ^ 1'b0 ;
  assign n26294 = n17247 ^ n8157 ^ 1'b0 ;
  assign n26295 = n708 & n2224 ;
  assign n26296 = n26295 ^ n4387 ^ 1'b0 ;
  assign n26297 = ~n11662 & n26296 ;
  assign n26298 = n26297 ^ n15680 ^ n14829 ;
  assign n26299 = ~n16479 & n25221 ;
  assign n26300 = n26299 ^ n24410 ^ 1'b0 ;
  assign n26301 = ( n17638 & n26298 ) | ( n17638 & ~n26300 ) | ( n26298 & ~n26300 ) ;
  assign n26302 = n12611 & ~n20603 ;
  assign n26303 = n16058 ^ n12515 ^ n6171 ;
  assign n26304 = n1217 & ~n26303 ;
  assign n26305 = ~n19797 & n26304 ;
  assign n26306 = n4569 | n9130 ;
  assign n26307 = n592 & ~n15479 ;
  assign n26308 = n7935 | n26307 ;
  assign n26309 = n14114 ^ n13384 ^ 1'b0 ;
  assign n26310 = n26308 | n26309 ;
  assign n26312 = n2622 & ~n12074 ;
  assign n26313 = n6202 & ~n26312 ;
  assign n26314 = n17168 & n26313 ;
  assign n26311 = n5539 & ~n21521 ;
  assign n26315 = n26314 ^ n26311 ^ 1'b0 ;
  assign n26316 = ~n1714 & n13762 ;
  assign n26317 = n9167 ^ n5722 ^ n498 ;
  assign n26318 = n26317 ^ n11657 ^ 1'b0 ;
  assign n26319 = n5177 ^ n4970 ^ n4447 ;
  assign n26320 = n16148 ^ n3682 ^ 1'b0 ;
  assign n26321 = n26319 & ~n26320 ;
  assign n26322 = n4065 | n7179 ;
  assign n26323 = n10470 & ~n26322 ;
  assign n26324 = ~n22923 & n26323 ;
  assign n26325 = n25702 & n26324 ;
  assign n26326 = n5278 & ~n22579 ;
  assign n26327 = ~n10899 & n26326 ;
  assign n26328 = n19399 & ~n26327 ;
  assign n26329 = n24391 ^ n8444 ^ 1'b0 ;
  assign n26330 = ~n14979 & n19722 ;
  assign n26331 = n14052 ^ n13452 ^ 1'b0 ;
  assign n26332 = n16801 ^ n1952 ^ 1'b0 ;
  assign n26333 = x163 & n10888 ;
  assign n26334 = n26333 ^ n25633 ^ 1'b0 ;
  assign n26335 = n5107 ^ n4391 ^ 1'b0 ;
  assign n26336 = ( ~n364 & n26334 ) | ( ~n364 & n26335 ) | ( n26334 & n26335 ) ;
  assign n26337 = ~n18221 & n26336 ;
  assign n26338 = ~n4642 & n16301 ;
  assign n26339 = ( n11529 & n12136 ) | ( n11529 & n19207 ) | ( n12136 & n19207 ) ;
  assign n26340 = ( x69 & n1682 ) | ( x69 & ~n26339 ) | ( n1682 & ~n26339 ) ;
  assign n26344 = n13602 ^ n6701 ^ n3195 ;
  assign n26341 = ( n3825 & n10988 ) | ( n3825 & ~n13184 ) | ( n10988 & ~n13184 ) ;
  assign n26342 = n13630 & n26341 ;
  assign n26343 = n7810 | n26342 ;
  assign n26345 = n26344 ^ n26343 ^ 1'b0 ;
  assign n26346 = ( n4011 & n26340 ) | ( n4011 & ~n26345 ) | ( n26340 & ~n26345 ) ;
  assign n26347 = n4210 & ~n12806 ;
  assign n26348 = ( n8717 & n15543 ) | ( n8717 & n26347 ) | ( n15543 & n26347 ) ;
  assign n26349 = ~n17520 & n18154 ;
  assign n26350 = n26349 ^ n23233 ^ 1'b0 ;
  assign n26351 = ~n19297 & n24418 ;
  assign n26352 = n26351 ^ n2552 ^ 1'b0 ;
  assign n26353 = n11069 | n15758 ;
  assign n26354 = n26353 ^ n16210 ^ 1'b0 ;
  assign n26355 = n10191 & ~n26354 ;
  assign n26356 = ~n547 & n26355 ;
  assign n26359 = ~n3918 & n10922 ;
  assign n26360 = ~n4830 & n26359 ;
  assign n26361 = ~n5951 & n24416 ;
  assign n26362 = n26360 & n26361 ;
  assign n26363 = n26362 ^ n3040 ^ 1'b0 ;
  assign n26364 = n21598 | n26363 ;
  assign n26357 = n1726 & ~n8391 ;
  assign n26358 = ~n5797 & n26357 ;
  assign n26365 = n26364 ^ n26358 ^ 1'b0 ;
  assign n26366 = n8214 ^ n3041 ^ 1'b0 ;
  assign n26367 = n9036 & n26366 ;
  assign n26368 = n21296 & ~n26367 ;
  assign n26369 = n25544 ^ n14122 ^ 1'b0 ;
  assign n26370 = n18396 ^ n922 ^ 1'b0 ;
  assign n26371 = n14584 ^ n2839 ^ 1'b0 ;
  assign n26372 = n2557 & ~n7579 ;
  assign n26373 = n26371 & ~n26372 ;
  assign n26374 = ~n12214 & n26373 ;
  assign n26375 = n8547 & n8860 ;
  assign n26376 = n8869 ^ n1802 ^ 1'b0 ;
  assign n26377 = n26376 ^ n19006 ^ 1'b0 ;
  assign n26378 = n16285 & n26377 ;
  assign n26379 = ( n6220 & n17752 ) | ( n6220 & n20693 ) | ( n17752 & n20693 ) ;
  assign n26380 = n26379 ^ n2916 ^ 1'b0 ;
  assign n26381 = n11759 ^ x25 ^ 1'b0 ;
  assign n26382 = n925 & n9912 ;
  assign n26383 = ~n925 & n26382 ;
  assign n26384 = n23485 ^ n16341 ^ 1'b0 ;
  assign n26385 = ~n26383 & n26384 ;
  assign n26386 = n23226 ^ n16987 ^ 1'b0 ;
  assign n26387 = x86 & n1866 ;
  assign n26388 = ~n4637 & n26387 ;
  assign n26389 = ( ~n394 & n16095 ) | ( ~n394 & n26388 ) | ( n16095 & n26388 ) ;
  assign n26390 = n26389 ^ n5420 ^ 1'b0 ;
  assign n26391 = n11529 & n25365 ;
  assign n26392 = n26391 ^ n11416 ^ 1'b0 ;
  assign n26393 = n2130 & n13845 ;
  assign n26394 = n11753 & ~n13364 ;
  assign n26395 = n13873 & n26394 ;
  assign n26400 = n5111 | n15608 ;
  assign n26401 = n14842 & n26400 ;
  assign n26396 = n1799 & ~n2789 ;
  assign n26397 = n26396 ^ n11178 ^ 1'b0 ;
  assign n26398 = n20172 | n26397 ;
  assign n26399 = n23810 | n26398 ;
  assign n26402 = n26401 ^ n26399 ^ 1'b0 ;
  assign n26403 = n7681 ^ n3142 ^ 1'b0 ;
  assign n26404 = n4198 & ~n26403 ;
  assign n26405 = n11458 & n13271 ;
  assign n26406 = n26405 ^ n23979 ^ n5029 ;
  assign n26407 = n5265 & n15773 ;
  assign n26408 = n26407 ^ n17721 ^ 1'b0 ;
  assign n26409 = n7686 ^ n3463 ^ 1'b0 ;
  assign n26410 = n4931 | n23786 ;
  assign n26411 = n26409 & ~n26410 ;
  assign n26412 = n15199 ^ n14240 ^ n5608 ;
  assign n26413 = n1901 & ~n2095 ;
  assign n26414 = n6395 & ~n8129 ;
  assign n26415 = ~n26413 & n26414 ;
  assign n26417 = n8424 ^ n1738 ^ 1'b0 ;
  assign n26418 = n10520 & ~n26417 ;
  assign n26419 = n9938 ^ n7569 ^ 1'b0 ;
  assign n26420 = ( n16214 & n26418 ) | ( n16214 & n26419 ) | ( n26418 & n26419 ) ;
  assign n26416 = n3627 | n16212 ;
  assign n26421 = n26420 ^ n26416 ^ 1'b0 ;
  assign n26423 = n4280 & ~n6483 ;
  assign n26424 = n26423 ^ n2711 ^ 1'b0 ;
  assign n26422 = n1671 & n15275 ;
  assign n26425 = n26424 ^ n26422 ^ 1'b0 ;
  assign n26426 = n23152 ^ n16612 ^ 1'b0 ;
  assign n26427 = n16480 & n26426 ;
  assign n26428 = n5034 | n14521 ;
  assign n26429 = x126 | n26428 ;
  assign n26430 = n15697 ^ n11924 ^ 1'b0 ;
  assign n26431 = ~n3898 & n26430 ;
  assign n26432 = n22378 ^ n20257 ^ 1'b0 ;
  assign n26433 = ~n26172 & n26432 ;
  assign n26434 = n8975 & n13271 ;
  assign n26435 = n14000 ^ x63 ^ 1'b0 ;
  assign n26436 = n7382 & ~n26435 ;
  assign n26437 = x13 & x199 ;
  assign n26438 = ~x199 & n26437 ;
  assign n26439 = n1023 & n1591 ;
  assign n26440 = ~n1591 & n26439 ;
  assign n26441 = n26438 & ~n26440 ;
  assign n26442 = n26436 & n26441 ;
  assign n26443 = ~n26436 & n26442 ;
  assign n26444 = n26443 ^ n22094 ^ 1'b0 ;
  assign n26445 = n10731 ^ x180 ^ 1'b0 ;
  assign n26446 = x244 & ~n22947 ;
  assign n26447 = n21766 & n26446 ;
  assign n26448 = n1360 | n3894 ;
  assign n26449 = n26448 ^ x243 ^ 1'b0 ;
  assign n26450 = n3028 & ~n26449 ;
  assign n26451 = n26450 ^ n9365 ^ 1'b0 ;
  assign n26452 = n1505 | n26451 ;
  assign n26453 = n12864 & ~n26452 ;
  assign n26454 = n26447 & n26453 ;
  assign n26456 = n1848 & n18770 ;
  assign n26457 = n26456 ^ n8914 ^ 1'b0 ;
  assign n26455 = n7361 | n9534 ;
  assign n26458 = n26457 ^ n26455 ^ 1'b0 ;
  assign n26460 = ~n6253 & n9984 ;
  assign n26461 = ~n1125 & n26460 ;
  assign n26459 = x36 & n10374 ;
  assign n26462 = n26461 ^ n26459 ^ 1'b0 ;
  assign n26463 = x129 & n25492 ;
  assign n26464 = n26462 | n26463 ;
  assign n26465 = ( n18862 & n20478 ) | ( n18862 & n22634 ) | ( n20478 & n22634 ) ;
  assign n26466 = n21712 | n22596 ;
  assign n26467 = n10316 & n13851 ;
  assign n26468 = ~n4869 & n26467 ;
  assign n26469 = ~n2687 & n26468 ;
  assign n26470 = n14206 ^ n10990 ^ n9215 ;
  assign n26471 = n26470 ^ n19805 ^ 1'b0 ;
  assign n26472 = ~n963 & n26471 ;
  assign n26473 = n1611 & n23044 ;
  assign n26474 = n6620 ^ n3989 ^ n3568 ;
  assign n26475 = n17722 ^ n1620 ^ 1'b0 ;
  assign n26476 = ( n4596 & ~n26474 ) | ( n4596 & n26475 ) | ( ~n26474 & n26475 ) ;
  assign n26477 = ~n13406 & n25334 ;
  assign n26478 = n25137 & n26477 ;
  assign n26481 = ( ~n6481 & n15500 ) | ( ~n6481 & n18248 ) | ( n15500 & n18248 ) ;
  assign n26479 = n6965 ^ n3729 ^ n850 ;
  assign n26480 = n26479 ^ n20245 ^ 1'b0 ;
  assign n26482 = n26481 ^ n26480 ^ 1'b0 ;
  assign n26483 = n8107 ^ n1129 ^ 1'b0 ;
  assign n26484 = n10674 | n26483 ;
  assign n26485 = n520 & ~n26484 ;
  assign n26486 = n26482 & ~n26485 ;
  assign n26487 = ~n24208 & n26486 ;
  assign n26488 = n18180 ^ n12290 ^ 1'b0 ;
  assign n26489 = n26488 ^ n11717 ^ 1'b0 ;
  assign n26490 = n2998 & ~n26489 ;
  assign n26491 = n784 & ~n1242 ;
  assign n26492 = n8632 | n11630 ;
  assign n26493 = n10248 | n22658 ;
  assign n26494 = n3291 & ~n26493 ;
  assign n26495 = n919 & ~n4593 ;
  assign n26496 = n26495 ^ n1086 ^ 1'b0 ;
  assign n26497 = ~n4906 & n26496 ;
  assign n26498 = ~n12030 & n21041 ;
  assign n26499 = ~n17635 & n26498 ;
  assign n26504 = n19919 ^ n5368 ^ 1'b0 ;
  assign n26500 = n2763 | n13765 ;
  assign n26501 = n3388 & ~n26500 ;
  assign n26502 = n26501 ^ n17701 ^ 1'b0 ;
  assign n26503 = ~n10251 & n26502 ;
  assign n26505 = n26504 ^ n26503 ^ 1'b0 ;
  assign n26506 = n26505 ^ n11623 ^ 1'b0 ;
  assign n26507 = n25137 ^ n9521 ^ 1'b0 ;
  assign n26508 = n8209 ^ n2514 ^ 1'b0 ;
  assign n26509 = n7365 & n22071 ;
  assign n26510 = ~n3067 & n11633 ;
  assign n26511 = ~n4659 & n26510 ;
  assign n26512 = n26511 ^ n13221 ^ n810 ;
  assign n26513 = n8308 | n26512 ;
  assign n26514 = ~n19934 & n26145 ;
  assign n26515 = ~n12625 & n26514 ;
  assign n26516 = n26515 ^ n1028 ^ 1'b0 ;
  assign n26517 = n2940 & ~n26516 ;
  assign n26518 = n2062 | n10599 ;
  assign n26519 = n11782 ^ n603 ^ 1'b0 ;
  assign n26520 = ( n2528 & ~n2653 ) | ( n2528 & n26519 ) | ( ~n2653 & n26519 ) ;
  assign n26521 = ( n7594 & n20833 ) | ( n7594 & n26520 ) | ( n20833 & n26520 ) ;
  assign n26522 = ~n4207 & n22723 ;
  assign n26523 = n26521 & n26522 ;
  assign n26524 = n25696 ^ n16025 ^ n6687 ;
  assign n26525 = n26524 ^ n2623 ^ 1'b0 ;
  assign n26526 = n25708 & ~n26525 ;
  assign n26527 = n2901 | n20443 ;
  assign n26528 = n466 & n5051 ;
  assign n26529 = ~n973 & n5309 ;
  assign n26530 = n23846 ^ n4821 ^ 1'b0 ;
  assign n26531 = n24655 & n26530 ;
  assign n26532 = ( ~n635 & n6069 ) | ( ~n635 & n6113 ) | ( n6069 & n6113 ) ;
  assign n26533 = ( n14758 & n17328 ) | ( n14758 & ~n26532 ) | ( n17328 & ~n26532 ) ;
  assign n26534 = n17544 ^ n7035 ^ 1'b0 ;
  assign n26535 = n15076 & n26534 ;
  assign n26536 = n26533 & n26535 ;
  assign n26537 = n26536 ^ n17753 ^ n513 ;
  assign n26538 = ~n1973 & n3121 ;
  assign n26539 = n26538 ^ n15070 ^ 1'b0 ;
  assign n26540 = n13827 | n26539 ;
  assign n26541 = n5459 | n26540 ;
  assign n26542 = n3667 | n26541 ;
  assign n26543 = n9207 ^ n1804 ^ 1'b0 ;
  assign n26544 = ~n4329 & n26543 ;
  assign n26545 = n26542 | n26544 ;
  assign n26546 = n12318 ^ n2008 ^ n1153 ;
  assign n26547 = ~n2271 & n7629 ;
  assign n26548 = n26546 & n26547 ;
  assign n26549 = n24973 | n26548 ;
  assign n26550 = n619 & ~n26549 ;
  assign n26551 = n3286 & ~n13228 ;
  assign n26552 = n6387 ^ n2065 ^ 1'b0 ;
  assign n26553 = n5596 & ~n26552 ;
  assign n26554 = n7624 & n24131 ;
  assign n26555 = n17114 | n26554 ;
  assign n26556 = n1611 | n4803 ;
  assign n26557 = n4981 & n21320 ;
  assign n26558 = n26557 ^ n10974 ^ 1'b0 ;
  assign n26559 = n26558 ^ n17038 ^ n270 ;
  assign n26560 = n19733 ^ n5350 ^ 1'b0 ;
  assign n26561 = n10425 ^ n2332 ^ 1'b0 ;
  assign n26562 = n26560 | n26561 ;
  assign n26563 = n19411 & ~n26562 ;
  assign n26564 = n26563 ^ n6017 ^ 1'b0 ;
  assign n26565 = n22709 ^ n6713 ^ 1'b0 ;
  assign n26566 = n6208 & ~n14146 ;
  assign n26567 = n26566 ^ n3736 ^ 1'b0 ;
  assign n26568 = n6402 & n13727 ;
  assign n26569 = n3419 ^ x199 ^ 1'b0 ;
  assign n26570 = ~n1124 & n5621 ;
  assign n26571 = ( n11291 & ~n21546 ) | ( n11291 & n26570 ) | ( ~n21546 & n26570 ) ;
  assign n26572 = n25135 ^ n13357 ^ 1'b0 ;
  assign n26573 = n4647 & ~n26572 ;
  assign n26574 = n3695 & n26573 ;
  assign n26575 = n8072 & n26574 ;
  assign n26576 = n8413 ^ n4065 ^ 1'b0 ;
  assign n26577 = ~n21901 & n26576 ;
  assign n26578 = ~n10241 & n22225 ;
  assign n26579 = n26578 ^ n15655 ^ 1'b0 ;
  assign n26580 = ~n3670 & n8517 ;
  assign n26581 = n13574 | n13863 ;
  assign n26582 = n18955 ^ n15109 ^ n4752 ;
  assign n26583 = n7613 ^ n1603 ^ 1'b0 ;
  assign n26584 = n4072 & n26583 ;
  assign n26588 = n2061 | n5729 ;
  assign n26585 = n9280 ^ n8041 ^ n3416 ;
  assign n26586 = n26585 ^ n2314 ^ n1610 ;
  assign n26587 = n11529 | n26586 ;
  assign n26589 = n26588 ^ n26587 ^ 1'b0 ;
  assign n26590 = ~n1067 & n7071 ;
  assign n26591 = n7303 & n26590 ;
  assign n26592 = n13149 | n26591 ;
  assign n26593 = n11057 ^ n2657 ^ 1'b0 ;
  assign n26594 = n26593 ^ n25671 ^ 1'b0 ;
  assign n26595 = n25053 | n26594 ;
  assign n26596 = ~n4896 & n8098 ;
  assign n26597 = n9065 & n26596 ;
  assign n26598 = n26597 ^ n1413 ^ 1'b0 ;
  assign n26599 = n10340 ^ n8119 ^ 1'b0 ;
  assign n26600 = n23690 & n26599 ;
  assign n26601 = ~n26598 & n26600 ;
  assign n26602 = ~n12725 & n16295 ;
  assign n26603 = n4541 | n26602 ;
  assign n26606 = n7300 & n18761 ;
  assign n26604 = n22644 ^ x45 ^ 1'b0 ;
  assign n26605 = n19098 | n26604 ;
  assign n26607 = n26606 ^ n26605 ^ n14514 ;
  assign n26608 = ~n8676 & n13814 ;
  assign n26609 = n4629 & ~n26608 ;
  assign n26610 = ( n19386 & n20510 ) | ( n19386 & n26609 ) | ( n20510 & n26609 ) ;
  assign n26611 = n24098 ^ n16388 ^ 1'b0 ;
  assign n26612 = ~n8371 & n9206 ;
  assign n26613 = ~n6315 & n15672 ;
  assign n26614 = n14711 & n26613 ;
  assign n26615 = n26614 ^ n2485 ^ 1'b0 ;
  assign n26616 = n7160 & ~n14526 ;
  assign n26617 = n8087 & ~n26616 ;
  assign n26618 = ~n10146 & n26617 ;
  assign n26619 = n24998 ^ n22591 ^ 1'b0 ;
  assign n26620 = n21084 & n26619 ;
  assign n26621 = n1744 & ~n19218 ;
  assign n26622 = n9961 & n23062 ;
  assign n26623 = n26622 ^ n15987 ^ 1'b0 ;
  assign n26624 = ~n419 & n16750 ;
  assign n26625 = n26624 ^ n12668 ^ 1'b0 ;
  assign n26626 = n8839 & ~n11833 ;
  assign n26627 = n26626 ^ n24775 ^ 1'b0 ;
  assign n26628 = n2172 & n24483 ;
  assign n26629 = n23156 & ~n26628 ;
  assign n26630 = n713 & ~n21436 ;
  assign n26631 = n7472 & n26630 ;
  assign n26632 = n8241 & ~n13377 ;
  assign n26633 = n16840 ^ n6496 ^ 1'b0 ;
  assign n26634 = n4840 | n13275 ;
  assign n26635 = n9711 ^ n1704 ^ 1'b0 ;
  assign n26636 = n4593 | n26635 ;
  assign n26637 = n5682 & n26636 ;
  assign n26638 = ~n4660 & n5592 ;
  assign n26639 = n26638 ^ n9919 ^ 1'b0 ;
  assign n26640 = n1039 & ~n10735 ;
  assign n26641 = n3158 & n7930 ;
  assign n26642 = ~n26640 & n26641 ;
  assign n26643 = n26639 | n26642 ;
  assign n26644 = n19185 | n26643 ;
  assign n26645 = n26644 ^ n18026 ^ 1'b0 ;
  assign n26646 = n9218 ^ n8236 ^ n5181 ;
  assign n26647 = n10268 | n10377 ;
  assign n26648 = n23164 ^ n11319 ^ 1'b0 ;
  assign n26649 = n26647 & n26648 ;
  assign n26650 = n24581 ^ n13610 ^ 1'b0 ;
  assign n26651 = n6502 | n26650 ;
  assign n26652 = n19052 ^ n16165 ^ 1'b0 ;
  assign n26653 = n18675 ^ n2161 ^ 1'b0 ;
  assign n26654 = ~n26652 & n26653 ;
  assign n26655 = ~n1605 & n26105 ;
  assign n26656 = n26655 ^ n3382 ^ 1'b0 ;
  assign n26657 = n15839 & ~n26656 ;
  assign n26658 = n26657 ^ n2622 ^ 1'b0 ;
  assign n26659 = ~n24717 & n26658 ;
  assign n26660 = n16588 ^ n5856 ^ 1'b0 ;
  assign n26661 = ~n4553 & n23907 ;
  assign n26662 = n26661 ^ n25294 ^ 1'b0 ;
  assign n26663 = ~n7443 & n15795 ;
  assign n26664 = n12815 | n20121 ;
  assign n26665 = n26664 ^ n1878 ^ 1'b0 ;
  assign n26666 = n21891 & n26665 ;
  assign n26667 = n9287 & n26666 ;
  assign n26668 = n5944 ^ n4316 ^ n3677 ;
  assign n26669 = n26668 ^ n23249 ^ 1'b0 ;
  assign n26670 = n9929 & n13828 ;
  assign n26671 = n26670 ^ n19990 ^ 1'b0 ;
  assign n26672 = n14440 & n26671 ;
  assign n26673 = n26672 ^ n9520 ^ 1'b0 ;
  assign n26674 = n1262 ^ n983 ^ 1'b0 ;
  assign n26675 = ~n5025 & n7685 ;
  assign n26676 = n26675 ^ n5825 ^ 1'b0 ;
  assign n26677 = n14663 | n26676 ;
  assign n26678 = n935 | n26677 ;
  assign n26679 = n26678 ^ n12013 ^ 1'b0 ;
  assign n26680 = ~n2047 & n16524 ;
  assign n26681 = n2047 & n26680 ;
  assign n26682 = n15858 & ~n26681 ;
  assign n26683 = ~n6104 & n26682 ;
  assign n26684 = n26683 ^ n10608 ^ 1'b0 ;
  assign n26685 = n16438 ^ n16320 ^ 1'b0 ;
  assign n26686 = n3458 ^ n3222 ^ 1'b0 ;
  assign n26687 = n26685 & n26686 ;
  assign n26688 = n17597 ^ n5232 ^ 1'b0 ;
  assign n26689 = n7584 & n7876 ;
  assign n26690 = n20450 ^ n4541 ^ 1'b0 ;
  assign n26691 = n26689 & n26690 ;
  assign n26692 = n25982 ^ n25616 ^ 1'b0 ;
  assign n26693 = n13829 & ~n17426 ;
  assign n26694 = ( n18649 & n23260 ) | ( n18649 & n26693 ) | ( n23260 & n26693 ) ;
  assign n26695 = ( n2932 & ~n5359 ) | ( n2932 & n9124 ) | ( ~n5359 & n9124 ) ;
  assign n26696 = n1330 & ~n26695 ;
  assign n26697 = n26696 ^ n16638 ^ 1'b0 ;
  assign n26698 = n8508 & n11659 ;
  assign n26699 = ~n1544 & n16429 ;
  assign n26700 = ~n1069 & n8622 ;
  assign n26701 = ~n13300 & n26700 ;
  assign n26702 = n14887 | n26701 ;
  assign n26703 = n26699 & ~n26702 ;
  assign n26704 = n14737 ^ n3233 ^ 1'b0 ;
  assign n26705 = n7507 | n26704 ;
  assign n26706 = ~n8883 & n23513 ;
  assign n26707 = n21720 ^ n14867 ^ 1'b0 ;
  assign n26708 = n18177 | n26707 ;
  assign n26709 = ~n14307 & n20578 ;
  assign n26710 = n26709 ^ n7107 ^ 1'b0 ;
  assign n26711 = n6998 & ~n11161 ;
  assign n26712 = ~n1903 & n26711 ;
  assign n26713 = n1124 & ~n18563 ;
  assign n26714 = n26713 ^ n2279 ^ 1'b0 ;
  assign n26715 = n8216 ^ n4579 ^ 1'b0 ;
  assign n26716 = ~n2730 & n26715 ;
  assign n26717 = n26716 ^ n7185 ^ n4525 ;
  assign n26718 = n6780 ^ n467 ^ 1'b0 ;
  assign n26719 = ( n7031 & n12233 ) | ( n7031 & n26718 ) | ( n12233 & n26718 ) ;
  assign n26720 = n3640 | n4883 ;
  assign n26721 = n26719 | n26720 ;
  assign n26722 = ~n369 & n26476 ;
  assign n26723 = n15540 | n17359 ;
  assign n26724 = n26723 ^ n14059 ^ n4222 ;
  assign n26725 = n14471 & ~n19551 ;
  assign n26726 = n3353 ^ n2900 ^ 1'b0 ;
  assign n26727 = n8291 & ~n26726 ;
  assign n26728 = ~n724 & n2250 ;
  assign n26729 = n26728 ^ n1023 ^ 1'b0 ;
  assign n26730 = n26729 ^ n20019 ^ 1'b0 ;
  assign n26731 = n26727 | n26730 ;
  assign n26732 = n672 | n26731 ;
  assign n26733 = n26732 ^ n7935 ^ 1'b0 ;
  assign n26734 = n992 | n14774 ;
  assign n26735 = n5248 | n26734 ;
  assign n26736 = n6202 & n9494 ;
  assign n26737 = n26736 ^ n16333 ^ 1'b0 ;
  assign n26738 = n5409 | n9324 ;
  assign n26739 = n10809 & ~n26738 ;
  assign n26740 = n22614 ^ n11728 ^ 1'b0 ;
  assign n26741 = n26740 ^ n16823 ^ 1'b0 ;
  assign n26742 = n2508 ^ n2078 ^ 1'b0 ;
  assign n26743 = ~n5156 & n12061 ;
  assign n26744 = n26742 & n26743 ;
  assign n26745 = n26744 ^ n14145 ^ 1'b0 ;
  assign n26746 = ~n25668 & n26745 ;
  assign n26747 = n26746 ^ n26639 ^ 1'b0 ;
  assign n26748 = n5407 & ~n26747 ;
  assign n26749 = n15798 | n26748 ;
  assign n26750 = n25297 ^ n11991 ^ n6106 ;
  assign n26756 = ~n12586 & n16403 ;
  assign n26757 = n26756 ^ n12074 ^ 1'b0 ;
  assign n26758 = n13908 ^ n12831 ^ n6599 ;
  assign n26759 = n26758 ^ n1481 ^ 1'b0 ;
  assign n26760 = ~n6220 & n26759 ;
  assign n26761 = n26760 ^ n23938 ^ 1'b0 ;
  assign n26762 = n26757 & ~n26761 ;
  assign n26751 = n26678 ^ n6452 ^ 1'b0 ;
  assign n26752 = ~n7386 & n26751 ;
  assign n26753 = n26752 ^ n5667 ^ 1'b0 ;
  assign n26754 = n14695 & ~n26753 ;
  assign n26755 = n10687 & n26754 ;
  assign n26763 = n26762 ^ n26755 ^ 1'b0 ;
  assign n26764 = ~n18392 & n19448 ;
  assign n26765 = n23068 & n26764 ;
  assign n26766 = n24319 ^ n20629 ^ 1'b0 ;
  assign n26767 = n19280 & n26766 ;
  assign n26768 = n8098 | n19006 ;
  assign n26769 = ~n17642 & n26768 ;
  assign n26770 = n26769 ^ n564 ^ 1'b0 ;
  assign n26771 = n17636 | n20503 ;
  assign n26772 = n26771 ^ n4554 ^ 1'b0 ;
  assign n26773 = n3683 & ~n26772 ;
  assign n26774 = n2755 | n14345 ;
  assign n26775 = n26774 ^ n5530 ^ 1'b0 ;
  assign n26776 = n4688 & n4881 ;
  assign n26777 = n20326 ^ n12239 ^ 1'b0 ;
  assign n26778 = n6576 & ~n26777 ;
  assign n26779 = n1570 | n11765 ;
  assign n26780 = n26779 ^ n23891 ^ n9216 ;
  assign n26781 = n6982 & n25708 ;
  assign n26782 = n4919 ^ n1111 ^ 1'b0 ;
  assign n26783 = n5840 | n8413 ;
  assign n26784 = n26783 ^ n8911 ^ 1'b0 ;
  assign n26785 = n26784 ^ n20141 ^ n5478 ;
  assign n26786 = n12863 ^ n11650 ^ 1'b0 ;
  assign n26787 = ( n1960 & ~n5471 ) | ( n1960 & n7964 ) | ( ~n5471 & n7964 ) ;
  assign n26788 = n26787 ^ n18096 ^ 1'b0 ;
  assign n26789 = ~n17517 & n26788 ;
  assign n26790 = n26789 ^ n3838 ^ 1'b0 ;
  assign n26791 = n1896 & n26790 ;
  assign n26792 = ~n518 & n26791 ;
  assign n26793 = n11072 & n25450 ;
  assign n26794 = ( ~n6151 & n8287 ) | ( ~n6151 & n24073 ) | ( n8287 & n24073 ) ;
  assign n26795 = ~n3114 & n6609 ;
  assign n26796 = ~n6609 & n26795 ;
  assign n26797 = ~n3582 & n26796 ;
  assign n26798 = n1098 & n26797 ;
  assign n26799 = n2564 & n26798 ;
  assign n26800 = ~n26794 & n26799 ;
  assign n26801 = n2929 & n17894 ;
  assign n26803 = n353 | n9334 ;
  assign n26804 = n26803 ^ n14912 ^ 1'b0 ;
  assign n26805 = n26804 ^ n15908 ^ 1'b0 ;
  assign n26806 = n5505 | n26805 ;
  assign n26802 = n14181 ^ n12491 ^ n10241 ;
  assign n26807 = n26806 ^ n26802 ^ 1'b0 ;
  assign n26808 = n26801 & n26807 ;
  assign n26812 = n4170 ^ n2343 ^ 1'b0 ;
  assign n26813 = n26812 ^ n15981 ^ 1'b0 ;
  assign n26809 = x179 & n2852 ;
  assign n26810 = ~n13198 & n26809 ;
  assign n26811 = n1153 & ~n26810 ;
  assign n26814 = n26813 ^ n26811 ^ 1'b0 ;
  assign n26815 = ~n2741 & n19736 ;
  assign n26816 = n6763 & n26815 ;
  assign n26817 = ~n17517 & n19656 ;
  assign n26819 = n19697 ^ n1619 ^ 1'b0 ;
  assign n26818 = n4066 ^ n564 ^ 1'b0 ;
  assign n26820 = n26819 ^ n26818 ^ n14911 ;
  assign n26821 = n15493 & n25857 ;
  assign n26822 = n26821 ^ n2590 ^ 1'b0 ;
  assign n26823 = n19886 | n26822 ;
  assign n26824 = n26823 ^ n4169 ^ 1'b0 ;
  assign n26825 = n9806 & ~n13584 ;
  assign n26826 = n11875 | n14342 ;
  assign n26827 = n26826 ^ n25680 ^ 1'b0 ;
  assign n26830 = ~n6615 & n10070 ;
  assign n26831 = n26830 ^ n1993 ^ 1'b0 ;
  assign n26828 = n11557 ^ n3926 ^ 1'b0 ;
  assign n26829 = n25598 & ~n26828 ;
  assign n26832 = n26831 ^ n26829 ^ 1'b0 ;
  assign n26833 = n7179 & n18532 ;
  assign n26834 = n3532 & n9411 ;
  assign n26835 = n26834 ^ n9922 ^ 1'b0 ;
  assign n26836 = n26833 | n26835 ;
  assign n26837 = n26836 ^ n11863 ^ n2945 ;
  assign n26838 = ( n4005 & ~n22252 ) | ( n4005 & n26837 ) | ( ~n22252 & n26837 ) ;
  assign n26839 = n25809 ^ n1180 ^ 1'b0 ;
  assign n26840 = n3684 & ~n26839 ;
  assign n26841 = n2830 & ~n3928 ;
  assign n26842 = n26841 ^ n24871 ^ 1'b0 ;
  assign n26843 = n1772 & ~n26842 ;
  assign n26844 = ~n997 & n1316 ;
  assign n26845 = n11253 | n16495 ;
  assign n26846 = n7855 & ~n26845 ;
  assign n26847 = n14202 ^ n625 ^ 1'b0 ;
  assign n26848 = ~n20770 & n26847 ;
  assign n26849 = n26848 ^ n22686 ^ 1'b0 ;
  assign n26851 = n18288 ^ n8804 ^ 1'b0 ;
  assign n26852 = n296 | n26851 ;
  assign n26850 = ~n8355 & n18891 ;
  assign n26853 = n26852 ^ n26850 ^ 1'b0 ;
  assign n26854 = n8733 & n12473 ;
  assign n26855 = n3055 & ~n5605 ;
  assign n26856 = n26855 ^ n22117 ^ 1'b0 ;
  assign n26857 = ~n2243 & n3887 ;
  assign n26858 = ~n6903 & n26857 ;
  assign n26859 = n24784 ^ n14661 ^ 1'b0 ;
  assign n26860 = ~n18169 & n26859 ;
  assign n26861 = n26858 & n26860 ;
  assign n26862 = n19085 ^ n12860 ^ 1'b0 ;
  assign n26863 = ~n10363 & n21029 ;
  assign n26864 = n9580 ^ n1958 ^ 1'b0 ;
  assign n26865 = n13071 & n26864 ;
  assign n26866 = ~n9740 & n26865 ;
  assign n26867 = n12754 ^ n4848 ^ 1'b0 ;
  assign n26868 = n6318 & ~n26867 ;
  assign n26869 = n9799 | n21965 ;
  assign n26870 = n26868 | n26869 ;
  assign n26871 = n10190 ^ n6367 ^ 1'b0 ;
  assign n26872 = n6950 & n26871 ;
  assign n26873 = ( n12375 & n13729 ) | ( n12375 & ~n23430 ) | ( n13729 & ~n23430 ) ;
  assign n26875 = n14708 & n16214 ;
  assign n26876 = n978 & n26875 ;
  assign n26874 = n6971 & n8580 ;
  assign n26877 = n26876 ^ n26874 ^ 1'b0 ;
  assign n26878 = n10336 & n10510 ;
  assign n26879 = n26878 ^ n1361 ^ 1'b0 ;
  assign n26880 = n12611 & n26879 ;
  assign n26881 = ~n3332 & n26880 ;
  assign n26882 = n26881 ^ n23382 ^ 1'b0 ;
  assign n26883 = n10133 | n26882 ;
  assign n26884 = n26056 ^ n24172 ^ 1'b0 ;
  assign n26885 = n9456 ^ n3823 ^ 1'b0 ;
  assign n26886 = ~n8508 & n15249 ;
  assign n26887 = n21688 & n26886 ;
  assign n26888 = n11554 & ~n25935 ;
  assign n26889 = n11374 & ~n13701 ;
  assign n26890 = n9746 & n26889 ;
  assign n26891 = n20220 ^ n830 ^ 1'b0 ;
  assign n26892 = n4417 & n26891 ;
  assign n26893 = n9753 ^ n6075 ^ n3928 ;
  assign n26894 = n23689 ^ n23205 ^ n3704 ;
  assign n26895 = n20244 ^ x196 ^ 1'b0 ;
  assign n26896 = n842 & ~n26895 ;
  assign n26897 = n2403 | n11592 ;
  assign n26898 = n16318 | n26897 ;
  assign n26899 = n8279 & n26898 ;
  assign n26900 = ~n26896 & n26899 ;
  assign n26901 = n2661 | n26900 ;
  assign n26902 = n5704 | n26901 ;
  assign n26903 = n5667 | n6395 ;
  assign n26904 = n7032 & n21050 ;
  assign n26905 = n26904 ^ n9540 ^ 1'b0 ;
  assign n26906 = n5695 & ~n9511 ;
  assign n26907 = n8978 ^ n4237 ^ 1'b0 ;
  assign n26908 = n26906 | n26907 ;
  assign n26909 = n15166 ^ n3435 ^ 1'b0 ;
  assign n26910 = n19540 ^ n17631 ^ n7674 ;
  assign n26911 = ~n4330 & n4603 ;
  assign n26912 = n11174 & n26911 ;
  assign n26913 = ~n4696 & n9237 ;
  assign n26914 = n4827 & n9288 ;
  assign n26915 = n26914 ^ n2679 ^ 1'b0 ;
  assign n26916 = n25908 ^ n16676 ^ n14207 ;
  assign n26917 = n8092 ^ n6182 ^ 1'b0 ;
  assign n26918 = n8604 & n26917 ;
  assign n26919 = ~n26916 & n26918 ;
  assign n26921 = n26585 ^ n13664 ^ 1'b0 ;
  assign n26922 = ~n6363 & n26921 ;
  assign n26920 = n8465 | n26858 ;
  assign n26923 = n26922 ^ n26920 ^ n4040 ;
  assign n26924 = n2146 & ~n2170 ;
  assign n26925 = n26924 ^ n10180 ^ 1'b0 ;
  assign n26926 = n26925 ^ n1137 ^ 1'b0 ;
  assign n26927 = x126 & ~n26926 ;
  assign n26928 = ~n26923 & n26927 ;
  assign n26929 = n8159 & ~n12070 ;
  assign n26930 = ~n13741 & n26929 ;
  assign n26931 = n19433 & ~n20853 ;
  assign n26932 = n26480 & n26931 ;
  assign n26933 = ~n26930 & n26932 ;
  assign n26935 = n3661 & ~n18081 ;
  assign n26934 = n7355 & ~n18259 ;
  assign n26936 = n26935 ^ n26934 ^ 1'b0 ;
  assign n26937 = n2472 & ~n15176 ;
  assign n26938 = ( n15090 & n18507 ) | ( n15090 & n19325 ) | ( n18507 & n19325 ) ;
  assign n26939 = ( n3160 & n17033 ) | ( n3160 & n21515 ) | ( n17033 & n21515 ) ;
  assign n26940 = n11290 | n12013 ;
  assign n26941 = n26940 ^ n17091 ^ 1'b0 ;
  assign n26942 = n22386 ^ n765 ^ 1'b0 ;
  assign n26943 = n987 & n24462 ;
  assign n26944 = ~n9526 & n26943 ;
  assign n26945 = n20405 ^ n16206 ^ 1'b0 ;
  assign n26946 = n3386 ^ n1220 ^ 1'b0 ;
  assign n26947 = n10276 & n26946 ;
  assign n26948 = n8546 & n14358 ;
  assign n26949 = n4442 & ~n5225 ;
  assign n26950 = n26949 ^ n9278 ^ 1'b0 ;
  assign n26951 = n1496 & n26950 ;
  assign n26952 = n14486 & n26951 ;
  assign n26953 = n4301 | n26952 ;
  assign n26954 = n9226 | n26953 ;
  assign n26955 = n20474 | n23893 ;
  assign n26956 = ( ~n18660 & n24615 ) | ( ~n18660 & n26955 ) | ( n24615 & n26955 ) ;
  assign n26957 = n10529 & n22857 ;
  assign n26958 = n13185 & n26957 ;
  assign n26959 = n2785 & n19784 ;
  assign n26960 = x212 ^ x154 ^ 1'b0 ;
  assign n26961 = n26959 | n26960 ;
  assign n26962 = n4589 & n16153 ;
  assign n26963 = n26962 ^ n16246 ^ 1'b0 ;
  assign n26964 = n16506 ^ n11659 ^ 1'b0 ;
  assign n26965 = n26964 ^ n3639 ^ 1'b0 ;
  assign n26966 = x107 | n7271 ;
  assign n26967 = n15091 ^ n6009 ^ 1'b0 ;
  assign n26968 = n15495 | n26967 ;
  assign n26969 = n4547 | n16595 ;
  assign n26970 = n12591 ^ n8627 ^ 1'b0 ;
  assign n26971 = n6159 & n26970 ;
  assign n26972 = ~n23883 & n26971 ;
  assign n26973 = ~n3790 & n10702 ;
  assign n26974 = n4300 & ~n8571 ;
  assign n26975 = ~n26973 & n26974 ;
  assign n26976 = n9352 & ~n26975 ;
  assign n26977 = n8722 & n26976 ;
  assign n26978 = n4204 | n18670 ;
  assign n26979 = x55 & ~n9091 ;
  assign n26980 = n7771 & n26979 ;
  assign n26981 = n26980 ^ n12554 ^ n585 ;
  assign n26982 = n13810 ^ n7056 ^ 1'b0 ;
  assign n26983 = n26982 ^ n13019 ^ 1'b0 ;
  assign n26984 = n11916 | n26983 ;
  assign n26985 = n20298 ^ n18391 ^ 1'b0 ;
  assign n26986 = ~n8233 & n26985 ;
  assign n26987 = n10920 & n26986 ;
  assign n26988 = ~n13546 & n19045 ;
  assign n26989 = n26988 ^ n9420 ^ 1'b0 ;
  assign n26990 = n26987 | n26989 ;
  assign n26991 = ~n4997 & n11586 ;
  assign n26992 = n26990 & n26991 ;
  assign n26994 = n2069 & n9070 ;
  assign n26995 = n26994 ^ n9695 ^ 1'b0 ;
  assign n26993 = ~n15153 & n19812 ;
  assign n26996 = n26995 ^ n26993 ^ 1'b0 ;
  assign n26997 = n19521 ^ n5962 ^ 1'b0 ;
  assign n26998 = n15744 & ~n15832 ;
  assign n26999 = n26998 ^ n8530 ^ 1'b0 ;
  assign n27000 = n830 & ~n3961 ;
  assign n27001 = n2085 | n17858 ;
  assign n27002 = n5110 & n14199 ;
  assign n27003 = n3133 & n9271 ;
  assign n27004 = ~n2730 & n3235 ;
  assign n27005 = ~n16396 & n27004 ;
  assign n27006 = ~n27003 & n27005 ;
  assign n27007 = n17609 ^ n6493 ^ n3023 ;
  assign n27008 = n1036 | n18563 ;
  assign n27009 = n16290 ^ n5426 ^ 1'b0 ;
  assign n27010 = n1494 & ~n27009 ;
  assign n27011 = n16926 | n27010 ;
  assign n27012 = n4919 & ~n15557 ;
  assign n27013 = n16061 ^ n11608 ^ 1'b0 ;
  assign n27014 = n2951 & n9886 ;
  assign n27015 = n27014 ^ n24061 ^ 1'b0 ;
  assign n27016 = n23854 & n25494 ;
  assign n27017 = x162 & n25094 ;
  assign n27018 = n27017 ^ n12332 ^ 1'b0 ;
  assign n27019 = n14371 & n14760 ;
  assign n27020 = n9705 ^ n2584 ^ 1'b0 ;
  assign n27021 = n4070 & ~n27020 ;
  assign n27022 = n27021 ^ n7493 ^ 1'b0 ;
  assign n27023 = n27022 ^ n4872 ^ 1'b0 ;
  assign n27024 = ~n27019 & n27023 ;
  assign n27025 = ~n15571 & n27024 ;
  assign n27026 = ~n6085 & n21602 ;
  assign n27027 = n3956 & n27026 ;
  assign n27028 = n3751 | n8033 ;
  assign n27029 = n2801 | n27028 ;
  assign n27030 = n27029 ^ n3999 ^ 1'b0 ;
  assign n27031 = n7976 & ~n11835 ;
  assign n27032 = ~n27030 & n27031 ;
  assign n27033 = n27032 ^ n2754 ^ 1'b0 ;
  assign n27034 = ( ~n6555 & n7810 ) | ( ~n6555 & n19038 ) | ( n7810 & n19038 ) ;
  assign n27035 = n27034 ^ n9573 ^ 1'b0 ;
  assign n27037 = n13177 ^ n10690 ^ 1'b0 ;
  assign n27038 = ~n9319 & n27037 ;
  assign n27036 = n18061 & ~n21861 ;
  assign n27039 = n27038 ^ n27036 ^ 1'b0 ;
  assign n27040 = n4706 & n10577 ;
  assign n27041 = ~n5340 & n27040 ;
  assign n27042 = n27041 ^ n9660 ^ 1'b0 ;
  assign n27043 = n7721 ^ n2202 ^ 1'b0 ;
  assign n27044 = n22910 ^ n12300 ^ 1'b0 ;
  assign n27045 = n11639 & n12247 ;
  assign n27046 = n21023 & n27045 ;
  assign n27047 = n3942 ^ n911 ^ 1'b0 ;
  assign n27048 = ~n5848 & n27047 ;
  assign n27049 = n14967 ^ n8861 ^ n3950 ;
  assign n27050 = n27048 & n27049 ;
  assign n27051 = n16379 | n17291 ;
  assign n27052 = n27051 ^ n20133 ^ 1'b0 ;
  assign n27053 = n6434 ^ n4547 ^ 1'b0 ;
  assign n27054 = n2426 & n5400 ;
  assign n27055 = n27054 ^ n8606 ^ 1'b0 ;
  assign n27056 = n3611 & n6149 ;
  assign n27057 = ( n18029 & ~n27055 ) | ( n18029 & n27056 ) | ( ~n27055 & n27056 ) ;
  assign n27058 = n11946 ^ n2116 ^ 1'b0 ;
  assign n27059 = n27058 ^ n25897 ^ 1'b0 ;
  assign n27060 = n15540 ^ n1898 ^ 1'b0 ;
  assign n27061 = n497 & ~n10452 ;
  assign n27062 = ( n7917 & n26768 ) | ( n7917 & ~n27061 ) | ( n26768 & ~n27061 ) ;
  assign n27063 = ( n7798 & n10350 ) | ( n7798 & n17861 ) | ( n10350 & n17861 ) ;
  assign n27064 = n22199 ^ n5954 ^ 1'b0 ;
  assign n27065 = n18727 ^ n9366 ^ 1'b0 ;
  assign n27066 = n16598 & n20308 ;
  assign n27067 = n27066 ^ n14752 ^ 1'b0 ;
  assign n27068 = n5130 | n21351 ;
  assign n27069 = ~n8450 & n21834 ;
  assign n27070 = n2396 & n27069 ;
  assign n27071 = n9700 ^ n3171 ^ 1'b0 ;
  assign n27072 = n27070 & n27071 ;
  assign n27073 = ~n5579 & n27072 ;
  assign n27074 = n3703 & n27073 ;
  assign n27075 = n11840 ^ n2477 ^ 1'b0 ;
  assign n27076 = n2925 & n16026 ;
  assign n27077 = n6199 | n27076 ;
  assign n27078 = n1766 & ~n27077 ;
  assign n27079 = n8018 | n27078 ;
  assign n27080 = ~n2165 & n18122 ;
  assign n27081 = n1221 & ~n19649 ;
  assign n27082 = n3677 & n27081 ;
  assign n27083 = n5864 & ~n8477 ;
  assign n27084 = n27083 ^ n24823 ^ 1'b0 ;
  assign n27085 = n26616 ^ n26508 ^ 1'b0 ;
  assign n27086 = ~n17054 & n27085 ;
  assign n27087 = n5891 & ~n14967 ;
  assign n27088 = n6495 & ~n20318 ;
  assign n27089 = n413 & n27088 ;
  assign n27090 = n20599 ^ n15668 ^ n3806 ;
  assign n27091 = ~n15285 & n19235 ;
  assign n27092 = n15076 ^ x196 ^ 1'b0 ;
  assign n27093 = n5498 & n23161 ;
  assign n27094 = n27093 ^ n13940 ^ 1'b0 ;
  assign n27095 = n15445 & ~n27094 ;
  assign n27096 = ( ~n4210 & n4914 ) | ( ~n4210 & n9713 ) | ( n4914 & n9713 ) ;
  assign n27097 = n10090 | n27096 ;
  assign n27098 = n11431 & ~n18841 ;
  assign n27099 = n27098 ^ n24981 ^ 1'b0 ;
  assign n27100 = n27099 ^ n11908 ^ 1'b0 ;
  assign n27101 = ( n4350 & n13513 ) | ( n4350 & ~n27100 ) | ( n13513 & ~n27100 ) ;
  assign n27102 = n13450 ^ n3293 ^ 1'b0 ;
  assign n27103 = n27102 ^ n2790 ^ n2649 ;
  assign n27104 = n20224 ^ n4287 ^ 1'b0 ;
  assign n27105 = n12318 & n15101 ;
  assign n27106 = n26119 & n27105 ;
  assign n27107 = n2319 & n4773 ;
  assign n27108 = ~n13779 & n27107 ;
  assign n27109 = n11636 ^ n2916 ^ 1'b0 ;
  assign n27110 = ~n3286 & n22718 ;
  assign n27111 = n4725 ^ x175 ^ 1'b0 ;
  assign n27112 = n716 | n27111 ;
  assign n27113 = ~n3461 & n21834 ;
  assign n27114 = n27112 & n27113 ;
  assign n27115 = n27114 ^ n20210 ^ 1'b0 ;
  assign n27116 = n15620 ^ n8466 ^ 1'b0 ;
  assign n27117 = n17864 & n27116 ;
  assign n27118 = n27117 ^ n15296 ^ 1'b0 ;
  assign n27122 = n11680 ^ n1964 ^ 1'b0 ;
  assign n27123 = ( n511 & ~n5456 ) | ( n511 & n27122 ) | ( ~n5456 & n27122 ) ;
  assign n27119 = ~n3217 & n8373 ;
  assign n27120 = ( x200 & ~n13954 ) | ( x200 & n27119 ) | ( ~n13954 & n27119 ) ;
  assign n27121 = ~n9496 & n27120 ;
  assign n27124 = n27123 ^ n27121 ^ 1'b0 ;
  assign n27125 = n13790 | n27124 ;
  assign n27126 = n16291 ^ n11314 ^ 1'b0 ;
  assign n27127 = x40 & n15809 ;
  assign n27128 = ~n15119 & n16674 ;
  assign n27129 = n22235 ^ n15654 ^ 1'b0 ;
  assign n27130 = n27128 & ~n27129 ;
  assign n27131 = n858 & ~n3432 ;
  assign n27132 = n27131 ^ n26911 ^ n22452 ;
  assign n27133 = n1251 | n23594 ;
  assign n27134 = n13725 ^ n9289 ^ 1'b0 ;
  assign n27135 = ~n1694 & n27134 ;
  assign n27136 = n27135 ^ n2316 ^ 1'b0 ;
  assign n27137 = n27133 & ~n27136 ;
  assign n27138 = n7132 & n11358 ;
  assign n27139 = n7646 & n16758 ;
  assign n27140 = ~n10817 & n27139 ;
  assign n27141 = n2666 | n27140 ;
  assign n27142 = n1534 | n1966 ;
  assign n27143 = ~n5525 & n9976 ;
  assign n27144 = n27143 ^ n17898 ^ 1'b0 ;
  assign n27145 = ~n1653 & n13301 ;
  assign n27146 = n6149 ^ n1490 ^ 1'b0 ;
  assign n27147 = n27146 ^ n12379 ^ 1'b0 ;
  assign n27148 = ~n1853 & n3613 ;
  assign n27149 = n3993 & n8224 ;
  assign n27150 = n27149 ^ n5797 ^ 1'b0 ;
  assign n27151 = n27150 ^ n21246 ^ 1'b0 ;
  assign n27152 = n27151 ^ n14847 ^ 1'b0 ;
  assign n27153 = n17938 | n27152 ;
  assign n27154 = n18693 ^ n3572 ^ 1'b0 ;
  assign n27155 = ~n7880 & n27154 ;
  assign n27156 = ~n5602 & n14457 ;
  assign n27157 = n27156 ^ n4498 ^ 1'b0 ;
  assign n27158 = ( n5851 & n18028 ) | ( n5851 & ~n27157 ) | ( n18028 & ~n27157 ) ;
  assign n27165 = n9788 ^ n2484 ^ n2110 ;
  assign n27166 = n27165 ^ n7581 ^ 1'b0 ;
  assign n27161 = n6157 ^ n2148 ^ 1'b0 ;
  assign n27162 = ~n10807 & n27161 ;
  assign n27163 = n27162 ^ n24071 ^ 1'b0 ;
  assign n27164 = n4542 | n27163 ;
  assign n27167 = n27166 ^ n27164 ^ n11435 ;
  assign n27159 = n5517 | n7893 ;
  assign n27160 = n20056 | n27159 ;
  assign n27168 = n27167 ^ n27160 ^ 1'b0 ;
  assign n27169 = n5581 | n15496 ;
  assign n27170 = n9976 ^ n5454 ^ 1'b0 ;
  assign n27171 = n7467 ^ x46 ^ 1'b0 ;
  assign n27172 = n15429 & ~n27171 ;
  assign n27173 = n5065 & ~n8966 ;
  assign n27174 = n11938 ^ n4481 ^ 1'b0 ;
  assign n27175 = n11291 & n27174 ;
  assign n27176 = n8322 & ~n17382 ;
  assign n27177 = n27176 ^ n4994 ^ 1'b0 ;
  assign n27178 = n5614 | n23148 ;
  assign n27179 = n19102 & ~n27178 ;
  assign n27180 = n27179 ^ n5293 ^ 1'b0 ;
  assign n27181 = n11699 ^ n9627 ^ 1'b0 ;
  assign n27182 = ~n8434 & n12264 ;
  assign n27183 = n23959 ^ n21068 ^ 1'b0 ;
  assign n27184 = n14562 | n27183 ;
  assign n27185 = n21863 ^ n2037 ^ 1'b0 ;
  assign n27186 = n10264 | n27185 ;
  assign n27187 = ( n880 & ~n8970 ) | ( n880 & n22084 ) | ( ~n8970 & n22084 ) ;
  assign n27188 = n327 | n11943 ;
  assign n27189 = n7596 & n27188 ;
  assign n27190 = n27189 ^ n1909 ^ 1'b0 ;
  assign n27191 = n23957 ^ n13862 ^ n7874 ;
  assign n27192 = n26352 ^ n5561 ^ 1'b0 ;
  assign n27193 = n21538 ^ n9463 ^ 1'b0 ;
  assign n27194 = n13610 & ~n27193 ;
  assign n27195 = n5307 & n13228 ;
  assign n27196 = n22619 ^ n6880 ^ 1'b0 ;
  assign n27197 = n7571 | n27196 ;
  assign n27198 = n27197 ^ n11433 ^ 1'b0 ;
  assign n27199 = n13774 & ~n27198 ;
  assign n27200 = ~n1914 & n3706 ;
  assign n27201 = ( n2335 & n13258 ) | ( n2335 & n18904 ) | ( n13258 & n18904 ) ;
  assign n27202 = ~n27200 & n27201 ;
  assign n27203 = n27202 ^ n18506 ^ 1'b0 ;
  assign n27204 = n21660 ^ n15472 ^ n1815 ;
  assign n27206 = n11229 & ~n12162 ;
  assign n27207 = n18178 & n27206 ;
  assign n27208 = n27207 ^ n4605 ^ 1'b0 ;
  assign n27205 = n671 & ~n17399 ;
  assign n27209 = n27208 ^ n27205 ^ 1'b0 ;
  assign n27210 = n22715 ^ n13406 ^ 1'b0 ;
  assign n27211 = n7165 | n27210 ;
  assign n27212 = n27211 ^ x93 ^ 1'b0 ;
  assign n27213 = n21262 & ~n27212 ;
  assign n27214 = n19488 | n25151 ;
  assign n27215 = n1172 | n9916 ;
  assign n27216 = n4036 | n27215 ;
  assign n27217 = n18296 ^ n5918 ^ 1'b0 ;
  assign n27218 = ~n4553 & n9525 ;
  assign n27219 = n27218 ^ n473 ^ 1'b0 ;
  assign n27220 = n8195 & ~n27219 ;
  assign n27221 = n27220 ^ n18315 ^ 1'b0 ;
  assign n27222 = n24644 & ~n27221 ;
  assign n27223 = n15577 ^ n13671 ^ 1'b0 ;
  assign n27224 = n3934 ^ x181 ^ 1'b0 ;
  assign n27225 = ( n6525 & n11684 ) | ( n6525 & n23177 ) | ( n11684 & n23177 ) ;
  assign n27226 = n19361 ^ n11981 ^ 1'b0 ;
  assign n27227 = n10982 ^ n6581 ^ 1'b0 ;
  assign n27228 = n22663 ^ n20174 ^ 1'b0 ;
  assign n27229 = n13051 & n27228 ;
  assign n27230 = n12878 ^ n908 ^ 1'b0 ;
  assign n27231 = n9016 & n27230 ;
  assign n27232 = ~n19940 & n27231 ;
  assign n27233 = n8030 ^ n2158 ^ 1'b0 ;
  assign n27234 = n5031 | n27233 ;
  assign n27235 = n27234 ^ n12953 ^ 1'b0 ;
  assign n27237 = n3577 & ~n7948 ;
  assign n27238 = ~n6896 & n27237 ;
  assign n27236 = ~n3351 & n10336 ;
  assign n27239 = n27238 ^ n27236 ^ 1'b0 ;
  assign n27240 = n9800 ^ n4964 ^ 1'b0 ;
  assign n27241 = n900 & n5190 ;
  assign n27242 = n27241 ^ n2199 ^ 1'b0 ;
  assign n27243 = ~n1736 & n27242 ;
  assign n27244 = n6983 | n11282 ;
  assign n27245 = n27243 & ~n27244 ;
  assign n27246 = n22824 ^ n11026 ^ 1'b0 ;
  assign n27247 = n8242 & ~n23285 ;
  assign n27248 = n27247 ^ n18776 ^ 1'b0 ;
  assign n27249 = n8079 ^ n6139 ^ 1'b0 ;
  assign n27250 = n4319 | n6348 ;
  assign n27251 = n27249 | n27250 ;
  assign n27255 = n2321 & n22572 ;
  assign n27254 = n7027 & n9724 ;
  assign n27256 = n27255 ^ n27254 ^ 1'b0 ;
  assign n27252 = n6477 ^ n4225 ^ 1'b0 ;
  assign n27253 = n3673 | n27252 ;
  assign n27257 = n27256 ^ n27253 ^ n5509 ;
  assign n27258 = n3892 | n15151 ;
  assign n27259 = n4123 & n9262 ;
  assign n27260 = n5671 ^ n5346 ^ 1'b0 ;
  assign n27261 = n4966 & n27260 ;
  assign n27262 = n8945 & ~n12939 ;
  assign n27263 = n27262 ^ n522 ^ 1'b0 ;
  assign n27264 = ( n9292 & ~n27261 ) | ( n9292 & n27263 ) | ( ~n27261 & n27263 ) ;
  assign n27265 = n13660 | n27264 ;
  assign n27266 = n23784 | n27265 ;
  assign n27267 = n6534 | n9285 ;
  assign n27268 = n6006 | n18801 ;
  assign n27269 = n4737 ^ n1466 ^ 1'b0 ;
  assign n27270 = n5847 | n27269 ;
  assign n27271 = n16820 ^ n6805 ^ 1'b0 ;
  assign n27272 = n6531 & ~n8700 ;
  assign n27273 = n27272 ^ n8771 ^ 1'b0 ;
  assign n27274 = ( n7089 & ~n12778 ) | ( n7089 & n21745 ) | ( ~n12778 & n21745 ) ;
  assign n27275 = n27274 ^ n5476 ^ 1'b0 ;
  assign n27276 = n8802 ^ n8246 ^ 1'b0 ;
  assign n27277 = ~n20752 & n27276 ;
  assign n27278 = n27277 ^ n17303 ^ 1'b0 ;
  assign n27279 = x105 & ~n26204 ;
  assign n27280 = n26738 ^ n9692 ^ n5604 ;
  assign n27281 = n27280 ^ n15741 ^ 1'b0 ;
  assign n27282 = n22667 ^ n3307 ^ n1453 ;
  assign n27283 = n25394 ^ n10381 ^ 1'b0 ;
  assign n27284 = ~n2911 & n27283 ;
  assign n27285 = n27284 ^ n16768 ^ 1'b0 ;
  assign n27286 = ~n15209 & n24491 ;
  assign n27287 = n7745 & n27286 ;
  assign n27288 = n12727 | n25829 ;
  assign n27289 = n27288 ^ n15104 ^ 1'b0 ;
  assign n27290 = n12787 ^ n8070 ^ 1'b0 ;
  assign n27291 = n7866 & n27290 ;
  assign n27292 = ~n7932 & n27291 ;
  assign n27293 = n13759 ^ n5398 ^ 1'b0 ;
  assign n27294 = ~n8678 & n16887 ;
  assign n27295 = ~n8302 & n27294 ;
  assign n27296 = n25584 ^ n16982 ^ 1'b0 ;
  assign n27297 = ~n3542 & n22041 ;
  assign n27298 = n2745 | n9753 ;
  assign n27299 = n4567 & n18385 ;
  assign n27300 = n27299 ^ n2061 ^ 1'b0 ;
  assign n27301 = n5587 ^ n1543 ^ 1'b0 ;
  assign n27302 = n27301 ^ n16502 ^ 1'b0 ;
  assign n27303 = ( n20648 & n27300 ) | ( n20648 & ~n27302 ) | ( n27300 & ~n27302 ) ;
  assign n27304 = n27303 ^ n14637 ^ 1'b0 ;
  assign n27305 = ~n1473 & n27304 ;
  assign n27306 = n27305 ^ n13398 ^ 1'b0 ;
  assign n27307 = n10499 ^ n4714 ^ n274 ;
  assign n27308 = n12649 & ~n27307 ;
  assign n27309 = n19022 ^ n274 ^ 1'b0 ;
  assign n27310 = ~n11081 & n27309 ;
  assign n27311 = ~n26357 & n27310 ;
  assign n27312 = ~n1505 & n2086 ;
  assign n27313 = n26327 & ~n27312 ;
  assign n27314 = n27313 ^ n8510 ^ 1'b0 ;
  assign n27315 = n27314 ^ n5988 ^ 1'b0 ;
  assign n27316 = n2706 ^ n2172 ^ 1'b0 ;
  assign n27317 = n27316 ^ n7549 ^ 1'b0 ;
  assign n27318 = n27317 ^ n22584 ^ 1'b0 ;
  assign n27319 = n10554 ^ n500 ^ 1'b0 ;
  assign n27323 = ~x143 & n6342 ;
  assign n27324 = n4042 & n27323 ;
  assign n27320 = ~n3393 & n14553 ;
  assign n27321 = n27320 ^ n17561 ^ 1'b0 ;
  assign n27322 = n4425 & ~n27321 ;
  assign n27325 = n27324 ^ n27322 ^ 1'b0 ;
  assign n27326 = n6739 & ~n14781 ;
  assign n27327 = n27326 ^ n3915 ^ 1'b0 ;
  assign n27328 = n7493 | n25680 ;
  assign n27329 = n27327 | n27328 ;
  assign n27330 = n27329 ^ n2549 ^ 1'b0 ;
  assign n27331 = n6506 ^ n2799 ^ 1'b0 ;
  assign n27332 = n3666 | n27331 ;
  assign n27333 = ~n4970 & n27332 ;
  assign n27334 = n16193 ^ n4585 ^ 1'b0 ;
  assign n27335 = ~n18543 & n27334 ;
  assign n27336 = ~n4096 & n27335 ;
  assign n27337 = n27336 ^ n19736 ^ 1'b0 ;
  assign n27338 = n16861 & n24160 ;
  assign n27339 = n1019 ^ n888 ^ 1'b0 ;
  assign n27340 = n25296 | n27339 ;
  assign n27341 = n19699 ^ n7769 ^ 1'b0 ;
  assign n27342 = n13370 & n27341 ;
  assign n27343 = ~n1197 & n27342 ;
  assign n27344 = n2472 & ~n4123 ;
  assign n27345 = n27343 & n27344 ;
  assign n27346 = n14765 ^ n9123 ^ 1'b0 ;
  assign n27347 = n8349 & ~n27346 ;
  assign n27348 = n27347 ^ n1232 ^ 1'b0 ;
  assign n27349 = ~n9540 & n18041 ;
  assign n27350 = n15491 ^ n12603 ^ n7279 ;
  assign n27351 = n17364 & ~n27350 ;
  assign n27352 = n21503 ^ n2830 ^ 1'b0 ;
  assign n27353 = n16527 ^ n14605 ^ 1'b0 ;
  assign n27354 = n27302 & n27353 ;
  assign n27355 = n27354 ^ n10501 ^ 1'b0 ;
  assign n27356 = ~n688 & n19046 ;
  assign n27357 = ~n19046 & n27356 ;
  assign n27358 = n1453 & ~n9267 ;
  assign n27359 = n9267 & n27358 ;
  assign n27360 = n5625 & n27359 ;
  assign n27361 = x91 & ~n11901 ;
  assign n27362 = n27361 ^ n9622 ^ 1'b0 ;
  assign n27363 = n27362 ^ n2101 ^ 1'b0 ;
  assign n27364 = ~n3932 & n27363 ;
  assign n27365 = n27360 & n27364 ;
  assign n27366 = n27365 ^ n17081 ^ 1'b0 ;
  assign n27367 = ~n27357 & n27366 ;
  assign n27372 = ( n2191 & ~n8192 ) | ( n2191 & n12870 ) | ( ~n8192 & n12870 ) ;
  assign n27369 = ~n6834 & n19045 ;
  assign n27370 = n27369 ^ n13789 ^ 1'b0 ;
  assign n27371 = n1231 & ~n27370 ;
  assign n27373 = n27372 ^ n27371 ^ 1'b0 ;
  assign n27374 = n13871 | n27373 ;
  assign n27375 = n27374 ^ n21546 ^ 1'b0 ;
  assign n27368 = ~n8190 & n12636 ;
  assign n27376 = n27375 ^ n27368 ^ 1'b0 ;
  assign n27377 = n26744 ^ n1577 ^ 1'b0 ;
  assign n27378 = ~n4593 & n27377 ;
  assign n27379 = n5322 & ~n22518 ;
  assign n27380 = n27379 ^ n2083 ^ 1'b0 ;
  assign n27381 = n7382 ^ n6789 ^ 1'b0 ;
  assign n27382 = n19634 | n27381 ;
  assign n27383 = n18551 | n27382 ;
  assign n27384 = ~n24678 & n25334 ;
  assign n27385 = n27384 ^ n16352 ^ 1'b0 ;
  assign n27386 = ~n9075 & n27385 ;
  assign n27387 = n21490 ^ n12078 ^ 1'b0 ;
  assign n27388 = ~n15555 & n24691 ;
  assign n27389 = n27388 ^ n1680 ^ 1'b0 ;
  assign n27390 = ~n27387 & n27389 ;
  assign n27391 = n1426 & n17911 ;
  assign n27392 = n1377 & n8722 ;
  assign n27394 = n8473 ^ n7061 ^ 1'b0 ;
  assign n27395 = ~n9024 & n27394 ;
  assign n27393 = n13624 ^ n9944 ^ 1'b0 ;
  assign n27396 = n27395 ^ n27393 ^ 1'b0 ;
  assign n27397 = ~n3837 & n26609 ;
  assign n27398 = n8957 | n13672 ;
  assign n27399 = n27397 & ~n27398 ;
  assign n27400 = ~n7053 & n21262 ;
  assign n27402 = n15802 ^ n9571 ^ 1'b0 ;
  assign n27401 = n14306 | n15889 ;
  assign n27403 = n27402 ^ n27401 ^ 1'b0 ;
  assign n27407 = n713 & n6679 ;
  assign n27408 = n13472 & n27407 ;
  assign n27409 = ~n9821 & n27408 ;
  assign n27404 = n8217 ^ n4520 ^ 1'b0 ;
  assign n27405 = x151 & ~n27404 ;
  assign n27406 = x221 & n27405 ;
  assign n27410 = n27409 ^ n27406 ^ n14109 ;
  assign n27411 = ~n3234 & n22442 ;
  assign n27412 = n10763 | n22957 ;
  assign n27413 = n27412 ^ n17114 ^ 1'b0 ;
  assign n27414 = ~n13048 & n14155 ;
  assign n27415 = n27414 ^ n13468 ^ 1'b0 ;
  assign n27419 = ~n3357 & n5476 ;
  assign n27420 = n27419 ^ n12953 ^ 1'b0 ;
  assign n27421 = n7275 & ~n18062 ;
  assign n27422 = ~n27420 & n27421 ;
  assign n27423 = n1903 & n10062 ;
  assign n27424 = n27423 ^ n2394 ^ 1'b0 ;
  assign n27425 = n27422 | n27424 ;
  assign n27416 = x109 | n14908 ;
  assign n27417 = n15387 | n15925 ;
  assign n27418 = n27416 & ~n27417 ;
  assign n27426 = n27425 ^ n27418 ^ 1'b0 ;
  assign n27427 = n12627 ^ n12603 ^ 1'b0 ;
  assign n27428 = n27427 ^ n20081 ^ 1'b0 ;
  assign n27429 = ~n27426 & n27428 ;
  assign n27430 = n11138 ^ n7676 ^ 1'b0 ;
  assign n27432 = n2223 | n7994 ;
  assign n27433 = n27432 ^ n2176 ^ 1'b0 ;
  assign n27431 = n3801 ^ n2559 ^ 1'b0 ;
  assign n27434 = n27433 ^ n27431 ^ n23111 ;
  assign n27435 = n8733 & n27434 ;
  assign n27436 = n4099 & n27435 ;
  assign n27438 = n477 | n19516 ;
  assign n27437 = n11367 & ~n20668 ;
  assign n27439 = n27438 ^ n27437 ^ 1'b0 ;
  assign n27440 = n12259 | n27439 ;
  assign n27441 = n13555 ^ n812 ^ 1'b0 ;
  assign n27442 = ~n7644 & n7966 ;
  assign n27443 = n935 & n27442 ;
  assign n27444 = n27443 ^ n3592 ^ 1'b0 ;
  assign n27445 = n6253 & n27444 ;
  assign n27446 = n9821 & ~n27445 ;
  assign n27447 = n10497 & n11344 ;
  assign n27448 = n13951 & n27447 ;
  assign n27449 = n14065 ^ n9742 ^ 1'b0 ;
  assign n27450 = ~n1545 & n4315 ;
  assign n27451 = n27449 & n27450 ;
  assign n27452 = n840 & n1822 ;
  assign n27453 = n13242 & ~n27452 ;
  assign n27454 = n27453 ^ n8816 ^ 1'b0 ;
  assign n27455 = ~n27451 & n27454 ;
  assign n27456 = n3928 & n27455 ;
  assign n27457 = n27456 ^ n19645 ^ 1'b0 ;
  assign n27458 = n1992 | n7000 ;
  assign n27459 = n3385 | n20238 ;
  assign n27460 = n22922 ^ n7587 ^ 1'b0 ;
  assign n27461 = n1494 & n27460 ;
  assign n27462 = n6402 ^ n4642 ^ 1'b0 ;
  assign n27463 = n8663 & n27462 ;
  assign n27464 = ~n4203 & n27463 ;
  assign n27465 = n1244 ^ n1125 ^ 1'b0 ;
  assign n27466 = n1344 & n27465 ;
  assign n27467 = ~n17960 & n20761 ;
  assign n27468 = n27467 ^ n7323 ^ 1'b0 ;
  assign n27472 = n19885 ^ x242 ^ 1'b0 ;
  assign n27469 = n3411 ^ n389 ^ 1'b0 ;
  assign n27470 = n10079 & ~n27469 ;
  assign n27471 = n18194 | n27470 ;
  assign n27473 = n27472 ^ n27471 ^ 1'b0 ;
  assign n27474 = n3222 ^ n2509 ^ x3 ;
  assign n27475 = n1841 & n27474 ;
  assign n27476 = n665 | n27475 ;
  assign n27477 = ~n755 & n12306 ;
  assign n27478 = ~n11450 & n27477 ;
  assign n27479 = n26195 ^ n19287 ^ n17548 ;
  assign n27480 = n20794 ^ n14711 ^ 1'b0 ;
  assign n27481 = n13610 & n27480 ;
  assign n27482 = n26787 & n27481 ;
  assign n27483 = n4730 & ~n22173 ;
  assign n27484 = n27483 ^ n18631 ^ 1'b0 ;
  assign n27485 = n5825 & ~n27484 ;
  assign n27486 = ~n5498 & n27485 ;
  assign n27487 = ~n6533 & n20330 ;
  assign n27488 = ~n12787 & n27487 ;
  assign n27489 = n5075 ^ n5036 ^ 1'b0 ;
  assign n27490 = n25980 | n27489 ;
  assign n27491 = ~n2072 & n2141 ;
  assign n27492 = n27491 ^ n8463 ^ 1'b0 ;
  assign n27493 = ~n10978 & n27492 ;
  assign n27494 = ~n16579 & n27493 ;
  assign n27495 = x251 & ~n27494 ;
  assign n27496 = n16803 & n27495 ;
  assign n27497 = n22739 ^ n3694 ^ 1'b0 ;
  assign n27498 = n13861 ^ n12356 ^ n11799 ;
  assign n27499 = n27498 ^ n26412 ^ n8523 ;
  assign n27500 = n20990 ^ n13292 ^ n6326 ;
  assign n27501 = n1634 & ~n22905 ;
  assign n27502 = n27501 ^ n4732 ^ 1'b0 ;
  assign n27503 = n9518 & ~n19986 ;
  assign n27504 = n4637 & n11164 ;
  assign n27505 = n4008 & n27504 ;
  assign n27506 = ~n432 & n3435 ;
  assign n27507 = n25657 ^ n20071 ^ 1'b0 ;
  assign n27508 = n8722 & ~n8832 ;
  assign n27509 = ( ~n276 & n8911 ) | ( ~n276 & n8921 ) | ( n8911 & n8921 ) ;
  assign n27510 = n27509 ^ n6269 ^ n1807 ;
  assign n27511 = n1699 | n2165 ;
  assign n27512 = n10731 ^ n6106 ^ 1'b0 ;
  assign n27513 = n13816 | n27512 ;
  assign n27514 = n20902 ^ n10733 ^ 1'b0 ;
  assign n27515 = n3041 | n6943 ;
  assign n27516 = n22316 | n27515 ;
  assign n27517 = n15028 ^ n11437 ^ 1'b0 ;
  assign n27518 = n20056 | n27517 ;
  assign n27519 = n21460 & ~n27518 ;
  assign n27520 = ( n1223 & ~n4846 ) | ( n1223 & n18053 ) | ( ~n4846 & n18053 ) ;
  assign n27521 = n1112 & n5815 ;
  assign n27522 = ~n17386 & n27521 ;
  assign n27523 = n6916 & ~n27522 ;
  assign n27524 = n25442 & ~n25660 ;
  assign n27525 = n13463 ^ n9428 ^ 1'b0 ;
  assign n27526 = n26379 & ~n27525 ;
  assign n27527 = n5051 ^ n1940 ^ 1'b0 ;
  assign n27528 = n3629 & ~n27527 ;
  assign n27529 = n9705 & ~n27528 ;
  assign n27530 = n27529 ^ n16044 ^ 1'b0 ;
  assign n27531 = n14562 & n23037 ;
  assign n27532 = ~n27530 & n27531 ;
  assign n27533 = n8620 | n19128 ;
  assign n27534 = n27533 ^ n23297 ^ 1'b0 ;
  assign n27535 = n26192 ^ n2069 ^ 1'b0 ;
  assign n27536 = n4562 | n10046 ;
  assign n27537 = n27536 ^ x231 ^ 1'b0 ;
  assign n27538 = n27537 ^ n7359 ^ 1'b0 ;
  assign n27539 = n16674 ^ n2013 ^ 1'b0 ;
  assign n27540 = n27539 ^ x31 ^ 1'b0 ;
  assign n27541 = n23852 & ~n27540 ;
  assign n27542 = ( ~n9670 & n16463 ) | ( ~n9670 & n27541 ) | ( n16463 & n27541 ) ;
  assign n27543 = n11320 ^ n2870 ^ 1'b0 ;
  assign n27544 = ~n2825 & n5626 ;
  assign n27545 = n27544 ^ n19158 ^ 1'b0 ;
  assign n27546 = n22551 ^ n5089 ^ n2076 ;
  assign n27547 = n13777 | n27546 ;
  assign n27548 = n27489 ^ n19952 ^ n4383 ;
  assign n27555 = n23012 ^ n16777 ^ 1'b0 ;
  assign n27556 = n11055 & ~n27555 ;
  assign n27549 = ~n2067 & n12275 ;
  assign n27550 = n1221 & n27549 ;
  assign n27551 = ~n27549 & n27550 ;
  assign n27552 = ~n5050 & n27551 ;
  assign n27553 = n15945 & ~n27552 ;
  assign n27554 = n15305 & ~n27553 ;
  assign n27557 = n27556 ^ n27554 ^ 1'b0 ;
  assign n27558 = ~n23369 & n25374 ;
  assign n27563 = ~n7120 & n18544 ;
  assign n27564 = n27563 ^ n15503 ^ 1'b0 ;
  assign n27559 = n1782 & n22743 ;
  assign n27560 = n20916 ^ n17456 ^ 1'b0 ;
  assign n27561 = x195 | n27560 ;
  assign n27562 = n27559 | n27561 ;
  assign n27565 = n27564 ^ n27562 ^ 1'b0 ;
  assign n27566 = n5416 & n13829 ;
  assign n27567 = n1961 & n27566 ;
  assign n27568 = n2502 | n4807 ;
  assign n27569 = n3157 | n27568 ;
  assign n27570 = n15633 & n27569 ;
  assign n27571 = n27570 ^ n8888 ^ 1'b0 ;
  assign n27572 = n24190 & n27571 ;
  assign n27573 = n4174 & ~n5725 ;
  assign n27574 = n7676 & n27573 ;
  assign n27575 = n14383 ^ n11494 ^ 1'b0 ;
  assign n27576 = n3344 | n27575 ;
  assign n27577 = n27576 ^ n8668 ^ 1'b0 ;
  assign n27578 = n2646 & ~n22313 ;
  assign n27579 = ~n4645 & n14363 ;
  assign n27580 = n27579 ^ n4694 ^ 1'b0 ;
  assign n27581 = ~n17161 & n27580 ;
  assign n27582 = n1611 & ~n27581 ;
  assign n27585 = n679 | n1193 ;
  assign n27586 = n679 & ~n27585 ;
  assign n27587 = x115 & ~n27586 ;
  assign n27583 = n2146 & ~n5546 ;
  assign n27584 = n5546 & n27583 ;
  assign n27588 = n27587 ^ n27584 ^ 1'b0 ;
  assign n27589 = n27588 ^ n6900 ^ 1'b0 ;
  assign n27590 = n5719 | n27589 ;
  assign n27591 = n13632 ^ n9210 ^ 1'b0 ;
  assign n27592 = n3645 ^ n765 ^ 1'b0 ;
  assign n27593 = n6745 & ~n25805 ;
  assign n27594 = n17258 ^ n3879 ^ 1'b0 ;
  assign n27595 = n27594 ^ n12514 ^ 1'b0 ;
  assign n27596 = n27120 ^ n8774 ^ 1'b0 ;
  assign n27597 = ~n15069 & n27596 ;
  assign n27598 = n8265 | n22718 ;
  assign n27599 = n14752 & ~n17552 ;
  assign n27600 = n16468 & ~n17448 ;
  assign n27601 = n3377 ^ n2058 ^ 1'b0 ;
  assign n27602 = n4348 | n27601 ;
  assign n27603 = n12746 & n27602 ;
  assign n27604 = ~n1695 & n6780 ;
  assign n27605 = n710 & ~n2835 ;
  assign n27606 = n27604 & n27605 ;
  assign n27607 = n5939 & ~n27606 ;
  assign n27608 = ~n16947 & n27607 ;
  assign n27609 = n27608 ^ n3755 ^ 1'b0 ;
  assign n27610 = n27603 | n27609 ;
  assign n27611 = n3974 & ~n15125 ;
  assign n27612 = n16061 & n27611 ;
  assign n27613 = ( n5243 & n6387 ) | ( n5243 & ~n15899 ) | ( n6387 & ~n15899 ) ;
  assign n27614 = ~n16615 & n27613 ;
  assign n27615 = n27614 ^ n22581 ^ 1'b0 ;
  assign n27616 = n27615 ^ n15316 ^ 1'b0 ;
  assign n27617 = n11941 & ~n27616 ;
  assign n27618 = n27612 & n27617 ;
  assign n27619 = ( ~n1696 & n15343 ) | ( ~n1696 & n22810 ) | ( n15343 & n22810 ) ;
  assign n27620 = n27619 ^ n4122 ^ 1'b0 ;
  assign n27621 = n12095 ^ n4771 ^ 1'b0 ;
  assign n27622 = n14823 ^ n7269 ^ 1'b0 ;
  assign n27623 = n2622 & n27622 ;
  assign n27624 = n16403 ^ n12630 ^ n4011 ;
  assign n27625 = n23022 ^ n2950 ^ 1'b0 ;
  assign n27626 = n13164 & n14843 ;
  assign n27627 = ~n13725 & n27626 ;
  assign n27628 = n16801 & n19535 ;
  assign n27629 = n10776 & n27628 ;
  assign n27630 = n27629 ^ n21786 ^ 1'b0 ;
  assign n27631 = n2722 & ~n2951 ;
  assign n27632 = n27631 ^ n3195 ^ 1'b0 ;
  assign n27634 = n6110 & ~n7966 ;
  assign n27633 = ~n12891 & n17867 ;
  assign n27635 = n27634 ^ n27633 ^ 1'b0 ;
  assign n27636 = n8276 ^ n7188 ^ x152 ;
  assign n27637 = n3432 | n15688 ;
  assign n27638 = ~n27636 & n27637 ;
  assign n27639 = n10516 ^ n6157 ^ n961 ;
  assign n27640 = n7617 ^ n2082 ^ 1'b0 ;
  assign n27641 = n27640 ^ n10559 ^ 1'b0 ;
  assign n27642 = n27639 | n27641 ;
  assign n27643 = n18246 ^ n13867 ^ 1'b0 ;
  assign n27644 = n12249 & n27643 ;
  assign n27647 = n4511 | n18210 ;
  assign n27648 = n13629 & ~n27647 ;
  assign n27645 = n4512 & n11342 ;
  assign n27646 = n7932 & n27645 ;
  assign n27649 = n27648 ^ n27646 ^ 1'b0 ;
  assign n27650 = n17010 & ~n21845 ;
  assign n27651 = n27649 & n27650 ;
  assign n27652 = n27651 ^ n1353 ^ 1'b0 ;
  assign n27653 = n24646 ^ n9006 ^ 1'b0 ;
  assign n27654 = n2400 & ~n27653 ;
  assign n27655 = n12041 & ~n27654 ;
  assign n27656 = n4899 & ~n26406 ;
  assign n27657 = n27656 ^ n15347 ^ 1'b0 ;
  assign n27658 = n12085 ^ n6674 ^ 1'b0 ;
  assign n27660 = n11891 & n15577 ;
  assign n27659 = ~n4848 & n5695 ;
  assign n27661 = n27660 ^ n27659 ^ 1'b0 ;
  assign n27662 = n12812 | n24920 ;
  assign n27663 = n27662 ^ n27197 ^ n16943 ;
  assign n27664 = n20267 | n27663 ;
  assign n27665 = ~n12162 & n27648 ;
  assign n27666 = n27665 ^ n2983 ^ 1'b0 ;
  assign n27667 = n27666 ^ n5255 ^ 1'b0 ;
  assign n27668 = n4026 & ~n9241 ;
  assign n27669 = ~n705 & n2172 ;
  assign n27670 = ~n2172 & n27669 ;
  assign n27671 = ~n24941 & n27670 ;
  assign n27672 = n3465 & n24691 ;
  assign n27673 = ~n4856 & n11355 ;
  assign n27674 = n14410 | n27673 ;
  assign n27675 = n27674 ^ n12298 ^ 1'b0 ;
  assign n27676 = n9110 | n27675 ;
  assign n27677 = n27672 & ~n27676 ;
  assign n27678 = n6454 ^ n3616 ^ 1'b0 ;
  assign n27679 = n11586 & n27678 ;
  assign n27680 = n27679 ^ n20108 ^ 1'b0 ;
  assign n27681 = n26378 ^ n328 ^ 1'b0 ;
  assign n27682 = n10648 & n27681 ;
  assign n27683 = n15814 ^ n395 ^ 1'b0 ;
  assign n27684 = n27682 & n27683 ;
  assign n27689 = n16545 ^ n836 ^ 1'b0 ;
  assign n27686 = n6166 & ~n8074 ;
  assign n27687 = n14521 & n27686 ;
  assign n27688 = n6655 | n27687 ;
  assign n27690 = n27689 ^ n27688 ^ 1'b0 ;
  assign n27685 = n11030 | n11665 ;
  assign n27691 = n27690 ^ n27685 ^ 1'b0 ;
  assign n27692 = n27691 ^ n8677 ^ 1'b0 ;
  assign n27693 = ~n13364 & n27692 ;
  assign n27694 = ~n5596 & n27693 ;
  assign n27695 = n26787 ^ n14756 ^ n3705 ;
  assign n27696 = n27695 ^ n26591 ^ n11871 ;
  assign n27697 = ~n5727 & n12096 ;
  assign n27698 = n27697 ^ n409 ^ 1'b0 ;
  assign n27699 = n27698 ^ n25960 ^ n8568 ;
  assign n27700 = n22888 ^ n14412 ^ 1'b0 ;
  assign n27701 = n5944 & n27700 ;
  assign n27702 = n27701 ^ n4146 ^ 1'b0 ;
  assign n27703 = n27699 & n27702 ;
  assign n27704 = n12930 | n27397 ;
  assign n27705 = n27704 ^ n23681 ^ 1'b0 ;
  assign n27706 = ~n9442 & n11941 ;
  assign n27707 = n27706 ^ n740 ^ 1'b0 ;
  assign n27708 = n27707 ^ n7963 ^ x159 ;
  assign n27709 = n11230 | n15738 ;
  assign n27710 = n27709 ^ n23833 ^ 1'b0 ;
  assign n27711 = n27708 & n27710 ;
  assign n27712 = n12112 ^ n8607 ^ n571 ;
  assign n27713 = n25682 & n27712 ;
  assign n27714 = n3190 ^ n2823 ^ 1'b0 ;
  assign n27715 = n3951 & n27714 ;
  assign n27716 = n1153 & n5401 ;
  assign n27717 = n27715 | n27716 ;
  assign n27718 = n17900 ^ n6873 ^ 1'b0 ;
  assign n27719 = n5455 & ~n7195 ;
  assign n27720 = n9391 ^ n6701 ^ 1'b0 ;
  assign n27721 = n19797 & n27720 ;
  assign n27722 = n7031 & n27721 ;
  assign n27723 = n27719 & n27722 ;
  assign n27724 = n6923 & ~n12138 ;
  assign n27725 = n27723 & n27724 ;
  assign n27726 = ~n12355 & n17073 ;
  assign n27727 = n14529 ^ n12148 ^ 1'b0 ;
  assign n27728 = ~n18766 & n27727 ;
  assign n27729 = n3588 | n18082 ;
  assign n27730 = n26407 ^ n6053 ^ 1'b0 ;
  assign n27731 = n8391 & ~n27730 ;
  assign n27732 = ~n2076 & n27731 ;
  assign n27733 = n3256 | n21899 ;
  assign n27734 = n27733 ^ n4855 ^ 1'b0 ;
  assign n27735 = n12614 ^ n5840 ^ 1'b0 ;
  assign n27736 = n4968 & ~n20168 ;
  assign n27737 = n10017 ^ n6394 ^ 1'b0 ;
  assign n27738 = n27737 ^ n9798 ^ 1'b0 ;
  assign n27739 = n3627 | n6274 ;
  assign n27740 = n24572 ^ n4090 ^ 1'b0 ;
  assign n27741 = n27739 | n27740 ;
  assign n27742 = n6788 ^ x198 ^ 1'b0 ;
  assign n27743 = n6398 & ~n27742 ;
  assign n27744 = ( ~n520 & n11067 ) | ( ~n520 & n27743 ) | ( n11067 & n27743 ) ;
  assign n27745 = n23983 ^ n17521 ^ 1'b0 ;
  assign n27746 = ~n8874 & n27745 ;
  assign n27755 = n4988 ^ n4128 ^ n2310 ;
  assign n27752 = n4343 & ~n6365 ;
  assign n27753 = n27752 ^ n3610 ^ 1'b0 ;
  assign n27754 = n16377 & ~n27753 ;
  assign n27756 = n27755 ^ n27754 ^ 1'b0 ;
  assign n27757 = ~n5893 & n27756 ;
  assign n27747 = n4123 ^ x118 ^ 1'b0 ;
  assign n27748 = ~n5018 & n27747 ;
  assign n27749 = n23560 & n27748 ;
  assign n27750 = n27749 ^ n1982 ^ 1'b0 ;
  assign n27751 = n12648 & n27750 ;
  assign n27758 = n27757 ^ n27751 ^ 1'b0 ;
  assign n27759 = n6252 ^ n905 ^ 1'b0 ;
  assign n27760 = n16390 | n27759 ;
  assign n27761 = n20826 & ~n23280 ;
  assign n27763 = ( n8763 & n9839 ) | ( n8763 & ~n11665 ) | ( n9839 & ~n11665 ) ;
  assign n27762 = n8278 & n18723 ;
  assign n27764 = n27763 ^ n27762 ^ 1'b0 ;
  assign n27765 = ~n4348 & n19830 ;
  assign n27766 = n27765 ^ x169 ^ 1'b0 ;
  assign n27767 = n27766 ^ n11541 ^ 1'b0 ;
  assign n27768 = n9007 & n27767 ;
  assign n27769 = n3099 & ~n8933 ;
  assign n27770 = ~n3099 & n27769 ;
  assign n27771 = n27770 ^ n14533 ^ 1'b0 ;
  assign n27772 = n4518 | n9385 ;
  assign n27773 = n4518 & ~n27772 ;
  assign n27774 = n27771 | n27773 ;
  assign n27775 = n1346 | n27774 ;
  assign n27776 = n27775 ^ n16679 ^ 1'b0 ;
  assign n27777 = n27768 & n27776 ;
  assign n27778 = n13839 | n14963 ;
  assign n27779 = n2331 | n27778 ;
  assign n27780 = n20006 & ~n22001 ;
  assign n27781 = ~n6284 & n8442 ;
  assign n27782 = n27781 ^ x173 ^ 1'b0 ;
  assign n27783 = n27782 ^ n1219 ^ 1'b0 ;
  assign n27784 = n4260 & n27783 ;
  assign n27785 = n12712 ^ n4784 ^ 1'b0 ;
  assign n27786 = ( n8009 & n25957 ) | ( n8009 & ~n27785 ) | ( n25957 & ~n27785 ) ;
  assign n27787 = n12611 ^ x151 ^ 1'b0 ;
  assign n27788 = n3400 ^ n2926 ^ 1'b0 ;
  assign n27789 = n2491 | n27788 ;
  assign n27790 = n1254 & n7800 ;
  assign n27791 = ( n1274 & n3966 ) | ( n1274 & ~n9728 ) | ( n3966 & ~n9728 ) ;
  assign n27792 = n27791 ^ n2595 ^ 1'b0 ;
  assign n27793 = n12006 & ~n17155 ;
  assign n27794 = n27793 ^ n14311 ^ 1'b0 ;
  assign n27795 = n27794 ^ n12133 ^ n6900 ;
  assign n27796 = n21748 ^ n1643 ^ 1'b0 ;
  assign n27797 = n27796 ^ n10616 ^ 1'b0 ;
  assign n27798 = n15178 ^ n4345 ^ 1'b0 ;
  assign n27799 = n3666 & ~n7120 ;
  assign n27800 = n1948 & n27799 ;
  assign n27801 = ~n11607 & n13131 ;
  assign n27802 = n27801 ^ n18493 ^ 1'b0 ;
  assign n27803 = n27800 | n27802 ;
  assign n27804 = n10467 ^ n6171 ^ 1'b0 ;
  assign n27805 = n4331 & ~n27804 ;
  assign n27806 = n14253 ^ n8632 ^ 1'b0 ;
  assign n27807 = n5871 ^ n2651 ^ n2496 ;
  assign n27808 = n7742 ^ n1086 ^ 1'b0 ;
  assign n27809 = n27808 ^ n3936 ^ n1262 ;
  assign n27810 = ~n4023 & n23156 ;
  assign n27811 = n27809 & n27810 ;
  assign n27812 = n19373 | n27811 ;
  assign n27813 = n15783 & ~n27812 ;
  assign n27814 = n20341 | n27813 ;
  assign n27815 = n27814 ^ x227 ^ 1'b0 ;
  assign n27816 = n6349 & ~n10041 ;
  assign n27817 = n11868 ^ n10474 ^ 1'b0 ;
  assign n27818 = n27816 & n27817 ;
  assign n27819 = n27818 ^ n15107 ^ 1'b0 ;
  assign n27820 = ~n12556 & n24658 ;
  assign n27821 = n27172 & n27820 ;
  assign n27822 = n27821 ^ n23128 ^ 1'b0 ;
  assign n27823 = n20868 ^ x104 ^ 1'b0 ;
  assign n27824 = n11367 & ~n27823 ;
  assign n27825 = n5619 | n10270 ;
  assign n27826 = n7739 | n27825 ;
  assign n27827 = n12501 & n27826 ;
  assign n27828 = ~n7961 & n8463 ;
  assign n27829 = ( n22297 & ~n26334 ) | ( n22297 & n27828 ) | ( ~n26334 & n27828 ) ;
  assign n27831 = n5951 | n6415 ;
  assign n27832 = n27831 ^ n24332 ^ 1'b0 ;
  assign n27830 = n8535 & ~n13085 ;
  assign n27833 = n27832 ^ n27830 ^ 1'b0 ;
  assign n27834 = n17965 ^ n2441 ^ x112 ;
  assign n27835 = n5076 & ~n10694 ;
  assign n27836 = ~n27834 & n27835 ;
  assign n27837 = n10363 ^ n1138 ^ 1'b0 ;
  assign n27838 = n15930 & ~n27837 ;
  assign n27839 = n17239 | n27838 ;
  assign n27841 = n12009 ^ n8391 ^ 1'b0 ;
  assign n27842 = n11116 & n27841 ;
  assign n27843 = ( n8751 & ~n12074 ) | ( n8751 & n27842 ) | ( ~n12074 & n27842 ) ;
  assign n27840 = n2216 | n15402 ;
  assign n27844 = n27843 ^ n27840 ^ 1'b0 ;
  assign n27845 = n27844 ^ n15405 ^ n2443 ;
  assign n27846 = n15481 ^ n14696 ^ 1'b0 ;
  assign n27847 = n27846 ^ n2812 ^ 1'b0 ;
  assign n27848 = n564 | n23099 ;
  assign n27849 = n9735 ^ n1730 ^ 1'b0 ;
  assign n27850 = ~n2719 & n17886 ;
  assign n27851 = n15608 & n27850 ;
  assign n27852 = n8415 ^ n5621 ^ 1'b0 ;
  assign n27853 = n5282 & n27852 ;
  assign n27854 = ~n7419 & n27853 ;
  assign n27855 = n2122 | n27719 ;
  assign n27856 = n25310 | n27855 ;
  assign n27857 = n27856 ^ n26466 ^ 1'b0 ;
  assign n27858 = ~n20783 & n27857 ;
  assign n27859 = n7107 & n11951 ;
  assign n27860 = n1701 & n27859 ;
  assign n27861 = n27860 ^ n5001 ^ 1'b0 ;
  assign n27862 = n1667 & n2998 ;
  assign n27863 = n21492 ^ n5458 ^ n3644 ;
  assign n27864 = n12468 & ~n18145 ;
  assign n27865 = n9735 ^ n8914 ^ n5392 ;
  assign n27866 = n20389 ^ n13355 ^ 1'b0 ;
  assign n27867 = n15713 ^ n2358 ^ 1'b0 ;
  assign n27868 = n27866 | n27867 ;
  assign n27869 = ~n13197 & n17254 ;
  assign n27874 = n4898 & ~n5758 ;
  assign n27875 = n27874 ^ n13828 ^ 1'b0 ;
  assign n27876 = n15779 & n27875 ;
  assign n27870 = n15636 ^ n10122 ^ n8201 ;
  assign n27871 = n27870 ^ n4921 ^ 1'b0 ;
  assign n27872 = n27871 ^ n2274 ^ 1'b0 ;
  assign n27873 = n8578 | n27872 ;
  assign n27877 = n27876 ^ n27873 ^ 1'b0 ;
  assign n27878 = n5917 & ~n20921 ;
  assign n27879 = n27878 ^ n19381 ^ 1'b0 ;
  assign n27881 = ~n5990 & n8112 ;
  assign n27882 = n27881 ^ n8880 ^ 1'b0 ;
  assign n27880 = n7930 & ~n27484 ;
  assign n27883 = n27882 ^ n27880 ^ 1'b0 ;
  assign n27884 = n20136 ^ n8444 ^ 1'b0 ;
  assign n27885 = n22596 | n27884 ;
  assign n27886 = n267 & n2481 ;
  assign n27887 = n13894 & n27886 ;
  assign n27888 = n2191 & n6464 ;
  assign n27889 = n27888 ^ n3539 ^ 1'b0 ;
  assign n27890 = n27739 ^ n11541 ^ 1'b0 ;
  assign n27891 = n27889 & n27890 ;
  assign n27892 = ~n1593 & n1680 ;
  assign n27893 = n27892 ^ n387 ^ 1'b0 ;
  assign n27894 = n2850 | n27893 ;
  assign n27895 = n25769 | n27894 ;
  assign n27896 = n2951 & ~n17443 ;
  assign n27897 = ~n27895 & n27896 ;
  assign n27898 = n11430 | n14505 ;
  assign n27899 = n13219 & ~n19785 ;
  assign n27900 = n27899 ^ n6553 ^ 1'b0 ;
  assign n27901 = ~n12383 & n27900 ;
  assign n27902 = n16106 & n27901 ;
  assign n27903 = n27898 & n27902 ;
  assign n27904 = n22024 | n27903 ;
  assign n27905 = n27904 ^ n3014 ^ 1'b0 ;
  assign n27906 = n22627 ^ n4076 ^ 1'b0 ;
  assign n27907 = n3942 & ~n27906 ;
  assign n27908 = n10918 & ~n15798 ;
  assign n27909 = n27908 ^ n14843 ^ 1'b0 ;
  assign n27910 = n7223 | n9603 ;
  assign n27911 = n27910 ^ n9456 ^ 1'b0 ;
  assign n27912 = n11655 & n27911 ;
  assign n27913 = n27912 ^ n19210 ^ 1'b0 ;
  assign n27914 = n8475 & n25259 ;
  assign n27915 = n9161 ^ n393 ^ 1'b0 ;
  assign n27916 = ~n3957 & n10339 ;
  assign n27917 = n9642 & ~n13604 ;
  assign n27918 = n14359 & n27917 ;
  assign n27919 = ~n16980 & n19026 ;
  assign n27920 = ~n5163 & n10044 ;
  assign n27921 = ~n17333 & n27920 ;
  assign n27922 = n19515 ^ n9423 ^ 1'b0 ;
  assign n27923 = n4733 ^ x72 ^ 1'b0 ;
  assign n27924 = ~n25512 & n27923 ;
  assign n27925 = n10996 & n27318 ;
  assign n27926 = n11323 & n15133 ;
  assign n27927 = n16983 & ~n27926 ;
  assign n27928 = x244 & ~n1458 ;
  assign n27929 = n27928 ^ n1439 ^ 1'b0 ;
  assign n27930 = n27929 ^ n2385 ^ 1'b0 ;
  assign n27931 = n8375 | n27930 ;
  assign n27932 = n1342 | n27931 ;
  assign n27933 = n14666 | n27932 ;
  assign n27934 = ~n12155 & n27933 ;
  assign n27935 = ~n27335 & n27934 ;
  assign n27936 = n16567 ^ n10907 ^ n10834 ;
  assign n27937 = ( n3407 & n9824 ) | ( n3407 & ~n27936 ) | ( n9824 & ~n27936 ) ;
  assign n27938 = ~n1593 & n8671 ;
  assign n27939 = n6582 & ~n27938 ;
  assign n27940 = n14622 & n27939 ;
  assign n27941 = n24502 ^ n19185 ^ 1'b0 ;
  assign n27942 = n13480 & n27941 ;
  assign n27943 = n27942 ^ n8337 ^ 1'b0 ;
  assign n27944 = n3931 & n27943 ;
  assign n27945 = ( ~n16003 & n27940 ) | ( ~n16003 & n27944 ) | ( n27940 & n27944 ) ;
  assign n27946 = n11147 ^ n6853 ^ 1'b0 ;
  assign n27947 = n5539 ^ n2528 ^ 1'b0 ;
  assign n27948 = n11137 & ~n12884 ;
  assign n27949 = n27948 ^ n15122 ^ 1'b0 ;
  assign n27950 = n17708 & n27949 ;
  assign n27951 = n27950 ^ n1536 ^ 1'b0 ;
  assign n27952 = ~x233 & n4714 ;
  assign n27953 = n8822 ^ n2022 ^ 1'b0 ;
  assign n27954 = n5134 & ~n24811 ;
  assign n27955 = n27954 ^ n20616 ^ 1'b0 ;
  assign n27956 = ~n23516 & n27955 ;
  assign n27957 = n13631 ^ n6749 ^ 1'b0 ;
  assign n27958 = ~n10988 & n27957 ;
  assign n27959 = n1760 & n27958 ;
  assign n27960 = n27959 ^ n8012 ^ 1'b0 ;
  assign n27961 = n4259 & n11271 ;
  assign n27962 = n27961 ^ n1474 ^ 1'b0 ;
  assign n27963 = ~n2223 & n27962 ;
  assign n27964 = n2223 & n27963 ;
  assign n27965 = n21658 & ~n27964 ;
  assign n27966 = n27965 ^ n9461 ^ 1'b0 ;
  assign n27967 = n20552 ^ n18904 ^ 1'b0 ;
  assign n27970 = n13626 & n23891 ;
  assign n27971 = n27970 ^ n24062 ^ n7511 ;
  assign n27968 = n1589 ^ n742 ^ 1'b0 ;
  assign n27969 = n2765 | n27968 ;
  assign n27972 = n27971 ^ n27969 ^ 1'b0 ;
  assign n27973 = n496 | n6877 ;
  assign n27974 = n27973 ^ n16753 ^ 1'b0 ;
  assign n27975 = n12161 & ~n13802 ;
  assign n27976 = ~n4827 & n27975 ;
  assign n27977 = n747 & n1869 ;
  assign n27978 = n1138 | n18794 ;
  assign n27979 = n6789 & ~n27978 ;
  assign n27980 = n1389 & ~n12765 ;
  assign n27981 = ~n27979 & n27980 ;
  assign n27983 = n9912 & ~n17773 ;
  assign n27984 = n2567 & n27983 ;
  assign n27982 = n5583 | n23348 ;
  assign n27985 = n27984 ^ n27982 ^ 1'b0 ;
  assign n27986 = n26825 | n27985 ;
  assign n27987 = n1223 | n15069 ;
  assign n27988 = ~n9132 & n16820 ;
  assign n27989 = n5363 ^ n1340 ^ 1'b0 ;
  assign n27990 = ~n2881 & n9549 ;
  assign n27991 = n1048 & n27990 ;
  assign n27992 = n3600 | n23022 ;
  assign n27993 = n12573 & ~n27992 ;
  assign n27994 = n2015 & n7467 ;
  assign n27995 = n27994 ^ n2688 ^ 1'b0 ;
  assign n27996 = n15549 ^ n12911 ^ x192 ;
  assign n27997 = n27996 ^ n1358 ^ 1'b0 ;
  assign n27998 = n27995 & n27997 ;
  assign n27999 = ~n611 & n1901 ;
  assign n28000 = n14048 | n18292 ;
  assign n28001 = n18535 ^ n1402 ^ 1'b0 ;
  assign n28002 = n407 | n28001 ;
  assign n28003 = ~n14546 & n20201 ;
  assign n28004 = n8311 & n28003 ;
  assign n28005 = n28004 ^ n2355 ^ 1'b0 ;
  assign n28006 = n9479 ^ n850 ^ 1'b0 ;
  assign n28007 = n3281 & ~n11398 ;
  assign n28008 = x14 | n2785 ;
  assign n28009 = ( n1799 & ~n4869 ) | ( n1799 & n7447 ) | ( ~n4869 & n7447 ) ;
  assign n28010 = n28009 ^ n19337 ^ 1'b0 ;
  assign n28011 = n6274 | n28010 ;
  assign n28012 = n1876 ^ n1328 ^ 1'b0 ;
  assign n28013 = n15301 ^ n10356 ^ n3567 ;
  assign n28014 = n6846 & n28013 ;
  assign n28015 = n4394 | n9329 ;
  assign n28016 = ~n13734 & n15622 ;
  assign n28017 = ~n4911 & n28016 ;
  assign n28018 = ~n17619 & n18059 ;
  assign n28019 = n28017 & n28018 ;
  assign n28020 = n24633 ^ n9362 ^ 1'b0 ;
  assign n28021 = ~n1317 & n9290 ;
  assign n28023 = ~n1770 & n13000 ;
  assign n28024 = n28023 ^ n17368 ^ 1'b0 ;
  assign n28022 = n1798 & ~n5338 ;
  assign n28025 = n28024 ^ n28022 ^ 1'b0 ;
  assign n28026 = n2936 & ~n16934 ;
  assign n28027 = n28026 ^ n19370 ^ 1'b0 ;
  assign n28028 = n7839 & n15389 ;
  assign n28036 = n1676 & n4286 ;
  assign n28029 = n2113 ^ n840 ^ 1'b0 ;
  assign n28030 = ~n18067 & n28029 ;
  assign n28031 = n14479 ^ n7810 ^ 1'b0 ;
  assign n28032 = n28030 & n28031 ;
  assign n28033 = n28032 ^ n11767 ^ n267 ;
  assign n28034 = n2504 & n28033 ;
  assign n28035 = n28034 ^ n23213 ^ 1'b0 ;
  assign n28037 = n28036 ^ n28035 ^ n1382 ;
  assign n28038 = n24625 ^ n12826 ^ 1'b0 ;
  assign n28039 = n4141 & n28038 ;
  assign n28040 = n10200 & ~n12681 ;
  assign n28041 = ~n26238 & n28040 ;
  assign n28042 = n1879 & ~n3736 ;
  assign n28043 = ~n8715 & n28042 ;
  assign n28044 = n28043 ^ n21109 ^ 1'b0 ;
  assign n28045 = n28041 | n28044 ;
  assign n28046 = n5937 & n10805 ;
  assign n28047 = ~n6429 & n28046 ;
  assign n28048 = n274 | n10157 ;
  assign n28049 = n28047 & ~n28048 ;
  assign n28050 = n28049 ^ n4009 ^ 1'b0 ;
  assign n28051 = x214 & ~n28050 ;
  assign n28052 = n17815 ^ n15343 ^ 1'b0 ;
  assign n28053 = n5532 & n28052 ;
  assign n28054 = n28053 ^ n3279 ^ 1'b0 ;
  assign n28055 = n3021 | n23019 ;
  assign n28056 = n11049 & ~n14967 ;
  assign n28057 = n14760 & n28056 ;
  assign n28058 = n28055 & n28057 ;
  assign n28059 = n28058 ^ n15492 ^ n10031 ;
  assign n28060 = n22113 ^ n18096 ^ n6533 ;
  assign n28061 = n28060 ^ n1447 ^ 1'b0 ;
  assign n28062 = n12628 | n28061 ;
  assign n28063 = n28062 ^ n10798 ^ 1'b0 ;
  assign n28064 = n12771 & n28063 ;
  assign n28065 = n9296 & n9911 ;
  assign n28067 = n5667 & n9237 ;
  assign n28066 = n14345 & ~n16728 ;
  assign n28068 = n28067 ^ n28066 ^ 1'b0 ;
  assign n28069 = n28068 ^ n22526 ^ 1'b0 ;
  assign n28070 = n13424 & n28069 ;
  assign n28071 = n13776 ^ n2924 ^ 1'b0 ;
  assign n28072 = n913 | n23779 ;
  assign n28073 = ~n28071 & n28072 ;
  assign n28074 = n28073 ^ n14249 ^ 1'b0 ;
  assign n28075 = n351 & ~n28074 ;
  assign n28076 = n28075 ^ n26828 ^ 1'b0 ;
  assign n28077 = n10111 & n14892 ;
  assign n28078 = n2868 & n28077 ;
  assign n28079 = n28078 ^ n6469 ^ 1'b0 ;
  assign n28080 = n794 & ~n28079 ;
  assign n28081 = n15999 ^ n3513 ^ 1'b0 ;
  assign n28082 = n13160 & ~n13573 ;
  assign n28083 = n5459 & ~n15131 ;
  assign n28084 = n28083 ^ n8072 ^ 1'b0 ;
  assign n28085 = n4937 & n28084 ;
  assign n28086 = ~n3542 & n28085 ;
  assign n28087 = n11589 | n28086 ;
  assign n28088 = n28087 ^ n260 ^ 1'b0 ;
  assign n28089 = n28088 ^ n20813 ^ 1'b0 ;
  assign n28092 = ~n3078 & n13390 ;
  assign n28093 = ~x30 & n28092 ;
  assign n28094 = n11901 ^ n8868 ^ 1'b0 ;
  assign n28095 = n28093 | n28094 ;
  assign n28096 = ( ~n928 & n21168 ) | ( ~n928 & n28095 ) | ( n21168 & n28095 ) ;
  assign n28090 = n1075 | n1413 ;
  assign n28091 = n11593 | n28090 ;
  assign n28097 = n28096 ^ n28091 ^ 1'b0 ;
  assign n28098 = ~n4568 & n7210 ;
  assign n28099 = ~n20096 & n28098 ;
  assign n28100 = ~n1177 & n12771 ;
  assign n28101 = n28100 ^ n3546 ^ 1'b0 ;
  assign n28102 = n19734 & ~n23547 ;
  assign n28103 = n28101 & n28102 ;
  assign n28104 = n13573 ^ n615 ^ 1'b0 ;
  assign n28105 = n2625 & n28104 ;
  assign n28106 = n6141 ^ n1841 ^ 1'b0 ;
  assign n28107 = n10988 ^ n2746 ^ 1'b0 ;
  assign n28108 = n10246 & ~n28107 ;
  assign n28109 = n17311 & n28108 ;
  assign n28110 = n25245 ^ n2142 ^ 1'b0 ;
  assign n28111 = n20829 | n25618 ;
  assign n28112 = n7462 | n28111 ;
  assign n28113 = ~n23607 & n28112 ;
  assign n28114 = n9009 & n28113 ;
  assign n28115 = n3131 & ~n5895 ;
  assign n28116 = n11127 & ~n28115 ;
  assign n28117 = n8501 | n16304 ;
  assign n28118 = n8916 & ~n28117 ;
  assign n28119 = n1851 | n12532 ;
  assign n28120 = n10279 | n28119 ;
  assign n28123 = n7223 & n17911 ;
  assign n28124 = ~n10988 & n11168 ;
  assign n28125 = n28123 & n28124 ;
  assign n28121 = x174 & n6782 ;
  assign n28122 = ~n8844 & n28121 ;
  assign n28126 = n28125 ^ n28122 ^ 1'b0 ;
  assign n28127 = n9967 & n13370 ;
  assign n28128 = n22784 | n27003 ;
  assign n28129 = n23255 | n28128 ;
  assign n28130 = ( ~n9268 & n15719 ) | ( ~n9268 & n28129 ) | ( n15719 & n28129 ) ;
  assign n28131 = n11951 ^ n9744 ^ 1'b0 ;
  assign n28132 = ~n27200 & n28131 ;
  assign n28133 = n4125 & n7241 ;
  assign n28134 = n5799 & n28133 ;
  assign n28135 = n23326 ^ n15946 ^ n7141 ;
  assign n28136 = n28135 ^ n25168 ^ 1'b0 ;
  assign n28138 = n2460 | n5608 ;
  assign n28137 = n10766 ^ n10241 ^ n4632 ;
  assign n28139 = n28138 ^ n28137 ^ 1'b0 ;
  assign n28140 = n15690 & ~n28139 ;
  assign n28141 = n10372 | n17695 ;
  assign n28142 = n28141 ^ n5879 ^ 1'b0 ;
  assign n28144 = n7099 & ~n11414 ;
  assign n28145 = ~n7099 & n28144 ;
  assign n28143 = n6429 & n12497 ;
  assign n28146 = n28145 ^ n28143 ^ 1'b0 ;
  assign n28147 = n28142 | n28146 ;
  assign n28148 = ~n14053 & n21701 ;
  assign n28149 = n27535 | n28148 ;
  assign n28150 = n14464 ^ n14350 ^ 1'b0 ;
  assign n28151 = n3823 & n28150 ;
  assign n28152 = n10264 ^ n5089 ^ n675 ;
  assign n28153 = n13912 ^ n4222 ^ 1'b0 ;
  assign n28154 = n4682 & ~n14247 ;
  assign n28155 = n13122 & n28154 ;
  assign n28156 = n21942 & ~n26634 ;
  assign n28157 = n19699 & n28156 ;
  assign n28158 = ( n3178 & n17012 ) | ( n3178 & ~n20688 ) | ( n17012 & ~n20688 ) ;
  assign n28159 = n6688 & ~n18133 ;
  assign n28160 = n1593 & n28159 ;
  assign n28161 = n6248 | n28160 ;
  assign n28162 = n15193 ^ n2297 ^ 1'b0 ;
  assign n28163 = ~n287 & n11040 ;
  assign n28164 = n28163 ^ n21261 ^ 1'b0 ;
  assign n28165 = ( n22201 & n28162 ) | ( n22201 & n28164 ) | ( n28162 & n28164 ) ;
  assign n28166 = n21484 & n28165 ;
  assign n28167 = n28166 ^ n6264 ^ 1'b0 ;
  assign n28168 = n5924 & n8165 ;
  assign n28169 = n22442 & ~n28168 ;
  assign n28170 = ~x45 & n28169 ;
  assign n28171 = n22570 | n28170 ;
  assign n28172 = x188 & ~n2121 ;
  assign n28173 = n28172 ^ x188 ^ 1'b0 ;
  assign n28174 = n17148 ^ n500 ^ 1'b0 ;
  assign n28175 = n1960 | n8630 ;
  assign n28176 = ~n8211 & n28175 ;
  assign n28177 = n12231 & ~n28176 ;
  assign n28178 = n1258 & n28177 ;
  assign n28179 = n3530 & n11276 ;
  assign n28180 = ~n12971 & n28179 ;
  assign n28181 = n28180 ^ n11609 ^ n7863 ;
  assign n28182 = n6318 ^ n5479 ^ 1'b0 ;
  assign n28183 = n13978 & n28182 ;
  assign n28184 = ~n10043 & n28183 ;
  assign n28185 = n28184 ^ n6817 ^ 1'b0 ;
  assign n28186 = n17809 ^ n6134 ^ 1'b0 ;
  assign n28187 = n13235 ^ n3386 ^ 1'b0 ;
  assign n28188 = n28186 & n28187 ;
  assign n28189 = n17638 & ~n28188 ;
  assign n28190 = n15104 & n18664 ;
  assign n28191 = n28190 ^ n2530 ^ 1'b0 ;
  assign n28192 = n15687 ^ n534 ^ 1'b0 ;
  assign n28193 = n872 | n17577 ;
  assign n28194 = n28193 ^ n4348 ^ 1'b0 ;
  assign n28195 = n27333 ^ n9928 ^ 1'b0 ;
  assign n28196 = n4598 & ~n28195 ;
  assign n28198 = n10129 | n14927 ;
  assign n28199 = n28198 ^ n2663 ^ 1'b0 ;
  assign n28197 = n3496 & n8947 ;
  assign n28200 = n28199 ^ n28197 ^ 1'b0 ;
  assign n28201 = n19486 & n28200 ;
  assign n28203 = x212 & n4123 ;
  assign n28202 = ~n779 & n18056 ;
  assign n28204 = n28203 ^ n28202 ^ 1'b0 ;
  assign n28205 = n28204 ^ n2706 ^ 1'b0 ;
  assign n28206 = n7365 & n28205 ;
  assign n28207 = n28206 ^ n7850 ^ 1'b0 ;
  assign n28208 = ~n12138 & n26626 ;
  assign n28209 = n22033 ^ n11203 ^ 1'b0 ;
  assign n28210 = n3362 & n28209 ;
  assign n28211 = n25512 ^ n4445 ^ 1'b0 ;
  assign n28212 = n3586 & ~n28211 ;
  assign n28213 = n28212 ^ n14114 ^ 1'b0 ;
  assign n28214 = n28213 ^ n14981 ^ n2119 ;
  assign n28215 = n11547 | n21497 ;
  assign n28216 = n12980 | n28215 ;
  assign n28217 = n2904 & n24041 ;
  assign n28218 = ~n28216 & n28217 ;
  assign n28219 = ~n28214 & n28218 ;
  assign n28220 = n10212 | n10897 ;
  assign n28221 = n28220 ^ n11610 ^ 1'b0 ;
  assign n28222 = ( n1125 & n5767 ) | ( n1125 & n8730 ) | ( n5767 & n8730 ) ;
  assign n28223 = n20463 & n28222 ;
  assign n28226 = ( ~n8678 & n11494 ) | ( ~n8678 & n14803 ) | ( n11494 & n14803 ) ;
  assign n28224 = n3290 | n15324 ;
  assign n28225 = n28224 ^ n22281 ^ 1'b0 ;
  assign n28227 = n28226 ^ n28225 ^ 1'b0 ;
  assign n28228 = ~n923 & n7967 ;
  assign n28229 = n2409 & ~n28228 ;
  assign n28230 = n28229 ^ n3075 ^ 1'b0 ;
  assign n28231 = ~n10532 & n28230 ;
  assign n28232 = n23202 ^ n20746 ^ 1'b0 ;
  assign n28233 = ~n1844 & n3747 ;
  assign n28234 = n1844 & n28233 ;
  assign n28235 = ~n1328 & n2570 ;
  assign n28236 = n28234 & n28235 ;
  assign n28237 = n1958 & ~n4593 ;
  assign n28238 = n28236 & n28237 ;
  assign n28239 = n1129 | n28238 ;
  assign n28240 = ~n22757 & n28239 ;
  assign n28241 = n28240 ^ n3511 ^ 1'b0 ;
  assign n28242 = n28241 ^ n4768 ^ 1'b0 ;
  assign n28243 = ( ~n14867 & n28232 ) | ( ~n14867 & n28242 ) | ( n28232 & n28242 ) ;
  assign n28244 = n7432 & n22303 ;
  assign n28245 = n11186 & n13245 ;
  assign n28246 = ~n19337 & n28245 ;
  assign n28247 = ~n8178 & n20747 ;
  assign n28248 = n28247 ^ n26128 ^ 1'b0 ;
  assign n28249 = n3770 ^ n1170 ^ 1'b0 ;
  assign n28250 = n5356 & n28249 ;
  assign n28251 = n26125 & n28250 ;
  assign n28252 = n28251 ^ n11118 ^ n10686 ;
  assign n28253 = ( n1874 & n9079 ) | ( n1874 & n25990 ) | ( n9079 & n25990 ) ;
  assign n28254 = n11191 & n14016 ;
  assign n28255 = ~n2116 & n28254 ;
  assign n28256 = n21579 & n28255 ;
  assign n28257 = n7844 & n8475 ;
  assign n28258 = n8968 & n28257 ;
  assign n28259 = ~n27658 & n28258 ;
  assign n28260 = n2306 | n14324 ;
  assign n28261 = n28260 ^ n738 ^ 1'b0 ;
  assign n28262 = ( x85 & ~n7630 ) | ( x85 & n13077 ) | ( ~n7630 & n13077 ) ;
  assign n28263 = n24276 ^ n14873 ^ 1'b0 ;
  assign n28264 = n5705 | n7771 ;
  assign n28265 = n28264 ^ n4055 ^ 1'b0 ;
  assign n28266 = ( n5142 & n21554 ) | ( n5142 & ~n28265 ) | ( n21554 & ~n28265 ) ;
  assign n28267 = n12552 ^ n2875 ^ 1'b0 ;
  assign n28268 = n10963 & ~n16059 ;
  assign n28269 = ( ~n7813 & n28267 ) | ( ~n7813 & n28268 ) | ( n28267 & n28268 ) ;
  assign n28270 = n18000 & ~n28269 ;
  assign n28271 = n23443 ^ n11950 ^ n3425 ;
  assign n28272 = n10296 & n28271 ;
  assign n28273 = ~n8981 & n28272 ;
  assign n28274 = n1660 & ~n28273 ;
  assign n28275 = n4458 | n12090 ;
  assign n28276 = n915 & ~n2077 ;
  assign n28277 = n1333 & ~n9758 ;
  assign n28278 = n10841 & ~n23794 ;
  assign n28279 = n2900 | n10139 ;
  assign n28284 = ~n13232 & n15137 ;
  assign n28280 = n7925 & ~n19923 ;
  assign n28281 = n9865 & n28280 ;
  assign n28282 = ( n1548 & n5939 ) | ( n1548 & ~n7966 ) | ( n5939 & ~n7966 ) ;
  assign n28283 = ~n28281 & n28282 ;
  assign n28285 = n28284 ^ n28283 ^ 1'b0 ;
  assign n28286 = ( ~n276 & n11816 ) | ( ~n276 & n26075 ) | ( n11816 & n26075 ) ;
  assign n28287 = n8943 ^ n3453 ^ 1'b0 ;
  assign n28288 = n27301 & ~n28287 ;
  assign n28289 = n28288 ^ n14317 ^ 1'b0 ;
  assign n28290 = n12553 & n28289 ;
  assign n28291 = ~n3624 & n28290 ;
  assign n28292 = n1170 | n22419 ;
  assign n28293 = n2024 | n9306 ;
  assign n28294 = n4117 & ~n16479 ;
  assign n28295 = n28294 ^ n20358 ^ 1'b0 ;
  assign n28296 = n3159 | n27666 ;
  assign n28297 = n12022 | n24297 ;
  assign n28299 = ~n9799 & n12485 ;
  assign n28300 = n12969 & n28299 ;
  assign n28301 = ~n12174 & n28300 ;
  assign n28298 = ~n6004 & n20858 ;
  assign n28302 = n28301 ^ n28298 ^ 1'b0 ;
  assign n28303 = n28302 ^ n11488 ^ n6272 ;
  assign n28304 = ~n15843 & n24476 ;
  assign n28305 = n28304 ^ n9742 ^ n6363 ;
  assign n28306 = ( n8219 & n20299 ) | ( n8219 & n28305 ) | ( n20299 & n28305 ) ;
  assign n28307 = n17267 ^ n9012 ^ 1'b0 ;
  assign n28308 = ~n8384 & n28307 ;
  assign n28309 = ~n28307 & n28308 ;
  assign n28310 = ~n2989 & n28309 ;
  assign n28311 = n10857 ^ n3114 ^ 1'b0 ;
  assign n28312 = n28310 & ~n28311 ;
  assign n28313 = n19464 & n28312 ;
  assign n28314 = ~n28312 & n28313 ;
  assign n28315 = n21881 ^ n2898 ^ 1'b0 ;
  assign n28316 = n10382 & ~n22697 ;
  assign n28317 = n23820 ^ n15866 ^ 1'b0 ;
  assign n28318 = n27405 ^ n4236 ^ 1'b0 ;
  assign n28319 = ~n10044 & n28318 ;
  assign n28320 = n28319 ^ n924 ^ 1'b0 ;
  assign n28321 = n5626 ^ n3954 ^ 1'b0 ;
  assign n28322 = n8243 & ~n11041 ;
  assign n28323 = ~n13216 & n28322 ;
  assign n28324 = ( n28320 & n28321 ) | ( n28320 & n28323 ) | ( n28321 & n28323 ) ;
  assign n28325 = ~n22821 & n27871 ;
  assign n28326 = ~n25381 & n28325 ;
  assign n28327 = n17951 ^ n6698 ^ 1'b0 ;
  assign n28328 = n274 | n7484 ;
  assign n28330 = n7455 ^ n1623 ^ 1'b0 ;
  assign n28329 = n4685 & ~n7238 ;
  assign n28331 = n28330 ^ n28329 ^ n17848 ;
  assign n28332 = n28331 ^ n23864 ^ n4111 ;
  assign n28335 = ~n8005 & n24332 ;
  assign n28336 = ~n9907 & n28335 ;
  assign n28333 = n7962 ^ n1638 ^ x149 ;
  assign n28334 = n23410 & n28333 ;
  assign n28337 = n28336 ^ n28334 ^ 1'b0 ;
  assign n28338 = n1593 & n4804 ;
  assign n28339 = n19433 & n28338 ;
  assign n28340 = n28339 ^ n17784 ^ 1'b0 ;
  assign n28341 = ~n1694 & n2904 ;
  assign n28342 = ~n5883 & n28341 ;
  assign n28343 = n28342 ^ n7174 ^ n4596 ;
  assign n28344 = n12201 | n28343 ;
  assign n28345 = ( n449 & n4512 ) | ( n449 & n7558 ) | ( n4512 & n7558 ) ;
  assign n28346 = n24809 ^ n3344 ^ 1'b0 ;
  assign n28347 = n28345 | n28346 ;
  assign n28348 = n28347 ^ n7879 ^ 1'b0 ;
  assign n28349 = n28348 ^ n10108 ^ 1'b0 ;
  assign n28350 = n28344 & ~n28349 ;
  assign n28351 = x6 & n1712 ;
  assign n28352 = n28351 ^ n7948 ^ n6966 ;
  assign n28353 = x226 & n1680 ;
  assign n28354 = n28353 ^ n6069 ^ 1'b0 ;
  assign n28355 = n2008 & n8198 ;
  assign n28356 = n26195 ^ n10509 ^ 1'b0 ;
  assign n28357 = ( n28354 & n28355 ) | ( n28354 & ~n28356 ) | ( n28355 & ~n28356 ) ;
  assign n28358 = n4375 & ~n9167 ;
  assign n28359 = ~n3124 & n4895 ;
  assign n28360 = ~n28358 & n28359 ;
  assign n28361 = n2924 | n10347 ;
  assign n28362 = n20229 & ~n28361 ;
  assign n28363 = n1220 & ~n4902 ;
  assign n28364 = n28363 ^ n1203 ^ 1'b0 ;
  assign n28365 = ~n22403 & n28364 ;
  assign n28366 = n28365 ^ n9110 ^ 1'b0 ;
  assign n28367 = n28362 & n28366 ;
  assign n28368 = n7179 | n18771 ;
  assign n28369 = n28368 ^ n10746 ^ 1'b0 ;
  assign n28370 = n3450 & n28369 ;
  assign n28371 = n16468 ^ n13779 ^ 1'b0 ;
  assign n28372 = n7449 & ~n28371 ;
  assign n28373 = n8136 ^ n3651 ^ 1'b0 ;
  assign n28374 = ~n26097 & n28373 ;
  assign n28375 = n20759 ^ n8564 ^ 1'b0 ;
  assign n28378 = n7738 ^ n7250 ^ 1'b0 ;
  assign n28379 = n3140 | n28378 ;
  assign n28376 = n13803 & ~n23957 ;
  assign n28377 = ~n23382 & n28376 ;
  assign n28380 = n28379 ^ n28377 ^ 1'b0 ;
  assign n28381 = ~n23075 & n28380 ;
  assign n28382 = n26861 ^ n4957 ^ 1'b0 ;
  assign n28383 = n6339 ^ n647 ^ 1'b0 ;
  assign n28384 = n16898 & n28383 ;
  assign n28385 = n28384 ^ n3253 ^ 1'b0 ;
  assign n28387 = n1935 & ~n17987 ;
  assign n28386 = ~n293 & n9930 ;
  assign n28388 = n28387 ^ n28386 ^ 1'b0 ;
  assign n28391 = ~n14294 & n17065 ;
  assign n28392 = n17578 & n18763 ;
  assign n28393 = n28391 & n28392 ;
  assign n28389 = n10666 | n17977 ;
  assign n28390 = n5379 & ~n28389 ;
  assign n28394 = n28393 ^ n28390 ^ x199 ;
  assign n28409 = n7815 ^ n7264 ^ 1'b0 ;
  assign n28396 = x25 & ~n1882 ;
  assign n28397 = n1882 & n28396 ;
  assign n28398 = n583 | n751 ;
  assign n28399 = n583 & ~n28398 ;
  assign n28400 = n3447 & ~n28399 ;
  assign n28401 = ~n3447 & n28400 ;
  assign n28402 = x69 & x211 ;
  assign n28403 = ~x211 & n28402 ;
  assign n28404 = ~n711 & n28403 ;
  assign n28405 = ~n348 & n28404 ;
  assign n28406 = ~n28404 & n28405 ;
  assign n28407 = n28401 | n28406 ;
  assign n28408 = n28397 & ~n28407 ;
  assign n28395 = n4745 ^ x207 ^ 1'b0 ;
  assign n28410 = n28409 ^ n28408 ^ n28395 ;
  assign n28411 = n3579 | n16096 ;
  assign n28412 = n28411 ^ n10172 ^ 1'b0 ;
  assign n28413 = n4603 & ~n11525 ;
  assign n28414 = n611 & n28413 ;
  assign n28415 = n1242 | n1775 ;
  assign n28416 = n1667 & ~n28415 ;
  assign n28417 = n729 & ~n28416 ;
  assign n28418 = n2291 & ~n4668 ;
  assign n28419 = n842 | n28418 ;
  assign n28420 = n4665 | n4821 ;
  assign n28421 = n16889 & ~n26247 ;
  assign n28422 = n18822 ^ n17954 ^ 1'b0 ;
  assign n28423 = n10247 & ~n16363 ;
  assign n28424 = n12842 | n28423 ;
  assign n28425 = n20360 ^ n2456 ^ 1'b0 ;
  assign n28426 = n28425 ^ n24310 ^ 1'b0 ;
  assign n28427 = ~n3826 & n28426 ;
  assign n28428 = n28424 & n28427 ;
  assign n28429 = n13285 ^ n973 ^ 1'b0 ;
  assign n28430 = n1010 & ~n28429 ;
  assign n28431 = n19543 ^ n18569 ^ 1'b0 ;
  assign n28432 = n18014 ^ n17926 ^ 1'b0 ;
  assign n28433 = n18910 & ~n28432 ;
  assign n28434 = n13163 | n14372 ;
  assign n28435 = n19458 ^ n6639 ^ 1'b0 ;
  assign n28436 = ~n28434 & n28435 ;
  assign n28437 = n1641 & ~n5920 ;
  assign n28438 = n15385 ^ n9742 ^ 1'b0 ;
  assign n28439 = n26868 ^ n22363 ^ 1'b0 ;
  assign n28440 = n20058 | n25775 ;
  assign n28441 = n2002 | n28440 ;
  assign n28442 = ~n8375 & n14708 ;
  assign n28443 = ~n7358 & n28442 ;
  assign n28444 = n18254 | n28443 ;
  assign n28446 = n15101 & ~n18350 ;
  assign n28445 = n22837 ^ n13521 ^ 1'b0 ;
  assign n28447 = n28446 ^ n28445 ^ 1'b0 ;
  assign n28448 = n5604 | n28447 ;
  assign n28450 = n611 | n19388 ;
  assign n28451 = n21676 | n28450 ;
  assign n28449 = n2328 & n4271 ;
  assign n28452 = n28451 ^ n28449 ^ 1'b0 ;
  assign n28453 = n10306 ^ n1680 ^ 1'b0 ;
  assign n28454 = n571 | n28453 ;
  assign n28455 = n28454 ^ n4114 ^ 1'b0 ;
  assign n28456 = n24887 ^ n7819 ^ 1'b0 ;
  assign n28457 = n9759 & ~n28456 ;
  assign n28458 = ~n17092 & n28457 ;
  assign n28459 = n18473 & ~n28458 ;
  assign n28460 = n8090 & n9623 ;
  assign n28461 = n28460 ^ n2023 ^ 1'b0 ;
  assign n28462 = n28459 | n28461 ;
  assign n28463 = n4950 & n15954 ;
  assign n28464 = n19496 ^ n16106 ^ 1'b0 ;
  assign n28465 = ~n13420 & n15884 ;
  assign n28466 = ~n28464 & n28465 ;
  assign n28467 = n28466 ^ n27539 ^ 1'b0 ;
  assign n28469 = n2819 & n5823 ;
  assign n28468 = ~n2492 & n7378 ;
  assign n28470 = n28469 ^ n28468 ^ 1'b0 ;
  assign n28471 = n7130 & n12398 ;
  assign n28472 = n3479 & n28471 ;
  assign n28473 = n16709 ^ n14784 ^ n9608 ;
  assign n28474 = ( n11450 & ~n28472 ) | ( n11450 & n28473 ) | ( ~n28472 & n28473 ) ;
  assign n28475 = n14101 ^ n9826 ^ 1'b0 ;
  assign n28476 = n14971 | n28475 ;
  assign n28477 = n24128 & ~n25696 ;
  assign n28478 = n1735 & n3839 ;
  assign n28479 = n17730 ^ n15644 ^ 1'b0 ;
  assign n28480 = ~n28478 & n28479 ;
  assign n28481 = x55 & n28480 ;
  assign n28482 = n1377 & ~n4815 ;
  assign n28483 = n4815 & n28482 ;
  assign n28484 = ~n3311 & n28483 ;
  assign n28485 = n28484 ^ n10582 ^ 1'b0 ;
  assign n28486 = ~n3721 & n28485 ;
  assign n28487 = n6260 | n28486 ;
  assign n28488 = n28487 ^ n5145 ^ 1'b0 ;
  assign n28489 = n28481 & ~n28488 ;
  assign n28490 = ~n14558 & n17477 ;
  assign n28491 = n3348 | n13277 ;
  assign n28492 = n28491 ^ n2058 ^ 1'b0 ;
  assign n28493 = n1851 & ~n28492 ;
  assign n28494 = n4888 & n8200 ;
  assign n28495 = ~n10189 & n20663 ;
  assign n28496 = n8043 | n28495 ;
  assign n28497 = n28496 ^ n16977 ^ 1'b0 ;
  assign n28498 = n2140 | n11773 ;
  assign n28499 = n28498 ^ n12812 ^ 1'b0 ;
  assign n28500 = ~n5362 & n28499 ;
  assign n28501 = n13135 & ~n15491 ;
  assign n28502 = ~n11492 & n15303 ;
  assign n28503 = n28464 ^ n24428 ^ 1'b0 ;
  assign n28504 = n28502 & n28503 ;
  assign n28505 = n9002 | n19810 ;
  assign n28506 = n22375 | n23273 ;
  assign n28507 = n969 & ~n28506 ;
  assign n28508 = n1803 & ~n5385 ;
  assign n28509 = ( n22879 & n24971 ) | ( n22879 & n28508 ) | ( n24971 & n28508 ) ;
  assign n28510 = n349 & ~n13779 ;
  assign n28511 = n5883 ^ n3034 ^ 1'b0 ;
  assign n28512 = n15273 & n28511 ;
  assign n28513 = n21126 | n28512 ;
  assign n28514 = n28513 ^ n11952 ^ 1'b0 ;
  assign n28515 = n17409 ^ n9065 ^ 1'b0 ;
  assign n28516 = n3769 & n28515 ;
  assign n28517 = ~n10781 & n28516 ;
  assign n28518 = n27564 & n28517 ;
  assign n28519 = ~n5608 & n15828 ;
  assign n28520 = ~n9067 & n28519 ;
  assign n28521 = n13435 & n28348 ;
  assign n28522 = ~n18285 & n28521 ;
  assign n28524 = n5812 & ~n8165 ;
  assign n28525 = n28524 ^ n498 ^ 1'b0 ;
  assign n28523 = ~n7223 & n19210 ;
  assign n28526 = n28525 ^ n28523 ^ 1'b0 ;
  assign n28527 = ( n2883 & n7398 ) | ( n2883 & ~n28526 ) | ( n7398 & ~n28526 ) ;
  assign n28528 = n18733 ^ n11815 ^ 1'b0 ;
  assign n28529 = n332 | n4327 ;
  assign n28530 = n28528 & ~n28529 ;
  assign n28531 = n28530 ^ n11496 ^ 1'b0 ;
  assign n28532 = n26349 | n28531 ;
  assign n28533 = n2426 | n2993 ;
  assign n28534 = n28533 ^ n1667 ^ 1'b0 ;
  assign n28535 = n19186 ^ n18387 ^ 1'b0 ;
  assign n28536 = ~n28534 & n28535 ;
  assign n28537 = n8058 & n28536 ;
  assign n28538 = n15883 | n28537 ;
  assign n28539 = n27826 & n28538 ;
  assign n28540 = n28539 ^ n24228 ^ 1'b0 ;
  assign n28541 = ~n12598 & n22307 ;
  assign n28542 = n28541 ^ n10717 ^ 1'b0 ;
  assign n28543 = ( n877 & n3449 ) | ( n877 & n9359 ) | ( n3449 & n9359 ) ;
  assign n28544 = n28543 ^ n1321 ^ 1'b0 ;
  assign n28545 = n28544 ^ n15533 ^ 1'b0 ;
  assign n28546 = ~n2065 & n4343 ;
  assign n28547 = n28546 ^ n12280 ^ 1'b0 ;
  assign n28548 = n4428 & ~n5127 ;
  assign n28549 = n4733 & n8471 ;
  assign n28550 = n525 & ~n1890 ;
  assign n28551 = n28550 ^ n4944 ^ n1796 ;
  assign n28552 = n28549 & n28551 ;
  assign n28553 = n28548 | n28552 ;
  assign n28554 = n628 & n2013 ;
  assign n28555 = ~n15366 & n22800 ;
  assign n28556 = ~x163 & n28555 ;
  assign n28557 = ~n2502 & n3606 ;
  assign n28558 = n2502 & n28557 ;
  assign n28559 = n9754 ^ n8184 ^ 1'b0 ;
  assign n28560 = n5667 & n28559 ;
  assign n28561 = n28560 ^ n11963 ^ 1'b0 ;
  assign n28562 = n3702 & n28561 ;
  assign n28563 = n432 & n28562 ;
  assign n28564 = n28563 ^ n28471 ^ 1'b0 ;
  assign n28565 = n6856 & ~n28564 ;
  assign n28566 = ( n9317 & n28558 ) | ( n9317 & n28565 ) | ( n28558 & n28565 ) ;
  assign n28567 = n6474 & n8466 ;
  assign n28568 = n12891 ^ n4268 ^ 1'b0 ;
  assign n28569 = n28567 | n28568 ;
  assign n28570 = ~n2301 & n12150 ;
  assign n28571 = n15572 & n28570 ;
  assign n28572 = n28571 ^ n7388 ^ 1'b0 ;
  assign n28573 = n25492 ^ n13266 ^ n8064 ;
  assign n28574 = n27343 & ~n28573 ;
  assign n28575 = n28574 ^ n27739 ^ 1'b0 ;
  assign n28576 = n12329 ^ n3174 ^ 1'b0 ;
  assign n28577 = n21660 | n28576 ;
  assign n28578 = ~x180 & n7839 ;
  assign n28579 = n4548 & ~n28578 ;
  assign n28580 = n28579 ^ n11384 ^ 1'b0 ;
  assign n28581 = ~n8072 & n28580 ;
  assign n28582 = n1819 & n5812 ;
  assign n28583 = n28582 ^ n4476 ^ 1'b0 ;
  assign n28586 = n618 | n9468 ;
  assign n28584 = n12989 & n14862 ;
  assign n28585 = n28584 ^ n12836 ^ 1'b0 ;
  assign n28587 = n28586 ^ n28585 ^ 1'b0 ;
  assign n28588 = n28587 ^ n10663 ^ 1'b0 ;
  assign n28589 = n12778 & n28588 ;
  assign n28590 = n28583 & n28589 ;
  assign n28591 = n22780 ^ n10552 ^ 1'b0 ;
  assign n28592 = n6358 ^ n1463 ^ 1'b0 ;
  assign n28593 = n28592 ^ n15086 ^ 1'b0 ;
  assign n28594 = n16334 & n28593 ;
  assign n28595 = n14544 ^ n12519 ^ 1'b0 ;
  assign n28596 = n25906 & ~n28595 ;
  assign n28597 = n17008 ^ n16579 ^ 1'b0 ;
  assign n28598 = n12441 & ~n28597 ;
  assign n28599 = n15117 ^ n998 ^ 1'b0 ;
  assign n28600 = ~n11965 & n28599 ;
  assign n28601 = n2569 & ~n7360 ;
  assign n28602 = n7784 & n28601 ;
  assign n28603 = n11542 ^ n1006 ^ 1'b0 ;
  assign n28604 = n3250 | n28603 ;
  assign n28605 = ( n8583 & n18434 ) | ( n8583 & n28604 ) | ( n18434 & n28604 ) ;
  assign n28606 = n28605 ^ n8309 ^ 1'b0 ;
  assign n28607 = n14787 & n28606 ;
  assign n28608 = n21739 ^ n1328 ^ 1'b0 ;
  assign n28609 = n20238 ^ n825 ^ 1'b0 ;
  assign n28610 = n14101 & ~n21240 ;
  assign n28611 = n28610 ^ n8999 ^ 1'b0 ;
  assign n28612 = ( ~n9413 & n14107 ) | ( ~n9413 & n28611 ) | ( n14107 & n28611 ) ;
  assign n28613 = ~n21513 & n28612 ;
  assign n28614 = n28613 ^ n10022 ^ 1'b0 ;
  assign n28615 = n1649 | n11245 ;
  assign n28616 = n17021 | n28615 ;
  assign n28617 = n5917 & n28616 ;
  assign n28618 = n1981 & n28617 ;
  assign n28619 = n15580 ^ n1475 ^ 1'b0 ;
  assign n28620 = n2366 & n28619 ;
  assign n28621 = n23155 & n28620 ;
  assign n28624 = n2942 ^ n723 ^ 1'b0 ;
  assign n28625 = ~n668 & n28624 ;
  assign n28622 = n4906 ^ n3088 ^ 1'b0 ;
  assign n28623 = n27559 | n28622 ;
  assign n28626 = n28625 ^ n28623 ^ 1'b0 ;
  assign n28627 = n6402 | n27307 ;
  assign n28628 = n3993 & n6881 ;
  assign n28629 = n28627 & n28628 ;
  assign n28630 = n15874 ^ n9289 ^ n375 ;
  assign n28631 = n5667 & ~n28630 ;
  assign n28632 = ( n5830 & n8352 ) | ( n5830 & n16271 ) | ( n8352 & n16271 ) ;
  assign n28633 = n17732 ^ n9321 ^ 1'b0 ;
  assign n28634 = n24039 & n28633 ;
  assign n28635 = n23449 | n28634 ;
  assign n28636 = ~n1613 & n7330 ;
  assign n28637 = n28636 ^ n19924 ^ n8359 ;
  assign n28638 = n17852 ^ n17071 ^ 1'b0 ;
  assign n28639 = n26420 & n28638 ;
  assign n28640 = n28639 ^ n7825 ^ 1'b0 ;
  assign n28641 = n17430 & n28640 ;
  assign n28642 = n1234 | n2075 ;
  assign n28643 = n847 | n28642 ;
  assign n28644 = n1255 | n5081 ;
  assign n28645 = n28643 | n28644 ;
  assign n28646 = n17929 | n28645 ;
  assign n28647 = n28646 ^ n826 ^ 1'b0 ;
  assign n28648 = n8077 & n16902 ;
  assign n28649 = n28648 ^ n14979 ^ 1'b0 ;
  assign n28650 = n4213 & ~n28649 ;
  assign n28651 = ~n4213 & n28650 ;
  assign n28652 = n12307 & n28651 ;
  assign n28653 = n28652 ^ n27198 ^ 1'b0 ;
  assign n28654 = n20527 ^ n3672 ^ 1'b0 ;
  assign n28655 = n21364 ^ n448 ^ 1'b0 ;
  assign n28656 = n5313 & n19210 ;
  assign n28657 = ~n28655 & n28656 ;
  assign n28658 = n17349 & ~n28657 ;
  assign n28659 = ~n2310 & n28658 ;
  assign n28660 = n28659 ^ n26716 ^ 1'b0 ;
  assign n28664 = n13016 & ~n16992 ;
  assign n28665 = n5505 & n28664 ;
  assign n28661 = n6648 & ~n11907 ;
  assign n28662 = n5420 & ~n17187 ;
  assign n28663 = n28661 | n28662 ;
  assign n28666 = n28665 ^ n28663 ^ 1'b0 ;
  assign n28667 = n2287 & ~n2743 ;
  assign n28668 = n28055 ^ n12201 ^ 1'b0 ;
  assign n28669 = n13771 | n23204 ;
  assign n28670 = n28669 ^ n18129 ^ 1'b0 ;
  assign n28677 = n3038 | n10675 ;
  assign n28678 = n3038 & ~n28677 ;
  assign n28679 = n1077 & n10986 ;
  assign n28680 = n28679 ^ n862 ^ 1'b0 ;
  assign n28681 = n28678 | n28680 ;
  assign n28682 = n28681 ^ n10258 ^ 1'b0 ;
  assign n28672 = n10512 ^ n638 ^ 1'b0 ;
  assign n28671 = x185 & n2430 ;
  assign n28673 = n28672 ^ n28671 ^ n16546 ;
  assign n28674 = n28673 ^ n27556 ^ 1'b0 ;
  assign n28675 = ~n23400 & n28674 ;
  assign n28676 = n23400 & n28675 ;
  assign n28683 = n28682 ^ n28676 ^ 1'b0 ;
  assign n28684 = ( x113 & ~n8676 ) | ( x113 & n15271 ) | ( ~n8676 & n15271 ) ;
  assign n28685 = n4584 ^ n848 ^ 1'b0 ;
  assign n28686 = n7822 ^ n3005 ^ 1'b0 ;
  assign n28687 = n3114 & n28686 ;
  assign n28688 = n28687 ^ n26344 ^ 1'b0 ;
  assign n28689 = ~n6719 & n8332 ;
  assign n28690 = ~n1678 & n28689 ;
  assign n28691 = n28690 ^ n3333 ^ 1'b0 ;
  assign n28692 = n28691 ^ n23880 ^ 1'b0 ;
  assign n28693 = ~n2776 & n16430 ;
  assign n28694 = ~n725 & n28693 ;
  assign n28695 = n1152 | n13267 ;
  assign n28696 = n18779 ^ x182 ^ 1'b0 ;
  assign n28697 = n28696 ^ n497 ^ 1'b0 ;
  assign n28698 = ( n2835 & ~n6046 ) | ( n2835 & n7597 ) | ( ~n6046 & n7597 ) ;
  assign n28699 = n28698 ^ n21837 ^ 1'b0 ;
  assign n28700 = n2396 & n28699 ;
  assign n28701 = n3371 & n18720 ;
  assign n28703 = n4148 & n11497 ;
  assign n28702 = ~n7707 & n9479 ;
  assign n28704 = n28703 ^ n28702 ^ 1'b0 ;
  assign n28705 = n9759 ^ n9357 ^ 1'b0 ;
  assign n28706 = n28705 ^ n21467 ^ 1'b0 ;
  assign n28707 = n8843 & ~n28706 ;
  assign n28708 = ~n4638 & n28707 ;
  assign n28709 = n21893 & n28708 ;
  assign n28714 = ~n2909 & n4479 ;
  assign n28712 = n2188 | n4896 ;
  assign n28713 = n28712 ^ n8169 ^ 1'b0 ;
  assign n28715 = n28714 ^ n28713 ^ n5988 ;
  assign n28710 = n6851 & ~n21088 ;
  assign n28711 = ~n9911 & n28710 ;
  assign n28716 = n28715 ^ n28711 ^ n25047 ;
  assign n28717 = n18453 ^ n14188 ^ 1'b0 ;
  assign n28718 = n14500 & ~n18453 ;
  assign n28719 = n28718 ^ n13905 ^ 1'b0 ;
  assign n28720 = ~n8323 & n13931 ;
  assign n28721 = ~n9022 & n28720 ;
  assign n28722 = n11963 & n24713 ;
  assign n28723 = ~n26069 & n28722 ;
  assign n28725 = n18164 ^ x181 ^ 1'b0 ;
  assign n28724 = n11790 & ~n14954 ;
  assign n28726 = n28725 ^ n28724 ^ 1'b0 ;
  assign n28727 = n19736 ^ n8224 ^ 1'b0 ;
  assign n28728 = n6481 | n14807 ;
  assign n28729 = n285 & ~n28728 ;
  assign n28730 = ~n3113 & n18637 ;
  assign n28731 = ~n4450 & n12146 ;
  assign n28732 = n28731 ^ n1101 ^ 1'b0 ;
  assign n28733 = n26501 | n28732 ;
  assign n28734 = n25062 ^ n6952 ^ 1'b0 ;
  assign n28735 = n5342 | n28734 ;
  assign n28736 = n4268 & n13813 ;
  assign n28737 = n28736 ^ n15759 ^ 1'b0 ;
  assign n28738 = ~n15191 & n23042 ;
  assign n28739 = n25897 ^ n10612 ^ 1'b0 ;
  assign n28740 = n17197 | n28739 ;
  assign n28741 = n3281 & ~n14767 ;
  assign n28742 = ~n9935 & n28741 ;
  assign n28743 = n5364 | n28742 ;
  assign n28744 = n3260 & n20640 ;
  assign n28745 = n7586 ^ n6281 ^ 1'b0 ;
  assign n28746 = n28745 ^ n16429 ^ n1819 ;
  assign n28747 = ( n12830 & n23376 ) | ( n12830 & ~n28746 ) | ( n23376 & ~n28746 ) ;
  assign n28748 = n23362 ^ n13372 ^ n10780 ;
  assign n28750 = n7501 & n26809 ;
  assign n28751 = n9190 & n28750 ;
  assign n28752 = n7617 | n28751 ;
  assign n28753 = n28752 ^ x138 ^ 1'b0 ;
  assign n28749 = n7749 & n20726 ;
  assign n28754 = n28753 ^ n28749 ^ 1'b0 ;
  assign n28755 = n21696 ^ n14990 ^ 1'b0 ;
  assign n28756 = n4838 & n28755 ;
  assign n28757 = n28756 ^ n27044 ^ 1'b0 ;
  assign n28758 = n9745 & ~n19983 ;
  assign n28759 = ~n27119 & n28758 ;
  assign n28760 = n2681 & n17858 ;
  assign n28761 = n28760 ^ n10593 ^ 1'b0 ;
  assign n28762 = ( n4958 & n5554 ) | ( n4958 & n28761 ) | ( n5554 & n28761 ) ;
  assign n28763 = n4755 & n7001 ;
  assign n28764 = ~n4755 & n28763 ;
  assign n28765 = n11488 & ~n28764 ;
  assign n28766 = ~n11488 & n28765 ;
  assign n28767 = n15775 ^ n12273 ^ 1'b0 ;
  assign n28768 = ~n28766 & n28767 ;
  assign n28769 = n1316 & ~n28768 ;
  assign n28770 = n4485 & n15547 ;
  assign n28771 = n15809 & ~n28770 ;
  assign n28772 = ( n10886 & n15602 ) | ( n10886 & ~n17505 ) | ( n15602 & ~n17505 ) ;
  assign n28773 = x137 & ~n26372 ;
  assign n28774 = n4520 & n19489 ;
  assign n28775 = n28774 ^ n26341 ^ 1'b0 ;
  assign n28776 = n14513 & ~n28775 ;
  assign n28777 = n19922 & n28776 ;
  assign n28778 = n28777 ^ n1738 ^ 1'b0 ;
  assign n28779 = ~n9210 & n28778 ;
  assign n28780 = n11997 ^ n10963 ^ 1'b0 ;
  assign n28781 = n13597 ^ n5021 ^ n1817 ;
  assign n28782 = n11526 | n28781 ;
  assign n28783 = n14479 | n28782 ;
  assign n28784 = n6106 & n8924 ;
  assign n28785 = n15065 & n26339 ;
  assign n28786 = n18034 ^ n2781 ^ 1'b0 ;
  assign n28787 = ~n2653 & n6506 ;
  assign n28788 = n874 | n11321 ;
  assign n28789 = n28788 ^ n21882 ^ 1'b0 ;
  assign n28790 = n7844 ^ n752 ^ 1'b0 ;
  assign n28791 = n28789 & ~n28790 ;
  assign n28792 = n7814 ^ n7165 ^ 1'b0 ;
  assign n28794 = n315 & n6906 ;
  assign n28795 = n5703 & ~n21218 ;
  assign n28796 = n28795 ^ n13258 ^ 1'b0 ;
  assign n28797 = n28794 & ~n28796 ;
  assign n28793 = ( n17484 & ~n19085 ) | ( n17484 & n24965 ) | ( ~n19085 & n24965 ) ;
  assign n28798 = n28797 ^ n28793 ^ 1'b0 ;
  assign n28799 = n14551 ^ n14256 ^ 1'b0 ;
  assign n28800 = n614 | n8134 ;
  assign n28801 = n17458 & ~n28800 ;
  assign n28802 = n3126 | n23780 ;
  assign n28803 = n27170 ^ n2178 ^ 1'b0 ;
  assign n28804 = ~n28802 & n28803 ;
  assign n28805 = n28804 ^ n6817 ^ 1'b0 ;
  assign n28806 = n3904 | n28805 ;
  assign n28807 = ~n21984 & n26233 ;
  assign n28811 = n25618 ^ n12664 ^ 1'b0 ;
  assign n28812 = ( n11186 & ~n13657 ) | ( n11186 & n16945 ) | ( ~n13657 & n16945 ) ;
  assign n28813 = n9256 ^ n9074 ^ 1'b0 ;
  assign n28814 = n10652 & ~n28813 ;
  assign n28815 = n28814 ^ n20628 ^ 1'b0 ;
  assign n28816 = n9027 & n28815 ;
  assign n28817 = ( ~n28811 & n28812 ) | ( ~n28811 & n28816 ) | ( n28812 & n28816 ) ;
  assign n28808 = n5242 | n22931 ;
  assign n28809 = n28808 ^ n15090 ^ 1'b0 ;
  assign n28810 = n24501 | n28809 ;
  assign n28818 = n28817 ^ n28810 ^ 1'b0 ;
  assign n28819 = n22837 ^ n1766 ^ 1'b0 ;
  assign n28820 = n2369 & ~n28819 ;
  assign n28821 = n28820 ^ n16822 ^ n8160 ;
  assign n28822 = n20108 ^ n19071 ^ 1'b0 ;
  assign n28823 = n25630 ^ n22929 ^ 1'b0 ;
  assign n28824 = n1832 & ~n28823 ;
  assign n28825 = n28824 ^ n25116 ^ 1'b0 ;
  assign n28826 = n15992 & ~n18453 ;
  assign n28827 = n15428 ^ n4204 ^ 1'b0 ;
  assign n28828 = n15647 ^ n2434 ^ 1'b0 ;
  assign n28829 = ~n6337 & n28828 ;
  assign n28830 = ( ~n366 & n5268 ) | ( ~n366 & n12218 ) | ( n5268 & n12218 ) ;
  assign n28831 = n6788 ^ n2063 ^ n716 ;
  assign n28832 = n28830 | n28831 ;
  assign n28833 = n28832 ^ n14582 ^ 1'b0 ;
  assign n28834 = n14572 ^ n9362 ^ 1'b0 ;
  assign n28835 = n11805 & n11936 ;
  assign n28836 = n28835 ^ n18611 ^ 1'b0 ;
  assign n28837 = ~n18426 & n22537 ;
  assign n28838 = n28837 ^ n4923 ^ n2130 ;
  assign n28839 = n13830 | n28838 ;
  assign n28840 = ( n11999 & ~n12848 ) | ( n11999 & n14580 ) | ( ~n12848 & n14580 ) ;
  assign n28841 = n6963 ^ n6062 ^ 1'b0 ;
  assign n28842 = n4705 & ~n28841 ;
  assign n28843 = ( n3839 & ~n15303 ) | ( n3839 & n28842 ) | ( ~n15303 & n28842 ) ;
  assign n28844 = n17718 ^ n2890 ^ 1'b0 ;
  assign n28845 = n18808 & ~n20224 ;
  assign n28846 = ~n7447 & n28586 ;
  assign n28847 = ~n11435 & n28846 ;
  assign n28848 = ~n10840 & n19328 ;
  assign n28849 = n1828 & n6442 ;
  assign n28850 = n7592 & n28849 ;
  assign n28851 = n20076 | n28850 ;
  assign n28852 = n14647 | n28851 ;
  assign n28853 = n5333 ^ n3962 ^ n367 ;
  assign n28854 = n28853 ^ n25407 ^ 1'b0 ;
  assign n28855 = n23596 ^ n7116 ^ 1'b0 ;
  assign n28856 = n8300 & ~n28855 ;
  assign n28857 = n23297 & n28856 ;
  assign n28858 = n23804 | n28857 ;
  assign n28860 = n5881 & n9944 ;
  assign n28861 = n28860 ^ n18420 ^ 1'b0 ;
  assign n28862 = n23646 | n28861 ;
  assign n28859 = n686 | n9056 ;
  assign n28863 = n28862 ^ n28859 ^ 1'b0 ;
  assign n28864 = n16675 & n25255 ;
  assign n28865 = n11447 ^ n5463 ^ 1'b0 ;
  assign n28866 = n14391 | n28865 ;
  assign n28867 = n9484 ^ x204 ^ 1'b0 ;
  assign n28868 = ( ~n5678 & n28866 ) | ( ~n5678 & n28867 ) | ( n28866 & n28867 ) ;
  assign n28869 = ( ~n1018 & n12871 ) | ( ~n1018 & n28868 ) | ( n12871 & n28868 ) ;
  assign n28870 = n24326 ^ n16857 ^ 1'b0 ;
  assign n28871 = ~n5798 & n12854 ;
  assign n28872 = n28871 ^ n27662 ^ 1'b0 ;
  assign n28873 = n10207 | n28872 ;
  assign n28874 = n4364 & n6529 ;
  assign n28875 = n18052 | n28874 ;
  assign n28876 = n28875 ^ n1744 ^ 1'b0 ;
  assign n28877 = n7306 & ~n8705 ;
  assign n28878 = n28877 ^ n21954 ^ n4714 ;
  assign n28879 = n28878 ^ n6164 ^ 1'b0 ;
  assign n28880 = n1309 & n10990 ;
  assign n28881 = n17149 ^ n15955 ^ 1'b0 ;
  assign n28882 = n28881 ^ n6803 ^ n3668 ;
  assign n28884 = n2970 | n23213 ;
  assign n28885 = n28884 ^ n2634 ^ 1'b0 ;
  assign n28883 = n3397 & ~n4639 ;
  assign n28886 = n28885 ^ n28883 ^ 1'b0 ;
  assign n28887 = n15880 & n28886 ;
  assign n28888 = n10250 ^ n6490 ^ 1'b0 ;
  assign n28889 = ~n24973 & n28888 ;
  assign n28890 = ~n6933 & n28889 ;
  assign n28891 = n28890 ^ n4563 ^ 1'b0 ;
  assign n28892 = ~n7271 & n11015 ;
  assign n28893 = ~n28891 & n28892 ;
  assign n28894 = n11592 ^ n4714 ^ 1'b0 ;
  assign n28895 = n4860 | n28894 ;
  assign n28896 = n4624 | n28895 ;
  assign n28897 = n28893 & ~n28896 ;
  assign n28898 = n17197 | n17794 ;
  assign n28899 = n8855 ^ n4676 ^ 1'b0 ;
  assign n28900 = n12690 | n28899 ;
  assign n28901 = n28900 ^ n3613 ^ 1'b0 ;
  assign n28902 = ~n4388 & n28901 ;
  assign n28903 = ~n7036 & n7848 ;
  assign n28904 = ~n466 & n2926 ;
  assign n28905 = ~n28903 & n28904 ;
  assign n28906 = n15311 & ~n28905 ;
  assign n28907 = ( n5173 & n17817 ) | ( n5173 & ~n28906 ) | ( n17817 & ~n28906 ) ;
  assign n28910 = n6805 ^ n6205 ^ n2436 ;
  assign n28908 = n1964 & ~n21696 ;
  assign n28909 = ~n6471 & n28908 ;
  assign n28911 = n28910 ^ n28909 ^ 1'b0 ;
  assign n28912 = n20298 ^ n6206 ^ 1'b0 ;
  assign n28913 = n7557 & ~n27739 ;
  assign n28914 = n4997 | n28913 ;
  assign n28915 = n23646 & ~n28914 ;
  assign n28916 = n20586 ^ n5065 ^ 1'b0 ;
  assign n28917 = n8234 | n28916 ;
  assign n28918 = n16391 ^ n10316 ^ 1'b0 ;
  assign n28919 = n27194 ^ n18277 ^ 1'b0 ;
  assign n28920 = n9193 ^ n4778 ^ 1'b0 ;
  assign n28921 = n11204 | n26495 ;
  assign n28922 = n20191 ^ n15902 ^ 1'b0 ;
  assign n28923 = ~n1992 & n28922 ;
  assign n28924 = n27899 ^ n13678 ^ 1'b0 ;
  assign n28925 = n6950 ^ n4374 ^ 1'b0 ;
  assign n28926 = n28925 ^ n14081 ^ 1'b0 ;
  assign n28927 = ( n24159 & ~n24805 ) | ( n24159 & n28926 ) | ( ~n24805 & n28926 ) ;
  assign n28928 = n10401 | n14956 ;
  assign n28929 = n25374 | n28928 ;
  assign n28930 = ~n7736 & n22810 ;
  assign n28931 = n20960 & ~n28930 ;
  assign n28932 = n21676 ^ n5598 ^ 1'b0 ;
  assign n28933 = n16977 ^ n12610 ^ 1'b0 ;
  assign n28934 = n20455 ^ n17979 ^ 1'b0 ;
  assign n28935 = n6286 & n22675 ;
  assign n28936 = n3588 & ~n5896 ;
  assign n28937 = ( n3012 & n15389 ) | ( n3012 & n28936 ) | ( n15389 & n28936 ) ;
  assign n28938 = n3513 | n28937 ;
  assign n28939 = n2724 & n7597 ;
  assign n28940 = ~n14048 & n18899 ;
  assign n28941 = n1522 & n2625 ;
  assign n28942 = n9747 & ~n28941 ;
  assign n28943 = n28942 ^ n9811 ^ n5812 ;
  assign n28944 = n1032 & n24644 ;
  assign n28945 = n407 ^ n291 ^ 1'b0 ;
  assign n28946 = n8645 & ~n28945 ;
  assign n28947 = n28946 ^ n10361 ^ 1'b0 ;
  assign n28948 = n13998 & n28947 ;
  assign n28949 = n28948 ^ n10443 ^ 1'b0 ;
  assign n28950 = ~n25002 & n28949 ;
  assign n28951 = n15315 & n27689 ;
  assign n28952 = n28951 ^ n13202 ^ 1'b0 ;
  assign n28953 = ( n6531 & n9063 ) | ( n6531 & ~n14688 ) | ( n9063 & ~n14688 ) ;
  assign n28954 = ~n17316 & n28953 ;
  assign n28955 = n20034 ^ n19379 ^ 1'b0 ;
  assign n28956 = n10914 ^ x184 ^ 1'b0 ;
  assign n28957 = n26409 & n28956 ;
  assign n28958 = n11564 & n14836 ;
  assign n28959 = n19417 ^ n3218 ^ 1'b0 ;
  assign n28960 = ~n5602 & n24375 ;
  assign n28961 = n14347 ^ n5619 ^ 1'b0 ;
  assign n28962 = n20392 | n28961 ;
  assign n28963 = n28960 & ~n28962 ;
  assign n28964 = n28963 ^ n15308 ^ 1'b0 ;
  assign n28965 = n22641 ^ n10768 ^ 1'b0 ;
  assign n28966 = n18056 & n28965 ;
  assign n28967 = n6957 | n15759 ;
  assign n28968 = n11737 & n15843 ;
  assign n28969 = n7022 & n14049 ;
  assign n28970 = n2655 & ~n5932 ;
  assign n28971 = n14437 ^ n997 ^ 1'b0 ;
  assign n28972 = ( n5646 & n28970 ) | ( n5646 & n28971 ) | ( n28970 & n28971 ) ;
  assign n28973 = n20910 | n25569 ;
  assign n28974 = n2394 | n5317 ;
  assign n28975 = n22123 & ~n28974 ;
  assign n28976 = n12622 | n28975 ;
  assign n28977 = n1730 | n28976 ;
  assign n28978 = n28977 ^ n10193 ^ 1'b0 ;
  assign n28979 = n17762 ^ n13221 ^ 1'b0 ;
  assign n28980 = n11763 | n28979 ;
  assign n28981 = n20358 | n28980 ;
  assign n28982 = n14655 ^ n1968 ^ 1'b0 ;
  assign n28983 = n491 | n28982 ;
  assign n28984 = n2164 | n28983 ;
  assign n28985 = x5 & n5058 ;
  assign n28986 = ~x5 & n28985 ;
  assign n28987 = n310 & ~n2681 ;
  assign n28988 = ~n310 & n28987 ;
  assign n28989 = n28986 | n28988 ;
  assign n28990 = ~n6413 & n8256 ;
  assign n28991 = ( ~n1615 & n9569 ) | ( ~n1615 & n28990 ) | ( n9569 & n28990 ) ;
  assign n28992 = n28991 ^ n28861 ^ n23690 ;
  assign n28993 = ( ~n4208 & n28989 ) | ( ~n4208 & n28992 ) | ( n28989 & n28992 ) ;
  assign n28994 = ~n17619 & n19503 ;
  assign n28995 = n992 & n28994 ;
  assign n28996 = n14526 & ~n27271 ;
  assign n28997 = n4721 & n14006 ;
  assign n28998 = n3690 & n8867 ;
  assign n28999 = n8198 ^ n6332 ^ 1'b0 ;
  assign n29000 = n28999 ^ n2953 ^ x54 ;
  assign n29001 = n28998 & ~n29000 ;
  assign n29002 = n16415 & ~n29001 ;
  assign n29003 = n12101 ^ n2097 ^ 1'b0 ;
  assign n29004 = n7579 | n15718 ;
  assign n29005 = ~n29003 & n29004 ;
  assign n29006 = n2073 ^ n575 ^ 1'b0 ;
  assign n29007 = ~n13098 & n29006 ;
  assign n29010 = n13171 ^ n11135 ^ 1'b0 ;
  assign n29008 = n11449 ^ n1905 ^ 1'b0 ;
  assign n29009 = n9105 & ~n29008 ;
  assign n29011 = n29010 ^ n29009 ^ n5066 ;
  assign n29012 = n28830 ^ n3431 ^ 1'b0 ;
  assign n29013 = n7674 | n29012 ;
  assign n29014 = n29011 & ~n29013 ;
  assign n29015 = ( n19195 & n29007 ) | ( n19195 & n29014 ) | ( n29007 & n29014 ) ;
  assign n29016 = x251 & ~n5496 ;
  assign n29017 = ~n24404 & n29016 ;
  assign n29018 = ~n2370 & n29017 ;
  assign n29019 = n3106 & n25577 ;
  assign n29020 = ~n6632 & n29019 ;
  assign n29021 = n9872 ^ n5442 ^ 1'b0 ;
  assign n29022 = x195 & n19671 ;
  assign n29023 = n8346 | n29022 ;
  assign n29024 = n11807 & n15850 ;
  assign n29025 = n5683 & n29024 ;
  assign n29026 = n29025 ^ n23208 ^ 1'b0 ;
  assign n29027 = n16545 & ~n29026 ;
  assign n29028 = n17811 ^ n14522 ^ n12238 ;
  assign n29029 = n29028 ^ n5168 ^ 1'b0 ;
  assign n29030 = n15543 ^ n943 ^ 1'b0 ;
  assign n29031 = x61 & ~n5278 ;
  assign n29032 = n8814 & ~n29031 ;
  assign n29033 = n20328 & n29032 ;
  assign n29034 = n29033 ^ n423 ^ 1'b0 ;
  assign n29035 = n10187 | n16430 ;
  assign n29036 = ~x92 & n15310 ;
  assign n29037 = n4634 & n7743 ;
  assign n29038 = n5587 & ~n8785 ;
  assign n29039 = n29038 ^ n7962 ^ 1'b0 ;
  assign n29040 = ( ~n7637 & n29037 ) | ( ~n7637 & n29039 ) | ( n29037 & n29039 ) ;
  assign n29041 = n6163 & ~n29040 ;
  assign n29042 = n5009 & n6193 ;
  assign n29043 = n5856 & n29042 ;
  assign n29044 = n29043 ^ n2580 ^ 1'b0 ;
  assign n29045 = x115 | n5859 ;
  assign n29046 = n2879 | n29045 ;
  assign n29047 = ~n1614 & n29046 ;
  assign n29048 = n19702 ^ n6687 ^ 1'b0 ;
  assign n29049 = n6157 & n29048 ;
  assign n29050 = ( n3805 & n9961 ) | ( n3805 & ~n29049 ) | ( n9961 & ~n29049 ) ;
  assign n29051 = ~n14389 & n29050 ;
  assign n29052 = n22707 & n25789 ;
  assign n29053 = n6206 & n14742 ;
  assign n29054 = n2613 & n29053 ;
  assign n29055 = ( n4222 & n23957 ) | ( n4222 & ~n29054 ) | ( n23957 & ~n29054 ) ;
  assign n29056 = n29055 ^ n14929 ^ n1307 ;
  assign n29057 = n29056 ^ n26128 ^ 1'b0 ;
  assign n29058 = ~n1544 & n4095 ;
  assign n29059 = ~n28409 & n29058 ;
  assign n29060 = n17238 | n26639 ;
  assign n29061 = n29059 & ~n29060 ;
  assign n29062 = n20633 | n29061 ;
  assign n29063 = n8414 & ~n10414 ;
  assign n29064 = n12646 & n29063 ;
  assign n29065 = n1437 & ~n12065 ;
  assign n29066 = n3790 | n29065 ;
  assign n29067 = x120 | n18528 ;
  assign n29068 = n6195 | n29067 ;
  assign n29069 = n23161 & ~n29068 ;
  assign n29070 = n5725 ^ n263 ^ 1'b0 ;
  assign n29071 = n22521 ^ n22327 ^ 1'b0 ;
  assign n29072 = n29070 | n29071 ;
  assign n29073 = ( n10120 & n13657 ) | ( n10120 & n20831 ) | ( n13657 & n20831 ) ;
  assign n29074 = ~n9202 & n13204 ;
  assign n29075 = n1884 & n3218 ;
  assign n29076 = n2817 & n29075 ;
  assign n29077 = n635 & n4323 ;
  assign n29078 = n5060 | n29077 ;
  assign n29079 = n3271 & n6701 ;
  assign n29080 = n29079 ^ n3271 ^ 1'b0 ;
  assign n29081 = n4589 & ~n21708 ;
  assign n29082 = n5069 | n19574 ;
  assign n29083 = n11608 | n29082 ;
  assign n29084 = n26312 & ~n29083 ;
  assign n29085 = n29081 & ~n29084 ;
  assign n29086 = ( ~n2775 & n6830 ) | ( ~n2775 & n20809 ) | ( n6830 & n20809 ) ;
  assign n29087 = n4269 ^ n1010 ^ 1'b0 ;
  assign n29088 = n8330 & ~n29087 ;
  assign n29090 = n2155 & ~n3139 ;
  assign n29091 = ~n1144 & n29090 ;
  assign n29089 = n15567 | n16851 ;
  assign n29092 = n29091 ^ n29089 ^ 1'b0 ;
  assign n29093 = n29088 | n29092 ;
  assign n29094 = n12339 | n19610 ;
  assign n29095 = n23636 & ~n29094 ;
  assign n29096 = ~n11735 & n12276 ;
  assign n29097 = n29096 ^ n28643 ^ 1'b0 ;
  assign n29099 = n15300 ^ n6527 ^ 1'b0 ;
  assign n29098 = n7197 & n19747 ;
  assign n29100 = n29099 ^ n29098 ^ 1'b0 ;
  assign n29101 = ~n29097 & n29100 ;
  assign n29102 = n4596 & ~n27569 ;
  assign n29103 = n14062 ^ n1160 ^ 1'b0 ;
  assign n29104 = n2545 & n29103 ;
  assign n29105 = n10174 & n15026 ;
  assign n29106 = n14565 ^ n12826 ^ 1'b0 ;
  assign n29107 = n16796 & n29106 ;
  assign n29108 = ~n1037 & n2946 ;
  assign n29109 = n22376 ^ n1237 ^ 1'b0 ;
  assign n29111 = n14559 | n24478 ;
  assign n29110 = n14111 ^ n6024 ^ 1'b0 ;
  assign n29112 = n29111 ^ n29110 ^ n10062 ;
  assign n29113 = n4166 | n16031 ;
  assign n29114 = n12515 | n29113 ;
  assign n29115 = n1137 | n12819 ;
  assign n29116 = n4642 & n29115 ;
  assign n29117 = n17577 ^ n6869 ^ n5523 ;
  assign n29118 = n26740 ^ n3213 ^ 1'b0 ;
  assign n29119 = n529 | n1915 ;
  assign n29120 = n29119 ^ n20644 ^ 1'b0 ;
  assign n29121 = ~n15080 & n29120 ;
  assign n29122 = n4449 & ~n13682 ;
  assign n29123 = ( n3382 & n4029 ) | ( n3382 & ~n29122 ) | ( n4029 & ~n29122 ) ;
  assign n29124 = n24781 ^ n6433 ^ 1'b0 ;
  assign n29125 = n20915 | n29124 ;
  assign n29126 = n3266 | n23346 ;
  assign n29127 = n19588 & ~n29126 ;
  assign n29128 = n22076 ^ n847 ^ 1'b0 ;
  assign n29129 = n6187 | n10663 ;
  assign n29130 = n29128 | n29129 ;
  assign n29131 = ~n25556 & n29130 ;
  assign n29132 = ~n8141 & n29131 ;
  assign n29133 = n21169 ^ n1820 ^ 1'b0 ;
  assign n29134 = ~n11551 & n22505 ;
  assign n29135 = ~n2704 & n29134 ;
  assign n29136 = n29135 ^ n23215 ^ 1'b0 ;
  assign n29137 = n20183 ^ n5752 ^ 1'b0 ;
  assign n29138 = n4124 | n29137 ;
  assign n29139 = n3231 & n19963 ;
  assign n29140 = n29139 ^ n23199 ^ 1'b0 ;
  assign n29141 = n7366 | n20625 ;
  assign n29142 = n1338 | n29141 ;
  assign n29143 = n6632 | n19335 ;
  assign n29144 = n23538 & ~n29143 ;
  assign n29148 = n12463 ^ n5773 ^ 1'b0 ;
  assign n29149 = ~n10864 & n29148 ;
  assign n29145 = n3682 & n16990 ;
  assign n29146 = n13962 & n29145 ;
  assign n29147 = ~n8250 & n29146 ;
  assign n29150 = n29149 ^ n29147 ^ n16145 ;
  assign n29151 = n1219 | n29150 ;
  assign n29152 = n29151 ^ n2924 ^ 1'b0 ;
  assign n29153 = n17457 ^ n4197 ^ 1'b0 ;
  assign n29154 = ~n7294 & n29153 ;
  assign n29155 = n5110 & n29154 ;
  assign n29156 = ( n3240 & n7791 ) | ( n3240 & n19559 ) | ( n7791 & n19559 ) ;
  assign n29157 = n10814 & n18756 ;
  assign n29158 = ~n6148 & n14533 ;
  assign n29159 = n6376 ^ n1838 ^ 1'b0 ;
  assign n29160 = n25462 | n29159 ;
  assign n29161 = n29160 ^ n17202 ^ 1'b0 ;
  assign n29164 = n11237 & ~n22740 ;
  assign n29162 = ( ~x107 & x150 ) | ( ~x107 & n5796 ) | ( x150 & n5796 ) ;
  assign n29163 = n10057 & n29162 ;
  assign n29165 = n29164 ^ n29163 ^ 1'b0 ;
  assign n29166 = n25206 ^ n9735 ^ 1'b0 ;
  assign n29167 = n7683 & ~n25327 ;
  assign n29168 = n29167 ^ n4441 ^ 1'b0 ;
  assign n29169 = n29168 ^ n10051 ^ 1'b0 ;
  assign n29170 = n11981 & n17199 ;
  assign n29171 = ~n6983 & n29170 ;
  assign n29172 = n9521 | n26508 ;
  assign n29173 = n29171 & ~n29172 ;
  assign n29174 = n675 & ~n12922 ;
  assign n29175 = n29174 ^ n9241 ^ 1'b0 ;
  assign n29176 = n3159 | n29175 ;
  assign n29177 = n29176 ^ n6005 ^ 1'b0 ;
  assign n29178 = ~n5009 & n12627 ;
  assign n29179 = n21057 ^ n17737 ^ 1'b0 ;
  assign n29180 = n4837 & n29179 ;
  assign n29181 = ~n22310 & n29180 ;
  assign n29182 = n16331 & n29181 ;
  assign n29183 = n7992 & n22028 ;
  assign n29184 = n29183 ^ n1121 ^ 1'b0 ;
  assign n29185 = n27472 ^ n13604 ^ 1'b0 ;
  assign n29186 = n12338 ^ n3465 ^ 1'b0 ;
  assign n29187 = ~n22527 & n29186 ;
  assign n29190 = n10857 & n20113 ;
  assign n29188 = ~n4154 & n10022 ;
  assign n29189 = n1219 & n29188 ;
  assign n29191 = n29190 ^ n29189 ^ 1'b0 ;
  assign n29192 = n5750 ^ n1495 ^ 1'b0 ;
  assign n29193 = n13327 & n29192 ;
  assign n29194 = n13225 & n29193 ;
  assign n29195 = n27382 ^ n20165 ^ 1'b0 ;
  assign n29196 = n4086 | n15730 ;
  assign n29197 = n3805 & ~n29196 ;
  assign n29198 = ~n6216 & n28684 ;
  assign n29200 = n1001 & ~n15504 ;
  assign n29201 = n15504 & n29200 ;
  assign n29199 = n930 & n10322 ;
  assign n29202 = n29201 ^ n29199 ^ 1'b0 ;
  assign n29203 = ( ~x50 & n7130 ) | ( ~x50 & n29202 ) | ( n7130 & n29202 ) ;
  assign n29204 = ( n22035 & n23678 ) | ( n22035 & ~n29203 ) | ( n23678 & ~n29203 ) ;
  assign n29205 = n9886 & ~n17054 ;
  assign n29206 = ~n2589 & n29205 ;
  assign n29207 = n20270 & ~n29206 ;
  assign n29208 = n18229 ^ n10240 ^ 1'b0 ;
  assign n29209 = n29208 ^ n26395 ^ 1'b0 ;
  assign n29210 = n4906 & ~n29209 ;
  assign n29211 = n29210 ^ n5342 ^ 1'b0 ;
  assign n29212 = n2509 & n3942 ;
  assign n29213 = ~n17974 & n29212 ;
  assign n29214 = n28614 ^ n4307 ^ 1'b0 ;
  assign n29215 = n6737 | n7521 ;
  assign n29216 = n23885 ^ n14150 ^ 1'b0 ;
  assign n29217 = n29215 | n29216 ;
  assign n29219 = n2403 | n3889 ;
  assign n29218 = n5402 & n17692 ;
  assign n29220 = n29219 ^ n29218 ^ 1'b0 ;
  assign n29221 = n29220 ^ n7173 ^ 1'b0 ;
  assign n29222 = n5713 & n29221 ;
  assign n29223 = n16521 & n29222 ;
  assign n29224 = n13803 ^ n6950 ^ 1'b0 ;
  assign n29225 = ( n5913 & n14067 ) | ( n5913 & ~n29224 ) | ( n14067 & ~n29224 ) ;
  assign n29226 = n15845 | n27347 ;
  assign n29227 = n11476 ^ n5392 ^ 1'b0 ;
  assign n29228 = ( ~n4970 & n11292 ) | ( ~n4970 & n29227 ) | ( n11292 & n29227 ) ;
  assign n29229 = n27750 & n29228 ;
  assign n29230 = ~n8333 & n29229 ;
  assign n29231 = n20855 ^ n8989 ^ 1'b0 ;
  assign n29232 = n29231 ^ n19308 ^ n4157 ;
  assign n29233 = n1077 & ~n15948 ;
  assign n29234 = n14589 & n29233 ;
  assign n29235 = ( n1259 & n12338 ) | ( n1259 & ~n29234 ) | ( n12338 & ~n29234 ) ;
  assign n29238 = n13767 & ~n18009 ;
  assign n29236 = ~n2397 & n2988 ;
  assign n29237 = ~n4181 & n29236 ;
  assign n29239 = n29238 ^ n29237 ^ 1'b0 ;
  assign n29240 = ~n1465 & n7624 ;
  assign n29241 = ~n29239 & n29240 ;
  assign n29242 = n29241 ^ n12054 ^ 1'b0 ;
  assign n29243 = ~n18915 & n29242 ;
  assign n29244 = ~n19777 & n29243 ;
  assign n29245 = ~n1384 & n6842 ;
  assign n29246 = n29244 & n29245 ;
  assign n29247 = n7329 ^ n5322 ^ 1'b0 ;
  assign n29248 = n14158 & n14614 ;
  assign n29249 = x146 & n2465 ;
  assign n29250 = n29249 ^ n882 ^ 1'b0 ;
  assign n29251 = ~n7586 & n29250 ;
  assign n29252 = n20536 ^ n8267 ^ 1'b0 ;
  assign n29253 = n9522 & ~n29252 ;
  assign n29254 = n29253 ^ n20435 ^ 1'b0 ;
  assign n29255 = n18196 ^ n7107 ^ 1'b0 ;
  assign n29256 = ~n3828 & n4515 ;
  assign n29257 = n10131 & n29256 ;
  assign n29258 = n3419 | n29257 ;
  assign n29259 = n29258 ^ n1634 ^ 1'b0 ;
  assign n29260 = n3702 & ~n4493 ;
  assign n29261 = n29260 ^ n1083 ^ 1'b0 ;
  assign n29262 = n29261 ^ n14767 ^ 1'b0 ;
  assign n29263 = ( n8874 & ~n9864 ) | ( n8874 & n21237 ) | ( ~n9864 & n21237 ) ;
  assign n29264 = n8994 ^ n7402 ^ 1'b0 ;
  assign n29265 = n29264 ^ n17758 ^ 1'b0 ;
  assign n29266 = ~n1864 & n29265 ;
  assign n29267 = n2694 | n11430 ;
  assign n29268 = ~n14352 & n18016 ;
  assign n29269 = n29267 & n29268 ;
  assign n29270 = n5771 | n29269 ;
  assign n29271 = n29270 ^ n8728 ^ 1'b0 ;
  assign n29272 = n1271 | n21485 ;
  assign n29273 = n29272 ^ n16356 ^ 1'b0 ;
  assign n29274 = ~n17457 & n29273 ;
  assign n29275 = n12070 ^ n3142 ^ 1'b0 ;
  assign n29276 = n5127 & n29275 ;
  assign n29277 = n5772 | n25637 ;
  assign n29279 = ~n2301 & n15357 ;
  assign n29278 = n3106 & n9515 ;
  assign n29280 = n29279 ^ n29278 ^ 1'b0 ;
  assign n29281 = n518 & n27799 ;
  assign n29282 = n29281 ^ n25715 ^ n7070 ;
  assign n29283 = n15719 & ~n29282 ;
  assign n29284 = n6391 & ~n19591 ;
  assign n29285 = ~n6186 & n29284 ;
  assign n29286 = n306 & ~n29285 ;
  assign n29287 = n11795 & n19529 ;
  assign n29288 = n23083 & n29287 ;
  assign n29289 = ( n8360 & n8694 ) | ( n8360 & ~n11990 ) | ( n8694 & ~n11990 ) ;
  assign n29290 = n27645 ^ n16986 ^ 1'b0 ;
  assign n29291 = n29289 | n29290 ;
  assign n29292 = n29291 ^ n2783 ^ 1'b0 ;
  assign n29293 = n1627 & ~n8391 ;
  assign n29294 = n29293 ^ n11389 ^ 1'b0 ;
  assign n29295 = n12143 ^ n6479 ^ 1'b0 ;
  assign n29296 = n10229 & n29295 ;
  assign n29297 = n5374 & n29296 ;
  assign n29298 = n27184 ^ n15765 ^ 1'b0 ;
  assign n29299 = n24934 ^ n18102 ^ 1'b0 ;
  assign n29300 = n24258 & n29299 ;
  assign n29301 = ~n10684 & n29300 ;
  assign n29302 = n22206 ^ n12958 ^ 1'b0 ;
  assign n29303 = n18796 & ~n24101 ;
  assign n29304 = n29303 ^ n26787 ^ n20631 ;
  assign n29305 = ( n2904 & n3496 ) | ( n2904 & n4499 ) | ( n3496 & n4499 ) ;
  assign n29306 = x176 | n14291 ;
  assign n29307 = n16035 ^ n1397 ^ 1'b0 ;
  assign n29308 = n19475 ^ n8219 ^ 1'b0 ;
  assign n29309 = n12732 ^ n2155 ^ 1'b0 ;
  assign n29310 = n28445 | n29309 ;
  assign n29311 = n9644 & n24431 ;
  assign n29312 = n4954 & n29311 ;
  assign n29316 = ( n938 & n1589 ) | ( n938 & n5783 ) | ( n1589 & n5783 ) ;
  assign n29317 = ~n9355 & n29316 ;
  assign n29318 = n29317 ^ n4640 ^ 1'b0 ;
  assign n29313 = n2489 | n8117 ;
  assign n29314 = n29313 ^ x80 ^ 1'b0 ;
  assign n29315 = n10218 & n29314 ;
  assign n29319 = n29318 ^ n29315 ^ 1'b0 ;
  assign n29320 = n29319 ^ n1344 ^ 1'b0 ;
  assign n29321 = n9413 | n17962 ;
  assign n29322 = n29321 ^ n5342 ^ 1'b0 ;
  assign n29324 = ( ~n12499 & n13580 ) | ( ~n12499 & n17526 ) | ( n13580 & n17526 ) ;
  assign n29323 = n4992 | n28623 ;
  assign n29325 = n29324 ^ n29323 ^ 1'b0 ;
  assign n29326 = n22181 ^ n20103 ^ 1'b0 ;
  assign n29327 = n26931 & n29326 ;
  assign n29328 = n29327 ^ n24281 ^ 1'b0 ;
  assign n29329 = n5623 ^ n5410 ^ 1'b0 ;
  assign n29330 = n22629 ^ n11692 ^ n8594 ;
  assign n29331 = ~n2193 & n12336 ;
  assign n29332 = n11467 & n29331 ;
  assign n29333 = ( ~n2861 & n20081 ) | ( ~n2861 & n29332 ) | ( n20081 & n29332 ) ;
  assign n29334 = n404 | n12782 ;
  assign n29335 = n24438 & n29334 ;
  assign n29336 = n5659 | n8619 ;
  assign n29337 = n26222 ^ n1378 ^ 1'b0 ;
  assign n29338 = n14415 ^ n7300 ^ n1855 ;
  assign n29339 = n19157 ^ n6327 ^ 1'b0 ;
  assign n29340 = ~n1276 & n14448 ;
  assign n29341 = ~n4951 & n29340 ;
  assign n29342 = n3726 ^ n1699 ^ 1'b0 ;
  assign n29343 = ~n29341 & n29342 ;
  assign n29344 = n23184 ^ n10674 ^ 1'b0 ;
  assign n29345 = n29286 & ~n29344 ;
  assign n29346 = n4066 | n13483 ;
  assign n29347 = ~n29286 & n29346 ;
  assign n29348 = n13110 ^ n649 ^ 1'b0 ;
  assign n29349 = ~n15889 & n27027 ;
  assign n29350 = ~n8234 & n29349 ;
  assign n29351 = ~n16681 & n18764 ;
  assign n29352 = n2925 & ~n16385 ;
  assign n29353 = n29352 ^ n19576 ^ n16018 ;
  assign n29354 = n16941 & n25958 ;
  assign n29355 = n29354 ^ n16810 ^ 1'b0 ;
  assign n29356 = ~n10805 & n15789 ;
  assign n29357 = n4458 ^ n3574 ^ 1'b0 ;
  assign n29358 = n27138 & n29357 ;
  assign n29359 = n2574 ^ n2431 ^ 1'b0 ;
  assign n29360 = ~n14128 & n29359 ;
  assign n29361 = n7257 & ~n10719 ;
  assign n29369 = x129 & n1486 ;
  assign n29370 = ~n3474 & n29369 ;
  assign n29371 = n5429 | n29370 ;
  assign n29372 = n29371 ^ n858 ^ 1'b0 ;
  assign n29373 = ~n20877 & n29372 ;
  assign n29374 = n29373 ^ n28232 ^ 1'b0 ;
  assign n29375 = n4737 | n29374 ;
  assign n29364 = n24967 ^ n15884 ^ 1'b0 ;
  assign n29365 = n12874 & n29364 ;
  assign n29366 = ~n12874 & n29365 ;
  assign n29362 = n6370 & ~n16336 ;
  assign n29363 = ~n3745 & n29362 ;
  assign n29367 = n29366 ^ n29363 ^ n14156 ;
  assign n29368 = ~n13571 & n29367 ;
  assign n29376 = n29375 ^ n29368 ^ 1'b0 ;
  assign n29377 = n14987 ^ n6817 ^ 1'b0 ;
  assign n29378 = n29377 ^ n7184 ^ 1'b0 ;
  assign n29379 = n14147 ^ n2469 ^ 1'b0 ;
  assign n29380 = n632 & n2980 ;
  assign n29381 = n29380 ^ n21812 ^ 1'b0 ;
  assign n29382 = n10840 | n29381 ;
  assign n29383 = ~n9560 & n14526 ;
  assign n29384 = ( n14807 & n16191 ) | ( n14807 & ~n18948 ) | ( n16191 & ~n18948 ) ;
  assign n29385 = ( n16953 & ~n21462 ) | ( n16953 & n29384 ) | ( ~n21462 & n29384 ) ;
  assign n29386 = n7489 | n29385 ;
  assign n29387 = n29383 & ~n29386 ;
  assign n29388 = n22845 ^ n634 ^ 1'b0 ;
  assign n29389 = n11863 | n29388 ;
  assign n29390 = ( ~x78 & n11386 ) | ( ~x78 & n17159 ) | ( n11386 & n17159 ) ;
  assign n29391 = x39 | n15952 ;
  assign n29392 = n20908 ^ n3494 ^ 1'b0 ;
  assign n29393 = n29392 ^ n6891 ^ n2047 ;
  assign n29394 = n29393 ^ n23091 ^ 1'b0 ;
  assign n29395 = n15877 ^ n12074 ^ 1'b0 ;
  assign n29396 = n2638 | n29395 ;
  assign n29397 = n7871 & ~n25109 ;
  assign n29398 = n29396 & n29397 ;
  assign n29399 = n10655 & ~n13695 ;
  assign n29400 = ~n26056 & n29399 ;
  assign n29401 = n29400 ^ n27201 ^ 1'b0 ;
  assign n29402 = n4527 | n6897 ;
  assign n29403 = n28226 ^ n14458 ^ 1'b0 ;
  assign n29404 = ~n12513 & n29403 ;
  assign n29405 = n29404 ^ n10363 ^ n466 ;
  assign n29406 = ~n1648 & n2331 ;
  assign n29407 = ~n14071 & n29406 ;
  assign n29408 = n26588 ^ n7660 ^ 1'b0 ;
  assign n29409 = x246 & n29408 ;
  assign n29410 = n29407 & n29409 ;
  assign n29411 = n11590 & ~n21428 ;
  assign n29413 = n13830 | n20776 ;
  assign n29414 = n6499 | n29413 ;
  assign n29412 = ~n16489 & n16549 ;
  assign n29415 = n29414 ^ n29412 ^ 1'b0 ;
  assign n29416 = n7013 ^ n6883 ^ 1'b0 ;
  assign n29417 = ~n6456 & n29416 ;
  assign n29418 = n20303 & ~n29417 ;
  assign n29419 = ~n11622 & n12226 ;
  assign n29420 = n18357 & ~n29419 ;
  assign n29421 = n4525 & ~n29420 ;
  assign n29422 = n24155 ^ n2845 ^ 1'b0 ;
  assign n29423 = ( n12242 & ~n13324 ) | ( n12242 & n24915 ) | ( ~n13324 & n24915 ) ;
  assign n29424 = ~n2602 & n14815 ;
  assign n29425 = n29423 & n29424 ;
  assign n29426 = n24372 ^ n13765 ^ n13338 ;
  assign n29427 = ~n13053 & n13429 ;
  assign n29428 = n4325 ^ n1189 ^ 1'b0 ;
  assign n29429 = n752 | n2139 ;
  assign n29430 = n2139 & ~n29429 ;
  assign n29431 = n749 & ~n29430 ;
  assign n29432 = n29430 & n29431 ;
  assign n29433 = n4225 | n29432 ;
  assign n29434 = n4225 & ~n29433 ;
  assign n29435 = n29434 ^ n19512 ^ 1'b0 ;
  assign n29436 = n12379 | n29435 ;
  assign n29437 = n29436 ^ n20381 ^ 1'b0 ;
  assign n29438 = n29428 | n29437 ;
  assign n29439 = ~n507 & n11563 ;
  assign n29440 = n29439 ^ n27220 ^ 1'b0 ;
  assign n29441 = n7251 & n17266 ;
  assign n29442 = n2844 & n29441 ;
  assign n29443 = n22349 | n23426 ;
  assign n29444 = n12625 & ~n13202 ;
  assign n29445 = n29444 ^ n28281 ^ n10395 ;
  assign n29446 = n29445 ^ n2487 ^ 1'b0 ;
  assign n29447 = n7838 | n11181 ;
  assign n29448 = ~n24063 & n29447 ;
  assign n29449 = n29448 ^ n11227 ^ 1'b0 ;
  assign n29450 = n7158 & n8023 ;
  assign n29451 = n23632 & n29450 ;
  assign n29452 = n29451 ^ n6937 ^ 1'b0 ;
  assign n29453 = ~n11336 & n12838 ;
  assign n29454 = n7791 & n29453 ;
  assign n29455 = n12585 & n29454 ;
  assign n29456 = n29455 ^ n3249 ^ 1'b0 ;
  assign n29457 = n5696 & ~n17430 ;
  assign n29458 = n18850 ^ n6307 ^ 1'b0 ;
  assign n29459 = n22726 | n29458 ;
  assign n29460 = n22522 ^ n4125 ^ 1'b0 ;
  assign n29461 = ~n18608 & n29460 ;
  assign n29462 = n675 & n13765 ;
  assign n29463 = n21881 ^ n17430 ^ 1'b0 ;
  assign n29464 = n2785 & n3133 ;
  assign n29465 = n16010 & ~n29464 ;
  assign n29466 = n7958 & ~n21428 ;
  assign n29467 = n5798 & n29466 ;
  assign n29468 = ~n485 & n22995 ;
  assign n29469 = n26606 & n29468 ;
  assign n29470 = n2443 & ~n25029 ;
  assign n29471 = ~n2443 & n29470 ;
  assign n29472 = n3223 & ~n10900 ;
  assign n29473 = n10900 & n29472 ;
  assign n29474 = n29473 ^ n12591 ^ n2956 ;
  assign n29475 = n7423 & ~n29474 ;
  assign n29476 = n29471 & n29475 ;
  assign n29477 = n15596 & n24633 ;
  assign n29478 = n2633 & n9009 ;
  assign n29479 = n9774 & n29478 ;
  assign n29480 = n7195 | n10402 ;
  assign n29481 = n29479 & n29480 ;
  assign n29482 = n28809 ^ n11650 ^ 1'b0 ;
  assign n29483 = ( ~n4770 & n10229 ) | ( ~n4770 & n29482 ) | ( n10229 & n29482 ) ;
  assign n29484 = n3622 | n17651 ;
  assign n29485 = n29484 ^ n6853 ^ 1'b0 ;
  assign n29486 = ~n771 & n10364 ;
  assign n29487 = n2167 & n29486 ;
  assign n29488 = n14767 ^ n12656 ^ 1'b0 ;
  assign n29489 = n8096 & n29488 ;
  assign n29490 = n4826 | n13958 ;
  assign n29491 = n13390 ^ n4142 ^ 1'b0 ;
  assign n29492 = n29490 | n29491 ;
  assign n29493 = n17858 & ~n25551 ;
  assign n29494 = n29493 ^ n1864 ^ 1'b0 ;
  assign n29495 = ~n20452 & n29494 ;
  assign n29496 = n10674 & n29495 ;
  assign n29497 = n8600 & n23625 ;
  assign n29498 = ( n3670 & n25580 ) | ( n3670 & ~n29497 ) | ( n25580 & ~n29497 ) ;
  assign n29499 = n11568 & ~n14463 ;
  assign n29500 = ~n20364 & n29499 ;
  assign n29501 = n29500 ^ n17957 ^ 1'b0 ;
  assign n29502 = ~n26093 & n29501 ;
  assign n29503 = n29502 ^ n26892 ^ 1'b0 ;
  assign n29504 = ~n18530 & n29503 ;
  assign n29505 = n6818 | n9362 ;
  assign n29506 = n29505 ^ n8406 ^ 1'b0 ;
  assign n29507 = ~n26906 & n29506 ;
  assign n29508 = ~n14693 & n23061 ;
  assign n29509 = n5775 ^ n2721 ^ 1'b0 ;
  assign n29510 = n29508 | n29509 ;
  assign n29511 = ~n23846 & n29510 ;
  assign n29512 = n279 & n29511 ;
  assign n29513 = ( n2428 & n3823 ) | ( n2428 & n7858 ) | ( n3823 & n7858 ) ;
  assign n29514 = n16560 ^ n6454 ^ 1'b0 ;
  assign n29515 = n2343 & n29514 ;
  assign n29516 = n9350 & ~n9859 ;
  assign n29517 = n3468 ^ x56 ^ 1'b0 ;
  assign n29518 = n29517 ^ n23094 ^ 1'b0 ;
  assign n29519 = n1508 & ~n6539 ;
  assign n29520 = n29519 ^ n7929 ^ 1'b0 ;
  assign n29521 = n11537 ^ n3380 ^ 1'b0 ;
  assign n29522 = n20028 & n29521 ;
  assign n29523 = n11181 & ~n22675 ;
  assign n29524 = ( n12789 & ~n13699 ) | ( n12789 & n29523 ) | ( ~n13699 & n29523 ) ;
  assign n29525 = ( ~n5859 & n16756 ) | ( ~n5859 & n22798 ) | ( n16756 & n22798 ) ;
  assign n29526 = ~n12802 & n14027 ;
  assign n29527 = n29526 ^ n18565 ^ 1'b0 ;
  assign n29529 = n15434 | n19009 ;
  assign n29528 = ~n714 & n23511 ;
  assign n29530 = n29529 ^ n29528 ^ 1'b0 ;
  assign n29531 = ~n3184 & n14890 ;
  assign n29532 = n12487 & n17383 ;
  assign n29533 = n29532 ^ n25971 ^ 1'b0 ;
  assign n29534 = n4938 & n10490 ;
  assign n29535 = ~n3260 & n24633 ;
  assign n29536 = n29535 ^ n17681 ^ 1'b0 ;
  assign n29537 = ( ~n4114 & n29534 ) | ( ~n4114 & n29536 ) | ( n29534 & n29536 ) ;
  assign n29538 = n12548 ^ n12294 ^ 1'b0 ;
  assign n29539 = ( n15213 & n15639 ) | ( n15213 & n29538 ) | ( n15639 & n29538 ) ;
  assign n29540 = n29539 ^ n3982 ^ 1'b0 ;
  assign n29541 = n9155 ^ n1610 ^ 1'b0 ;
  assign n29542 = ~n883 & n29541 ;
  assign n29543 = ~n17752 & n29542 ;
  assign n29544 = n29543 ^ n10001 ^ 1'b0 ;
  assign n29545 = ( n479 & n3230 ) | ( n479 & n19529 ) | ( n3230 & n19529 ) ;
  assign n29546 = n5554 ^ n5124 ^ 1'b0 ;
  assign n29547 = n29546 ^ n3690 ^ 1'b0 ;
  assign n29548 = n9100 & n20877 ;
  assign n29549 = n9433 ^ n6202 ^ 1'b0 ;
  assign n29552 = ( n893 & n2400 ) | ( n893 & n3856 ) | ( n2400 & n3856 ) ;
  assign n29550 = n6106 & n11804 ;
  assign n29551 = n29550 ^ n10262 ^ 1'b0 ;
  assign n29553 = n29552 ^ n29551 ^ 1'b0 ;
  assign n29554 = n1983 & ~n10530 ;
  assign n29555 = n29554 ^ n7702 ^ 1'b0 ;
  assign n29556 = n11560 & ~n18658 ;
  assign n29557 = ~n12839 & n29556 ;
  assign n29558 = n6333 & n18828 ;
  assign n29559 = n29558 ^ n3486 ^ 1'b0 ;
  assign n29560 = n24182 & ~n29559 ;
  assign n29561 = n20243 ^ n7416 ^ 1'b0 ;
  assign n29565 = n21858 ^ n6873 ^ 1'b0 ;
  assign n29566 = n3760 | n9096 ;
  assign n29567 = n29565 & ~n29566 ;
  assign n29568 = n29567 ^ n17741 ^ 1'b0 ;
  assign n29569 = n29568 ^ n6581 ^ 1'b0 ;
  assign n29562 = ~n2482 & n7932 ;
  assign n29563 = n18092 & n23562 ;
  assign n29564 = n29562 & n29563 ;
  assign n29570 = n29569 ^ n29564 ^ n5581 ;
  assign n29571 = n7397 ^ n7195 ^ 1'b0 ;
  assign n29572 = n21860 ^ n8880 ^ 1'b0 ;
  assign n29573 = n9582 & n29572 ;
  assign n29574 = ~n4360 & n23451 ;
  assign n29575 = ~n29573 & n29574 ;
  assign n29576 = n29571 & n29575 ;
  assign n29577 = n6386 | n24038 ;
  assign n29578 = ( ~n9610 & n9758 ) | ( ~n9610 & n26449 ) | ( n9758 & n26449 ) ;
  assign n29579 = n29578 ^ n19959 ^ n11414 ;
  assign n29580 = n5182 & ~n29579 ;
  assign n29581 = ~n3346 & n29580 ;
  assign n29582 = n29577 & n29581 ;
  assign n29583 = n9669 | n14025 ;
  assign n29584 = n14025 & ~n29583 ;
  assign n29585 = n10673 ^ n8153 ^ 1'b0 ;
  assign n29586 = n8781 & ~n29585 ;
  assign n29588 = n5806 | n11437 ;
  assign n29589 = ~n5363 & n29588 ;
  assign n29587 = n6510 | n7839 ;
  assign n29590 = n29589 ^ n29587 ^ 1'b0 ;
  assign n29591 = n20485 & n29590 ;
  assign n29592 = ~n2127 & n19037 ;
  assign n29593 = n1784 & n7002 ;
  assign n29594 = n11640 & ~n29593 ;
  assign n29595 = n29594 ^ n21521 ^ 1'b0 ;
  assign n29596 = n29595 ^ n1695 ^ n1404 ;
  assign n29597 = n262 & ~n21282 ;
  assign n29598 = n29597 ^ n15577 ^ 1'b0 ;
  assign n29599 = n5772 & n14895 ;
  assign n29600 = n25319 & n29599 ;
  assign n29601 = n24648 ^ n20420 ^ 1'b0 ;
  assign n29602 = ~n5183 & n29601 ;
  assign n29603 = ~n5534 & n29602 ;
  assign n29604 = n29603 ^ n15877 ^ 1'b0 ;
  assign n29605 = ~n8733 & n13042 ;
  assign n29606 = n18938 | n29605 ;
  assign n29607 = n29604 & ~n29606 ;
  assign n29608 = n20761 ^ n16297 ^ 1'b0 ;
  assign n29609 = n3223 & n29608 ;
  assign n29610 = n9767 & ~n22443 ;
  assign n29611 = n8782 ^ n5885 ^ 1'b0 ;
  assign n29612 = n7580 ^ n6265 ^ 1'b0 ;
  assign n29613 = n6984 ^ n4905 ^ 1'b0 ;
  assign n29614 = n12247 | n29613 ;
  assign n29615 = n29614 ^ n569 ^ 1'b0 ;
  assign n29616 = n3413 ^ n2411 ^ 1'b0 ;
  assign n29617 = n9045 | n29616 ;
  assign n29618 = n7340 & ~n29617 ;
  assign n29619 = n2252 & n18472 ;
  assign n29620 = ( n2579 & n2825 ) | ( n2579 & ~n11730 ) | ( n2825 & ~n11730 ) ;
  assign n29621 = n1279 | n2268 ;
  assign n29622 = n2529 & ~n15721 ;
  assign n29623 = ~n1839 & n29622 ;
  assign n29624 = n8868 & ~n29623 ;
  assign n29625 = n29621 & n29624 ;
  assign n29626 = n29625 ^ n19466 ^ n5192 ;
  assign n29627 = n13880 ^ n2004 ^ 1'b0 ;
  assign n29628 = ~n18005 & n29627 ;
  assign n29629 = n29628 ^ n4325 ^ 1'b0 ;
  assign n29630 = n19988 ^ n682 ^ 1'b0 ;
  assign n29631 = n4337 & n12116 ;
  assign n29632 = ~n19285 & n29631 ;
  assign n29633 = n814 & n29632 ;
  assign n29637 = n3754 ^ n1442 ^ 1'b0 ;
  assign n29638 = n4566 & n29637 ;
  assign n29634 = n12733 ^ n1635 ^ 1'b0 ;
  assign n29635 = ~n27076 & n29634 ;
  assign n29636 = n16322 & n29635 ;
  assign n29639 = n29638 ^ n29636 ^ 1'b0 ;
  assign n29640 = n29566 ^ n2897 ^ 1'b0 ;
  assign n29641 = n29640 ^ n21713 ^ n13189 ;
  assign n29642 = n3814 & n26736 ;
  assign n29643 = n13761 ^ n943 ^ 1'b0 ;
  assign n29644 = n21626 ^ n15614 ^ 1'b0 ;
  assign n29645 = n3221 | n29644 ;
  assign n29646 = n4827 ^ n2712 ^ 1'b0 ;
  assign n29647 = n24391 ^ n22542 ^ 1'b0 ;
  assign n29648 = n23641 & ~n29647 ;
  assign n29649 = n2262 & ~n4488 ;
  assign n29650 = n29649 ^ n22812 ^ 1'b0 ;
  assign n29651 = n8423 ^ n2988 ^ 1'b0 ;
  assign n29652 = n29651 ^ n16393 ^ 1'b0 ;
  assign n29653 = n4150 | n29652 ;
  assign n29654 = n10372 ^ n3701 ^ 1'b0 ;
  assign n29655 = n4299 | n29654 ;
  assign n29656 = x181 & ~n16385 ;
  assign n29657 = n29656 ^ n13275 ^ 1'b0 ;
  assign n29658 = n9821 ^ n9267 ^ 1'b0 ;
  assign n29659 = n2030 & ~n5195 ;
  assign n29660 = n29659 ^ n14059 ^ 1'b0 ;
  assign n29661 = n29306 ^ n19967 ^ 1'b0 ;
  assign n29662 = n29660 | n29661 ;
  assign n29663 = n8391 ^ n2153 ^ 1'b0 ;
  assign n29664 = n6659 | n10167 ;
  assign n29665 = x40 & ~n267 ;
  assign n29666 = n4460 | n13437 ;
  assign n29667 = n262 | n6564 ;
  assign n29668 = n12354 | n29667 ;
  assign n29669 = ~n1583 & n27466 ;
  assign n29670 = n29669 ^ n28321 ^ 1'b0 ;
  assign n29671 = n6587 ^ n2104 ^ 1'b0 ;
  assign n29672 = n2383 | n7745 ;
  assign n29673 = n29672 ^ n14237 ^ 1'b0 ;
  assign n29674 = n2282 & ~n20291 ;
  assign n29675 = n29673 & n29674 ;
  assign n29676 = n25440 ^ n14376 ^ n10588 ;
  assign n29677 = n29401 & n29676 ;
  assign n29678 = n29675 & n29677 ;
  assign n29679 = n24353 ^ n7872 ^ 1'b0 ;
  assign n29680 = n14522 & ~n29679 ;
  assign n29681 = ~n15825 & n20284 ;
  assign n29682 = n10085 & n22427 ;
  assign n29683 = n12450 | n19222 ;
  assign n29684 = n4447 | n29683 ;
  assign n29685 = n8087 & n26265 ;
  assign n29686 = n19244 & n29685 ;
  assign n29687 = n22028 ^ n18771 ^ 1'b0 ;
  assign n29688 = n29686 | n29687 ;
  assign n29689 = n29688 ^ n10296 ^ 1'b0 ;
  assign n29690 = n9934 | n29689 ;
  assign n29691 = n5714 & n21720 ;
  assign n29692 = n2360 & n11128 ;
  assign n29693 = n4649 ^ n3420 ^ n2736 ;
  assign n29694 = ~n24454 & n29693 ;
  assign n29695 = n2366 & ~n14486 ;
  assign n29696 = n29695 ^ n10706 ^ 1'b0 ;
  assign n29697 = ~n9788 & n12764 ;
  assign n29698 = n29696 & n29697 ;
  assign n29699 = n294 & ~n10711 ;
  assign n29700 = ~n5455 & n29699 ;
  assign n29701 = n13097 & n28116 ;
  assign n29702 = n29701 ^ n15571 ^ 1'b0 ;
  assign n29703 = ( n4088 & n20604 ) | ( n4088 & ~n25094 ) | ( n20604 & ~n25094 ) ;
  assign n29704 = n7987 & ~n17827 ;
  assign n29705 = n28955 ^ x99 ^ 1'b0 ;
  assign n29706 = ~n14060 & n27347 ;
  assign n29707 = n12297 & n29706 ;
  assign n29708 = n28112 ^ n24889 ^ 1'b0 ;
  assign n29709 = n7670 ^ n2803 ^ 1'b0 ;
  assign n29710 = n18339 | n29709 ;
  assign n29711 = x24 & n24825 ;
  assign n29712 = n9303 ^ n5961 ^ 1'b0 ;
  assign n29713 = ~n6701 & n29712 ;
  assign n29714 = n20696 ^ n701 ^ 1'b0 ;
  assign n29715 = ~n15689 & n29714 ;
  assign n29716 = n29715 ^ n2399 ^ 1'b0 ;
  assign n29717 = n8503 & ~n29716 ;
  assign n29718 = n13661 & ~n14491 ;
  assign n29719 = x21 & n6701 ;
  assign n29720 = n29719 ^ n16628 ^ 1'b0 ;
  assign n29721 = n6648 & ~n9511 ;
  assign n29722 = n19267 & n29721 ;
  assign n29723 = n28564 ^ n7360 ^ 1'b0 ;
  assign n29724 = ( n8814 & n25023 ) | ( n8814 & n29693 ) | ( n25023 & n29693 ) ;
  assign n29725 = n22604 ^ n12708 ^ 1'b0 ;
  assign n29726 = n13686 ^ n6921 ^ 1'b0 ;
  assign n29727 = n24996 & ~n29726 ;
  assign n29728 = ~n28499 & n29727 ;
  assign n29729 = n8882 & n23049 ;
  assign n29730 = n29728 & n29729 ;
  assign n29731 = n5596 ^ n1522 ^ 1'b0 ;
  assign n29732 = ~n1551 & n29731 ;
  assign n29733 = x89 | n17503 ;
  assign n29734 = ~n21473 & n29733 ;
  assign n29735 = n29732 & n29734 ;
  assign n29736 = n29735 ^ n15647 ^ 1'b0 ;
  assign n29737 = n2774 & n23864 ;
  assign n29738 = n29737 ^ n28925 ^ 1'b0 ;
  assign n29739 = n13654 | n16042 ;
  assign n29740 = n29739 ^ n24862 ^ 1'b0 ;
  assign n29741 = n17430 ^ n6069 ^ 1'b0 ;
  assign n29742 = n4293 & ~n5665 ;
  assign n29743 = n23024 ^ n716 ^ 1'b0 ;
  assign n29744 = n15178 ^ n12430 ^ 1'b0 ;
  assign n29745 = n2182 & ~n15213 ;
  assign n29746 = n1603 | n14152 ;
  assign n29747 = n29745 | n29746 ;
  assign n29748 = n29553 ^ n20486 ^ n4503 ;
  assign n29749 = n11566 ^ n1121 ^ 1'b0 ;
  assign n29750 = n7404 & n29749 ;
  assign n29751 = n29750 ^ n9841 ^ 1'b0 ;
  assign n29752 = n7840 & n29751 ;
  assign n29753 = n3400 | n21169 ;
  assign n29754 = n9313 & ~n29753 ;
  assign n29755 = n4097 | n6928 ;
  assign n29756 = ~n16233 & n29755 ;
  assign n29758 = n1474 & ~n1772 ;
  assign n29757 = n9053 ^ n8403 ^ n3272 ;
  assign n29759 = n29758 ^ n29757 ^ 1'b0 ;
  assign n29760 = n29756 & n29759 ;
  assign n29761 = ~n10353 & n29760 ;
  assign n29762 = ( n29752 & ~n29754 ) | ( n29752 & n29761 ) | ( ~n29754 & n29761 ) ;
  assign n29763 = n4185 | n5785 ;
  assign n29764 = n6716 | n14974 ;
  assign n29765 = n11070 | n29764 ;
  assign n29766 = ~n1851 & n4300 ;
  assign n29767 = n29766 ^ x214 ^ 1'b0 ;
  assign n29768 = n537 & n7714 ;
  assign n29769 = ~n16090 & n29768 ;
  assign n29770 = n29767 & n29769 ;
  assign n29771 = n4520 ^ n547 ^ 1'b0 ;
  assign n29772 = ~n29770 & n29771 ;
  assign n29773 = ( n3957 & n8556 ) | ( n3957 & n10059 ) | ( n8556 & n10059 ) ;
  assign n29774 = n12783 & n29773 ;
  assign n29775 = n29774 ^ n26005 ^ 1'b0 ;
  assign n29776 = n29775 ^ n21963 ^ 1'b0 ;
  assign n29777 = n2311 & n24056 ;
  assign n29778 = ( n20023 & n20105 ) | ( n20023 & n26192 ) | ( n20105 & n26192 ) ;
  assign n29779 = ~n10377 & n13905 ;
  assign n29780 = ~n819 & n16674 ;
  assign n29781 = n20585 & n29780 ;
  assign n29782 = n29781 ^ n5130 ^ 1'b0 ;
  assign n29783 = ( n5806 & n12542 ) | ( n5806 & ~n29782 ) | ( n12542 & ~n29782 ) ;
  assign n29784 = ~n2883 & n29783 ;
  assign n29785 = n29784 ^ n1738 ^ 1'b0 ;
  assign n29786 = n6246 ^ n2375 ^ 1'b0 ;
  assign n29787 = n1437 | n29786 ;
  assign n29788 = n11841 ^ n7757 ^ n6659 ;
  assign n29789 = n20832 | n29788 ;
  assign n29790 = n29789 ^ n20291 ^ 1'b0 ;
  assign n29791 = ~n714 & n7685 ;
  assign n29792 = n29791 ^ n8094 ^ 1'b0 ;
  assign n29793 = n1186 & n29792 ;
  assign n29794 = n29793 ^ n12856 ^ n5028 ;
  assign n29795 = n15479 & n27362 ;
  assign n29796 = ~n7923 & n29795 ;
  assign n29797 = n4740 & ~n5535 ;
  assign n29798 = n9009 & n10622 ;
  assign n29799 = n15812 ^ n5535 ^ 1'b0 ;
  assign n29800 = ~n29798 & n29799 ;
  assign n29801 = ~n1891 & n20521 ;
  assign n29802 = n8015 & n29801 ;
  assign n29803 = n3594 & ~n5047 ;
  assign n29804 = n29803 ^ n2506 ^ 1'b0 ;
  assign n29805 = n3864 & ~n20287 ;
  assign n29806 = n29805 ^ n10666 ^ 1'b0 ;
  assign n29807 = ~n7374 & n13031 ;
  assign n29808 = n29807 ^ n11185 ^ 1'b0 ;
  assign n29809 = n4733 & n7240 ;
  assign n29810 = n14490 ^ x148 ^ 1'b0 ;
  assign n29811 = n9801 & ~n29810 ;
  assign n29812 = n29811 ^ n3500 ^ n2998 ;
  assign n29813 = ( ~n9051 & n12595 ) | ( ~n9051 & n17303 ) | ( n12595 & n17303 ) ;
  assign n29814 = n15617 ^ n3450 ^ 1'b0 ;
  assign n29815 = ~n13424 & n18028 ;
  assign n29816 = n6255 & ~n25219 ;
  assign n29817 = n10437 & n19465 ;
  assign n29818 = n10722 | n25981 ;
  assign n29819 = n29817 & ~n29818 ;
  assign n29820 = n7379 | n17226 ;
  assign n29821 = n29820 ^ n24869 ^ 1'b0 ;
  assign n29825 = n7143 ^ n3529 ^ 1'b0 ;
  assign n29826 = n9574 | n29825 ;
  assign n29822 = ~n752 & n9157 ;
  assign n29823 = ~x159 & n29822 ;
  assign n29824 = n11653 & ~n29823 ;
  assign n29827 = n29826 ^ n29824 ^ 1'b0 ;
  assign n29828 = n16810 ^ n9951 ^ 1'b0 ;
  assign n29829 = n14191 | n29828 ;
  assign n29830 = n29829 ^ n17239 ^ 1'b0 ;
  assign n29831 = ~n1721 & n17490 ;
  assign n29832 = n3819 | n8602 ;
  assign n29833 = n1051 & ~n29832 ;
  assign n29834 = n8353 ^ n4256 ^ 1'b0 ;
  assign n29835 = n29834 ^ n28325 ^ 1'b0 ;
  assign n29836 = n3342 & n6202 ;
  assign n29837 = n2891 & n29836 ;
  assign n29838 = ~x80 & n7395 ;
  assign n29839 = ~n5958 & n29838 ;
  assign n29840 = ~n29837 & n29839 ;
  assign n29841 = n20594 & n29840 ;
  assign n29842 = n20616 | n27069 ;
  assign n29843 = ~n9735 & n15337 ;
  assign n29844 = ~n5139 & n15276 ;
  assign n29845 = ~n18728 & n29844 ;
  assign n29846 = n29845 ^ n16660 ^ n10754 ;
  assign n29847 = n8522 & ~n29846 ;
  assign n29848 = n23579 ^ n5320 ^ n4616 ;
  assign n29849 = ~n3850 & n10534 ;
  assign n29850 = n29849 ^ n16796 ^ 1'b0 ;
  assign n29851 = n29850 ^ n25055 ^ n15674 ;
  assign n29852 = n29851 ^ n24869 ^ 1'b0 ;
  assign n29853 = n3494 | n11719 ;
  assign n29854 = n13239 & n19325 ;
  assign n29855 = n29853 & n29854 ;
  assign n29856 = n845 | n14341 ;
  assign n29857 = n6977 & ~n29856 ;
  assign n29858 = n23003 & n29857 ;
  assign n29859 = n25454 ^ n14527 ^ 1'b0 ;
  assign n29860 = n29858 | n29859 ;
  assign n29861 = n15160 ^ n4198 ^ 1'b0 ;
  assign n29862 = n15427 | n19871 ;
  assign n29863 = n5273 & ~n15204 ;
  assign n29864 = n4637 ^ n1021 ^ 1'b0 ;
  assign n29865 = n18026 & ~n29864 ;
  assign n29866 = n29865 ^ n13316 ^ 1'b0 ;
  assign n29867 = n7676 ^ n1422 ^ 1'b0 ;
  assign n29868 = n3145 & n29867 ;
  assign n29869 = n19504 ^ n1880 ^ 1'b0 ;
  assign n29870 = n29837 | n29869 ;
  assign n29871 = n10817 ^ n2392 ^ 1'b0 ;
  assign n29872 = n4906 & ~n29871 ;
  assign n29873 = n23802 ^ n9076 ^ n1255 ;
  assign n29874 = n3189 & ~n6872 ;
  assign n29875 = n29874 ^ n10353 ^ 1'b0 ;
  assign n29876 = n688 & n29061 ;
  assign n29877 = n19364 ^ n17378 ^ 1'b0 ;
  assign n29879 = n3736 | n3830 ;
  assign n29880 = n3830 & ~n29879 ;
  assign n29881 = n29880 ^ n3670 ^ 1'b0 ;
  assign n29882 = n4931 & ~n29881 ;
  assign n29878 = n988 & n1462 ;
  assign n29883 = n29882 ^ n29878 ^ n16576 ;
  assign n29884 = n1807 & ~n9431 ;
  assign n29885 = n29884 ^ n22800 ^ n8180 ;
  assign n29886 = x82 | n8786 ;
  assign n29887 = n7990 ^ n7683 ^ 1'b0 ;
  assign n29888 = n29886 & ~n29887 ;
  assign n29889 = n2875 & n15387 ;
  assign n29890 = n4685 | n6155 ;
  assign n29891 = ~n10849 & n14507 ;
  assign n29892 = n4237 & ~n29891 ;
  assign n29893 = ~n15998 & n29892 ;
  assign n29894 = n5479 ^ n3328 ^ 1'b0 ;
  assign n29895 = x145 & n10194 ;
  assign n29896 = ~n14138 & n20759 ;
  assign n29897 = ~n29895 & n29896 ;
  assign n29898 = n4922 & ~n10236 ;
  assign n29899 = n19084 & n29898 ;
  assign n29900 = n1175 & ~n29899 ;
  assign n29903 = n5010 ^ n2301 ^ 1'b0 ;
  assign n29901 = n3210 | n4388 ;
  assign n29902 = n14315 & ~n29901 ;
  assign n29904 = n29903 ^ n29902 ^ n7061 ;
  assign n29905 = ( n12469 & n14768 ) | ( n12469 & n29904 ) | ( n14768 & n29904 ) ;
  assign n29906 = n18922 ^ n8781 ^ 1'b0 ;
  assign n29907 = n8336 & ~n25152 ;
  assign n29908 = n29906 & n29907 ;
  assign n29909 = n3262 & n17589 ;
  assign n29910 = n1665 | n20138 ;
  assign n29911 = n29910 ^ n19733 ^ 1'b0 ;
  assign n29912 = n15652 & n29911 ;
  assign n29913 = n2286 & ~n29912 ;
  assign n29914 = n12246 & n26667 ;
  assign n29915 = n5509 & ~n10974 ;
  assign n29916 = n1910 & n29915 ;
  assign n29917 = ~n11705 & n29916 ;
  assign n29918 = n29917 ^ n13981 ^ n9806 ;
  assign n29919 = ~n3335 & n19561 ;
  assign n29920 = n25296 ^ n9710 ^ n8254 ;
  assign n29921 = ( n29918 & n29919 ) | ( n29918 & n29920 ) | ( n29919 & n29920 ) ;
  assign n29922 = ( ~n7220 & n8052 ) | ( ~n7220 & n17114 ) | ( n8052 & n17114 ) ;
  assign n29923 = n29922 ^ n9676 ^ n5690 ;
  assign n29924 = n10714 | n28936 ;
  assign n29925 = n29924 ^ n8465 ^ 1'b0 ;
  assign n29926 = n2383 & ~n27185 ;
  assign n29927 = n29926 ^ n11941 ^ 1'b0 ;
  assign n29928 = n9674 | n19955 ;
  assign n29929 = n29928 ^ n15351 ^ 1'b0 ;
  assign n29932 = ~n3344 & n11030 ;
  assign n29930 = n9722 ^ n7285 ^ n3030 ;
  assign n29931 = ~n15874 & n29930 ;
  assign n29933 = n29932 ^ n29931 ^ 1'b0 ;
  assign n29934 = n3494 | n6506 ;
  assign n29935 = n29934 ^ x241 ^ 1'b0 ;
  assign n29936 = n17811 & n29935 ;
  assign n29937 = n21523 ^ n2638 ^ 1'b0 ;
  assign n29938 = n7070 | n8587 ;
  assign n29939 = n19460 & ~n29938 ;
  assign n29940 = n2568 & ~n29939 ;
  assign n29941 = n29940 ^ n19575 ^ 1'b0 ;
  assign n29942 = ~n4815 & n26418 ;
  assign n29943 = n29942 ^ n12854 ^ 1'b0 ;
  assign n29944 = n14708 ^ n4993 ^ 1'b0 ;
  assign n29945 = n2191 & ~n29944 ;
  assign n29946 = n28125 ^ n11680 ^ 1'b0 ;
  assign n29947 = n29945 & ~n29946 ;
  assign n29948 = ~n5383 & n6433 ;
  assign n29949 = n29948 ^ n353 ^ 1'b0 ;
  assign n29950 = n14364 & ~n29949 ;
  assign n29951 = n11850 | n13503 ;
  assign n29952 = n29951 ^ n19318 ^ 1'b0 ;
  assign n29953 = n20089 & n21655 ;
  assign n29954 = n26418 ^ n15304 ^ 1'b0 ;
  assign n29955 = ~n3772 & n29954 ;
  assign n29959 = n12894 & n15812 ;
  assign n29956 = ~n3899 & n4828 ;
  assign n29957 = n3266 | n29956 ;
  assign n29958 = n29957 ^ x6 ^ 1'b0 ;
  assign n29960 = n29959 ^ n29958 ^ 1'b0 ;
  assign n29961 = n2307 & ~n5604 ;
  assign n29962 = ~n13757 & n29961 ;
  assign n29963 = n3590 | n11626 ;
  assign n29964 = n29963 ^ n6496 ^ 1'b0 ;
  assign n29965 = n27637 & n29964 ;
  assign n29968 = ~n1981 & n12452 ;
  assign n29969 = n25604 & n29968 ;
  assign n29966 = n8927 | n14897 ;
  assign n29967 = n2868 & ~n29966 ;
  assign n29970 = n29969 ^ n29967 ^ 1'b0 ;
  assign n29971 = n13193 ^ n6387 ^ 1'b0 ;
  assign n29972 = n3947 & n29971 ;
  assign n29973 = n29972 ^ n8738 ^ 1'b0 ;
  assign n29974 = n8899 | n29973 ;
  assign n29975 = n29974 ^ n7385 ^ 1'b0 ;
  assign n29976 = n18741 & n29975 ;
  assign n29977 = n29976 ^ n18859 ^ 1'b0 ;
  assign n29978 = n20818 & n29977 ;
  assign n29979 = n906 & ~n13080 ;
  assign n29980 = n29785 & n29979 ;
  assign n29981 = ~n14059 & n29980 ;
  assign n29982 = n18133 ^ n17824 ^ 1'b0 ;
  assign n29983 = n12610 | n27828 ;
  assign n29984 = n22973 | n29983 ;
  assign n29985 = n4852 & n28635 ;
  assign n29986 = n29985 ^ n3873 ^ 1'b0 ;
  assign n29987 = n18822 & n20435 ;
  assign n29988 = ~n13976 & n29987 ;
  assign n29989 = n12892 & ~n17592 ;
  assign n29990 = n29989 ^ n372 ^ 1'b0 ;
  assign n29991 = n4669 & n29990 ;
  assign n29992 = n29988 & n29991 ;
  assign n29993 = n14526 ^ n13317 ^ 1'b0 ;
  assign n29994 = n17818 & ~n29993 ;
  assign n29995 = n5975 ^ n4511 ^ 1'b0 ;
  assign n29996 = ~n1891 & n29995 ;
  assign n29997 = ( ~n10442 & n23475 ) | ( ~n10442 & n29996 ) | ( n23475 & n29996 ) ;
  assign n29998 = n3601 & n22586 ;
  assign n29999 = n29998 ^ n2004 ^ 1'b0 ;
  assign n30000 = n15161 & ~n19529 ;
  assign n30001 = n19080 | n21168 ;
  assign n30002 = n4260 & n7513 ;
  assign n30003 = ~n6686 & n30002 ;
  assign n30004 = n8820 | n30003 ;
  assign n30005 = n30001 | n30004 ;
  assign n30006 = n26347 ^ n7761 ^ 1'b0 ;
  assign n30007 = n24132 ^ n10012 ^ 1'b0 ;
  assign n30008 = ~n4619 & n7558 ;
  assign n30009 = n30008 ^ n2223 ^ 1'b0 ;
  assign n30010 = n4632 | n30009 ;
  assign n30011 = n23854 & n30010 ;
  assign n30012 = ~n9543 & n11775 ;
  assign n30013 = n30012 ^ n3349 ^ 1'b0 ;
  assign n30015 = n8071 & n11285 ;
  assign n30014 = n13650 | n25745 ;
  assign n30016 = n30015 ^ n30014 ^ 1'b0 ;
  assign n30017 = n8522 & ~n16695 ;
  assign n30018 = ~n15053 & n30017 ;
  assign n30019 = ( ~n4381 & n12896 ) | ( ~n4381 & n30018 ) | ( n12896 & n30018 ) ;
  assign n30020 = n3593 & ~n8401 ;
  assign n30021 = n13176 ^ n12807 ^ 1'b0 ;
  assign n30022 = n1196 | n30021 ;
  assign n30023 = n4834 ^ n2641 ^ 1'b0 ;
  assign n30024 = ~n22493 & n22787 ;
  assign n30025 = n5330 & n6713 ;
  assign n30026 = n21129 | n30025 ;
  assign n30028 = n3055 | n14944 ;
  assign n30029 = n6036 | n30028 ;
  assign n30027 = n9205 & n9934 ;
  assign n30030 = n30029 ^ n30027 ^ 1'b0 ;
  assign n30031 = ~n8129 & n9192 ;
  assign n30032 = n28942 & n30031 ;
  assign n30033 = n13888 & ~n17974 ;
  assign n30034 = ~x249 & n30033 ;
  assign n30035 = n14285 & n23065 ;
  assign n30036 = n30035 ^ n11895 ^ 1'b0 ;
  assign n30037 = n19755 ^ n14497 ^ 1'b0 ;
  assign n30038 = n24852 ^ n16147 ^ x100 ;
  assign n30039 = n2715 | n4078 ;
  assign n30040 = n21034 & n30039 ;
  assign n30041 = ~n23369 & n30040 ;
  assign n30042 = n17707 ^ n1672 ^ 1'b0 ;
  assign n30043 = n30042 ^ n3899 ^ 1'b0 ;
  assign n30044 = n10950 & ~n30043 ;
  assign n30045 = n14291 | n30044 ;
  assign n30046 = n1101 | n10570 ;
  assign n30047 = n2493 & ~n7903 ;
  assign n30048 = n20896 ^ n4509 ^ n453 ;
  assign n30049 = n30048 ^ n417 ^ 1'b0 ;
  assign n30050 = ~n4574 & n30049 ;
  assign n30051 = n7243 ^ n708 ^ 1'b0 ;
  assign n30052 = n23133 & ~n30051 ;
  assign n30053 = n30052 ^ n4571 ^ 1'b0 ;
  assign n30054 = n23065 & ~n30053 ;
  assign n30056 = ( n453 & n812 ) | ( n453 & ~n7066 ) | ( n812 & ~n7066 ) ;
  assign n30055 = ~n12802 & n23751 ;
  assign n30057 = n30056 ^ n30055 ^ n24931 ;
  assign n30058 = ( n7170 & n17252 ) | ( n7170 & ~n30057 ) | ( n17252 & ~n30057 ) ;
  assign n30059 = n3383 & n4025 ;
  assign n30060 = n6567 | n30059 ;
  assign n30061 = n30060 ^ n5402 ^ 1'b0 ;
  assign n30062 = n30061 ^ n3549 ^ 1'b0 ;
  assign n30063 = n27757 ^ n4608 ^ 1'b0 ;
  assign n30064 = n293 & n4145 ;
  assign n30065 = n30064 ^ n8616 ^ 1'b0 ;
  assign n30066 = n10071 | n30065 ;
  assign n30067 = n11653 & n26450 ;
  assign n30071 = n4013 & ~n8457 ;
  assign n30072 = ~n4013 & n30071 ;
  assign n30073 = n30072 ^ n7301 ^ 1'b0 ;
  assign n30068 = n3760 & ~n13530 ;
  assign n30069 = n13530 & n30068 ;
  assign n30070 = n30069 ^ n21320 ^ 1'b0 ;
  assign n30074 = n30073 ^ n30070 ^ 1'b0 ;
  assign n30075 = ~n13047 & n30074 ;
  assign n30076 = n30075 ^ n21965 ^ 1'b0 ;
  assign n30077 = n20933 & ~n30076 ;
  assign n30078 = n14699 ^ n5452 ^ 1'b0 ;
  assign n30079 = n30078 ^ n17263 ^ 1'b0 ;
  assign n30080 = n5853 & n7329 ;
  assign n30081 = ~x175 & n11297 ;
  assign n30082 = ( n8058 & n30080 ) | ( n8058 & n30081 ) | ( n30080 & n30081 ) ;
  assign n30083 = n8344 ^ n1389 ^ 1'b0 ;
  assign n30084 = ~n6006 & n16109 ;
  assign n30085 = n22467 ^ n19837 ^ 1'b0 ;
  assign n30086 = n30084 & ~n30085 ;
  assign n30087 = n5410 & n29277 ;
  assign n30088 = n30087 ^ x227 ^ 1'b0 ;
  assign n30089 = n11756 ^ n3240 ^ 1'b0 ;
  assign n30090 = n22467 & n30089 ;
  assign n30091 = n1180 & ~n15366 ;
  assign n30092 = n30091 ^ n25107 ^ 1'b0 ;
  assign n30093 = n10575 | n29693 ;
  assign n30094 = n5453 | n30093 ;
  assign n30095 = n30094 ^ n27104 ^ 1'b0 ;
  assign n30096 = n25084 ^ n15299 ^ 1'b0 ;
  assign n30097 = n22228 ^ n12574 ^ 1'b0 ;
  assign n30099 = n18420 ^ n11297 ^ 1'b0 ;
  assign n30098 = n1690 | n25091 ;
  assign n30100 = n30099 ^ n30098 ^ 1'b0 ;
  assign n30102 = n3400 ^ n3246 ^ 1'b0 ;
  assign n30103 = n5525 | n30102 ;
  assign n30101 = x61 & ~n5005 ;
  assign n30104 = n30103 ^ n30101 ^ 1'b0 ;
  assign n30105 = n30104 ^ n8344 ^ 1'b0 ;
  assign n30106 = n18256 & ~n18415 ;
  assign n30107 = n4603 ^ n997 ^ 1'b0 ;
  assign n30108 = n12911 & ~n30107 ;
  assign n30109 = n18476 & ~n30108 ;
  assign n30110 = n1989 ^ n966 ^ 1'b0 ;
  assign n30111 = n12650 & ~n14538 ;
  assign n30112 = n2750 & ~n30111 ;
  assign n30113 = n14861 & n30112 ;
  assign n30114 = n10182 & ~n19469 ;
  assign n30115 = ~n256 & n7914 ;
  assign n30116 = n19682 & n30115 ;
  assign n30117 = ( n872 & n27739 ) | ( n872 & ~n30116 ) | ( n27739 & ~n30116 ) ;
  assign n30118 = n27003 ^ n15432 ^ 1'b0 ;
  assign n30119 = ~n9777 & n30118 ;
  assign n30120 = n5511 | n21347 ;
  assign n30121 = n30120 ^ n5579 ^ 1'b0 ;
  assign n30122 = n7914 & ~n30121 ;
  assign n30123 = n27470 | n30122 ;
  assign n30124 = n30123 ^ n6771 ^ 1'b0 ;
  assign n30125 = n23640 & ~n30124 ;
  assign n30126 = n917 & n15076 ;
  assign n30127 = n30126 ^ n2286 ^ 1'b0 ;
  assign n30128 = n23632 ^ n16882 ^ n15774 ;
  assign n30129 = n9777 ^ n8772 ^ 1'b0 ;
  assign n30130 = n3309 & n4603 ;
  assign n30131 = ~n4433 & n11204 ;
  assign n30132 = n25348 & n30131 ;
  assign n30133 = n27603 ^ n20108 ^ n7476 ;
  assign n30134 = ~n17678 & n30133 ;
  assign n30135 = ~n624 & n1738 ;
  assign n30136 = n30135 ^ n8112 ^ 1'b0 ;
  assign n30137 = n14967 | n30136 ;
  assign n30138 = n30137 ^ n9440 ^ 1'b0 ;
  assign n30139 = n29031 ^ n19554 ^ 1'b0 ;
  assign n30140 = n30139 ^ n24849 ^ 1'b0 ;
  assign n30141 = n5095 | n9627 ;
  assign n30142 = n5459 | n30141 ;
  assign n30143 = n16758 & ~n20776 ;
  assign n30144 = n8175 & n30143 ;
  assign n30145 = n30144 ^ n11860 ^ 1'b0 ;
  assign n30146 = n5135 & n7903 ;
  assign n30147 = n1774 & n24208 ;
  assign n30148 = ( n3809 & ~n30146 ) | ( n3809 & n30147 ) | ( ~n30146 & n30147 ) ;
  assign n30149 = n15894 ^ n11875 ^ 1'b0 ;
  assign n30150 = ~n4056 & n12486 ;
  assign n30151 = n8603 & ~n12574 ;
  assign n30152 = n30151 ^ n14312 ^ 1'b0 ;
  assign n30153 = n4381 | n30152 ;
  assign n30154 = ~n4258 & n6864 ;
  assign n30155 = n30154 ^ n1517 ^ 1'b0 ;
  assign n30156 = n6579 & n20696 ;
  assign n30157 = n2988 & n30156 ;
  assign n30158 = n30157 ^ n18725 ^ n12670 ;
  assign n30159 = n22824 ^ n11917 ^ n1891 ;
  assign n30160 = n10852 | n30159 ;
  assign n30161 = n30122 ^ n4069 ^ 1'b0 ;
  assign n30162 = n4260 & n24462 ;
  assign n30163 = n22303 & n30162 ;
  assign n30164 = n10649 | n16228 ;
  assign n30165 = n30164 ^ n18873 ^ 1'b0 ;
  assign n30166 = n7811 | n21757 ;
  assign n30167 = n30166 ^ n8112 ^ 1'b0 ;
  assign n30168 = n3515 | n30167 ;
  assign n30169 = n25633 & ~n26658 ;
  assign n30170 = n9844 | n24920 ;
  assign n30171 = n2809 & ~n30170 ;
  assign n30172 = n1628 & ~n30171 ;
  assign n30173 = n13466 ^ n2164 ^ 1'b0 ;
  assign n30174 = n16257 & ~n30173 ;
  assign n30175 = ~n21347 & n29118 ;
  assign n30176 = ~n30174 & n30175 ;
  assign n30177 = n26488 ^ n779 ^ 1'b0 ;
  assign n30178 = n18549 & ~n30177 ;
  assign n30179 = n12559 ^ n8289 ^ 1'b0 ;
  assign n30180 = n30178 & n30179 ;
  assign n30181 = n9912 ^ n2268 ^ 1'b0 ;
  assign n30182 = n23056 ^ n19132 ^ 1'b0 ;
  assign n30183 = ~n8463 & n9532 ;
  assign n30184 = n6075 & n30183 ;
  assign n30185 = n30184 ^ n3657 ^ 1'b0 ;
  assign n30186 = n5051 & ~n15485 ;
  assign n30187 = n17628 | n25977 ;
  assign n30188 = n15028 | n15395 ;
  assign n30189 = n30187 | n30188 ;
  assign n30190 = ( ~n2120 & n10331 ) | ( ~n2120 & n25088 ) | ( n10331 & n25088 ) ;
  assign n30191 = n30190 ^ n10175 ^ 1'b0 ;
  assign n30192 = n30191 ^ n14939 ^ 1'b0 ;
  assign n30193 = ~n11961 & n30192 ;
  assign n30194 = n30193 ^ n3037 ^ 1'b0 ;
  assign n30195 = n2873 | n3815 ;
  assign n30196 = n1042 & n27882 ;
  assign n30197 = n24246 ^ n7484 ^ 1'b0 ;
  assign n30198 = n5607 & ~n10527 ;
  assign n30199 = ~n2747 & n24807 ;
  assign n30200 = n2848 ^ n1351 ^ 1'b0 ;
  assign n30201 = n19690 ^ n18525 ^ 1'b0 ;
  assign n30202 = n19617 | n30201 ;
  assign n30203 = ( n21650 & n30200 ) | ( n21650 & ~n30202 ) | ( n30200 & ~n30202 ) ;
  assign n30204 = n30203 ^ n23586 ^ 1'b0 ;
  assign n30205 = n858 & n12937 ;
  assign n30206 = n28120 ^ n5118 ^ 1'b0 ;
  assign n30207 = n2450 & n30206 ;
  assign n30208 = n30207 ^ n14202 ^ 1'b0 ;
  assign n30209 = n30205 & n30208 ;
  assign n30210 = n7223 & ~n23800 ;
  assign n30211 = n6075 & n28910 ;
  assign n30212 = n10174 & n28833 ;
  assign n30213 = ~n4608 & n30212 ;
  assign n30214 = n21507 & n24137 ;
  assign n30215 = ~n10903 & n30214 ;
  assign n30216 = n2868 & n4306 ;
  assign n30217 = ~n14499 & n30216 ;
  assign n30218 = n30001 & ~n30217 ;
  assign n30219 = n20744 ^ n15104 ^ n12631 ;
  assign n30220 = ( ~n15277 & n24816 ) | ( ~n15277 & n30219 ) | ( n24816 & n30219 ) ;
  assign n30221 = n18754 ^ n6036 ^ 1'b0 ;
  assign n30222 = n13765 & ~n30221 ;
  assign n30223 = n11605 & n30222 ;
  assign n30224 = ~n8147 & n30223 ;
  assign n30225 = n3685 ^ n1763 ^ 1'b0 ;
  assign n30226 = n4610 & ~n30225 ;
  assign n30227 = n6339 & n19241 ;
  assign n30228 = n2870 & n30227 ;
  assign n30229 = x132 & ~n4484 ;
  assign n30230 = n30228 & n30229 ;
  assign n30231 = n30226 & ~n30230 ;
  assign n30232 = n30231 ^ n22931 ^ 1'b0 ;
  assign n30233 = n2167 & n5180 ;
  assign n30234 = n30233 ^ x54 ^ 1'b0 ;
  assign n30235 = n30234 ^ n15787 ^ n7157 ;
  assign n30236 = n1254 & n20644 ;
  assign n30237 = n1492 | n30236 ;
  assign n30238 = n25400 ^ n7405 ^ 1'b0 ;
  assign n30239 = n2206 & ~n30238 ;
  assign n30240 = n22266 ^ n16416 ^ 1'b0 ;
  assign n30241 = n16920 | n20526 ;
  assign n30242 = ( n2544 & n2701 ) | ( n2544 & ~n15834 ) | ( n2701 & ~n15834 ) ;
  assign n30243 = n7789 ^ n5541 ^ 1'b0 ;
  assign n30244 = n1894 & n16723 ;
  assign n30245 = ~n30243 & n30244 ;
  assign n30246 = n28874 | n30245 ;
  assign n30247 = n25866 ^ n7273 ^ 1'b0 ;
  assign n30248 = ~n24646 & n30247 ;
  assign n30249 = n29785 & ~n30248 ;
  assign n30250 = n30249 ^ n1561 ^ 1'b0 ;
  assign n30251 = ~n1276 & n4410 ;
  assign n30252 = n30251 ^ n4894 ^ 1'b0 ;
  assign n30253 = n1832 & n30252 ;
  assign n30254 = n699 | n3483 ;
  assign n30255 = ~n5649 & n14117 ;
  assign n30256 = ( n2063 & n3207 ) | ( n2063 & ~n30255 ) | ( n3207 & ~n30255 ) ;
  assign n30257 = x155 & ~n30256 ;
  assign n30258 = n30257 ^ n13339 ^ 1'b0 ;
  assign n30259 = n27832 ^ n15765 ^ 1'b0 ;
  assign n30260 = x178 & n30259 ;
  assign n30261 = n12573 & ~n16291 ;
  assign n30262 = n15429 & ~n18340 ;
  assign n30263 = n30261 & n30262 ;
  assign n30265 = n16505 ^ n2674 ^ 1'b0 ;
  assign n30266 = n22523 & n30265 ;
  assign n30267 = n8276 & n30266 ;
  assign n30264 = n4878 | n9850 ;
  assign n30268 = n30267 ^ n30264 ^ 1'b0 ;
  assign n30269 = ~n2920 & n24851 ;
  assign n30270 = ~n30268 & n30269 ;
  assign n30271 = n466 | n22079 ;
  assign n30272 = n30271 ^ n2319 ^ 1'b0 ;
  assign n30273 = n9177 & ~n30272 ;
  assign n30274 = n8373 & n16947 ;
  assign n30275 = n30274 ^ n5354 ^ 1'b0 ;
  assign n30276 = n13424 & ~n30275 ;
  assign n30277 = n2526 & n22636 ;
  assign n30278 = n11909 & ~n29997 ;
  assign n30279 = ~n12767 & n30278 ;
  assign n30280 = n21462 ^ n13303 ^ 1'b0 ;
  assign n30281 = ( ~n14755 & n23683 ) | ( ~n14755 & n24937 ) | ( n23683 & n24937 ) ;
  assign n30282 = n9611 | n27921 ;
  assign n30283 = n30282 ^ n29861 ^ 1'b0 ;
  assign n30284 = n2192 | n12058 ;
  assign n30285 = n11840 | n30284 ;
  assign n30286 = n16167 & n30285 ;
  assign n30287 = n30286 ^ n29154 ^ 1'b0 ;
  assign n30288 = n11856 & n30287 ;
  assign n30289 = n26349 & n28092 ;
  assign n30290 = n13742 ^ n10487 ^ n8195 ;
  assign n30291 = n29221 ^ n11253 ^ n5088 ;
  assign n30292 = ~n20989 & n28055 ;
  assign n30293 = n15811 ^ n8912 ^ 1'b0 ;
  assign n30294 = n2785 & ~n30293 ;
  assign n30295 = n18742 ^ n4265 ^ 1'b0 ;
  assign n30296 = n15070 & n30295 ;
  assign n30297 = ( ~n1508 & n18026 ) | ( ~n1508 & n28017 ) | ( n18026 & n28017 ) ;
  assign n30298 = n30296 & ~n30297 ;
  assign n30301 = n25731 ^ n13911 ^ 1'b0 ;
  assign n30299 = ~n6273 & n7805 ;
  assign n30300 = n30299 ^ n9701 ^ 1'b0 ;
  assign n30302 = n30301 ^ n30300 ^ 1'b0 ;
  assign n30303 = n20336 & n30302 ;
  assign n30304 = n18141 ^ n3119 ^ 1'b0 ;
  assign n30305 = n30303 & n30304 ;
  assign n30306 = n826 & n2283 ;
  assign n30307 = n9252 & n30306 ;
  assign n30308 = n18313 | n30307 ;
  assign n30309 = n30308 ^ n8964 ^ 1'b0 ;
  assign n30310 = n11014 ^ n5749 ^ 1'b0 ;
  assign n30311 = n8837 ^ n7303 ^ 1'b0 ;
  assign n30313 = n16104 ^ n4310 ^ n2866 ;
  assign n30312 = ~n15498 & n16877 ;
  assign n30314 = n30313 ^ n30312 ^ 1'b0 ;
  assign n30322 = ~n1667 & n7737 ;
  assign n30323 = n1667 & n30322 ;
  assign n30324 = ~n7276 & n30323 ;
  assign n30325 = ~n3186 & n30324 ;
  assign n30326 = n3186 & n30325 ;
  assign n30315 = n4881 | n8864 ;
  assign n30316 = n4113 & ~n7786 ;
  assign n30317 = n7786 & n30316 ;
  assign n30318 = n3829 & ~n30317 ;
  assign n30319 = ~n3829 & n30318 ;
  assign n30320 = n28263 & ~n30319 ;
  assign n30321 = ~n30315 & n30320 ;
  assign n30327 = n30326 ^ n30321 ^ 1'b0 ;
  assign n30328 = n19970 ^ n12679 ^ n8609 ;
  assign n30330 = ( x120 & n5605 ) | ( x120 & n10364 ) | ( n5605 & n10364 ) ;
  assign n30329 = n10925 & n20416 ;
  assign n30331 = n30330 ^ n30329 ^ 1'b0 ;
  assign n30332 = ~n30328 & n30331 ;
  assign n30333 = n30332 ^ n9853 ^ 1'b0 ;
  assign n30334 = n13181 ^ n1665 ^ 1'b0 ;
  assign n30335 = x89 | n5851 ;
  assign n30336 = n9889 & ~n30335 ;
  assign n30337 = n29544 & ~n30336 ;
  assign n30338 = n3709 | n4988 ;
  assign n30339 = ~n4268 & n10894 ;
  assign n30340 = ~n25029 & n30339 ;
  assign n30341 = ~n2907 & n30340 ;
  assign n30342 = n13459 ^ n4557 ^ 1'b0 ;
  assign n30346 = n15073 & n23757 ;
  assign n30347 = n30346 ^ n15155 ^ 1'b0 ;
  assign n30348 = n4929 & ~n30347 ;
  assign n30349 = n30348 ^ n6668 ^ 1'b0 ;
  assign n30350 = n9628 & ~n30349 ;
  assign n30343 = n13894 ^ n9443 ^ 1'b0 ;
  assign n30344 = n2521 | n30343 ;
  assign n30345 = n3671 | n30344 ;
  assign n30351 = n30350 ^ n30345 ^ 1'b0 ;
  assign n30352 = ( x86 & n17546 ) | ( x86 & ~n28058 ) | ( n17546 & ~n28058 ) ;
  assign n30353 = n7332 ^ n890 ^ n516 ;
  assign n30354 = n30353 ^ n14534 ^ 1'b0 ;
  assign n30355 = n3944 & n30354 ;
  assign n30356 = n25566 ^ n24627 ^ 1'b0 ;
  assign n30357 = n30355 & ~n30356 ;
  assign n30358 = n30357 ^ n9800 ^ 1'b0 ;
  assign n30359 = n5218 & ~n7778 ;
  assign n30360 = n30359 ^ n11035 ^ 1'b0 ;
  assign n30361 = ~n733 & n24967 ;
  assign n30362 = n11183 & n30361 ;
  assign n30363 = n30362 ^ n20864 ^ 1'b0 ;
  assign n30364 = n8397 & n30363 ;
  assign n30365 = n10957 | n30364 ;
  assign n30366 = n30360 | n30365 ;
  assign n30367 = n10711 ^ n4132 ^ 1'b0 ;
  assign n30368 = n28286 | n30367 ;
  assign n30369 = n30368 ^ n16885 ^ 1'b0 ;
  assign n30370 = n25600 ^ n22548 ^ 1'b0 ;
  assign n30371 = n11834 & ~n30370 ;
  assign n30372 = n10666 ^ n8984 ^ 1'b0 ;
  assign n30373 = n30372 ^ n10354 ^ 1'b0 ;
  assign n30374 = n30371 | n30373 ;
  assign n30375 = n25467 ^ n6045 ^ n4255 ;
  assign n30376 = n29861 ^ n2354 ^ 1'b0 ;
  assign n30377 = n30375 & n30376 ;
  assign n30378 = n4317 & ~n23342 ;
  assign n30379 = n30378 ^ n6313 ^ 1'b0 ;
  assign n30380 = n3256 | n30379 ;
  assign n30381 = n12170 | n30380 ;
  assign n30382 = n20519 ^ x116 ^ 1'b0 ;
  assign n30383 = n30382 ^ n25332 ^ n15327 ;
  assign n30384 = n11672 & ~n15783 ;
  assign n30385 = n30384 ^ n23866 ^ 1'b0 ;
  assign n30386 = ( ~n9628 & n21014 ) | ( ~n9628 & n30385 ) | ( n21014 & n30385 ) ;
  assign n30387 = n8182 & n25255 ;
  assign n30388 = ~n22440 & n30387 ;
  assign n30389 = n3243 | n16042 ;
  assign n30390 = n17355 & ~n30389 ;
  assign n30391 = ~n6965 & n13521 ;
  assign n30392 = ~n3707 & n30391 ;
  assign n30393 = n1322 & ~n7347 ;
  assign n30394 = n8133 ^ n7266 ^ 1'b0 ;
  assign n30395 = ~n15122 & n29403 ;
  assign n30396 = n2192 & n6337 ;
  assign n30397 = n30396 ^ n4524 ^ 1'b0 ;
  assign n30398 = n13697 | n18240 ;
  assign n30399 = n30397 | n30398 ;
  assign n30400 = n24731 ^ n16330 ^ n14630 ;
  assign n30401 = n30399 | n30400 ;
  assign n30403 = ~n2613 & n16255 ;
  assign n30402 = n1278 & ~n13240 ;
  assign n30404 = n30403 ^ n30402 ^ 1'b0 ;
  assign n30405 = n6661 & n30404 ;
  assign n30406 = n30405 ^ n4911 ^ 1'b0 ;
  assign n30407 = n26207 ^ n14458 ^ 1'b0 ;
  assign n30408 = n25737 | n30407 ;
  assign n30410 = n12720 | n12837 ;
  assign n30409 = n4922 & n5333 ;
  assign n30411 = n30410 ^ n30409 ^ 1'b0 ;
  assign n30412 = ~n18922 & n30411 ;
  assign n30413 = n5293 ^ n4428 ^ 1'b0 ;
  assign n30414 = ~n697 & n30413 ;
  assign n30415 = n30414 ^ n8868 ^ 1'b0 ;
  assign n30416 = n30412 & n30415 ;
  assign n30417 = n15135 | n24071 ;
  assign n30418 = n2972 & ~n23285 ;
  assign n30419 = n30418 ^ n12848 ^ n11523 ;
  assign n30420 = n4710 & ~n11377 ;
  assign n30421 = n29396 & n30420 ;
  assign n30422 = n30421 ^ n5799 ^ 1'b0 ;
  assign n30424 = n8354 & n10984 ;
  assign n30423 = n2801 | n11628 ;
  assign n30425 = n30424 ^ n30423 ^ 1'b0 ;
  assign n30426 = n21285 ^ n9501 ^ 1'b0 ;
  assign n30427 = n30425 | n30426 ;
  assign n30428 = n6590 & n24963 ;
  assign n30429 = n5429 | n30428 ;
  assign n30430 = n30429 ^ n24498 ^ 1'b0 ;
  assign n30431 = n10557 ^ n8463 ^ n4453 ;
  assign n30432 = ~n10947 & n30431 ;
  assign n30433 = n4608 & ~n8432 ;
  assign n30434 = n30433 ^ n24000 ^ 1'b0 ;
  assign n30435 = n1149 | n7473 ;
  assign n30436 = n13456 & ~n30435 ;
  assign n30437 = n30434 & ~n30436 ;
  assign n30438 = n24985 ^ n6456 ^ 1'b0 ;
  assign n30439 = n15004 | n24449 ;
  assign n30440 = n18250 ^ n13259 ^ 1'b0 ;
  assign n30441 = n10831 & n30440 ;
  assign n30442 = n30441 ^ n1867 ^ 1'b0 ;
  assign n30443 = ~n9239 & n11883 ;
  assign n30444 = n8951 ^ n7736 ^ 1'b0 ;
  assign n30445 = n30444 ^ n12544 ^ 1'b0 ;
  assign n30446 = ~n30443 & n30445 ;
  assign n30447 = n14415 ^ n14224 ^ 1'b0 ;
  assign n30448 = n1894 | n30447 ;
  assign n30449 = n3734 & n30448 ;
  assign n30450 = n28268 ^ n20351 ^ 1'b0 ;
  assign n30451 = n14218 ^ n10826 ^ 1'b0 ;
  assign n30452 = n17782 & n30451 ;
  assign n30453 = n11118 & ~n23563 ;
  assign n30454 = n8690 ^ x108 ^ 1'b0 ;
  assign n30455 = n3515 & n3962 ;
  assign n30456 = ~n10822 & n30455 ;
  assign n30457 = n30454 & n30456 ;
  assign n30458 = ~n15896 & n25109 ;
  assign n30459 = ~n5525 & n30458 ;
  assign n30460 = n30459 ^ n18472 ^ 1'b0 ;
  assign n30461 = n10905 & ~n30460 ;
  assign n30462 = ~n2624 & n30461 ;
  assign n30463 = ~n2271 & n13384 ;
  assign n30464 = n7662 | n14800 ;
  assign n30465 = n8112 & ~n30464 ;
  assign n30466 = ~n10765 & n30465 ;
  assign n30467 = n5293 & n21741 ;
  assign n30468 = n30467 ^ n23334 ^ 1'b0 ;
  assign n30469 = n25952 ^ n8664 ^ 1'b0 ;
  assign n30470 = n12514 & n30469 ;
  assign n30472 = n12677 & n17474 ;
  assign n30473 = n30472 ^ n11936 ^ 1'b0 ;
  assign n30474 = ~n20225 & n30473 ;
  assign n30471 = x3 & ~n24454 ;
  assign n30475 = n30474 ^ n30471 ^ 1'b0 ;
  assign n30476 = n5811 & n30475 ;
  assign n30477 = ~n5379 & n14053 ;
  assign n30478 = n1741 & n30477 ;
  assign n30479 = n30478 ^ n10416 ^ 1'b0 ;
  assign n30480 = n3863 & n30479 ;
  assign n30482 = ~n4744 & n7872 ;
  assign n30481 = n8295 & ~n17910 ;
  assign n30483 = n30482 ^ n30481 ^ 1'b0 ;
  assign n30485 = n13630 ^ n8976 ^ 1'b0 ;
  assign n30486 = n9655 & ~n30485 ;
  assign n30487 = n2508 ^ n2396 ^ 1'b0 ;
  assign n30488 = n14890 & ~n30487 ;
  assign n30489 = ~n30486 & n30488 ;
  assign n30484 = ~n5509 & n15930 ;
  assign n30490 = n30489 ^ n30484 ^ 1'b0 ;
  assign n30491 = ~n30483 & n30490 ;
  assign n30492 = n522 | n29011 ;
  assign n30493 = n28316 & ~n30492 ;
  assign n30494 = ~n1545 & n8838 ;
  assign n30495 = n30494 ^ n4547 ^ 1'b0 ;
  assign n30496 = ~n4994 & n30495 ;
  assign n30497 = n30496 ^ n1371 ^ 1'b0 ;
  assign n30498 = ~n9651 & n30497 ;
  assign n30499 = n26644 ^ n26449 ^ 1'b0 ;
  assign n30500 = n16038 ^ n7966 ^ x240 ;
  assign n30504 = n8974 & ~n10598 ;
  assign n30505 = n30504 ^ n1568 ^ 1'b0 ;
  assign n30506 = n1462 & ~n30505 ;
  assign n30507 = n30506 ^ n29709 ^ 1'b0 ;
  assign n30501 = ~n11041 & n17551 ;
  assign n30502 = ~n10477 & n30501 ;
  assign n30503 = n20423 | n30502 ;
  assign n30508 = n30507 ^ n30503 ^ n27133 ;
  assign n30509 = ~n2774 & n15787 ;
  assign n30510 = ~n1105 & n8888 ;
  assign n30511 = n17555 & n30510 ;
  assign n30512 = n14128 ^ n9912 ^ 1'b0 ;
  assign n30513 = n13860 & ~n30512 ;
  assign n30514 = n25802 ^ n2901 ^ 1'b0 ;
  assign n30515 = n26338 ^ n19230 ^ n8414 ;
  assign n30516 = ~n906 & n14553 ;
  assign n30517 = n12029 ^ n5118 ^ 1'b0 ;
  assign n30518 = ~n9213 & n30517 ;
  assign n30519 = ( n1782 & ~n15549 ) | ( n1782 & n29098 ) | ( ~n15549 & n29098 ) ;
  assign n30520 = n9663 & n14479 ;
  assign n30521 = ~n30519 & n30520 ;
  assign n30522 = n19529 ^ n8144 ^ 1'b0 ;
  assign n30523 = n904 & n24288 ;
  assign n30524 = n11015 & n30523 ;
  assign n30525 = n13266 ^ n8639 ^ 1'b0 ;
  assign n30526 = n30525 ^ n13426 ^ 1'b0 ;
  assign n30527 = n1371 & n28344 ;
  assign n30528 = n20249 & n30527 ;
  assign n30529 = n22170 ^ n13545 ^ 1'b0 ;
  assign n30530 = n9813 | n21851 ;
  assign n30531 = n30530 ^ n20251 ^ 1'b0 ;
  assign n30532 = n5999 & n30531 ;
  assign n30533 = x10 & n1462 ;
  assign n30534 = n30533 ^ n20480 ^ 1'b0 ;
  assign n30535 = n2102 ^ x102 ^ 1'b0 ;
  assign n30536 = n13463 ^ n2326 ^ 1'b0 ;
  assign n30537 = n30535 & n30536 ;
  assign n30538 = n30537 ^ n6985 ^ 1'b0 ;
  assign n30539 = n18485 ^ n579 ^ 1'b0 ;
  assign n30540 = x132 | n8125 ;
  assign n30541 = ~n11206 & n30540 ;
  assign n30542 = ~n25968 & n30541 ;
  assign n30543 = n5122 & ~n27828 ;
  assign n30544 = n26836 ^ n7147 ^ 1'b0 ;
  assign n30545 = n18715 & n30544 ;
  assign n30546 = n16104 ^ n9215 ^ 1'b0 ;
  assign n30547 = ~n14965 & n30546 ;
  assign n30548 = n16181 ^ n2455 ^ 1'b0 ;
  assign n30549 = n2345 | n9529 ;
  assign n30550 = n7602 | n30549 ;
  assign n30551 = n30550 ^ n15726 ^ n15107 ;
  assign n30552 = n11149 ^ n4835 ^ x248 ;
  assign n30553 = n29179 ^ n24816 ^ n11750 ;
  assign n30554 = n30553 ^ n26539 ^ 1'b0 ;
  assign n30555 = n25122 ^ n17458 ^ 1'b0 ;
  assign n30556 = n9721 | n18804 ;
  assign n30557 = n27081 & ~n30556 ;
  assign n30558 = n29533 ^ n22010 ^ 1'b0 ;
  assign n30559 = n23560 & ~n30558 ;
  assign n30560 = ( n15285 & n22944 ) | ( n15285 & ~n28416 ) | ( n22944 & ~n28416 ) ;
  assign n30561 = n5549 & n13129 ;
  assign n30562 = n23761 & n30561 ;
  assign n30563 = n29215 ^ n9753 ^ 1'b0 ;
  assign n30564 = n26860 & n30563 ;
  assign n30565 = ~n4864 & n22053 ;
  assign n30566 = ~n3714 & n30565 ;
  assign n30567 = n19045 ^ n8058 ^ 1'b0 ;
  assign n30568 = n8816 & n30567 ;
  assign n30569 = n30566 & n30568 ;
  assign n30571 = n14916 & ~n25809 ;
  assign n30570 = n23424 | n25753 ;
  assign n30572 = n30571 ^ n30570 ^ 1'b0 ;
  assign n30573 = n2813 & ~n30572 ;
  assign n30574 = ~n17252 & n27475 ;
  assign n30575 = n3158 & n30574 ;
  assign n30576 = n19106 ^ n12557 ^ 1'b0 ;
  assign n30577 = n12673 | n30576 ;
  assign n30578 = n8683 & ~n30577 ;
  assign n30579 = n306 | n22053 ;
  assign n30580 = n9976 ^ n2409 ^ 1'b0 ;
  assign n30581 = n8728 | n27312 ;
  assign n30582 = n2062 & n2434 ;
  assign n30583 = ~n3146 & n30582 ;
  assign n30584 = n30581 | n30583 ;
  assign n30585 = n4672 & ~n30584 ;
  assign n30586 = n10858 ^ n7366 ^ 1'b0 ;
  assign n30587 = n5686 & n30586 ;
  assign n30588 = n30587 ^ n8011 ^ 1'b0 ;
  assign n30589 = n13649 & n30588 ;
  assign n30590 = n13524 & ~n30589 ;
  assign n30593 = n17965 ^ n9173 ^ 1'b0 ;
  assign n30594 = n18306 | n30593 ;
  assign n30591 = n20134 & ~n23733 ;
  assign n30592 = n30591 ^ n15457 ^ 1'b0 ;
  assign n30595 = n30594 ^ n30592 ^ 1'b0 ;
  assign n30596 = n5443 ^ n1177 ^ 1'b0 ;
  assign n30597 = ~n25334 & n30596 ;
  assign n30598 = n1734 & n6495 ;
  assign n30599 = n7306 & n30598 ;
  assign n30600 = n13807 | n30599 ;
  assign n30601 = n30600 ^ n14235 ^ 1'b0 ;
  assign n30602 = n17635 & n28142 ;
  assign n30603 = n6793 | n8956 ;
  assign n30604 = n3180 ^ n505 ^ 1'b0 ;
  assign n30605 = ~n2203 & n30604 ;
  assign n30606 = n30605 ^ n17386 ^ 1'b0 ;
  assign n30607 = ~n25494 & n30606 ;
  assign n30608 = n29860 ^ x143 ^ 1'b0 ;
  assign n30609 = n4943 ^ n1547 ^ 1'b0 ;
  assign n30610 = n7307 & n30609 ;
  assign n30611 = ( n1968 & ~n9693 ) | ( n1968 & n27826 ) | ( ~n9693 & n27826 ) ;
  assign n30612 = ~n15046 & n30611 ;
  assign n30613 = n4230 & n7002 ;
  assign n30614 = ~n5690 & n30613 ;
  assign n30615 = n24715 ^ n22673 ^ 1'b0 ;
  assign n30616 = ~n23114 & n30615 ;
  assign n30618 = n3329 ^ n1508 ^ 1'b0 ;
  assign n30617 = n8278 & ~n11891 ;
  assign n30619 = n30618 ^ n30617 ^ 1'b0 ;
  assign n30620 = n30619 ^ n22982 ^ n2216 ;
  assign n30621 = n1851 & n27799 ;
  assign n30622 = n7444 | n30621 ;
  assign n30623 = n5062 ^ n4004 ^ 1'b0 ;
  assign n30624 = n14122 & ~n24073 ;
  assign n30625 = ~x0 & n30624 ;
  assign n30626 = n2297 | n26613 ;
  assign n30627 = n15576 & n30626 ;
  assign n30628 = n9892 | n17284 ;
  assign n30629 = n18952 & n30628 ;
  assign n30630 = ~n30627 & n30629 ;
  assign n30631 = n6844 ^ n2301 ^ 1'b0 ;
  assign n30632 = ~n11470 & n11506 ;
  assign n30633 = n30631 & n30632 ;
  assign n30634 = n1568 & n13539 ;
  assign n30635 = n30634 ^ n11496 ^ 1'b0 ;
  assign n30636 = n27818 ^ n455 ^ 1'b0 ;
  assign n30637 = n30635 | n30636 ;
  assign n30638 = ~n1250 & n13664 ;
  assign n30639 = n30638 ^ n5529 ^ 1'b0 ;
  assign n30640 = n9632 & ~n21749 ;
  assign n30641 = ( n4421 & n30639 ) | ( n4421 & ~n30640 ) | ( n30639 & ~n30640 ) ;
  assign n30642 = n9319 | n11539 ;
  assign n30643 = ~n13941 & n16348 ;
  assign n30644 = n30643 ^ n7285 ^ 1'b0 ;
  assign n30645 = n30642 & n30644 ;
  assign n30646 = n29257 ^ n21841 ^ n8308 ;
  assign n30647 = n15692 ^ n6624 ^ 1'b0 ;
  assign n30648 = ~n825 & n30647 ;
  assign n30649 = n5767 & n30648 ;
  assign n30650 = ( n1623 & ~n2594 ) | ( n1623 & n30649 ) | ( ~n2594 & n30649 ) ;
  assign n30651 = n24897 ^ n3481 ^ 1'b0 ;
  assign n30652 = n6739 & n30651 ;
  assign n30653 = n2691 & n14234 ;
  assign n30654 = n30653 ^ n4131 ^ 1'b0 ;
  assign n30655 = ~n22032 & n30654 ;
  assign n30656 = n19581 & ~n29713 ;
  assign n30657 = n14311 ^ n1738 ^ 1'b0 ;
  assign n30658 = n24290 & n30657 ;
  assign n30662 = n2702 | n5742 ;
  assign n30663 = n3451 & ~n30662 ;
  assign n30660 = n15652 ^ n4966 ^ 1'b0 ;
  assign n30659 = n6888 | n24703 ;
  assign n30661 = n30660 ^ n30659 ^ 1'b0 ;
  assign n30664 = n30663 ^ n30661 ^ 1'b0 ;
  assign n30665 = n28374 ^ n18875 ^ 1'b0 ;
  assign n30666 = ( n5209 & n10657 ) | ( n5209 & n30665 ) | ( n10657 & n30665 ) ;
  assign n30667 = n13710 ^ n4953 ^ 1'b0 ;
  assign n30668 = ~n6912 & n16771 ;
  assign n30669 = ( n22609 & n28597 ) | ( n22609 & ~n30668 ) | ( n28597 & ~n30668 ) ;
  assign n30670 = n2687 | n30669 ;
  assign n30671 = ~n1160 & n7375 ;
  assign n30672 = n25420 | n30671 ;
  assign n30673 = n24506 ^ n7109 ^ 1'b0 ;
  assign n30674 = ( n2338 & n3367 ) | ( n2338 & n15515 ) | ( n3367 & n15515 ) ;
  assign n30675 = x82 | x141 ;
  assign n30676 = ~n30674 & n30675 ;
  assign n30677 = n7602 ^ n5779 ^ 1'b0 ;
  assign n30678 = n6689 & n30677 ;
  assign n30679 = n17610 & n30678 ;
  assign n30680 = n30679 ^ n9612 ^ 1'b0 ;
  assign n30681 = n8333 ^ n2103 ^ 1'b0 ;
  assign n30682 = x114 & x237 ;
  assign n30683 = ~x114 & n30682 ;
  assign n30684 = n1586 | n4399 ;
  assign n30685 = n1586 & ~n30684 ;
  assign n30686 = n589 | n1078 ;
  assign n30687 = n1078 & ~n30686 ;
  assign n30688 = n30685 | n30687 ;
  assign n30689 = n30683 & ~n30688 ;
  assign n30690 = n1684 & ~n1968 ;
  assign n30691 = ~n1684 & n30690 ;
  assign n30692 = n7397 & ~n30691 ;
  assign n30693 = ~n17606 & n30692 ;
  assign n30694 = n30689 & n30693 ;
  assign n30695 = ~n2841 & n8360 ;
  assign n30696 = n15504 & n30695 ;
  assign n30697 = n1828 & ~n30696 ;
  assign n30698 = n30697 ^ n4595 ^ 1'b0 ;
  assign n30699 = n18725 & ~n30698 ;
  assign n30700 = n18244 ^ n886 ^ 1'b0 ;
  assign n30701 = ~n7825 & n30700 ;
  assign n30702 = n25053 ^ n14736 ^ 1'b0 ;
  assign n30703 = n7089 & n30702 ;
  assign n30704 = n799 & n30703 ;
  assign n30705 = ( x100 & ~n5184 ) | ( x100 & n14677 ) | ( ~n5184 & n14677 ) ;
  assign n30706 = n425 & n9389 ;
  assign n30707 = n4753 & n19275 ;
  assign n30708 = n25580 ^ n17264 ^ n6075 ;
  assign n30709 = n22614 | n24922 ;
  assign n30710 = n30709 ^ n5344 ^ 1'b0 ;
  assign n30713 = n458 & ~n5214 ;
  assign n30714 = ~n7061 & n30713 ;
  assign n30711 = n6989 ^ n6794 ^ 1'b0 ;
  assign n30712 = ~n13283 & n30711 ;
  assign n30715 = n30714 ^ n30712 ^ 1'b0 ;
  assign n30716 = n19634 ^ n17562 ^ 1'b0 ;
  assign n30717 = n2770 | n30716 ;
  assign n30718 = n27853 ^ n24131 ^ 1'b0 ;
  assign n30719 = n30717 | n30718 ;
  assign n30720 = n4309 & n11747 ;
  assign n30721 = n21965 & n28426 ;
  assign n30722 = n1055 & n11599 ;
  assign n30723 = n8578 & n30722 ;
  assign n30724 = n1295 | n2296 ;
  assign n30725 = n30724 ^ n17285 ^ 1'b0 ;
  assign n30726 = ( n6357 & ~n30723 ) | ( n6357 & n30725 ) | ( ~n30723 & n30725 ) ;
  assign n30727 = n30721 & ~n30726 ;
  assign n30728 = ~n4288 & n6453 ;
  assign n30729 = n30728 ^ n8133 ^ 1'b0 ;
  assign n30730 = ~n6620 & n23630 ;
  assign n30731 = ~n30729 & n30730 ;
  assign n30732 = n22874 ^ n7939 ^ 1'b0 ;
  assign n30733 = n17572 ^ n5971 ^ 1'b0 ;
  assign n30734 = n5091 & ~n30733 ;
  assign n30735 = n17360 ^ n11153 ^ 1'b0 ;
  assign n30736 = ~n3911 & n30735 ;
  assign n30737 = n15278 | n28970 ;
  assign n30738 = ~n7491 & n7631 ;
  assign n30739 = n4218 ^ x242 ^ 1'b0 ;
  assign n30740 = n3121 & ~n30739 ;
  assign n30741 = n5311 | n10880 ;
  assign n30742 = n11367 & n19714 ;
  assign n30743 = n30742 ^ n8260 ^ 1'b0 ;
  assign n30744 = ( n1360 & ~n14311 ) | ( n1360 & n26736 ) | ( ~n14311 & n26736 ) ;
  assign n30745 = n12167 | n17364 ;
  assign n30746 = n17872 ^ n9276 ^ n6582 ;
  assign n30747 = n6291 & n30490 ;
  assign n30748 = n25377 ^ n17114 ^ 1'b0 ;
  assign n30749 = n9522 & ~n22935 ;
  assign n30750 = n30749 ^ n13070 ^ 1'b0 ;
  assign n30751 = n16322 | n25579 ;
  assign n30752 = n6621 & ~n17074 ;
  assign n30753 = n30751 & n30752 ;
  assign n30754 = n6722 | n9529 ;
  assign n30755 = n9516 ^ n3996 ^ 1'b0 ;
  assign n30756 = n4195 & ~n30755 ;
  assign n30757 = n30756 ^ n30245 ^ 1'b0 ;
  assign n30758 = n30754 & n30757 ;
  assign n30759 = n30758 ^ n19752 ^ 1'b0 ;
  assign n30760 = n4597 & ~n19812 ;
  assign n30761 = ~n13064 & n30760 ;
  assign n30762 = n30761 ^ n20044 ^ 1'b0 ;
  assign n30763 = n15950 ^ n10889 ^ 1'b0 ;
  assign n30764 = n12502 & ~n30763 ;
  assign n30765 = n3855 & n20373 ;
  assign n30766 = x171 | n755 ;
  assign n30767 = ( ~n28461 & n30765 ) | ( ~n28461 & n30766 ) | ( n30765 & n30766 ) ;
  assign n30768 = n1633 | n16177 ;
  assign n30769 = n30768 ^ n8107 ^ 1'b0 ;
  assign n30770 = n2634 & ~n30769 ;
  assign n30771 = n12320 ^ n5398 ^ 1'b0 ;
  assign n30772 = n9429 & ~n18703 ;
  assign n30773 = n347 & n30772 ;
  assign n30774 = ~n8303 & n30773 ;
  assign n30775 = n14652 & n22601 ;
  assign n30776 = n30775 ^ n3481 ^ 1'b0 ;
  assign n30777 = ~n10663 & n16710 ;
  assign n30778 = n2920 & n30777 ;
  assign n30779 = ~n21391 & n30778 ;
  assign n30780 = ~n7496 & n30779 ;
  assign n30781 = n30780 ^ n20442 ^ n11627 ;
  assign n30782 = n30781 ^ n2301 ^ 1'b0 ;
  assign n30783 = n2657 | n24082 ;
  assign n30784 = n14568 ^ n3494 ^ 1'b0 ;
  assign n30785 = n30784 ^ n28167 ^ 1'b0 ;
  assign n30786 = n9704 & ~n21240 ;
  assign n30787 = n30786 ^ n464 ^ 1'b0 ;
  assign n30788 = n30787 ^ n18718 ^ 1'b0 ;
  assign n30789 = n18248 ^ n1271 ^ 1'b0 ;
  assign n30790 = n400 & n1690 ;
  assign n30791 = n838 & ~n7179 ;
  assign n30792 = n30791 ^ n15102 ^ 1'b0 ;
  assign n30793 = n30790 & n30792 ;
  assign n30794 = n23610 | n29675 ;
  assign n30795 = n30794 ^ n22236 ^ 1'b0 ;
  assign n30796 = n24809 ^ n18383 ^ n17872 ;
  assign n30797 = n20279 ^ x96 ^ 1'b0 ;
  assign n30798 = n8868 & n30797 ;
  assign n30799 = n5309 & n30798 ;
  assign n30800 = n10506 ^ n2693 ^ 1'b0 ;
  assign n30801 = n30799 & ~n30800 ;
  assign n30802 = ~n2096 & n22252 ;
  assign n30803 = n30802 ^ n7130 ^ 1'b0 ;
  assign n30804 = ~n27639 & n30803 ;
  assign n30805 = n30804 ^ n17812 ^ 1'b0 ;
  assign n30806 = n16363 & n16505 ;
  assign n30807 = n30806 ^ n2321 ^ 1'b0 ;
  assign n30808 = n4501 & n11330 ;
  assign n30809 = n22829 | n30808 ;
  assign n30810 = n719 & n15680 ;
  assign n30811 = n12725 ^ n11549 ^ n9761 ;
  assign n30812 = n30811 ^ n3678 ^ 1'b0 ;
  assign n30813 = n14714 & ~n30812 ;
  assign n30814 = ~n17747 & n30813 ;
  assign n30815 = ( ~n5127 & n30810 ) | ( ~n5127 & n30814 ) | ( n30810 & n30814 ) ;
  assign n30816 = ( ~n1254 & n2501 ) | ( ~n1254 & n30815 ) | ( n2501 & n30815 ) ;
  assign n30817 = n13082 ^ n12168 ^ 1'b0 ;
  assign n30818 = ~n9068 & n30817 ;
  assign n30819 = n30818 ^ n18554 ^ 1'b0 ;
  assign n30820 = n5186 ^ n4315 ^ 1'b0 ;
  assign n30821 = n12876 ^ n9722 ^ 1'b0 ;
  assign n30822 = n30821 ^ n8679 ^ 1'b0 ;
  assign n30823 = n372 | n30822 ;
  assign n30824 = n23869 ^ n23196 ^ 1'b0 ;
  assign n30825 = n19435 & n22394 ;
  assign n30826 = n8440 | n18927 ;
  assign n30827 = n14754 & n28839 ;
  assign n30828 = ~n4860 & n16812 ;
  assign n30829 = ~n2821 & n30828 ;
  assign n30830 = n7170 | n30829 ;
  assign n30834 = ~n1116 & n30410 ;
  assign n30831 = n13668 ^ n3594 ^ 1'b0 ;
  assign n30832 = n11072 | n30831 ;
  assign n30833 = n21054 | n30832 ;
  assign n30835 = n30834 ^ n30833 ^ 1'b0 ;
  assign n30836 = n24781 ^ n23683 ^ n21445 ;
  assign n30837 = n14680 ^ n10490 ^ 1'b0 ;
  assign n30838 = ( n1596 & ~n15950 ) | ( n1596 & n30837 ) | ( ~n15950 & n30837 ) ;
  assign n30839 = n3744 & ~n13636 ;
  assign n30840 = ~n1123 & n30839 ;
  assign n30841 = n30840 ^ n5188 ^ 1'b0 ;
  assign n30842 = n4113 & ~n30841 ;
  assign n30843 = n6398 & ~n17758 ;
  assign n30844 = n30842 & n30843 ;
  assign n30845 = ~n11353 & n21967 ;
  assign n30846 = n3408 & n30845 ;
  assign n30847 = n3416 & ~n30846 ;
  assign n30848 = n3775 & n4565 ;
  assign n30849 = n22825 ^ n14175 ^ 1'b0 ;
  assign n30850 = n25255 ^ n14794 ^ n14595 ;
  assign n30851 = n4718 ^ n3483 ^ 1'b0 ;
  assign n30852 = n5772 & ~n30851 ;
  assign n30853 = n3028 | n7536 ;
  assign n30854 = n27874 ^ n26006 ^ 1'b0 ;
  assign n30855 = n30853 | n30854 ;
  assign n30856 = n26890 | n30855 ;
  assign n30857 = n30852 | n30856 ;
  assign n30858 = n13964 | n19564 ;
  assign n30859 = n30858 ^ n17415 ^ 1'b0 ;
  assign n30860 = n18122 & n19271 ;
  assign n30861 = n30860 ^ n25518 ^ 1'b0 ;
  assign n30862 = n8722 | n9345 ;
  assign n30863 = n30862 ^ n25628 ^ 1'b0 ;
  assign n30864 = n6496 ^ n2868 ^ 1'b0 ;
  assign n30865 = n7507 | n30864 ;
  assign n30866 = ~n13060 & n30865 ;
  assign n30867 = n30866 ^ n6031 ^ 1'b0 ;
  assign n30868 = n7467 & ~n22039 ;
  assign n30869 = n30868 ^ n19553 ^ 1'b0 ;
  assign n30872 = n8785 ^ n8309 ^ 1'b0 ;
  assign n30873 = n10399 | n30872 ;
  assign n30874 = n4011 | n30873 ;
  assign n30870 = n7109 ^ n1859 ^ 1'b0 ;
  assign n30871 = n10512 & ~n30870 ;
  assign n30875 = n30874 ^ n30871 ^ 1'b0 ;
  assign n30876 = n349 | n12982 ;
  assign n30877 = n1561 & n10973 ;
  assign n30878 = ~n1561 & n30877 ;
  assign n30879 = n3474 | n4088 ;
  assign n30880 = n3474 & ~n30879 ;
  assign n30881 = ~x195 & n30880 ;
  assign n30882 = n30881 ^ n5775 ^ 1'b0 ;
  assign n30883 = x24 & x232 ;
  assign n30884 = ~x24 & n30883 ;
  assign n30885 = x161 & n3601 ;
  assign n30886 = ~n3601 & n30885 ;
  assign n30887 = n3152 & ~n30886 ;
  assign n30888 = n30884 & n30887 ;
  assign n30889 = n30882 | n30888 ;
  assign n30890 = n30882 & ~n30889 ;
  assign n30891 = n5622 & ~n30890 ;
  assign n30892 = ~n5622 & n30891 ;
  assign n30893 = n30878 | n30892 ;
  assign n30894 = n30878 & ~n30893 ;
  assign n30895 = n6585 | n11665 ;
  assign n30896 = n30894 & ~n30895 ;
  assign n30897 = n1733 | n14306 ;
  assign n30898 = n30896 & ~n30897 ;
  assign n30899 = n883 | n1583 ;
  assign n30900 = n1583 & ~n30899 ;
  assign n30901 = n7723 & ~n30900 ;
  assign n30902 = ~n7723 & n30901 ;
  assign n30903 = n30902 ^ n4516 ^ 1'b0 ;
  assign n30904 = n30898 | n30903 ;
  assign n30905 = n30898 & ~n30904 ;
  assign n30906 = n9609 & ~n21863 ;
  assign n30907 = ~n9609 & n30906 ;
  assign n30908 = n1077 & ~n17373 ;
  assign n30909 = n30907 & n30908 ;
  assign n30910 = n17120 | n30909 ;
  assign n30911 = n30905 & ~n30910 ;
  assign n30912 = n17794 ^ n4512 ^ 1'b0 ;
  assign n30913 = n23864 & ~n30912 ;
  assign n30914 = n10096 ^ n8873 ^ 1'b0 ;
  assign n30915 = n18904 | n30914 ;
  assign n30916 = n3956 | n30915 ;
  assign n30919 = n18307 ^ n7634 ^ 1'b0 ;
  assign n30920 = n4195 ^ n2037 ^ 1'b0 ;
  assign n30921 = n25405 & n30920 ;
  assign n30922 = ( n29088 & n30919 ) | ( n29088 & ~n30921 ) | ( n30919 & ~n30921 ) ;
  assign n30917 = n7651 ^ n6868 ^ n6154 ;
  assign n30918 = ~n5579 & n30917 ;
  assign n30923 = n30922 ^ n30918 ^ n16410 ;
  assign n30924 = n13266 ^ n676 ^ 1'b0 ;
  assign n30925 = n1356 & ~n30924 ;
  assign n30926 = n13762 | n22610 ;
  assign n30927 = n25977 | n30926 ;
  assign n30928 = n24347 ^ n1424 ^ 1'b0 ;
  assign n30929 = n12652 | n24914 ;
  assign n30930 = n24835 ^ n13969 ^ 1'b0 ;
  assign n30931 = n30929 | n30930 ;
  assign n30932 = n12517 ^ n3296 ^ 1'b0 ;
  assign n30933 = x176 & n30932 ;
  assign n30934 = n14462 & ~n30933 ;
  assign n30935 = n4575 & n8073 ;
  assign n30936 = n30935 ^ n9987 ^ 1'b0 ;
  assign n30937 = n14066 ^ n10336 ^ n10155 ;
  assign n30938 = n3149 & ~n10886 ;
  assign n30939 = n26307 & n30938 ;
  assign n30940 = n5498 ^ n2872 ^ n2039 ;
  assign n30941 = ~n17330 & n30940 ;
  assign n30942 = n16438 & ~n19229 ;
  assign n30943 = n15896 | n24148 ;
  assign n30944 = n25043 & ~n30943 ;
  assign n30945 = n24015 | n28329 ;
  assign n30946 = n16693 ^ n14532 ^ 1'b0 ;
  assign n30947 = n9595 ^ n1051 ^ 1'b0 ;
  assign n30948 = ~n10731 & n22714 ;
  assign n30949 = n30947 & n30948 ;
  assign n30950 = n18195 & ~n30949 ;
  assign n30951 = n22156 ^ n16866 ^ n2870 ;
  assign n30952 = n16412 & ~n30412 ;
  assign n30953 = n3546 & n21879 ;
  assign n30954 = n3316 | n30953 ;
  assign n30955 = n4521 & ~n30954 ;
  assign n30956 = n14181 ^ n11576 ^ 1'b0 ;
  assign n30957 = n3747 & ~n5442 ;
  assign n30958 = n30957 ^ n6532 ^ 1'b0 ;
  assign n30959 = n23244 & n30958 ;
  assign n30960 = n30959 ^ n9515 ^ 1'b0 ;
  assign n30961 = n19704 ^ n6846 ^ 1'b0 ;
  assign n30962 = ( n10072 & n15138 ) | ( n10072 & ~n30961 ) | ( n15138 & ~n30961 ) ;
  assign n30963 = n703 & n7784 ;
  assign n30964 = ~n1274 & n28761 ;
  assign n30965 = n26381 & ~n30964 ;
  assign n30966 = n30965 ^ n16066 ^ 1'b0 ;
  assign n30967 = n11838 ^ n3561 ^ 1'b0 ;
  assign n30968 = ~n30092 & n30967 ;
  assign n30969 = n7205 & ~n29136 ;
  assign n30970 = ~n1208 & n5280 ;
  assign n30971 = n14172 & n30970 ;
  assign n30972 = n30971 ^ n16129 ^ 1'b0 ;
  assign n30973 = ~n29286 & n30972 ;
  assign n30979 = n406 & ~n12538 ;
  assign n30980 = n22709 & n30979 ;
  assign n30975 = n7895 ^ n1705 ^ 1'b0 ;
  assign n30976 = ~n2881 & n30975 ;
  assign n30977 = ( n985 & ~n16947 ) | ( n985 & n30976 ) | ( ~n16947 & n30976 ) ;
  assign n30974 = n10120 & n11585 ;
  assign n30978 = n30977 ^ n30974 ^ 1'b0 ;
  assign n30981 = n30980 ^ n30978 ^ n11872 ;
  assign n30982 = ~n13958 & n30981 ;
  assign n30983 = n16679 & ~n26836 ;
  assign n30984 = ( ~n5065 & n7646 ) | ( ~n5065 & n29838 ) | ( n7646 & n29838 ) ;
  assign n30985 = n21035 | n30984 ;
  assign n30986 = n30985 ^ n23422 ^ 1'b0 ;
  assign n30987 = n6636 & n11743 ;
  assign n30988 = n30987 ^ n17238 ^ 1'b0 ;
  assign n30989 = n16280 | n30988 ;
  assign n30990 = n21191 ^ n18041 ^ n7624 ;
  assign n30991 = n5686 & ~n28636 ;
  assign n30992 = n30991 ^ n27489 ^ n3923 ;
  assign n30993 = ~n340 & n1501 ;
  assign n30994 = n340 & n30993 ;
  assign n30995 = n1486 | n30994 ;
  assign n30996 = n15018 & n21781 ;
  assign n30997 = n30996 ^ n30592 ^ 1'b0 ;
  assign n30998 = n25413 ^ n14335 ^ 1'b0 ;
  assign n30999 = n4988 & n30998 ;
  assign n31000 = n3190 & ~n12569 ;
  assign n31001 = n7097 & ~n26588 ;
  assign n31002 = n31001 ^ n6499 ^ 1'b0 ;
  assign n31003 = n31000 & ~n31002 ;
  assign n31004 = ~n30999 & n31003 ;
  assign n31005 = n25229 ^ n11162 ^ 1'b0 ;
  assign n31006 = n11751 ^ n7415 ^ n2096 ;
  assign n31007 = ~n24887 & n28627 ;
  assign n31008 = n13803 & ~n31007 ;
  assign n31009 = n31008 ^ n6257 ^ 1'b0 ;
  assign n31010 = n14794 & n31009 ;
  assign n31011 = n31010 ^ n11274 ^ n7984 ;
  assign n31012 = ~n7292 & n14428 ;
  assign n31013 = n11730 ^ n8363 ^ 1'b0 ;
  assign n31014 = n31012 | n31013 ;
  assign n31015 = n2841 & n4770 ;
  assign n31016 = n31015 ^ n28009 ^ 1'b0 ;
  assign n31017 = n3474 | n31016 ;
  assign n31018 = n7716 | n13412 ;
  assign n31019 = n6483 ^ n1738 ^ 1'b0 ;
  assign n31020 = n31019 ^ n13412 ^ 1'b0 ;
  assign n31021 = n29660 ^ n5272 ^ 1'b0 ;
  assign n31022 = n23844 ^ n6785 ^ n436 ;
  assign n31023 = ~n1490 & n4794 ;
  assign n31024 = n15544 ^ n4493 ^ 1'b0 ;
  assign n31025 = n25898 ^ n6994 ^ 1'b0 ;
  assign n31026 = n9921 ^ n6679 ^ 1'b0 ;
  assign n31027 = n11442 & n31026 ;
  assign n31028 = n31027 ^ n16146 ^ n2640 ;
  assign n31029 = n4977 ^ n3904 ^ 1'b0 ;
  assign n31030 = n10077 ^ n7972 ^ 1'b0 ;
  assign n31031 = n4562 ^ n710 ^ 1'b0 ;
  assign n31032 = n31031 ^ n29539 ^ 1'b0 ;
  assign n31033 = ~n2378 & n31032 ;
  assign n31034 = n26630 ^ n2746 ^ 1'b0 ;
  assign n31035 = n17308 & ~n31034 ;
  assign n31036 = n18356 ^ n12313 ^ n2092 ;
  assign n31037 = n16252 ^ n5056 ^ 1'b0 ;
  assign n31038 = n31036 & ~n31037 ;
  assign n31039 = n1664 ^ n772 ^ 1'b0 ;
  assign n31040 = n28940 ^ n7620 ^ 1'b0 ;
  assign n31041 = n2963 & ~n9839 ;
  assign n31042 = ~n2657 & n31041 ;
  assign n31043 = n19098 ^ n13401 ^ 1'b0 ;
  assign n31044 = n11155 & n31043 ;
  assign n31045 = n27380 & n31044 ;
  assign n31046 = n15300 ^ n11732 ^ 1'b0 ;
  assign n31047 = n29616 | n31046 ;
  assign n31048 = n4970 ^ n759 ^ 1'b0 ;
  assign n31049 = n31048 ^ n22096 ^ n5365 ;
  assign n31050 = n16822 & n29052 ;
  assign n31051 = n6854 ^ n643 ^ 1'b0 ;
  assign n31052 = n31051 ^ n22015 ^ n353 ;
  assign n31053 = n31052 ^ n11034 ^ 1'b0 ;
  assign n31054 = n3348 ^ n1894 ^ 1'b0 ;
  assign n31055 = ~n13832 & n31054 ;
  assign n31056 = n5400 & ~n7173 ;
  assign n31057 = n2098 & n31056 ;
  assign n31058 = n6254 & n31057 ;
  assign n31059 = n4040 ^ n2224 ^ 1'b0 ;
  assign n31060 = ~n21660 & n31059 ;
  assign n31061 = n5132 | n31060 ;
  assign n31062 = ( ~n11449 & n25652 ) | ( ~n11449 & n31061 ) | ( n25652 & n31061 ) ;
  assign n31065 = n10526 ^ n4509 ^ 1'b0 ;
  assign n31066 = ~n12515 & n31065 ;
  assign n31063 = n11508 ^ n4638 ^ 1'b0 ;
  assign n31064 = n4105 & ~n31063 ;
  assign n31067 = n31066 ^ n31064 ^ 1'b0 ;
  assign n31068 = n19758 & n21808 ;
  assign n31069 = n20259 | n27680 ;
  assign n31070 = n31069 ^ n13773 ^ 1'b0 ;
  assign n31071 = ~n13767 & n28561 ;
  assign n31072 = ~n18081 & n31071 ;
  assign n31073 = n11647 ^ n6620 ^ 1'b0 ;
  assign n31075 = n14376 ^ n8419 ^ 1'b0 ;
  assign n31074 = n1749 & ~n3494 ;
  assign n31076 = n31075 ^ n31074 ^ n25426 ;
  assign n31077 = n400 | n2875 ;
  assign n31078 = n8758 | n28756 ;
  assign n31079 = n4995 | n14444 ;
  assign n31080 = n13090 & n31079 ;
  assign n31081 = n1219 & ~n22960 ;
  assign n31082 = ( n3901 & n9753 ) | ( n3901 & ~n14114 ) | ( n9753 & ~n14114 ) ;
  assign n31083 = n8390 | n10820 ;
  assign n31084 = ~n9548 & n31083 ;
  assign n31085 = n31084 ^ n9098 ^ 1'b0 ;
  assign n31086 = n31082 & n31085 ;
  assign n31087 = ~n4876 & n17967 ;
  assign n31088 = n12274 & ~n31087 ;
  assign n31089 = n31088 ^ n2953 ^ 1'b0 ;
  assign n31090 = n25300 ^ n14698 ^ 1'b0 ;
  assign n31091 = n8884 ^ n4266 ^ 1'b0 ;
  assign n31092 = n31090 | n31091 ;
  assign n31093 = n31092 ^ n3777 ^ 1'b0 ;
  assign n31094 = n2959 & n31093 ;
  assign n31095 = n31094 ^ n26836 ^ 1'b0 ;
  assign n31096 = n5497 & n17654 ;
  assign n31097 = n16548 ^ n11118 ^ 1'b0 ;
  assign n31098 = n21497 ^ n13268 ^ 1'b0 ;
  assign n31099 = n29712 & n31098 ;
  assign n31100 = n27728 ^ n1968 ^ 1'b0 ;
  assign n31101 = n8835 & ~n31100 ;
  assign n31102 = ( n1810 & ~n2574 ) | ( n1810 & n20181 ) | ( ~n2574 & n20181 ) ;
  assign n31103 = n16560 ^ n14105 ^ 1'b0 ;
  assign n31104 = n31102 & n31103 ;
  assign n31105 = n10709 & ~n16618 ;
  assign n31106 = n15061 & n17053 ;
  assign n31107 = n642 & n31106 ;
  assign n31108 = n13362 ^ n7418 ^ 1'b0 ;
  assign n31109 = ~n15895 & n23079 ;
  assign n31110 = n31108 & n31109 ;
  assign n31111 = ~n2274 & n31110 ;
  assign n31112 = n31111 ^ n23881 ^ 1'b0 ;
  assign n31113 = n31107 | n31112 ;
  assign n31114 = n11713 | n19102 ;
  assign n31115 = ~n2178 & n3670 ;
  assign n31116 = n13482 & n31115 ;
  assign n31117 = n6075 | n19424 ;
  assign n31118 = n31116 & ~n31117 ;
  assign n31119 = n30961 ^ n26176 ^ 1'b0 ;
  assign n31120 = n498 | n20699 ;
  assign n31121 = n19372 | n31120 ;
  assign n31122 = n7757 & ~n18053 ;
  assign n31123 = n7693 ^ n5962 ^ 1'b0 ;
  assign n31124 = ~n842 & n12943 ;
  assign n31125 = n31124 ^ n7347 ^ 1'b0 ;
  assign n31126 = n3714 | n31125 ;
  assign n31127 = ( ~n7862 & n9365 ) | ( ~n7862 & n20716 ) | ( n9365 & n20716 ) ;
  assign n31128 = n27624 ^ n15051 ^ 1'b0 ;
  assign n31129 = n2689 & n31128 ;
  assign n31130 = n5121 | n17229 ;
  assign n31131 = n31130 ^ n26175 ^ 1'b0 ;
  assign n31132 = n18098 | n31131 ;
  assign n31133 = n13337 ^ x159 ^ 1'b0 ;
  assign n31134 = ~n26315 & n31133 ;
  assign n31135 = n7109 & ~n7634 ;
  assign n31136 = n31135 ^ n7975 ^ 1'b0 ;
  assign n31137 = n11508 ^ n2177 ^ 1'b0 ;
  assign n31138 = n5061 & n31137 ;
  assign n31139 = ~n6440 & n31138 ;
  assign n31140 = ~n31136 & n31139 ;
  assign n31141 = n30802 ^ n13931 ^ 1'b0 ;
  assign n31142 = ~n13353 & n31141 ;
  assign n31143 = n20977 ^ n19365 ^ 1'b0 ;
  assign n31144 = n20709 & n31143 ;
  assign n31145 = n16606 ^ n9243 ^ 1'b0 ;
  assign n31146 = n23701 ^ n19788 ^ 1'b0 ;
  assign n31147 = n12611 & n15857 ;
  assign n31148 = n31147 ^ n24453 ^ 1'b0 ;
  assign n31149 = n24632 ^ n19050 ^ 1'b0 ;
  assign n31150 = ~n3195 & n31149 ;
  assign n31151 = n27447 ^ n8246 ^ 1'b0 ;
  assign n31152 = n24169 ^ n10884 ^ 1'b0 ;
  assign n31153 = n31152 ^ n1330 ^ 1'b0 ;
  assign n31154 = n31153 ^ n8722 ^ 1'b0 ;
  assign n31155 = n7874 ^ n3698 ^ 1'b0 ;
  assign n31156 = n15551 & n26544 ;
  assign n31157 = n31155 & n31156 ;
  assign n31158 = n3155 & ~n31157 ;
  assign n31159 = n10359 ^ n2137 ^ 1'b0 ;
  assign n31160 = n9767 & ~n31159 ;
  assign n31161 = n31160 ^ n7876 ^ 1'b0 ;
  assign n31162 = n14030 ^ n12364 ^ 1'b0 ;
  assign n31163 = n2369 & ~n31162 ;
  assign n31164 = n3760 & ~n17009 ;
  assign n31165 = ~n8281 & n31164 ;
  assign n31166 = n21877 ^ n18396 ^ 1'b0 ;
  assign n31167 = n13420 & ~n31166 ;
  assign n31168 = n8153 & n31167 ;
  assign n31169 = x190 & ~n2099 ;
  assign n31170 = ~n15434 & n31169 ;
  assign n31171 = n31170 ^ n4615 ^ 1'b0 ;
  assign n31172 = n18768 & ~n25266 ;
  assign n31173 = ~n404 & n21801 ;
  assign n31175 = n10135 ^ n10075 ^ 1'b0 ;
  assign n31176 = ~n14080 & n31175 ;
  assign n31174 = n21887 ^ n579 ^ 1'b0 ;
  assign n31177 = n31176 ^ n31174 ^ n16679 ;
  assign n31178 = n5132 ^ n2799 ^ 1'b0 ;
  assign n31180 = n8564 ^ n7814 ^ 1'b0 ;
  assign n31179 = n8997 & ~n26125 ;
  assign n31181 = n31180 ^ n31179 ^ 1'b0 ;
  assign n31182 = n8936 ^ n415 ^ 1'b0 ;
  assign n31183 = n31182 ^ n26347 ^ 1'b0 ;
  assign n31184 = n9698 | n31183 ;
  assign n31185 = ~n9218 & n21234 ;
  assign n31186 = ~n466 & n21479 ;
  assign n31187 = ~n30385 & n31186 ;
  assign n31191 = n15227 ^ n1590 ^ 1'b0 ;
  assign n31192 = ~n4719 & n31191 ;
  assign n31193 = ~n22675 & n31192 ;
  assign n31194 = n6805 & n31193 ;
  assign n31188 = n9130 ^ n2230 ^ 1'b0 ;
  assign n31189 = n31188 ^ n7999 ^ 1'b0 ;
  assign n31190 = n24586 & ~n31189 ;
  assign n31195 = n31194 ^ n31190 ^ 1'b0 ;
  assign n31196 = n6144 & n15196 ;
  assign n31197 = n27872 ^ n3485 ^ 1'b0 ;
  assign n31198 = n31196 & ~n31197 ;
  assign n31199 = n31198 ^ n24013 ^ 1'b0 ;
  assign n31200 = n16363 & n31199 ;
  assign n31201 = ~n25187 & n31200 ;
  assign n31202 = n12873 ^ n9886 ^ 1'b0 ;
  assign n31203 = n10934 & n31202 ;
  assign n31204 = n7148 & n31203 ;
  assign n31205 = n31204 ^ n25935 ^ 1'b0 ;
  assign n31206 = n31205 ^ n3059 ^ 1'b0 ;
  assign n31207 = n10385 ^ n2418 ^ 1'b0 ;
  assign n31208 = n15176 | n31207 ;
  assign n31209 = n2413 & n31208 ;
  assign n31210 = n4562 ^ n613 ^ 1'b0 ;
  assign n31211 = ( n9275 & ~n14994 ) | ( n9275 & n24484 ) | ( ~n14994 & n24484 ) ;
  assign n31212 = n13805 ^ n5616 ^ 1'b0 ;
  assign n31213 = n31211 & n31212 ;
  assign n31214 = n24443 ^ n11253 ^ n542 ;
  assign n31215 = n6931 | n22582 ;
  assign n31216 = n14371 & ~n31215 ;
  assign n31217 = ~n8642 & n26097 ;
  assign n31218 = ~n4241 & n31217 ;
  assign n31219 = n30751 | n31218 ;
  assign n31220 = n31219 ^ n21560 ^ 1'b0 ;
  assign n31222 = n8133 | n10763 ;
  assign n31223 = n31222 ^ n12878 ^ 1'b0 ;
  assign n31221 = n4693 & ~n10382 ;
  assign n31224 = n31223 ^ n31221 ^ 1'b0 ;
  assign n31225 = n15514 & ~n16105 ;
  assign n31226 = n31225 ^ n473 ^ 1'b0 ;
  assign n31227 = n13742 ^ n6826 ^ 1'b0 ;
  assign n31228 = n27485 & ~n31227 ;
  assign n31229 = n2256 & ~n31228 ;
  assign n31230 = n31226 & n31229 ;
  assign n31231 = n994 | n12955 ;
  assign n31232 = n9649 & ~n31231 ;
  assign n31235 = n7036 ^ n2559 ^ 1'b0 ;
  assign n31236 = n13119 & ~n31235 ;
  assign n31233 = x15 & n1170 ;
  assign n31234 = n6818 | n31233 ;
  assign n31237 = n31236 ^ n31234 ^ 1'b0 ;
  assign n31238 = n21038 & n28014 ;
  assign n31239 = n20637 | n29256 ;
  assign n31240 = ~n18242 & n30431 ;
  assign n31241 = n31240 ^ n19026 ^ 1'b0 ;
  assign n31242 = n18770 & n22882 ;
  assign n31243 = ~n6166 & n31242 ;
  assign n31244 = n5780 | n6066 ;
  assign n31245 = n20201 ^ n9912 ^ n8103 ;
  assign n31246 = n31245 ^ n14505 ^ 1'b0 ;
  assign n31247 = n3674 ^ n1240 ^ 1'b0 ;
  assign n31248 = ( n1981 & n13630 ) | ( n1981 & n25255 ) | ( n13630 & n25255 ) ;
  assign n31249 = n20631 | n21191 ;
  assign n31250 = n7710 & ~n31249 ;
  assign n31251 = n31250 ^ n28722 ^ n2540 ;
  assign n31252 = n11137 ^ n9200 ^ 1'b0 ;
  assign n31253 = n5081 | n31252 ;
  assign n31254 = ( n10309 & n18390 ) | ( n10309 & n19595 ) | ( n18390 & n19595 ) ;
  assign n31255 = n31254 ^ n16296 ^ 1'b0 ;
  assign n31256 = n31253 | n31255 ;
  assign n31257 = n7848 & ~n15730 ;
  assign n31258 = ~n5132 & n17107 ;
  assign n31259 = ~n22754 & n31258 ;
  assign n31260 = x116 & ~n8328 ;
  assign n31261 = n14818 & ~n19983 ;
  assign n31262 = ( n11799 & n31260 ) | ( n11799 & n31261 ) | ( n31260 & n31261 ) ;
  assign n31263 = n19788 ^ n11544 ^ 1'b0 ;
  assign n31264 = n12513 ^ n12258 ^ 1'b0 ;
  assign n31265 = n10290 | n31264 ;
  assign n31266 = n17091 | n31265 ;
  assign n31267 = n31266 ^ n844 ^ 1'b0 ;
  assign n31268 = n23541 & n31267 ;
  assign n31269 = n9746 ^ n8762 ^ 1'b0 ;
  assign n31270 = ~n7813 & n31269 ;
  assign n31271 = n14567 & n17903 ;
  assign n31272 = n4621 ^ n2471 ^ 1'b0 ;
  assign n31273 = n31271 & ~n31272 ;
  assign n31274 = n11976 | n31273 ;
  assign n31275 = n4370 | n10316 ;
  assign n31276 = n31275 ^ n25152 ^ 1'b0 ;
  assign n31277 = n26481 | n30362 ;
  assign n31278 = ~n13042 & n31277 ;
  assign n31279 = n856 & n31278 ;
  assign n31280 = ( n606 & ~n6963 ) | ( n606 & n18268 ) | ( ~n6963 & n18268 ) ;
  assign n31281 = n462 | n31280 ;
  assign n31282 = n16280 & ~n31281 ;
  assign n31283 = ~n8391 & n31282 ;
  assign n31284 = ~n6354 & n9921 ;
  assign n31285 = n14470 & n31284 ;
  assign n31286 = n27621 | n27806 ;
  assign n31287 = n31285 & ~n31286 ;
  assign n31289 = n18108 ^ n2916 ^ 1'b0 ;
  assign n31290 = n19897 & ~n31289 ;
  assign n31288 = n1428 & ~n3172 ;
  assign n31291 = n31290 ^ n31288 ^ 1'b0 ;
  assign n31292 = n27284 ^ n17442 ^ n14125 ;
  assign n31293 = n24773 ^ n11689 ^ 1'b0 ;
  assign n31294 = n19159 & ~n31293 ;
  assign n31295 = n29208 & n31294 ;
  assign n31296 = n15730 ^ n9432 ^ 1'b0 ;
  assign n31297 = ~n2995 & n31296 ;
  assign n31298 = n13668 ^ n9438 ^ n5450 ;
  assign n31299 = n6522 & n31298 ;
  assign n31300 = n3022 & ~n7675 ;
  assign n31301 = ~n7855 & n13565 ;
  assign n31302 = n23537 ^ n22724 ^ 1'b0 ;
  assign n31303 = n9276 | n19885 ;
  assign n31304 = n4325 ^ n2918 ^ 1'b0 ;
  assign n31305 = n31303 | n31304 ;
  assign n31306 = n3372 | n31305 ;
  assign n31307 = n16104 & n23447 ;
  assign n31308 = n28021 ^ n19819 ^ 1'b0 ;
  assign n31309 = n31308 ^ n16020 ^ 1'b0 ;
  assign n31310 = n16618 | n31309 ;
  assign n31311 = n18938 | n23683 ;
  assign n31312 = n18899 | n31311 ;
  assign n31313 = n2782 | n8555 ;
  assign n31314 = n2231 | n31313 ;
  assign n31315 = n31314 ^ n15214 ^ 1'b0 ;
  assign n31316 = n20494 & n31315 ;
  assign n31317 = n937 & ~n20183 ;
  assign n31318 = ~n15012 & n31317 ;
  assign n31321 = n10682 | n23794 ;
  assign n31322 = n15449 & ~n31321 ;
  assign n31319 = n13701 | n27927 ;
  assign n31320 = n31319 ^ n31083 ^ 1'b0 ;
  assign n31323 = n31322 ^ n31320 ^ 1'b0 ;
  assign n31324 = n19440 & n30023 ;
  assign n31325 = n31324 ^ n8704 ^ 1'b0 ;
  assign n31326 = n20913 | n31325 ;
  assign n31327 = n3564 & n17903 ;
  assign n31328 = n31327 ^ x119 ^ 1'b0 ;
  assign n31329 = n15271 & n31328 ;
  assign n31330 = n16783 ^ n16273 ^ 1'b0 ;
  assign n31331 = n30556 | n31330 ;
  assign n31332 = n7571 & n11574 ;
  assign n31333 = ~n29643 & n31332 ;
  assign n31334 = n19986 & n29853 ;
  assign n31337 = n12612 ^ n2722 ^ 1'b0 ;
  assign n31336 = n13468 ^ n9454 ^ 1'b0 ;
  assign n31335 = n11514 | n13297 ;
  assign n31338 = n31337 ^ n31336 ^ n31335 ;
  assign n31339 = n18674 ^ n18071 ^ 1'b0 ;
  assign n31340 = n26902 & n31339 ;
  assign n31341 = n5406 & ~n12802 ;
  assign n31342 = ~n7183 & n8098 ;
  assign n31343 = n7742 & n31342 ;
  assign n31344 = n31343 ^ x209 ^ 1'b0 ;
  assign n31345 = n19162 | n31344 ;
  assign n31346 = n14158 | n31345 ;
  assign n31347 = n31346 ^ n5413 ^ 1'b0 ;
  assign n31348 = ~n6226 & n19471 ;
  assign n31349 = n31348 ^ n20516 ^ 1'b0 ;
  assign n31350 = n20647 ^ n11684 ^ 1'b0 ;
  assign n31351 = ~n16171 & n18922 ;
  assign n31352 = n10374 ^ n1130 ^ 1'b0 ;
  assign n31353 = n11593 | n31352 ;
  assign n31354 = n31353 ^ n20596 ^ 1'b0 ;
  assign n31355 = ( n6138 & n23184 ) | ( n6138 & ~n29768 ) | ( n23184 & ~n29768 ) ;
  assign n31356 = ~n30738 & n31355 ;
  assign n31357 = n13343 & n19160 ;
  assign n31358 = n31357 ^ n12519 ^ 1'b0 ;
  assign n31359 = ( ~n12740 & n17139 ) | ( ~n12740 & n25603 ) | ( n17139 & n25603 ) ;
  assign n31360 = n22740 | n27995 ;
  assign n31361 = n16327 ^ n9509 ^ 1'b0 ;
  assign n31362 = n22003 | n26447 ;
  assign n31363 = n13523 & ~n31362 ;
  assign n31364 = n8425 ^ n5836 ^ 1'b0 ;
  assign n31365 = n924 & ~n25249 ;
  assign n31366 = n22303 ^ n5195 ^ n4541 ;
  assign n31367 = n20140 ^ n5893 ^ 1'b0 ;
  assign n31368 = n7260 & n7792 ;
  assign n31369 = n16764 & ~n31368 ;
  assign n31370 = n23753 | n31369 ;
  assign n31371 = n8322 | n31370 ;
  assign n31372 = n31371 ^ n2883 ^ 1'b0 ;
  assign n31373 = n9788 & ~n20753 ;
  assign n31374 = n31373 ^ n3904 ^ 1'b0 ;
  assign n31377 = n4821 | n15560 ;
  assign n31378 = n31377 ^ n5648 ^ 1'b0 ;
  assign n31375 = n12854 | n18703 ;
  assign n31376 = n5004 & n31375 ;
  assign n31379 = n31378 ^ n31376 ^ n19889 ;
  assign n31380 = n3957 & n28674 ;
  assign n31381 = ~n4356 & n9779 ;
  assign n31382 = ~n3235 & n31381 ;
  assign n31383 = n7876 & n15027 ;
  assign n31384 = n31382 & n31383 ;
  assign n31385 = n31384 ^ n15010 ^ 1'b0 ;
  assign n31386 = ~n1465 & n19068 ;
  assign n31387 = n31385 & n31386 ;
  assign n31388 = ~n9366 & n24633 ;
  assign n31389 = ( n7632 & n9839 ) | ( n7632 & ~n18933 ) | ( n9839 & ~n18933 ) ;
  assign n31390 = n5076 & n5529 ;
  assign n31391 = n31390 ^ n24921 ^ 1'b0 ;
  assign n31392 = n2209 & n20364 ;
  assign n31393 = n7577 | n17888 ;
  assign n31394 = n31393 ^ n2424 ^ 1'b0 ;
  assign n31395 = n2746 & n19134 ;
  assign n31396 = n31395 ^ n9560 ^ 1'b0 ;
  assign n31397 = n8116 & ~n31396 ;
  assign n31398 = n31394 & n31397 ;
  assign n31399 = n18094 ^ n16042 ^ 1'b0 ;
  assign n31400 = n6571 ^ n705 ^ 1'b0 ;
  assign n31401 = n21347 ^ n2907 ^ 1'b0 ;
  assign n31402 = n12260 | n16178 ;
  assign n31403 = n31298 | n31402 ;
  assign n31404 = x229 | n22783 ;
  assign n31405 = ~n5582 & n29277 ;
  assign n31406 = n31405 ^ n10437 ^ 1'b0 ;
  assign n31407 = ( n12014 & n13075 ) | ( n12014 & n21802 ) | ( n13075 & n21802 ) ;
  assign n31408 = n22305 ^ n10934 ^ 1'b0 ;
  assign n31409 = n31407 & ~n31408 ;
  assign n31410 = n31409 ^ n1321 ^ 1'b0 ;
  assign n31411 = n17458 ^ n12398 ^ n1746 ;
  assign n31412 = n20566 ^ n2230 ^ 1'b0 ;
  assign n31413 = n18631 & ~n28201 ;
  assign n31414 = ~n13668 & n31413 ;
  assign n31415 = ~n3291 & n8807 ;
  assign n31416 = n30283 ^ n4649 ^ 1'b0 ;
  assign n31417 = n21169 ^ n3416 ^ 1'b0 ;
  assign n31418 = n30412 ^ n3973 ^ 1'b0 ;
  assign n31419 = n31418 ^ n6177 ^ n3019 ;
  assign n31420 = ( n12975 & ~n21131 ) | ( n12975 & n31419 ) | ( ~n21131 & n31419 ) ;
  assign n31421 = n11458 & n16967 ;
  assign n31422 = n7361 ^ n4782 ^ 1'b0 ;
  assign n31423 = n7798 & n31422 ;
  assign n31424 = n14758 & n19188 ;
  assign n31425 = n1583 & n31424 ;
  assign n31426 = n31425 ^ n10674 ^ 1'b0 ;
  assign n31427 = n31423 & n31426 ;
  assign n31428 = n6109 | n29128 ;
  assign n31429 = n2622 & ~n21601 ;
  assign n31430 = n31429 ^ n19201 ^ 1'b0 ;
  assign n31431 = ~n908 & n4053 ;
  assign n31432 = n10253 & ~n31431 ;
  assign n31433 = n31432 ^ n13360 ^ 1'b0 ;
  assign n31434 = n14887 ^ n12081 ^ 1'b0 ;
  assign n31435 = n31434 ^ n13221 ^ n970 ;
  assign n31436 = ~n13611 & n24691 ;
  assign n31437 = ( n3382 & n12449 ) | ( n3382 & n25680 ) | ( n12449 & n25680 ) ;
  assign n31438 = n30403 ^ n4387 ^ 1'b0 ;
  assign n31439 = n31437 & ~n31438 ;
  assign n31441 = n8994 | n27744 ;
  assign n31440 = n3744 | n29625 ;
  assign n31442 = n31441 ^ n31440 ^ 1'b0 ;
  assign n31443 = ~n14218 & n15492 ;
  assign n31444 = n1859 | n31443 ;
  assign n31446 = n2120 ^ n1078 ^ 1'b0 ;
  assign n31445 = x159 & n9191 ;
  assign n31447 = n31446 ^ n31445 ^ 1'b0 ;
  assign n31448 = n31447 ^ n29546 ^ 1'b0 ;
  assign n31449 = ~n8347 & n31448 ;
  assign n31450 = n11271 ^ n4844 ^ 1'b0 ;
  assign n31451 = n21467 ^ n19284 ^ 1'b0 ;
  assign n31452 = ~n11043 & n31451 ;
  assign n31453 = n30003 ^ n4557 ^ 1'b0 ;
  assign n31455 = n27639 ^ n2813 ^ 1'b0 ;
  assign n31454 = n9605 | n23055 ;
  assign n31456 = n31455 ^ n31454 ^ 1'b0 ;
  assign n31457 = n2335 ^ n1994 ^ 1'b0 ;
  assign n31458 = n28653 & ~n31457 ;
  assign n31459 = n20148 & n31458 ;
  assign n31460 = n2609 & n31459 ;
  assign n31461 = n15697 ^ n9385 ^ 1'b0 ;
  assign n31462 = n5758 | n31461 ;
  assign n31463 = n18320 | n21766 ;
  assign n31464 = n31463 ^ n13811 ^ 1'b0 ;
  assign n31465 = n453 & n17984 ;
  assign n31466 = ~n2992 & n31465 ;
  assign n31467 = ~n6268 & n31466 ;
  assign n31468 = n31467 ^ n21588 ^ 1'b0 ;
  assign n31469 = x34 & n31468 ;
  assign n31470 = n28956 ^ n11195 ^ 1'b0 ;
  assign n31471 = n16308 & n31470 ;
  assign n31472 = ~n25421 & n31471 ;
  assign n31473 = n13578 ^ n3155 ^ 1'b0 ;
  assign n31474 = n31472 & n31473 ;
  assign n31476 = n28256 ^ n2679 ^ 1'b0 ;
  assign n31478 = n3610 & n16026 ;
  assign n31479 = ~n3850 & n31478 ;
  assign n31477 = n4037 & ~n14844 ;
  assign n31480 = n31479 ^ n31477 ^ n14381 ;
  assign n31481 = n31476 & n31480 ;
  assign n31475 = n1129 & n9509 ;
  assign n31482 = n31481 ^ n31475 ^ 1'b0 ;
  assign n31483 = n10168 ^ n3214 ^ 1'b0 ;
  assign n31484 = ~n6746 & n10401 ;
  assign n31485 = n31484 ^ n11687 ^ 1'b0 ;
  assign n31486 = ~n15363 & n31485 ;
  assign n31487 = n31486 ^ n5598 ^ 1'b0 ;
  assign n31488 = n1606 ^ x167 ^ 1'b0 ;
  assign n31489 = ~n1557 & n22800 ;
  assign n31490 = n10237 ^ n8064 ^ 1'b0 ;
  assign n31491 = n3685 & ~n31490 ;
  assign n31492 = n29665 ^ n6632 ^ 1'b0 ;
  assign n31493 = ~n14010 & n31492 ;
  assign n31494 = n8930 & n14890 ;
  assign n31495 = n31494 ^ n4610 ^ 1'b0 ;
  assign n31496 = n31495 ^ n11794 ^ n11253 ;
  assign n31497 = n18933 & ~n31057 ;
  assign n31498 = ( n3656 & n14703 ) | ( n3656 & ~n17700 ) | ( n14703 & ~n17700 ) ;
  assign n31499 = n31498 ^ n19441 ^ 1'b0 ;
  assign n31500 = n4565 & n31499 ;
  assign n31502 = ~n23653 & n28761 ;
  assign n31501 = n17669 | n27162 ;
  assign n31503 = n31502 ^ n31501 ^ 1'b0 ;
  assign n31504 = n24390 ^ n3742 ^ 1'b0 ;
  assign n31505 = ~n21846 & n31504 ;
  assign n31509 = ( n2815 & ~n12058 ) | ( n2815 & n19437 ) | ( ~n12058 & n19437 ) ;
  assign n31506 = n18314 ^ n5512 ^ 1'b0 ;
  assign n31507 = n5705 | n31506 ;
  assign n31508 = n367 & ~n31507 ;
  assign n31510 = n31509 ^ n31508 ^ 1'b0 ;
  assign n31511 = ( n18110 & n19471 ) | ( n18110 & ~n30230 ) | ( n19471 & ~n30230 ) ;
  assign n31512 = ~n14787 & n18016 ;
  assign n31513 = n21401 ^ x107 ^ 1'b0 ;
  assign n31514 = n8862 ^ n5282 ^ 1'b0 ;
  assign n31515 = n3734 & n7989 ;
  assign n31516 = n1006 & ~n12894 ;
  assign n31517 = ~n3155 & n23508 ;
  assign n31518 = n31517 ^ n7964 ^ 1'b0 ;
  assign n31519 = ~n1114 & n31518 ;
  assign n31520 = n24702 ^ n15973 ^ 1'b0 ;
  assign n31521 = n2903 & n6661 ;
  assign n31522 = n31520 & n31521 ;
  assign n31523 = n15640 ^ n3768 ^ 1'b0 ;
  assign n31524 = n9701 ^ n5031 ^ 1'b0 ;
  assign n31525 = n17483 ^ n2366 ^ 1'b0 ;
  assign n31526 = n31524 & n31525 ;
  assign n31527 = ~n23145 & n31526 ;
  assign n31528 = n31527 ^ n10402 ^ 1'b0 ;
  assign n31529 = n3447 & n5988 ;
  assign n31530 = n31529 ^ n11843 ^ 1'b0 ;
  assign n31531 = ~n9451 & n14816 ;
  assign n31532 = n14669 | n16301 ;
  assign n31533 = n6772 & n16562 ;
  assign n31534 = n31532 & n31533 ;
  assign n31535 = n4307 & n5467 ;
  assign n31536 = n9173 & n15906 ;
  assign n31537 = n18348 ^ n13255 ^ 1'b0 ;
  assign n31538 = n12727 & n31537 ;
  assign n31539 = n16687 & n23800 ;
  assign n31540 = n29207 ^ n14984 ^ 1'b0 ;
  assign n31541 = n4169 ^ n2397 ^ 1'b0 ;
  assign n31542 = n7880 | n15831 ;
  assign n31543 = ~n15491 & n31542 ;
  assign n31544 = n13077 & n28605 ;
  assign n31545 = ~n7510 & n31544 ;
  assign n31546 = n31545 ^ n6979 ^ 1'b0 ;
  assign n31547 = n5511 | n31546 ;
  assign n31548 = n7319 & ~n7672 ;
  assign n31549 = n31548 ^ n15565 ^ 1'b0 ;
  assign n31550 = n571 | n2595 ;
  assign n31551 = n31549 & n31550 ;
  assign n31552 = ~n14466 & n23904 ;
  assign n31553 = n8103 & ~n14578 ;
  assign n31554 = n7187 & n9577 ;
  assign n31555 = ~x106 & n31554 ;
  assign n31556 = ( n1100 & n19416 ) | ( n1100 & n31555 ) | ( n19416 & n31555 ) ;
  assign n31557 = n8770 & ~n16525 ;
  assign n31558 = n17789 ^ n7605 ^ 1'b0 ;
  assign n31559 = ~n9855 & n31558 ;
  assign n31560 = n24263 & ~n31559 ;
  assign n31561 = n6783 & ~n31560 ;
  assign n31562 = n31561 ^ n18750 ^ 1'b0 ;
  assign n31563 = n28856 & ~n31562 ;
  assign n31564 = ~n1135 & n10368 ;
  assign n31565 = n23372 & ~n31564 ;
  assign n31566 = n5890 & n16791 ;
  assign n31567 = n31566 ^ n31116 ^ 1'b0 ;
  assign n31568 = n18756 ^ n4803 ^ 1'b0 ;
  assign n31569 = x163 | n16803 ;
  assign n31570 = n31569 ^ n22490 ^ n5500 ;
  assign n31571 = n10880 & ~n12892 ;
  assign n31572 = n935 & n14968 ;
  assign n31573 = n20314 & n30439 ;
  assign n31574 = n31572 & n31573 ;
  assign n31575 = ~n3757 & n31000 ;
  assign n31578 = n4649 | n19665 ;
  assign n31579 = n3755 | n31578 ;
  assign n31576 = ~n2058 & n3959 ;
  assign n31577 = n31576 ^ n22139 ^ 1'b0 ;
  assign n31580 = n31579 ^ n31577 ^ n27974 ;
  assign n31581 = n9022 & ~n9132 ;
  assign n31582 = n9132 & n31581 ;
  assign n31583 = n31582 ^ n14218 ^ 1'b0 ;
  assign n31587 = n1051 | n17397 ;
  assign n31588 = n17397 & ~n31587 ;
  assign n31584 = n23249 ^ n10976 ^ n8241 ;
  assign n31585 = n17901 & ~n31584 ;
  assign n31586 = n31585 ^ n3210 ^ 1'b0 ;
  assign n31589 = n31588 ^ n31586 ^ 1'b0 ;
  assign n31590 = ( n10068 & ~n31583 ) | ( n10068 & n31589 ) | ( ~n31583 & n31589 ) ;
  assign n31591 = n3861 | n14795 ;
  assign n31592 = n31591 ^ n4803 ^ 1'b0 ;
  assign n31593 = n12764 & n31592 ;
  assign n31594 = ~n4252 & n31593 ;
  assign n31595 = n31594 ^ n26960 ^ 1'b0 ;
  assign n31596 = ~n18658 & n24484 ;
  assign n31597 = n21250 | n29595 ;
  assign n31599 = n364 | n1398 ;
  assign n31600 = n31599 ^ n2098 ^ 1'b0 ;
  assign n31598 = x134 & n10746 ;
  assign n31601 = n31600 ^ n31598 ^ 1'b0 ;
  assign n31602 = n31597 & ~n31601 ;
  assign n31603 = n31602 ^ n18433 ^ n6027 ;
  assign n31604 = n13364 ^ n757 ^ 1'b0 ;
  assign n31605 = n1512 ^ n1245 ^ 1'b0 ;
  assign n31607 = n1103 | n4775 ;
  assign n31608 = n8519 | n8847 ;
  assign n31609 = n31607 & ~n31608 ;
  assign n31606 = n11366 | n11935 ;
  assign n31610 = n31609 ^ n31606 ^ 1'b0 ;
  assign n31611 = n31610 ^ n2651 ^ 1'b0 ;
  assign n31612 = ~n23238 & n31611 ;
  assign n31613 = n2900 | n23381 ;
  assign n31614 = n31613 ^ n6726 ^ 1'b0 ;
  assign n31615 = n2164 & n20389 ;
  assign n31616 = ~x14 & n31615 ;
  assign n31617 = n29700 ^ n12389 ^ 1'b0 ;
  assign n31618 = ~n31616 & n31617 ;
  assign n31619 = n4083 | n14089 ;
  assign n31620 = n31619 ^ n1432 ^ 1'b0 ;
  assign n31621 = ( ~x0 & n4652 ) | ( ~x0 & n31620 ) | ( n4652 & n31620 ) ;
  assign n31622 = n17283 ^ n12943 ^ n12712 ;
  assign n31623 = n6537 ^ n1738 ^ 1'b0 ;
  assign n31624 = n17260 | n31623 ;
  assign n31625 = n4865 & n31025 ;
  assign n31626 = n31625 ^ n28325 ^ 1'b0 ;
  assign n31628 = n23128 ^ n11331 ^ 1'b0 ;
  assign n31627 = n20487 & ~n29033 ;
  assign n31629 = n31628 ^ n31627 ^ 1'b0 ;
  assign n31630 = n30957 ^ n5728 ^ 1'b0 ;
  assign n31631 = n8131 ^ n4076 ^ 1'b0 ;
  assign n31632 = n31630 & n31631 ;
  assign n31633 = ~n16237 & n25326 ;
  assign n31634 = n31633 ^ n13610 ^ 1'b0 ;
  assign n31635 = n7486 & n10845 ;
  assign n31636 = n31356 ^ n1468 ^ 1'b0 ;
  assign n31637 = n1884 | n31636 ;
  assign n31638 = n2889 & ~n8927 ;
  assign n31639 = n24615 & n31638 ;
  assign n31642 = n2785 & ~n21814 ;
  assign n31643 = n31642 ^ n8094 ^ 1'b0 ;
  assign n31640 = n14540 ^ n10941 ^ 1'b0 ;
  assign n31641 = n29425 | n31640 ;
  assign n31644 = n31643 ^ n31641 ^ 1'b0 ;
  assign n31645 = ( n8819 & ~n10878 ) | ( n8819 & n15929 ) | ( ~n10878 & n15929 ) ;
  assign n31646 = ~n16433 & n20972 ;
  assign n31647 = ( n31273 & n31645 ) | ( n31273 & ~n31646 ) | ( n31645 & ~n31646 ) ;
  assign n31648 = n24043 | n31647 ;
  assign n31649 = n4739 ^ n2086 ^ 1'b0 ;
  assign n31650 = n31649 ^ n5101 ^ n2355 ;
  assign n31651 = n1064 & ~n27141 ;
  assign n31652 = n27086 ^ n15015 ^ 1'b0 ;
  assign n31653 = n27727 ^ n23164 ^ 1'b0 ;
  assign n31654 = n9833 & ~n18388 ;
  assign n31655 = n31654 ^ n12782 ^ 1'b0 ;
  assign n31656 = n16404 ^ n13863 ^ 1'b0 ;
  assign n31657 = n22278 & ~n31656 ;
  assign n31658 = n23560 ^ n14297 ^ n7419 ;
  assign n31659 = ~n5210 & n9957 ;
  assign n31660 = n17193 ^ n2439 ^ 1'b0 ;
  assign n31661 = n9850 ^ n6812 ^ 1'b0 ;
  assign n31667 = ~n3134 & n11578 ;
  assign n31668 = n31667 ^ n2602 ^ 1'b0 ;
  assign n31666 = ~n1491 & n6414 ;
  assign n31669 = n31668 ^ n31666 ^ 1'b0 ;
  assign n31664 = n19837 ^ n3904 ^ n320 ;
  assign n31662 = ( ~n5669 & n10180 ) | ( ~n5669 & n14038 ) | ( n10180 & n14038 ) ;
  assign n31663 = n3233 & n31662 ;
  assign n31665 = n31664 ^ n31663 ^ 1'b0 ;
  assign n31670 = n31669 ^ n31665 ^ 1'b0 ;
  assign n31671 = n24831 ^ n14115 ^ 1'b0 ;
  assign n31672 = ~n2477 & n20336 ;
  assign n31673 = n3263 | n10331 ;
  assign n31674 = n13666 & n31673 ;
  assign n31675 = ~n5276 & n31674 ;
  assign n31676 = n7811 | n31675 ;
  assign n31677 = n7109 & ~n31676 ;
  assign n31678 = ~n10689 & n14360 ;
  assign n31679 = n6004 & n31678 ;
  assign n31680 = ~n31677 & n31679 ;
  assign n31681 = ~n13133 & n15779 ;
  assign n31682 = n31681 ^ n24005 ^ 1'b0 ;
  assign n31683 = ( n15713 & ~n19504 ) | ( n15713 & n31682 ) | ( ~n19504 & n31682 ) ;
  assign n31684 = n21488 ^ n1856 ^ 1'b0 ;
  assign n31685 = n11057 & n31684 ;
  assign n31686 = n29750 ^ n2951 ^ n1979 ;
  assign n31687 = n31686 ^ n24840 ^ 1'b0 ;
  assign n31688 = n5811 | n31687 ;
  assign n31689 = n31688 ^ n21538 ^ 1'b0 ;
  assign n31690 = n11029 ^ n3460 ^ 1'b0 ;
  assign n31691 = ~n2020 & n31690 ;
  assign n31692 = ~n15015 & n31691 ;
  assign n31693 = n22044 | n31692 ;
  assign n31694 = n2823 & n6977 ;
  assign n31695 = n31694 ^ n21901 ^ 1'b0 ;
  assign n31696 = n8300 & n14575 ;
  assign n31697 = ( n5496 & n17768 ) | ( n5496 & n19988 ) | ( n17768 & n19988 ) ;
  assign n31699 = n4449 & n8963 ;
  assign n31700 = n7545 & n31699 ;
  assign n31698 = n13839 | n19784 ;
  assign n31701 = n31700 ^ n31698 ^ 1'b0 ;
  assign n31702 = ( ~x137 & n31697 ) | ( ~x137 & n31701 ) | ( n31697 & n31701 ) ;
  assign n31703 = n1707 | n11511 ;
  assign n31704 = n1707 & ~n31703 ;
  assign n31705 = n22632 & ~n31704 ;
  assign n31706 = n13454 ^ x151 ^ 1'b0 ;
  assign n31707 = n2045 & ~n9336 ;
  assign n31708 = n9853 & n31707 ;
  assign n31709 = n19650 ^ n8202 ^ 1'b0 ;
  assign n31710 = n30027 & ~n31709 ;
  assign n31711 = n12553 & n20505 ;
  assign n31712 = n31711 ^ n4512 ^ 1'b0 ;
  assign n31713 = n20566 ^ n12244 ^ 1'b0 ;
  assign n31714 = ~n264 & n2279 ;
  assign n31715 = n22833 & n30146 ;
  assign n31716 = n2172 & n13960 ;
  assign n31717 = n2368 | n4222 ;
  assign n31718 = x222 | n31717 ;
  assign n31719 = n5912 | n31718 ;
  assign n31720 = n11733 & n12040 ;
  assign n31721 = n31720 ^ n3067 ^ 1'b0 ;
  assign n31722 = n9202 & n29307 ;
  assign n31723 = n31721 & n31722 ;
  assign n31724 = n11450 & n11589 ;
  assign n31725 = ~n5101 & n31724 ;
  assign n31726 = n31725 ^ n7170 ^ 1'b0 ;
  assign n31727 = n28673 ^ n18043 ^ n11087 ;
  assign n31728 = n31727 ^ n14288 ^ 1'b0 ;
  assign n31729 = n22955 | n31728 ;
  assign n31730 = n11292 & n11843 ;
  assign n31731 = n3050 | n25208 ;
  assign n31732 = n10506 | n31731 ;
  assign n31733 = n944 ^ n287 ^ 1'b0 ;
  assign n31734 = n9105 & n31733 ;
  assign n31735 = ~n9512 & n31734 ;
  assign n31736 = n4916 ^ n3938 ^ 1'b0 ;
  assign n31737 = ~n3588 & n31736 ;
  assign n31738 = n31735 & ~n31737 ;
  assign n31739 = n31738 ^ n13562 ^ 1'b0 ;
  assign n31742 = n4198 | n6072 ;
  assign n31743 = n31742 ^ n1851 ^ 1'b0 ;
  assign n31740 = n27003 | n27647 ;
  assign n31741 = n31740 ^ n24660 ^ 1'b0 ;
  assign n31744 = n31743 ^ n31741 ^ n11413 ;
  assign n31745 = n19413 ^ n957 ^ 1'b0 ;
  assign n31746 = n8558 & n8978 ;
  assign n31747 = n31746 ^ n5619 ^ 1'b0 ;
  assign n31748 = n12246 & ~n31747 ;
  assign n31749 = n370 | n10694 ;
  assign n31750 = n3216 | n31749 ;
  assign n31751 = n8857 ^ n1400 ^ 1'b0 ;
  assign n31752 = n15662 | n30076 ;
  assign n31753 = n5675 & ~n31752 ;
  assign n31754 = n8165 | n16649 ;
  assign n31755 = n11130 | n31754 ;
  assign n31756 = n31755 ^ n28910 ^ 1'b0 ;
  assign n31757 = n6345 ^ n3686 ^ 1'b0 ;
  assign n31758 = n6421 | n31757 ;
  assign n31761 = n961 & n9829 ;
  assign n31759 = n3799 & n5509 ;
  assign n31760 = n31759 ^ n6333 ^ 1'b0 ;
  assign n31762 = n31761 ^ n31760 ^ 1'b0 ;
  assign n31763 = n9959 & n31762 ;
  assign n31764 = n1238 & n10248 ;
  assign n31765 = ~n21114 & n31764 ;
  assign n31766 = n10404 | n30848 ;
  assign n31767 = n4084 | n26398 ;
  assign n31768 = n31767 ^ n16893 ^ 1'b0 ;
  assign n31769 = ~n1763 & n31768 ;
  assign n31770 = ( n256 & ~n13402 ) | ( n256 & n28199 ) | ( ~n13402 & n28199 ) ;
  assign n31771 = n31770 ^ n26056 ^ 1'b0 ;
  assign n31772 = ( ~n3491 & n19533 ) | ( ~n3491 & n27070 ) | ( n19533 & n27070 ) ;
  assign n31773 = n20191 & ~n31586 ;
  assign n31774 = ~n17763 & n31773 ;
  assign n31775 = ~n5298 & n29502 ;
  assign n31776 = n31775 ^ n21696 ^ 1'b0 ;
  assign n31777 = n13668 ^ n7332 ^ 1'b0 ;
  assign n31778 = n23635 | n31777 ;
  assign n31779 = n25470 | n31778 ;
  assign n31780 = n13586 ^ n10905 ^ 1'b0 ;
  assign n31781 = n8612 & ~n31780 ;
  assign n31782 = n20918 ^ n2282 ^ 1'b0 ;
  assign n31783 = n16348 | n31782 ;
  assign n31784 = n31783 ^ n4548 ^ 1'b0 ;
  assign n31785 = n15955 | n31784 ;
  assign n31786 = n9649 ^ n5700 ^ 1'b0 ;
  assign n31787 = ~n19983 & n31786 ;
  assign n31788 = n26280 ^ n6387 ^ 1'b0 ;
  assign n31789 = n31787 & n31788 ;
  assign n31790 = ( n407 & n5664 ) | ( n407 & ~n31789 ) | ( n5664 & ~n31789 ) ;
  assign n31791 = ~n31785 & n31790 ;
  assign n31792 = n10062 ^ n7482 ^ n6119 ;
  assign n31793 = n25805 ^ n15723 ^ 1'b0 ;
  assign n31794 = n8289 ^ n4739 ^ 1'b0 ;
  assign n31795 = ~n11016 & n31794 ;
  assign n31796 = n3034 ^ n2929 ^ 1'b0 ;
  assign n31797 = n1387 & n31796 ;
  assign n31798 = ~n16471 & n18557 ;
  assign n31799 = ~n31797 & n31798 ;
  assign n31800 = n7154 & n10650 ;
  assign n31801 = n19357 & n31800 ;
  assign n31802 = n17692 & ~n31801 ;
  assign n31803 = n11963 & n31802 ;
  assign n31804 = ~n8219 & n14276 ;
  assign n31805 = n31804 ^ n342 ^ 1'b0 ;
  assign n31806 = n906 & n31805 ;
  assign n31807 = n31806 ^ n6722 ^ 1'b0 ;
  assign n31808 = n31807 ^ n20830 ^ 1'b0 ;
  assign n31809 = n11479 | n12734 ;
  assign n31810 = n5218 | n31809 ;
  assign n31811 = n31810 ^ n17417 ^ 1'b0 ;
  assign n31812 = n24601 ^ n11462 ^ 1'b0 ;
  assign n31813 = ~n2203 & n28005 ;
  assign n31814 = n31813 ^ n23539 ^ n5446 ;
  assign n31815 = n31812 & n31814 ;
  assign n31816 = n15484 ^ n6854 ^ 1'b0 ;
  assign n31817 = n22366 & ~n31816 ;
  assign n31818 = n759 & ~n31817 ;
  assign n31819 = n1541 ^ n984 ^ 1'b0 ;
  assign n31820 = n26570 & ~n31819 ;
  assign n31823 = n5257 & n6741 ;
  assign n31824 = n11170 ^ n5582 ^ 1'b0 ;
  assign n31825 = n31823 & n31824 ;
  assign n31821 = n4128 ^ n1004 ^ 1'b0 ;
  assign n31822 = n1510 & n31821 ;
  assign n31826 = n31825 ^ n31822 ^ 1'b0 ;
  assign n31827 = n2213 & ~n10118 ;
  assign n31828 = n31827 ^ n5565 ^ 1'b0 ;
  assign n31829 = ~x196 & n2622 ;
  assign n31830 = ( n18307 & n31828 ) | ( n18307 & ~n31829 ) | ( n31828 & ~n31829 ) ;
  assign n31831 = n21447 ^ n2424 ^ 1'b0 ;
  assign n31832 = n31831 ^ n18110 ^ n6373 ;
  assign n31833 = n16044 & n28703 ;
  assign n31834 = n31833 ^ n23372 ^ 1'b0 ;
  assign n31835 = n22225 & ~n31834 ;
  assign n31836 = n16709 ^ n16073 ^ n10056 ;
  assign n31839 = n5942 | n15445 ;
  assign n31840 = n5942 & ~n31839 ;
  assign n31841 = n17638 & ~n21890 ;
  assign n31842 = n31840 & n31841 ;
  assign n31837 = n4313 & ~n15946 ;
  assign n31838 = n15946 & n31837 ;
  assign n31843 = n31842 ^ n31838 ^ n7464 ;
  assign n31844 = n31843 ^ n9526 ^ 1'b0 ;
  assign n31845 = ~n31836 & n31844 ;
  assign n31846 = ~n9322 & n31845 ;
  assign n31847 = n31846 ^ n13099 ^ 1'b0 ;
  assign n31848 = n29397 ^ n22339 ^ 1'b0 ;
  assign n31850 = n19496 | n23682 ;
  assign n31849 = ~n9749 & n30619 ;
  assign n31851 = n31850 ^ n31849 ^ 1'b0 ;
  assign n31852 = n22347 ^ n4685 ^ n1772 ;
  assign n31853 = n20688 & ~n25445 ;
  assign n31854 = n31852 & n31853 ;
  assign n31858 = n12940 | n16952 ;
  assign n31855 = n9227 ^ n7054 ^ 1'b0 ;
  assign n31856 = n387 | n31855 ;
  assign n31857 = n31856 ^ n5020 ^ 1'b0 ;
  assign n31859 = n31858 ^ n31857 ^ n24889 ;
  assign n31860 = ~n9260 & n14936 ;
  assign n31861 = ( n7035 & ~n14367 ) | ( n7035 & n15304 ) | ( ~n14367 & n15304 ) ;
  assign n31862 = n31860 | n31861 ;
  assign n31863 = n3966 & n22053 ;
  assign n31864 = n14969 ^ n7222 ^ n2919 ;
  assign n31865 = n31864 ^ n13448 ^ 1'b0 ;
  assign n31866 = ~n15336 & n31865 ;
  assign n31867 = n31866 ^ n18110 ^ 1'b0 ;
  assign n31868 = n1482 | n31867 ;
  assign n31869 = ~n9241 & n18104 ;
  assign n31870 = n31869 ^ n20320 ^ 1'b0 ;
  assign n31871 = n31870 ^ n14312 ^ 1'b0 ;
  assign n31872 = n31871 ^ n22658 ^ 1'b0 ;
  assign n31873 = n24201 | n25057 ;
  assign n31874 = n2593 & ~n31873 ;
  assign n31875 = n23755 ^ n9665 ^ 1'b0 ;
  assign n31876 = n19250 & n31875 ;
  assign n31877 = n11877 & n31876 ;
  assign n31878 = n20903 ^ n799 ^ 1'b0 ;
  assign n31879 = n22193 ^ n7239 ^ 1'b0 ;
  assign n31880 = n14970 ^ n2082 ^ 1'b0 ;
  assign n31881 = n18459 | n31880 ;
  assign n31882 = n25866 ^ n7583 ^ n1835 ;
  assign n31883 = n31882 ^ n23911 ^ 1'b0 ;
  assign n31884 = n2589 & n16898 ;
  assign n31885 = ~n12871 & n31884 ;
  assign n31886 = n26285 | n31885 ;
  assign n31887 = n31886 ^ n3410 ^ 1'b0 ;
  assign n31888 = ~n26046 & n28804 ;
  assign n31889 = n31888 ^ n26654 ^ 1'b0 ;
  assign n31890 = n18747 ^ n16355 ^ 1'b0 ;
  assign n31891 = n21879 & ~n23423 ;
  assign n31892 = n1605 | n31891 ;
  assign n31893 = n31890 & ~n31892 ;
  assign n31894 = ~n4051 & n9476 ;
  assign n31895 = n31894 ^ n1367 ^ 1'b0 ;
  assign n31896 = n13743 | n23859 ;
  assign n31897 = n30440 ^ n25400 ^ n18457 ;
  assign n31898 = n28092 ^ n10280 ^ 1'b0 ;
  assign n31899 = n5038 ^ n619 ^ 1'b0 ;
  assign n31900 = n11071 & n13439 ;
  assign n31901 = ~n606 & n8990 ;
  assign n31902 = ~n9509 & n31901 ;
  assign n31903 = n15135 | n31902 ;
  assign n31904 = n31903 ^ n5931 ^ 1'b0 ;
  assign n31905 = n9048 ^ n6522 ^ 1'b0 ;
  assign n31906 = n3362 & ~n31905 ;
  assign n31907 = n31906 ^ n9365 ^ 1'b0 ;
  assign n31908 = n22758 | n31907 ;
  assign n31909 = n31908 ^ n21831 ^ 1'b0 ;
  assign n31910 = ~n812 & n7693 ;
  assign n31911 = n31910 ^ n20347 ^ 1'b0 ;
  assign n31912 = n31911 ^ n2239 ^ 1'b0 ;
  assign n31913 = n24136 ^ n7871 ^ 1'b0 ;
  assign n31914 = ~n14747 & n31913 ;
  assign n31915 = n5119 | n31914 ;
  assign n31916 = n25543 ^ n3279 ^ 1'b0 ;
  assign n31920 = n23287 ^ n2232 ^ 1'b0 ;
  assign n31917 = n15967 | n25858 ;
  assign n31918 = n26510 | n31917 ;
  assign n31919 = n3190 & n31918 ;
  assign n31921 = n31920 ^ n31919 ^ 1'b0 ;
  assign n31922 = ~n2395 & n4125 ;
  assign n31923 = ~n16869 & n31922 ;
  assign n31924 = n31923 ^ n13518 ^ 1'b0 ;
  assign n31925 = ~n9773 & n31924 ;
  assign n31926 = ( n9479 & ~n31921 ) | ( n9479 & n31925 ) | ( ~n31921 & n31925 ) ;
  assign n31927 = n932 | n9447 ;
  assign n31928 = n31927 ^ n6171 ^ 1'b0 ;
  assign n31929 = n22026 ^ n2370 ^ 1'b0 ;
  assign n31930 = n18361 ^ n8626 ^ 1'b0 ;
  assign n31931 = n3560 & ~n31930 ;
  assign n31933 = n2433 & n7989 ;
  assign n31932 = ~n8517 & n9642 ;
  assign n31934 = n31933 ^ n31932 ^ 1'b0 ;
  assign n31935 = n26171 ^ n21528 ^ n5186 ;
  assign n31945 = n28084 ^ x70 ^ 1'b0 ;
  assign n31946 = n1002 | n31945 ;
  assign n31947 = n4554 & ~n31946 ;
  assign n31938 = n7199 | n9045 ;
  assign n31939 = n31938 ^ n3655 ^ 1'b0 ;
  assign n31937 = n12595 & n26746 ;
  assign n31940 = n31939 ^ n31937 ^ 1'b0 ;
  assign n31936 = n17251 | n24293 ;
  assign n31941 = n31940 ^ n31936 ^ 1'b0 ;
  assign n31942 = n1543 & ~n31941 ;
  assign n31943 = n31942 ^ n10616 ^ 1'b0 ;
  assign n31944 = n26000 & ~n31943 ;
  assign n31948 = n31947 ^ n31944 ^ 1'b0 ;
  assign n31949 = n2228 | n19482 ;
  assign n31950 = n688 & ~n31949 ;
  assign n31951 = n31950 ^ x122 ^ 1'b0 ;
  assign n31952 = n1532 ^ n751 ^ 1'b0 ;
  assign n31953 = n31951 & n31952 ;
  assign n31954 = n3298 & n20449 ;
  assign n31955 = n5442 | n27102 ;
  assign n31956 = n20699 & ~n31955 ;
  assign n31957 = n9451 | n31956 ;
  assign n31958 = n18002 | n20826 ;
  assign n31959 = n26285 ^ n12704 ^ 1'b0 ;
  assign n31960 = n31958 & ~n31959 ;
  assign n31961 = n19974 ^ n13370 ^ 1'b0 ;
  assign n31962 = n9736 & ~n16352 ;
  assign n31963 = n31962 ^ n18182 ^ 1'b0 ;
  assign n31964 = ~n998 & n7061 ;
  assign n31965 = ~x150 & n31964 ;
  assign n31966 = n6173 & ~n31965 ;
  assign n31967 = n31966 ^ n4218 ^ 1'b0 ;
  assign n31968 = n9934 & n31967 ;
  assign n31969 = n10950 ^ x82 ^ 1'b0 ;
  assign n31970 = ~n3210 & n31969 ;
  assign n31971 = n2301 & ~n31970 ;
  assign n31972 = n1943 & ~n8395 ;
  assign n31973 = ~n2550 & n31972 ;
  assign n31974 = ~n3656 & n8974 ;
  assign n31975 = n31973 & n31974 ;
  assign n31976 = n24745 & ~n31975 ;
  assign n31977 = n5076 ^ n2739 ^ 1'b0 ;
  assign n31978 = ~n1048 & n15854 ;
  assign n31979 = n12520 | n17448 ;
  assign n31980 = n2924 & ~n31979 ;
  assign n31981 = n17883 ^ n7600 ^ 1'b0 ;
  assign n31982 = n19022 | n20406 ;
  assign n31983 = n21162 ^ n7111 ^ 1'b0 ;
  assign n31984 = ~n2829 & n31983 ;
  assign n31985 = n31984 ^ n21322 ^ 1'b0 ;
  assign n31986 = n7578 & ~n11121 ;
  assign n31987 = n31986 ^ n708 ^ 1'b0 ;
  assign n31988 = n31987 ^ n20332 ^ n4974 ;
  assign n31989 = n31988 ^ n1094 ^ 1'b0 ;
  assign n31990 = n4793 & n20456 ;
  assign n31991 = ~n786 & n20967 ;
  assign n31992 = n31990 & n31991 ;
  assign n31993 = n28874 ^ n8430 ^ 1'b0 ;
  assign n31994 = n30729 ^ n5404 ^ 1'b0 ;
  assign n31995 = n11333 ^ n6897 ^ 1'b0 ;
  assign n31996 = n7264 & ~n16857 ;
  assign n31997 = ( ~n16019 & n31995 ) | ( ~n16019 & n31996 ) | ( n31995 & n31996 ) ;
  assign n31998 = n14994 | n23683 ;
  assign n31999 = n31998 ^ n1293 ^ 1'b0 ;
  assign n32000 = n6027 ^ n2580 ^ 1'b0 ;
  assign n32001 = n5590 & ~n21812 ;
  assign n32003 = x23 & ~n274 ;
  assign n32002 = n8305 ^ n6236 ^ n3640 ;
  assign n32004 = n32003 ^ n32002 ^ 1'b0 ;
  assign n32005 = ( n7513 & ~n19102 ) | ( n7513 & n23457 ) | ( ~n19102 & n23457 ) ;
  assign n32006 = n296 & ~n12218 ;
  assign n32007 = n24848 ^ n4317 ^ 1'b0 ;
  assign n32008 = ~n2936 & n32007 ;
  assign n32009 = ( n2167 & n16252 ) | ( n2167 & n20821 ) | ( n16252 & n20821 ) ;
  assign n32010 = n287 & n22119 ;
  assign n32011 = n32010 ^ x105 ^ 1'b0 ;
  assign n32012 = n1086 | n14124 ;
  assign n32013 = n15676 & ~n32012 ;
  assign n32014 = n32013 ^ n3435 ^ 1'b0 ;
  assign n32015 = ~n5097 & n7248 ;
  assign n32016 = n12856 & n32015 ;
  assign n32017 = n23091 | n32016 ;
  assign n32018 = n32017 ^ n16264 ^ 1'b0 ;
  assign n32019 = x45 & ~n10387 ;
  assign n32020 = n32019 ^ n9654 ^ 1'b0 ;
  assign n32021 = ~n12516 & n16153 ;
  assign n32022 = n32020 & n32021 ;
  assign n32024 = x17 & ~n3109 ;
  assign n32023 = x45 & ~n21171 ;
  assign n32025 = n32024 ^ n32023 ^ 1'b0 ;
  assign n32026 = n4501 & ~n32025 ;
  assign n32027 = n13689 ^ n4916 ^ 1'b0 ;
  assign n32028 = n11147 & ~n14198 ;
  assign n32029 = n994 | n18346 ;
  assign n32030 = ~n20507 & n32029 ;
  assign n32031 = n6394 ^ n1545 ^ 1'b0 ;
  assign n32032 = n1342 & n32031 ;
  assign n32033 = n2904 ^ n1134 ^ 1'b0 ;
  assign n32034 = ~n7562 & n32033 ;
  assign n32035 = n2369 & n32034 ;
  assign n32036 = n18277 & n32035 ;
  assign n32037 = n7116 & ~n32036 ;
  assign n32038 = ~n14717 & n32037 ;
  assign n32043 = n10152 ^ n3786 ^ 1'b0 ;
  assign n32039 = ~n10711 & n10785 ;
  assign n32040 = ( n11137 & ~n20566 ) | ( n11137 & n32039 ) | ( ~n20566 & n32039 ) ;
  assign n32041 = n32040 ^ n12904 ^ 1'b0 ;
  assign n32042 = n7724 & ~n32041 ;
  assign n32044 = n32043 ^ n32042 ^ 1'b0 ;
  assign n32045 = n3326 & n6765 ;
  assign n32046 = n4254 & n18321 ;
  assign n32047 = n32045 & n32046 ;
  assign n32048 = n3468 & n32047 ;
  assign n32049 = ~n3419 & n23248 ;
  assign n32050 = ~n11147 & n32049 ;
  assign n32051 = n5582 | n32050 ;
  assign n32052 = n20543 | n32051 ;
  assign n32053 = n14590 ^ n9317 ^ n6822 ;
  assign n32054 = n9036 & ~n9821 ;
  assign n32055 = ~n4638 & n32054 ;
  assign n32056 = n32055 ^ n9727 ^ n2062 ;
  assign n32057 = n17081 ^ n1474 ^ 1'b0 ;
  assign n32058 = n9195 ^ n2986 ^ 1'b0 ;
  assign n32059 = ~n27094 & n32058 ;
  assign n32060 = n15818 & ~n25990 ;
  assign n32061 = n19819 & n32060 ;
  assign n32062 = n29033 ^ n5208 ^ 1'b0 ;
  assign n32063 = n32062 ^ n29793 ^ n14732 ;
  assign n32064 = n9529 ^ n2244 ^ 1'b0 ;
  assign n32065 = n8866 | n32064 ;
  assign n32066 = n7986 & ~n25008 ;
  assign n32067 = n32066 ^ n22425 ^ 1'b0 ;
  assign n32068 = n19690 ^ n16403 ^ 1'b0 ;
  assign n32069 = n2301 & n32068 ;
  assign n32070 = ~n6339 & n15709 ;
  assign n32071 = n32070 ^ n23865 ^ 1'b0 ;
  assign n32072 = n27328 ^ n15761 ^ 1'b0 ;
  assign n32073 = n6984 & n32072 ;
  assign n32074 = n15428 | n21590 ;
  assign n32075 = n542 & ~n32074 ;
  assign n32076 = n5282 & n14696 ;
  assign n32077 = n5391 & n26397 ;
  assign n32078 = x63 & ~n5626 ;
  assign n32079 = n10179 ^ n3845 ^ 1'b0 ;
  assign n32080 = n11381 ^ n9890 ^ n4567 ;
  assign n32081 = n1442 ^ n1269 ^ 1'b0 ;
  assign n32082 = ~n15465 & n32081 ;
  assign n32083 = n32082 ^ n18742 ^ 1'b0 ;
  assign n32084 = n4878 | n6957 ;
  assign n32085 = n32084 ^ n7308 ^ 1'b0 ;
  assign n32086 = n4638 & n32085 ;
  assign n32087 = n32086 ^ n13693 ^ 1'b0 ;
  assign n32088 = n12677 & ~n15162 ;
  assign n32089 = n32087 & n32088 ;
  assign n32090 = n1621 & n3312 ;
  assign n32091 = ~n24311 & n32090 ;
  assign n32092 = n13688 ^ n5393 ^ 1'b0 ;
  assign n32093 = n19528 ^ n2736 ^ 1'b0 ;
  assign n32094 = n8976 & n32093 ;
  assign n32095 = n18865 & ~n32094 ;
  assign n32096 = n2954 | n16461 ;
  assign n32097 = n2743 | n32096 ;
  assign n32098 = n10258 ^ n7842 ^ 1'b0 ;
  assign n32099 = ~n24974 & n32098 ;
  assign n32100 = ~n3329 & n32099 ;
  assign n32101 = n22037 | n32100 ;
  assign n32102 = n32101 ^ n1262 ^ 1'b0 ;
  assign n32103 = ~n1387 & n4432 ;
  assign n32104 = n32103 ^ n28671 ^ 1'b0 ;
  assign n32105 = ~n4379 & n5237 ;
  assign n32106 = n32105 ^ n9569 ^ 1'b0 ;
  assign n32107 = n2332 | n32106 ;
  assign n32108 = n32107 ^ n9982 ^ n1439 ;
  assign n32109 = n32108 ^ n14873 ^ 1'b0 ;
  assign n32111 = ~n6083 & n11934 ;
  assign n32110 = n2602 | n6479 ;
  assign n32112 = n32111 ^ n32110 ^ 1'b0 ;
  assign n32113 = n11316 | n12418 ;
  assign n32114 = n32113 ^ n15709 ^ 1'b0 ;
  assign n32115 = ~n26194 & n32114 ;
  assign n32116 = n4420 & ~n13124 ;
  assign n32117 = n32116 ^ n24502 ^ n7066 ;
  assign n32118 = n14440 | n32117 ;
  assign n32119 = n32118 ^ n17836 ^ 1'b0 ;
  assign n32120 = n32115 & ~n32119 ;
  assign n32121 = n10044 ^ n6121 ^ 1'b0 ;
  assign n32122 = n27116 ^ n8523 ^ 1'b0 ;
  assign n32123 = ~n32121 & n32122 ;
  assign n32124 = n11450 ^ n5142 ^ 1'b0 ;
  assign n32125 = n32124 ^ n11605 ^ 1'b0 ;
  assign n32126 = ~n2096 & n32125 ;
  assign n32127 = n15273 & ~n31297 ;
  assign n32128 = n14329 & n32127 ;
  assign n32129 = n10743 & n18477 ;
  assign n32130 = n5322 & n8952 ;
  assign n32131 = ~n5242 & n20181 ;
  assign n32132 = n32131 ^ n20012 ^ 1'b0 ;
  assign n32133 = n32130 & ~n32132 ;
  assign n32134 = n25965 & n27059 ;
  assign n32135 = n32134 ^ n24996 ^ 1'b0 ;
  assign n32136 = n25512 ^ n9745 ^ 1'b0 ;
  assign n32137 = n31025 & ~n32136 ;
  assign n32138 = n2926 & n5934 ;
  assign n32139 = ~n9835 & n9984 ;
  assign n32140 = ~n32138 & n32139 ;
  assign n32141 = n4900 & n5457 ;
  assign n32142 = ( n744 & ~n4240 ) | ( n744 & n32141 ) | ( ~n4240 & n32141 ) ;
  assign n32143 = n32142 ^ n8740 ^ 1'b0 ;
  assign n32144 = n421 & ~n3277 ;
  assign n32145 = n32144 ^ n2269 ^ 1'b0 ;
  assign n32147 = ( n2900 & ~n13283 ) | ( n2900 & n19695 ) | ( ~n13283 & n19695 ) ;
  assign n32146 = n4795 | n29267 ;
  assign n32148 = n32147 ^ n32146 ^ 1'b0 ;
  assign n32149 = ~n32145 & n32148 ;
  assign n32150 = n6022 & n7902 ;
  assign n32151 = n32150 ^ n19819 ^ n19695 ;
  assign n32152 = n8603 & n32151 ;
  assign n32153 = n32152 ^ n15611 ^ 1'b0 ;
  assign n32154 = n11106 ^ n1667 ^ 1'b0 ;
  assign n32155 = n8907 & n26132 ;
  assign n32156 = n32155 ^ n21541 ^ 1'b0 ;
  assign n32157 = ~n32154 & n32156 ;
  assign n32158 = ~n17556 & n20095 ;
  assign n32159 = n5941 & ~n32158 ;
  assign n32160 = n32159 ^ n11191 ^ 1'b0 ;
  assign n32161 = n661 | n4069 ;
  assign n32162 = n2007 | n32161 ;
  assign n32163 = n30207 ^ n4169 ^ 1'b0 ;
  assign n32164 = n32162 & n32163 ;
  assign n32165 = n14597 | n22824 ;
  assign n32166 = n20995 | n27114 ;
  assign n32167 = n26319 | n32166 ;
  assign n32168 = n32167 ^ n22800 ^ n21843 ;
  assign n32169 = n26204 ^ n6224 ^ x2 ;
  assign n32170 = n26908 | n32169 ;
  assign n32171 = n6385 | n32170 ;
  assign n32172 = n32170 & ~n32171 ;
  assign n32173 = ( ~n3419 & n29204 ) | ( ~n3419 & n32172 ) | ( n29204 & n32172 ) ;
  assign n32174 = n9587 ^ n7573 ^ 1'b0 ;
  assign n32175 = ~n835 & n8133 ;
  assign n32176 = n8004 & ~n32175 ;
  assign n32177 = n32174 & n32176 ;
  assign n32178 = n9004 ^ n274 ^ 1'b0 ;
  assign n32179 = n7849 ^ n1506 ^ 1'b0 ;
  assign n32180 = n3290 ^ x32 ^ 1'b0 ;
  assign n32181 = n32180 ^ n26562 ^ n6131 ;
  assign n32183 = ( n10146 & n11512 ) | ( n10146 & ~n23362 ) | ( n11512 & ~n23362 ) ;
  assign n32184 = n9745 ^ n4874 ^ 1'b0 ;
  assign n32185 = ( ~n8915 & n32183 ) | ( ~n8915 & n32184 ) | ( n32183 & n32184 ) ;
  assign n32182 = n4741 & n7101 ;
  assign n32186 = n32185 ^ n32182 ^ n12621 ;
  assign n32187 = n28543 ^ n3150 ^ 1'b0 ;
  assign n32188 = n675 & ~n953 ;
  assign n32189 = ~x226 & n32188 ;
  assign n32190 = n14016 & n17663 ;
  assign n32191 = ~n30166 & n32190 ;
  assign n32192 = n25650 ^ n12754 ^ 1'b0 ;
  assign n32193 = ~n2691 & n25682 ;
  assign n32194 = n1439 & ~n32193 ;
  assign n32195 = n13888 & ~n32194 ;
  assign n32196 = n32195 ^ n6080 ^ 1'b0 ;
  assign n32197 = n18029 ^ n1815 ^ 1'b0 ;
  assign n32198 = n25973 ^ n22719 ^ 1'b0 ;
  assign n32199 = ( n11234 & n17918 ) | ( n11234 & n32198 ) | ( n17918 & n32198 ) ;
  assign n32200 = n4720 ^ n3368 ^ 1'b0 ;
  assign n32201 = x134 & ~n32200 ;
  assign n32202 = n11976 & ~n13607 ;
  assign n32203 = n10684 & ~n32202 ;
  assign n32204 = n9659 & ~n27482 ;
  assign n32205 = n4659 | n25409 ;
  assign n32206 = ( ~n21072 & n23862 ) | ( ~n21072 & n32205 ) | ( n23862 & n32205 ) ;
  assign n32207 = n2736 & ~n4875 ;
  assign n32208 = n4875 & n32207 ;
  assign n32209 = n32208 ^ n5074 ^ 1'b0 ;
  assign n32210 = ~n779 & n19758 ;
  assign n32211 = n27238 & n32210 ;
  assign n32212 = n32209 & ~n32211 ;
  assign n32213 = n21371 ^ n12338 ^ 1'b0 ;
  assign n32214 = n25383 ^ n15821 ^ 1'b0 ;
  assign n32215 = n6619 | n32214 ;
  assign n32216 = n23031 ^ n9294 ^ 1'b0 ;
  assign n32217 = n2887 & ~n32216 ;
  assign n32218 = ~n2745 & n18013 ;
  assign n32219 = ~n9094 & n32218 ;
  assign n32220 = n32219 ^ n1633 ^ 1'b0 ;
  assign n32221 = n742 & ~n8688 ;
  assign n32222 = ~n29565 & n32221 ;
  assign n32223 = ( n6437 & ~n16038 ) | ( n6437 & n32222 ) | ( ~n16038 & n32222 ) ;
  assign n32224 = n16784 | n19788 ;
  assign n32225 = n30192 ^ n7941 ^ 1'b0 ;
  assign n32226 = ( n2199 & ~n16384 ) | ( n2199 & n24816 ) | ( ~n16384 & n24816 ) ;
  assign n32227 = n32226 ^ n15518 ^ 1'b0 ;
  assign n32228 = n518 & ~n32227 ;
  assign n32229 = n25023 & n32228 ;
  assign n32230 = n1878 & n31836 ;
  assign n32231 = n17392 ^ n5461 ^ n1725 ;
  assign n32232 = ~n11862 & n32231 ;
  assign n32233 = ~n24053 & n32232 ;
  assign n32234 = n6681 & n32233 ;
  assign n32235 = n19568 ^ n8815 ^ 1'b0 ;
  assign n32236 = n25827 & ~n32235 ;
  assign n32237 = n6797 & n19368 ;
  assign n32238 = n10092 & n32237 ;
  assign n32239 = ~n6551 & n7187 ;
  assign n32240 = n32239 ^ n11803 ^ 1'b0 ;
  assign n32241 = n16030 ^ n9090 ^ 1'b0 ;
  assign n32242 = n19383 & ~n32241 ;
  assign n32243 = n10030 & ~n29138 ;
  assign n32244 = n11127 & ~n15798 ;
  assign n32245 = n32244 ^ n6582 ^ 1'b0 ;
  assign n32246 = n5836 ^ n5425 ^ 1'b0 ;
  assign n32247 = n497 | n32246 ;
  assign n32248 = n2697 & n9327 ;
  assign n32249 = n6854 & n32248 ;
  assign n32250 = n28802 & n32249 ;
  assign n32251 = x143 & n6200 ;
  assign n32252 = n29390 ^ n1696 ^ 1'b0 ;
  assign n32253 = n32251 | n32252 ;
  assign n32254 = n19271 & n23118 ;
  assign n32255 = n904 & n10041 ;
  assign n32256 = n13268 & n32255 ;
  assign n32257 = ~n23872 & n30464 ;
  assign n32258 = n24139 & ~n32257 ;
  assign n32259 = ~n20905 & n29573 ;
  assign n32260 = n32259 ^ n17126 ^ 1'b0 ;
  assign n32261 = ( n12332 & n13678 ) | ( n12332 & ~n20292 ) | ( n13678 & ~n20292 ) ;
  assign n32262 = ~n4003 & n11669 ;
  assign n32263 = n32262 ^ n4159 ^ 1'b0 ;
  assign n32264 = n32263 ^ n6337 ^ 1'b0 ;
  assign n32265 = n4306 & ~n32264 ;
  assign n32266 = ~n1575 & n5470 ;
  assign n32267 = n32266 ^ n20388 ^ 1'b0 ;
  assign n32268 = n32267 ^ n31830 ^ 1'b0 ;
  assign n32269 = n2889 ^ x14 ^ 1'b0 ;
  assign n32270 = n11377 | n11725 ;
  assign n32271 = n32270 ^ n25359 ^ 1'b0 ;
  assign n32272 = n10608 ^ n5864 ^ 1'b0 ;
  assign n32273 = ~n2325 & n3942 ;
  assign n32274 = n32273 ^ n15042 ^ 1'b0 ;
  assign n32275 = n29445 ^ n16892 ^ 1'b0 ;
  assign n32276 = n20629 & n32275 ;
  assign n32277 = n7704 | n7890 ;
  assign n32278 = n1589 & n6358 ;
  assign n32279 = ~n17051 & n32278 ;
  assign n32280 = n27604 & n32279 ;
  assign n32281 = n13562 ^ n10847 ^ 1'b0 ;
  assign n32282 = ( n4025 & n4261 ) | ( n4025 & n32281 ) | ( n4261 & n32281 ) ;
  assign n32283 = n32282 ^ n15579 ^ n10807 ;
  assign n32284 = n15178 & ~n23152 ;
  assign n32285 = n5815 | n8943 ;
  assign n32286 = n20653 & n32285 ;
  assign n32287 = ~n24440 & n32286 ;
  assign n32288 = n7791 & ~n30545 ;
  assign n32290 = n5385 ^ n5050 ^ 1'b0 ;
  assign n32289 = n6793 | n10290 ;
  assign n32291 = n32290 ^ n32289 ^ 1'b0 ;
  assign n32292 = n1714 | n20389 ;
  assign n32293 = n15795 & n32292 ;
  assign n32294 = n25544 ^ n1048 ^ 1'b0 ;
  assign n32295 = n322 & n32294 ;
  assign n32296 = n23180 ^ n14036 ^ 1'b0 ;
  assign n32298 = n1813 ^ n599 ^ 1'b0 ;
  assign n32299 = n1385 | n32298 ;
  assign n32297 = n5540 & n17763 ;
  assign n32300 = n32299 ^ n32297 ^ 1'b0 ;
  assign n32301 = n32300 ^ n5560 ^ 1'b0 ;
  assign n32302 = n5959 & ~n30525 ;
  assign n32303 = n32302 ^ n320 ^ 1'b0 ;
  assign n32304 = n865 | n4005 ;
  assign n32305 = n32304 ^ n2372 ^ 1'b0 ;
  assign n32306 = n1737 & n9930 ;
  assign n32307 = n7757 | n32306 ;
  assign n32308 = ~n4263 & n25049 ;
  assign n32309 = ~n8499 & n32308 ;
  assign n32310 = n14994 ^ n3726 ^ 1'b0 ;
  assign n32311 = n3432 & ~n32310 ;
  assign n32312 = n9447 | n32311 ;
  assign n32313 = n27663 ^ n19644 ^ 1'b0 ;
  assign n32314 = n18563 | n32313 ;
  assign n32315 = ~n978 & n20375 ;
  assign n32316 = n978 & n32315 ;
  assign n32317 = n15004 ^ n4524 ^ 1'b0 ;
  assign n32318 = n14919 | n32317 ;
  assign n32319 = n3291 & n29846 ;
  assign n32320 = n21944 ^ n4799 ^ n3302 ;
  assign n32321 = n6008 | n31376 ;
  assign n32322 = n32321 ^ n27332 ^ 1'b0 ;
  assign n32323 = ~n6409 & n20845 ;
  assign n32324 = n17707 & n32323 ;
  assign n32325 = ~n4380 & n28856 ;
  assign n32326 = n16506 ^ n5709 ^ 1'b0 ;
  assign n32327 = n4123 & ~n13187 ;
  assign n32328 = n32327 ^ n32111 ^ 1'b0 ;
  assign n32329 = n32328 ^ n23597 ^ n11494 ;
  assign n32330 = n30261 ^ n3210 ^ 1'b0 ;
  assign n32331 = n32330 ^ n25763 ^ 1'b0 ;
  assign n32332 = n21428 | n32331 ;
  assign n32333 = n25104 ^ n4701 ^ 1'b0 ;
  assign n32334 = n6943 & n27480 ;
  assign n32336 = n12280 ^ n305 ^ 1'b0 ;
  assign n32337 = n32336 ^ n18385 ^ 1'b0 ;
  assign n32338 = n4181 ^ n983 ^ 1'b0 ;
  assign n32339 = n32337 & ~n32338 ;
  assign n32335 = ~n851 & n16404 ;
  assign n32340 = n32339 ^ n32335 ^ 1'b0 ;
  assign n32341 = n1977 & ~n2600 ;
  assign n32342 = n2600 & n32341 ;
  assign n32343 = n32342 ^ n6920 ^ 1'b0 ;
  assign n32344 = n3936 & ~n4775 ;
  assign n32345 = n4775 & n32344 ;
  assign n32346 = n1219 | n32345 ;
  assign n32347 = n32343 | n32346 ;
  assign n32348 = ~n3424 & n18933 ;
  assign n32349 = n32348 ^ n12612 ^ 1'b0 ;
  assign n32350 = ( ~n18254 & n32347 ) | ( ~n18254 & n32349 ) | ( n32347 & n32349 ) ;
  assign n32351 = n9699 & ~n13693 ;
  assign n32352 = n32351 ^ n4941 ^ 1'b0 ;
  assign n32353 = n6547 ^ n2542 ^ 1'b0 ;
  assign n32354 = n6812 & ~n32353 ;
  assign n32355 = ~n9448 & n28698 ;
  assign n32356 = n8138 | n15042 ;
  assign n32357 = ~n1489 & n5792 ;
  assign n32358 = n6357 | n32357 ;
  assign n32359 = n27418 ^ n8991 ^ 1'b0 ;
  assign n32360 = n7385 | n25755 ;
  assign n32361 = n14456 & n16923 ;
  assign n32363 = n5075 & ~n17653 ;
  assign n32362 = ( n7799 & ~n13950 ) | ( n7799 & n15056 ) | ( ~n13950 & n15056 ) ;
  assign n32364 = n32363 ^ n32362 ^ 1'b0 ;
  assign n32365 = n2995 | n32364 ;
  assign n32366 = n32365 ^ n6033 ^ 1'b0 ;
  assign n32367 = ~n6112 & n19390 ;
  assign n32368 = n15582 | n20305 ;
  assign n32369 = n32368 ^ n11412 ^ 1'b0 ;
  assign n32371 = n10803 ^ n7873 ^ 1'b0 ;
  assign n32372 = ~n23938 & n32371 ;
  assign n32370 = n9489 & n18549 ;
  assign n32373 = n32372 ^ n32370 ^ 1'b0 ;
  assign n32374 = n27639 ^ n5385 ^ 1'b0 ;
  assign n32375 = n3007 ^ n739 ^ 1'b0 ;
  assign n32376 = n5402 & n6765 ;
  assign n32377 = n32376 ^ n12648 ^ 1'b0 ;
  assign n32378 = n27409 ^ n21479 ^ n16018 ;
  assign n32379 = n23253 | n32378 ;
  assign n32380 = n11976 ^ n3633 ^ n1165 ;
  assign n32381 = ~n888 & n32380 ;
  assign n32382 = n24300 ^ n8882 ^ 1'b0 ;
  assign n32383 = n21050 ^ n16975 ^ 1'b0 ;
  assign n32386 = n22539 & ~n22669 ;
  assign n32387 = n22669 & n32386 ;
  assign n32388 = n32387 ^ n10905 ^ 1'b0 ;
  assign n32389 = n4374 | n32388 ;
  assign n32384 = n3967 ^ n3925 ^ 1'b0 ;
  assign n32385 = ~n2142 & n32384 ;
  assign n32390 = n32389 ^ n32385 ^ 1'b0 ;
  assign n32391 = n28815 ^ n6254 ^ 1'b0 ;
  assign n32392 = n32391 ^ n3172 ^ 1'b0 ;
  assign n32393 = n26992 & ~n32392 ;
  assign n32394 = n14911 | n26841 ;
  assign n32395 = n32394 ^ n4730 ^ 1'b0 ;
  assign n32396 = ( ~n2106 & n26925 ) | ( ~n2106 & n32395 ) | ( n26925 & n32395 ) ;
  assign n32397 = n2165 | n13162 ;
  assign n32398 = n32397 ^ n1738 ^ 1'b0 ;
  assign n32399 = n6734 | n8189 ;
  assign n32400 = n16545 | n32399 ;
  assign n32401 = n27198 & n27945 ;
  assign n32402 = ~n32400 & n32401 ;
  assign n32403 = n11439 & ~n15301 ;
  assign n32404 = n32402 & n32403 ;
  assign n32405 = n22041 ^ n8275 ^ 1'b0 ;
  assign n32406 = n29750 & ~n32405 ;
  assign n32407 = n14760 ^ n4871 ^ 1'b0 ;
  assign n32408 = n32406 & n32407 ;
  assign n32410 = ( n1032 & ~n4611 ) | ( n1032 & n7964 ) | ( ~n4611 & n7964 ) ;
  assign n32409 = n1870 & n14562 ;
  assign n32411 = n32410 ^ n32409 ^ 1'b0 ;
  assign n32412 = n19235 ^ n13761 ^ n8277 ;
  assign n32413 = ~n4753 & n22303 ;
  assign n32414 = n32413 ^ n4060 ^ 1'b0 ;
  assign n32415 = n19369 & n27973 ;
  assign n32416 = ( n3075 & ~n18392 ) | ( n3075 & n28512 ) | ( ~n18392 & n28512 ) ;
  assign n32417 = n11946 ^ n7381 ^ 1'b0 ;
  assign n32418 = n13104 ^ x82 ^ 1'b0 ;
  assign n32419 = n3357 | n32418 ;
  assign n32420 = n12933 ^ n3360 ^ 1'b0 ;
  assign n32421 = ~n19948 & n32420 ;
  assign n32422 = n4192 ^ n3100 ^ 1'b0 ;
  assign n32423 = n32422 ^ n6450 ^ 1'b0 ;
  assign n32424 = n31205 ^ n15264 ^ 1'b0 ;
  assign n32425 = n23983 & ~n31604 ;
  assign n32426 = n32425 ^ n25768 ^ 1'b0 ;
  assign n32427 = n1315 | n32426 ;
  assign n32428 = n24128 ^ n7035 ^ 1'b0 ;
  assign n32431 = n13759 ^ n10596 ^ n6163 ;
  assign n32432 = ~n12709 & n32431 ;
  assign n32433 = n4968 & n32432 ;
  assign n32429 = ~n879 & n12703 ;
  assign n32430 = n32429 ^ n18319 ^ 1'b0 ;
  assign n32434 = n32433 ^ n32430 ^ n12733 ;
  assign n32436 = n4388 | n11628 ;
  assign n32437 = n12789 | n32436 ;
  assign n32435 = n3195 & n16427 ;
  assign n32438 = n32437 ^ n32435 ^ 1'b0 ;
  assign n32439 = n27687 & ~n29236 ;
  assign n32440 = n8943 | n22033 ;
  assign n32441 = n19983 ^ n11253 ^ n6616 ;
  assign n32442 = ~n22480 & n29162 ;
  assign n32443 = n32442 ^ n14988 ^ 1'b0 ;
  assign n32444 = n24173 ^ n9072 ^ 1'b0 ;
  assign n32445 = n15871 ^ n14408 ^ n4637 ;
  assign n32446 = n21318 ^ n3588 ^ 1'b0 ;
  assign n32447 = n11766 & n14376 ;
  assign n32448 = ~n27506 & n28634 ;
  assign n32449 = n1688 & ~n2646 ;
  assign n32450 = n32449 ^ n16428 ^ 1'b0 ;
  assign n32451 = ~n32107 & n32450 ;
  assign n32452 = n32451 ^ n6401 ^ 1'b0 ;
  assign n32453 = n19979 ^ n2582 ^ 1'b0 ;
  assign n32454 = n14272 ^ n13108 ^ 1'b0 ;
  assign n32455 = ~n6274 & n32454 ;
  assign n32456 = n32455 ^ n3437 ^ 1'b0 ;
  assign n32457 = n4733 & n32456 ;
  assign n32458 = n32457 ^ n3868 ^ 1'b0 ;
  assign n32459 = n946 & ~n9380 ;
  assign n32460 = n14652 & n28096 ;
  assign n32461 = n759 | n1556 ;
  assign n32462 = n32461 ^ n6689 ^ n5586 ;
  assign n32463 = n7882 & n32462 ;
  assign n32464 = n29696 & n32463 ;
  assign n32465 = n32464 ^ n9770 ^ 1'b0 ;
  assign n32466 = ~n21364 & n32465 ;
  assign n32467 = n32466 ^ n17902 ^ 1'b0 ;
  assign n32468 = n9353 ^ n8784 ^ 1'b0 ;
  assign n32469 = n2259 & ~n3975 ;
  assign n32470 = n32468 & n32469 ;
  assign n32471 = x208 & n32057 ;
  assign n32472 = n32470 & n32471 ;
  assign n32473 = ~n11751 & n25276 ;
  assign n32474 = n9775 ^ n6437 ^ 1'b0 ;
  assign n32475 = n4426 | n13121 ;
  assign n32476 = n18959 | n32475 ;
  assign n32477 = n1612 & ~n10356 ;
  assign n32478 = ~n19515 & n32477 ;
  assign n32480 = n12226 ^ n8529 ^ 1'b0 ;
  assign n32481 = x46 & n32480 ;
  assign n32479 = ~n12894 & n17545 ;
  assign n32482 = n32481 ^ n32479 ^ 1'b0 ;
  assign n32483 = n13163 | n29736 ;
  assign n32484 = n25174 & ~n32483 ;
  assign n32485 = n3837 & n20407 ;
  assign n32486 = n1130 | n32485 ;
  assign n32487 = n2514 & ~n32486 ;
  assign n32488 = n10609 | n12913 ;
  assign n32489 = n6378 & ~n32488 ;
  assign n32490 = n4045 | n32489 ;
  assign n32491 = ( n25755 & n30136 ) | ( n25755 & ~n32490 ) | ( n30136 & ~n32490 ) ;
  assign n32492 = n17336 ^ n3758 ^ 1'b0 ;
  assign n32493 = n22971 ^ n13305 ^ 1'b0 ;
  assign n32494 = n7702 & n32493 ;
  assign n32495 = ~n13418 & n17444 ;
  assign n32496 = n6749 & n14379 ;
  assign n32497 = n9608 | n27307 ;
  assign n32498 = n7797 | n32497 ;
  assign n32499 = ( n8067 & n32496 ) | ( n8067 & n32498 ) | ( n32496 & n32498 ) ;
  assign n32500 = n32499 ^ n19947 ^ 1'b0 ;
  assign n32501 = n9241 & ~n32500 ;
  assign n32502 = n4083 | n32501 ;
  assign n32504 = n860 | n12508 ;
  assign n32505 = n32504 ^ n15619 ^ 1'b0 ;
  assign n32506 = n25374 & n32505 ;
  assign n32507 = n32506 ^ n2477 ^ 1'b0 ;
  assign n32503 = n5561 & n26844 ;
  assign n32508 = n32507 ^ n32503 ^ 1'b0 ;
  assign n32509 = ~n4042 & n12911 ;
  assign n32510 = ~n9333 & n32509 ;
  assign n32511 = n28101 ^ n8066 ^ 1'b0 ;
  assign n32512 = n18410 | n21926 ;
  assign n32513 = n32511 | n32512 ;
  assign n32514 = n9028 | n13951 ;
  assign n32515 = n26342 & ~n32514 ;
  assign n32516 = n16018 ^ n4004 ^ 1'b0 ;
  assign n32517 = n16303 & ~n32516 ;
  assign n32518 = n9994 | n13741 ;
  assign n32519 = ~n18268 & n27029 ;
  assign n32520 = n32519 ^ n10520 ^ 1'b0 ;
  assign n32521 = ~n10706 & n32520 ;
  assign n32525 = n9502 | n14433 ;
  assign n32526 = n11935 & ~n32525 ;
  assign n32527 = ~n19373 & n32526 ;
  assign n32528 = n32527 ^ n10710 ^ 1'b0 ;
  assign n32522 = n11662 & n23947 ;
  assign n32523 = n32522 ^ n27639 ^ 1'b0 ;
  assign n32524 = n10352 & n32523 ;
  assign n32529 = n32528 ^ n32524 ^ 1'b0 ;
  assign n32530 = n8353 | n27166 ;
  assign n32531 = n32530 ^ n11754 ^ 1'b0 ;
  assign n32532 = n13896 & ~n26391 ;
  assign n32533 = n361 & n27146 ;
  assign n32534 = ~n22467 & n32533 ;
  assign n32535 = n24483 ^ n13809 ^ 1'b0 ;
  assign n32536 = n5639 ^ n2332 ^ 1'b0 ;
  assign n32537 = n32535 | n32536 ;
  assign n32538 = n28204 & ~n32537 ;
  assign n32539 = n26640 ^ n6412 ^ 1'b0 ;
  assign n32540 = n4206 | n9898 ;
  assign n32541 = n31111 & ~n32540 ;
  assign n32542 = ~x102 & n27201 ;
  assign n32543 = n27606 ^ n12361 ^ n3058 ;
  assign n32544 = n363 | n2065 ;
  assign n32545 = n32544 ^ n1554 ^ 1'b0 ;
  assign n32546 = n29852 & ~n32545 ;
  assign n32547 = n2400 | n4404 ;
  assign n32548 = n32547 ^ n1664 ^ 1'b0 ;
  assign n32549 = n32548 ^ n6402 ^ 1'b0 ;
  assign n32550 = n21391 | n32549 ;
  assign n32551 = n2999 & n26699 ;
  assign n32552 = n30298 & ~n32551 ;
  assign n32553 = n32550 & n32552 ;
  assign n32554 = n1925 | n12802 ;
  assign n32555 = n4605 ^ n4198 ^ 1'b0 ;
  assign n32556 = n32554 | n32555 ;
  assign n32557 = n31883 | n32556 ;
  assign n32558 = n6436 ^ n796 ^ 1'b0 ;
  assign n32559 = n29962 ^ n27173 ^ n22523 ;
  assign n32560 = n23974 | n25923 ;
  assign n32561 = n2286 | n13574 ;
  assign n32562 = n32121 & ~n32561 ;
  assign n32563 = ~n4010 & n6061 ;
  assign n32564 = n17911 | n20469 ;
  assign n32565 = n32563 & ~n32564 ;
  assign n32566 = n3906 ^ n3546 ^ 1'b0 ;
  assign n32567 = n25535 ^ n17635 ^ 1'b0 ;
  assign n32570 = n7379 ^ n1878 ^ 1'b0 ;
  assign n32571 = n5101 & n32570 ;
  assign n32568 = n5087 & n26089 ;
  assign n32569 = n11909 & ~n32568 ;
  assign n32572 = n32571 ^ n32569 ^ 1'b0 ;
  assign n32573 = n28777 & n29808 ;
  assign n32574 = n18278 ^ n6357 ^ 1'b0 ;
  assign n32575 = ~n9992 & n32574 ;
  assign n32576 = n32575 ^ n27768 ^ 1'b0 ;
  assign n32577 = n23784 ^ n11148 ^ 1'b0 ;
  assign n32578 = n14392 & ~n32577 ;
  assign n32579 = n21801 ^ n4370 ^ 1'b0 ;
  assign n32580 = n12665 | n32579 ;
  assign n32581 = n4546 & n32580 ;
  assign n32582 = n2170 | n9971 ;
  assign n32583 = n19439 | n25940 ;
  assign n32584 = n3505 | n32583 ;
  assign n32585 = ~n28570 & n32584 ;
  assign n32586 = n32582 | n32585 ;
  assign n32587 = x129 & n11692 ;
  assign n32588 = n32587 ^ n2665 ^ 1'b0 ;
  assign n32589 = n8909 ^ n4508 ^ 1'b0 ;
  assign n32590 = n3127 & n32589 ;
  assign n32591 = ( n12176 & ~n32588 ) | ( n12176 & n32590 ) | ( ~n32588 & n32590 ) ;
  assign n32592 = n32591 ^ n21712 ^ 1'b0 ;
  assign n32593 = n32592 ^ n18490 ^ n12865 ;
  assign n32594 = n21757 ^ n18482 ^ 1'b0 ;
  assign n32595 = n6168 & n8322 ;
  assign n32596 = ~n28872 & n32595 ;
  assign n32597 = n4174 & ~n23516 ;
  assign n32598 = n1552 & n32597 ;
  assign n32599 = n1335 & n7641 ;
  assign n32600 = n32598 & n32599 ;
  assign n32601 = n7016 | n8880 ;
  assign n32602 = n3837 & ~n32601 ;
  assign n32603 = n1981 ^ n922 ^ 1'b0 ;
  assign n32604 = ~n22487 & n32603 ;
  assign n32605 = n632 & ~n1422 ;
  assign n32606 = n11151 & n32605 ;
  assign n32607 = ~n6888 & n16058 ;
  assign n32608 = ~n9191 & n32607 ;
  assign n32609 = n1664 | n14281 ;
  assign n32610 = n32609 ^ x46 ^ 1'b0 ;
  assign n32611 = n9541 & n32610 ;
  assign n32612 = n32611 ^ n6230 ^ 1'b0 ;
  assign n32613 = n4300 & n5292 ;
  assign n32614 = n32613 ^ n2511 ^ 1'b0 ;
  assign n32615 = n32614 ^ n5648 ^ n4066 ;
  assign n32616 = n19491 & ~n21610 ;
  assign n32618 = n5507 & ~n11134 ;
  assign n32617 = n7586 ^ n2414 ^ n608 ;
  assign n32619 = n32618 ^ n32617 ^ 1'b0 ;
  assign n32620 = n21306 ^ n12612 ^ n2325 ;
  assign n32621 = n32620 ^ n15271 ^ 1'b0 ;
  assign n32622 = n27509 & n32621 ;
  assign n32623 = ~n5195 & n5284 ;
  assign n32624 = n32623 ^ n13521 ^ 1'b0 ;
  assign n32625 = n763 & n18597 ;
  assign n32626 = n32625 ^ n836 ^ 1'b0 ;
  assign n32627 = n32624 & n32626 ;
  assign n32628 = n3679 | n9458 ;
  assign n32629 = n1694 | n2215 ;
  assign n32630 = x157 | n32629 ;
  assign n32631 = n13275 & n17093 ;
  assign n32632 = n27794 & n32631 ;
  assign n32633 = n6272 | n16928 ;
  assign n32634 = n8950 & ~n13435 ;
  assign n32635 = n5664 & n9204 ;
  assign n32636 = ~n5664 & n32635 ;
  assign n32637 = n6751 & ~n32636 ;
  assign n32638 = ~n6751 & n32637 ;
  assign n32639 = n32638 ^ n21050 ^ n3070 ;
  assign n32640 = n32639 ^ n30344 ^ n7066 ;
  assign n32641 = n24132 ^ n11936 ^ 1'b0 ;
  assign n32642 = n2255 | n32641 ;
  assign n32643 = n7478 & ~n22921 ;
  assign n32644 = n32643 ^ n19050 ^ 1'b0 ;
  assign n32645 = n1322 & ~n13812 ;
  assign n32646 = n32645 ^ n12242 ^ 1'b0 ;
  assign n32647 = n6608 | n32646 ;
  assign n32648 = n13127 ^ n8485 ^ 1'b0 ;
  assign n32649 = n7677 & n32648 ;
  assign n32650 = n32649 ^ n1647 ^ 1'b0 ;
  assign n32651 = ( n4621 & ~n10134 ) | ( n4621 & n24172 ) | ( ~n10134 & n24172 ) ;
  assign n32652 = n22060 & n32651 ;
  assign n32653 = n2585 & n32652 ;
  assign n32654 = n4260 & n15555 ;
  assign n32655 = ~n14978 & n32654 ;
  assign n32656 = n32655 ^ n20406 ^ 1'b0 ;
  assign n32657 = n5802 & ~n17494 ;
  assign n32658 = n13953 & n23003 ;
  assign n32659 = n14117 ^ n6654 ^ 1'b0 ;
  assign n32660 = n18597 & ~n32659 ;
  assign n32661 = n30766 ^ n17122 ^ 1'b0 ;
  assign n32662 = ( n11469 & n13993 ) | ( n11469 & ~n32661 ) | ( n13993 & ~n32661 ) ;
  assign n32663 = n32660 | n32662 ;
  assign n32664 = n5429 | n31693 ;
  assign n32665 = ~n1067 & n9072 ;
  assign n32666 = n1508 & ~n20818 ;
  assign n32668 = n5690 & n9262 ;
  assign n32667 = n763 & ~n6236 ;
  assign n32669 = n32668 ^ n32667 ^ 1'b0 ;
  assign n32670 = n7405 ^ n5630 ^ 1'b0 ;
  assign n32671 = ~n14497 & n32670 ;
  assign n32672 = n32669 & n32671 ;
  assign n32673 = ~n2719 & n4562 ;
  assign n32674 = ~n32672 & n32673 ;
  assign n32675 = n2699 & n4589 ;
  assign n32676 = n8844 & n32675 ;
  assign n32677 = n12815 | n18533 ;
  assign n32678 = n32677 ^ n3486 ^ 1'b0 ;
  assign n32679 = n32678 ^ n1929 ^ 1'b0 ;
  assign n32680 = n30648 ^ n7161 ^ 1'b0 ;
  assign n32681 = ~n5600 & n32680 ;
  assign n32682 = n5245 | n25402 ;
  assign n32683 = ~n24214 & n32682 ;
  assign n32684 = n32683 ^ n24749 ^ 1'b0 ;
  assign n32685 = x169 & ~n4921 ;
  assign n32686 = ~n5948 & n32685 ;
  assign n32687 = ~n9977 & n31236 ;
  assign n32688 = n32686 & n32687 ;
  assign n32689 = n12953 ^ n3754 ^ 1'b0 ;
  assign n32690 = ~n4905 & n32689 ;
  assign n32691 = n26727 | n31957 ;
  assign n32692 = n32691 ^ n16225 ^ 1'b0 ;
  assign n32693 = n8744 | n11394 ;
  assign n32694 = n23264 ^ n2304 ^ 1'b0 ;
  assign n32695 = n25499 | n32694 ;
  assign n32696 = n21222 ^ n4303 ^ 1'b0 ;
  assign n32697 = n18568 ^ n2041 ^ 1'b0 ;
  assign n32698 = n25002 | n32697 ;
  assign n32699 = n13034 ^ n6097 ^ 1'b0 ;
  assign n32700 = n6920 & ~n32699 ;
  assign n32701 = n32700 ^ n7159 ^ 1'b0 ;
  assign n32702 = ~n31943 & n32701 ;
  assign n32703 = n19744 & n26810 ;
  assign n32704 = n21712 ^ n2015 ^ 1'b0 ;
  assign n32705 = n1346 & n32704 ;
  assign n32706 = ( ~n24070 & n32703 ) | ( ~n24070 & n32705 ) | ( n32703 & n32705 ) ;
  assign n32707 = ~n10746 & n26877 ;
  assign n32708 = n32707 ^ n9037 ^ 1'b0 ;
  assign n32709 = n3529 ^ n1347 ^ 1'b0 ;
  assign n32710 = ~n5025 & n32709 ;
  assign n32711 = n10803 | n16533 ;
  assign n32712 = n20579 & ~n32711 ;
  assign n32713 = x167 & n11435 ;
  assign n32714 = ~n11435 & n32713 ;
  assign n32715 = n3417 & ~n32714 ;
  assign n32716 = n32714 & n32715 ;
  assign n32719 = n12122 & n23678 ;
  assign n32717 = ( n1183 & n4472 ) | ( n1183 & ~n18019 ) | ( n4472 & ~n18019 ) ;
  assign n32718 = n18830 & n32717 ;
  assign n32720 = n32719 ^ n32718 ^ 1'b0 ;
  assign n32721 = n26504 ^ n12638 ^ 1'b0 ;
  assign n32722 = n17272 ^ n14730 ^ n11297 ;
  assign n32723 = n26498 ^ n25729 ^ 1'b0 ;
  assign n32724 = n10165 & ~n32723 ;
  assign n32725 = n19336 ^ n8763 ^ 1'b0 ;
  assign n32726 = n7871 ^ n7638 ^ 1'b0 ;
  assign n32727 = n14000 | n32726 ;
  assign n32728 = n32727 ^ n14619 ^ 1'b0 ;
  assign n32729 = n6254 & n32728 ;
  assign n32730 = ( n9720 & n12504 ) | ( n9720 & n32729 ) | ( n12504 & n32729 ) ;
  assign n32731 = n20358 | n32730 ;
  assign n32732 = n10149 ^ n759 ^ 1'b0 ;
  assign n32733 = n5437 ^ n1049 ^ 1'b0 ;
  assign n32734 = n32733 ^ n400 ^ 1'b0 ;
  assign n32735 = ~n32732 & n32734 ;
  assign n32736 = n2622 & ~n2819 ;
  assign n32737 = n13892 & n14666 ;
  assign n32738 = ~n978 & n1447 ;
  assign n32739 = n8302 & ~n32738 ;
  assign n32740 = n32739 ^ n20665 ^ 1'b0 ;
  assign n32741 = n12487 & n19299 ;
  assign n32742 = n32741 ^ n8816 ^ 1'b0 ;
  assign n32743 = n1503 & ~n5368 ;
  assign n32744 = n15852 ^ n5659 ^ 1'b0 ;
  assign n32745 = n30157 ^ n14869 ^ 1'b0 ;
  assign n32746 = n32744 | n32745 ;
  assign n32747 = n28481 ^ n2113 ^ 1'b0 ;
  assign n32748 = n20589 | n32747 ;
  assign n32751 = n1379 & n7187 ;
  assign n32749 = n17765 | n21999 ;
  assign n32750 = n32749 ^ n13387 ^ 1'b0 ;
  assign n32752 = n32751 ^ n32750 ^ 1'b0 ;
  assign n32753 = n9024 ^ n8034 ^ 1'b0 ;
  assign n32754 = n32753 ^ n21701 ^ 1'b0 ;
  assign n32755 = n12052 | n24810 ;
  assign n32756 = n4333 & n23613 ;
  assign n32757 = ( ~n2756 & n6753 ) | ( ~n2756 & n9638 ) | ( n6753 & n9638 ) ;
  assign n32758 = ~n13952 & n32757 ;
  assign n32759 = n32758 ^ n12303 ^ 1'b0 ;
  assign n32760 = n20470 ^ n17238 ^ 1'b0 ;
  assign n32761 = n32759 & n32760 ;
  assign n32762 = n17960 ^ n13162 ^ n9470 ;
  assign n32763 = ( n10191 & n19534 ) | ( n10191 & n32762 ) | ( n19534 & n32762 ) ;
  assign n32764 = ( n6655 & ~n8659 ) | ( n6655 & n17273 ) | ( ~n8659 & n17273 ) ;
  assign n32765 = n20817 ^ n5675 ^ 1'b0 ;
  assign n32766 = n1534 & ~n32765 ;
  assign n32767 = ~n12138 & n14141 ;
  assign n32768 = ~x105 & n32767 ;
  assign n32769 = n4315 & ~n32768 ;
  assign n32770 = n7196 & ~n9196 ;
  assign n32771 = ~n12033 & n32770 ;
  assign n32772 = n25650 ^ n1909 ^ 1'b0 ;
  assign n32773 = n12381 ^ n3246 ^ 1'b0 ;
  assign n32774 = ~n9004 & n32773 ;
  assign n32775 = n3679 & ~n4953 ;
  assign n32776 = ~n12861 & n32775 ;
  assign n32777 = ( n992 & n32774 ) | ( n992 & ~n32776 ) | ( n32774 & ~n32776 ) ;
  assign n32778 = ~n1014 & n4279 ;
  assign n32779 = n16307 & n17631 ;
  assign n32780 = n1874 & n32779 ;
  assign n32781 = n30865 & ~n32780 ;
  assign n32782 = ~n32778 & n32781 ;
  assign n32783 = n26876 & ~n32782 ;
  assign n32785 = n22343 ^ n8098 ^ 1'b0 ;
  assign n32786 = ~n31303 & n32785 ;
  assign n32784 = n5150 & ~n5909 ;
  assign n32787 = n32786 ^ n32784 ^ x119 ;
  assign n32790 = n23205 ^ n14470 ^ 1'b0 ;
  assign n32791 = n20915 | n32790 ;
  assign n32788 = ( n1844 & ~n4610 ) | ( n1844 & n7200 ) | ( ~n4610 & n7200 ) ;
  assign n32789 = n5308 | n32788 ;
  assign n32792 = n32791 ^ n32789 ^ 1'b0 ;
  assign n32793 = ~n1879 & n15648 ;
  assign n32794 = n17543 | n30631 ;
  assign n32795 = n9100 & ~n20284 ;
  assign n32796 = n7948 | n32795 ;
  assign n32797 = n32796 ^ n14532 ^ 1'b0 ;
  assign n32798 = n986 & n14335 ;
  assign n32799 = n28168 & n32798 ;
  assign n32803 = n19953 ^ n8260 ^ 1'b0 ;
  assign n32804 = x236 & ~n32803 ;
  assign n32805 = n14730 & n32804 ;
  assign n32800 = n8606 & n14304 ;
  assign n32801 = n12655 & ~n32800 ;
  assign n32802 = n11617 & n32801 ;
  assign n32806 = n32805 ^ n32802 ^ 1'b0 ;
  assign n32807 = ~n649 & n8224 ;
  assign n32808 = n268 & n10079 ;
  assign n32809 = n32807 & ~n32808 ;
  assign n32810 = ~n3249 & n8659 ;
  assign n32811 = n32810 ^ n3348 ^ 1'b0 ;
  assign n32812 = n4090 & n11570 ;
  assign n32813 = ~n9857 & n32812 ;
  assign n32814 = n11840 & ~n32813 ;
  assign n32815 = n5364 & n29099 ;
  assign n32816 = ~n14930 & n32815 ;
  assign n32817 = ~n26272 & n27811 ;
  assign n32818 = ~n14677 & n17573 ;
  assign n32819 = ~n12892 & n32818 ;
  assign n32820 = ~n6357 & n12064 ;
  assign n32821 = n32820 ^ n3640 ^ 1'b0 ;
  assign n32822 = n12807 | n19211 ;
  assign n32823 = n30242 & ~n32822 ;
  assign n32824 = ( n32819 & ~n32821 ) | ( n32819 & n32823 ) | ( ~n32821 & n32823 ) ;
  assign n32825 = n21007 ^ n11040 ^ 1'b0 ;
  assign n32826 = ~n32824 & n32825 ;
  assign n32827 = n5014 | n23163 ;
  assign n32828 = n3423 & ~n24715 ;
  assign n32829 = n14514 & n32828 ;
  assign n32830 = n32829 ^ n27150 ^ n1982 ;
  assign n32833 = n19524 & n25327 ;
  assign n32831 = n7731 & n19817 ;
  assign n32832 = n32831 ^ n18397 ^ 1'b0 ;
  assign n32834 = n32833 ^ n32832 ^ 1'b0 ;
  assign n32835 = n31367 ^ n2544 ^ 1'b0 ;
  assign n32836 = n32834 & n32835 ;
  assign n32837 = n19030 & n26824 ;
  assign n32838 = n21521 ^ n10179 ^ 1'b0 ;
  assign n32839 = ~n9438 & n13888 ;
  assign n32840 = ~n23410 & n32839 ;
  assign n32841 = x249 & ~n14259 ;
  assign n32842 = ~n1371 & n7596 ;
  assign n32843 = n10317 | n14522 ;
  assign n32844 = x192 & n10776 ;
  assign n32845 = x129 & ~n23400 ;
  assign n32846 = n15571 & n32845 ;
  assign n32847 = n32846 ^ n31622 ^ 1'b0 ;
  assign n32850 = n12720 ^ n3055 ^ n585 ;
  assign n32848 = n1635 & n24192 ;
  assign n32849 = n32848 ^ n17877 ^ 1'b0 ;
  assign n32851 = n32850 ^ n32849 ^ n13664 ;
  assign n32852 = n13934 ^ n11196 ^ 1'b0 ;
  assign n32853 = n1784 & n32852 ;
  assign n32854 = ~n7061 & n32853 ;
  assign n32855 = n32854 ^ n6619 ^ n5208 ;
  assign n32857 = n25724 ^ n4964 ^ 1'b0 ;
  assign n32856 = n1004 & ~n21391 ;
  assign n32858 = n32857 ^ n32856 ^ 1'b0 ;
  assign n32859 = n21629 & n32858 ;
  assign n32860 = n11473 & ~n18848 ;
  assign n32861 = n13976 ^ n10407 ^ 1'b0 ;
  assign n32862 = n8277 & ~n32861 ;
  assign n32863 = ~n4244 & n32862 ;
  assign n32864 = n28745 & n32863 ;
  assign n32865 = n19492 & n26074 ;
  assign n32866 = n6646 ^ n1482 ^ 1'b0 ;
  assign n32867 = n16243 & ~n32866 ;
  assign n32868 = n12262 | n32867 ;
  assign n32869 = n13781 & ~n27355 ;
  assign n32870 = n419 & n32869 ;
  assign n32871 = n32870 ^ n12245 ^ 1'b0 ;
  assign n32872 = ~n32868 & n32871 ;
  assign n32873 = n20630 ^ n16989 ^ 1'b0 ;
  assign n32874 = n12473 & ~n32873 ;
  assign n32875 = n1931 & n18725 ;
  assign n32876 = ~n32874 & n32875 ;
  assign n32877 = n14598 & n16120 ;
  assign n32878 = n32877 ^ n17646 ^ 1'b0 ;
  assign n32879 = ( ~n12982 & n17895 ) | ( ~n12982 & n32878 ) | ( n17895 & n32878 ) ;
  assign n32880 = n1335 & ~n32879 ;
  assign n32881 = n32880 ^ n4128 ^ 1'b0 ;
  assign n32882 = n7579 & ~n29949 ;
  assign n32883 = n22732 ^ n13531 ^ n2128 ;
  assign n32884 = n32883 ^ n14800 ^ 1'b0 ;
  assign n32885 = n15290 ^ n1656 ^ 1'b0 ;
  assign n32886 = n32884 & n32885 ;
  assign n32887 = ~n1864 & n16893 ;
  assign n32888 = n15912 & n32887 ;
  assign n32889 = n13670 ^ n13496 ^ 1'b0 ;
  assign n32890 = n25593 | n32889 ;
  assign n32891 = n12044 & n24809 ;
  assign n32892 = n8114 | n15347 ;
  assign n32893 = ~n22044 & n28807 ;
  assign n32894 = n32893 ^ n19006 ^ 1'b0 ;
  assign n32895 = n13419 | n31870 ;
  assign n32896 = n29396 & ~n32895 ;
  assign n32899 = n7096 & ~n7467 ;
  assign n32897 = n9053 | n9206 ;
  assign n32898 = n4442 & ~n32897 ;
  assign n32900 = n32899 ^ n32898 ^ 1'b0 ;
  assign n32901 = ~n8951 & n17406 ;
  assign n32902 = n32901 ^ n17858 ^ 1'b0 ;
  assign n32903 = n8572 ^ n4108 ^ 1'b0 ;
  assign n32904 = n16431 | n32903 ;
  assign n32905 = n32904 ^ n18633 ^ 1'b0 ;
  assign n32906 = x57 & n5121 ;
  assign n32907 = ~n11969 & n18450 ;
  assign n32908 = ~n19491 & n32907 ;
  assign n32909 = n32908 ^ n5728 ^ 1'b0 ;
  assign n32910 = n1138 & n32909 ;
  assign n32911 = n2400 & n8087 ;
  assign n32912 = n6182 & n32911 ;
  assign n32913 = n10295 & n17518 ;
  assign n32914 = n32913 ^ n689 ^ 1'b0 ;
  assign n32915 = n3305 & ~n32914 ;
  assign n32916 = ~n23113 & n32915 ;
  assign n32917 = n2772 & ~n32916 ;
  assign n32918 = n17433 ^ n3258 ^ 1'b0 ;
  assign n32919 = ~n8907 & n9955 ;
  assign n32920 = ~n2267 & n32919 ;
  assign n32921 = n6891 & ~n7117 ;
  assign n32922 = n5095 & ~n32921 ;
  assign n32923 = n7458 & ~n7542 ;
  assign n32924 = n7240 & n32923 ;
  assign n32925 = n20083 & ~n32924 ;
  assign n32926 = n32925 ^ n676 ^ 1'b0 ;
  assign n32927 = ~n4033 & n32028 ;
  assign n32928 = n23383 ^ n22170 ^ 1'b0 ;
  assign n32929 = n32927 | n32928 ;
  assign n32930 = n9083 & ~n12080 ;
  assign n32931 = n14533 | n21461 ;
  assign n32932 = n32931 ^ n13313 ^ 1'b0 ;
  assign n32933 = ~n4542 & n9110 ;
  assign n32934 = n15783 ^ n1508 ^ 1'b0 ;
  assign n32935 = n32933 & ~n32934 ;
  assign n32936 = n30205 & ~n32935 ;
  assign n32937 = n27372 ^ n4637 ^ n2163 ;
  assign n32938 = n17847 ^ n11114 ^ n9436 ;
  assign n32939 = n431 & ~n1775 ;
  assign n32940 = n32939 ^ n842 ^ 1'b0 ;
  assign n32941 = n32940 ^ n4766 ^ 1'b0 ;
  assign n32942 = x129 & ~n32941 ;
  assign n32943 = n22975 ^ n5482 ^ 1'b0 ;
  assign n32944 = n507 | n32943 ;
  assign n32945 = n6337 ^ n4241 ^ 1'b0 ;
  assign n32946 = n6062 | n32945 ;
  assign n32947 = n7914 | n32946 ;
  assign n32948 = n22625 ^ n1264 ^ 1'b0 ;
  assign n32949 = n6781 | n20291 ;
  assign n32950 = n24371 ^ n3419 ^ 1'b0 ;
  assign n32951 = n25344 ^ n14727 ^ 1'b0 ;
  assign n32953 = n1014 | n19783 ;
  assign n32954 = n25399 & ~n32953 ;
  assign n32952 = n14556 ^ n2466 ^ 1'b0 ;
  assign n32955 = n32954 ^ n32952 ^ 1'b0 ;
  assign n32956 = n11950 & n32955 ;
  assign n32957 = n32956 ^ n18759 ^ 1'b0 ;
  assign n32958 = n10144 ^ n8143 ^ 1'b0 ;
  assign n32959 = n20994 ^ n5009 ^ 1'b0 ;
  assign n32960 = n10529 & ~n27234 ;
  assign n32961 = ~n6233 & n32960 ;
  assign n32962 = ~n1824 & n30160 ;
  assign n32963 = n27327 & n32962 ;
  assign n32964 = n2801 ^ n2464 ^ 1'b0 ;
  assign n32965 = n29146 | n32964 ;
  assign n32966 = n17417 & n27891 ;
  assign n32967 = n1185 & n32966 ;
  assign n32968 = n3692 | n32967 ;
  assign n32969 = n9167 | n19037 ;
  assign n32970 = n32969 ^ n5118 ^ 1'b0 ;
  assign n32971 = n17458 | n32970 ;
  assign n32973 = n11392 ^ n5980 ^ 1'b0 ;
  assign n32974 = n11167 & n32973 ;
  assign n32975 = ( n3920 & ~n3966 ) | ( n3920 & n32974 ) | ( ~n3966 & n32974 ) ;
  assign n32972 = ~n4117 & n32285 ;
  assign n32976 = n32975 ^ n32972 ^ 1'b0 ;
  assign n32977 = n8369 | n12335 ;
  assign n32978 = n32977 ^ n3050 ^ 1'b0 ;
  assign n32979 = n18700 ^ n2663 ^ 1'b0 ;
  assign n32980 = n6349 & ~n9216 ;
  assign n32981 = n10217 ^ n5685 ^ 1'b0 ;
  assign n32982 = n32980 & ~n32981 ;
  assign n32983 = n32982 ^ n5816 ^ 1'b0 ;
  assign n32984 = n18288 | n32983 ;
  assign n32985 = ~n12593 & n14859 ;
  assign n32986 = n24324 ^ n6376 ^ n4207 ;
  assign n32987 = ~n6389 & n16701 ;
  assign n32988 = n15338 & n32987 ;
  assign n32989 = n13315 | n32988 ;
  assign n32990 = n32989 ^ n6270 ^ 1'b0 ;
  assign n32991 = n25659 ^ n2477 ^ 1'b0 ;
  assign n32992 = n32991 ^ n16196 ^ 1'b0 ;
  assign n32993 = n32990 | n32992 ;
  assign n32994 = n32993 ^ n2675 ^ 1'b0 ;
  assign n32995 = n2268 & ~n15904 ;
  assign n32996 = ~n2611 & n5767 ;
  assign n32997 = n32996 ^ n21340 ^ 1'b0 ;
  assign n32998 = n32422 | n32997 ;
  assign n32999 = n10529 ^ n1353 ^ 1'b0 ;
  assign n33000 = n29255 & n32999 ;
  assign n33001 = n33000 ^ n10182 ^ 1'b0 ;
  assign n33002 = ~n3498 & n8280 ;
  assign n33003 = n4852 & n33002 ;
  assign n33004 = n7716 & n33003 ;
  assign n33005 = n6684 | n12066 ;
  assign n33006 = n8129 ^ n7768 ^ 1'b0 ;
  assign n33007 = n24851 ^ n1424 ^ 1'b0 ;
  assign n33008 = n33006 | n33007 ;
  assign n33009 = n33008 ^ n3749 ^ 1'b0 ;
  assign n33010 = ~n33005 & n33009 ;
  assign n33011 = n33010 ^ n17609 ^ 1'b0 ;
  assign n33012 = n16788 & n33011 ;
  assign n33013 = n28006 ^ n16612 ^ 1'b0 ;
  assign n33014 = ( n9218 & n33012 ) | ( n9218 & ~n33013 ) | ( n33012 & ~n33013 ) ;
  assign n33015 = n2685 & ~n33014 ;
  assign n33016 = n33015 ^ n16686 ^ 1'b0 ;
  assign n33017 = ( n14653 & n15471 ) | ( n14653 & ~n19333 ) | ( n15471 & ~n19333 ) ;
  assign n33018 = n4551 ^ n1298 ^ 1'b0 ;
  assign n33019 = n20399 ^ n16481 ^ n6600 ;
  assign n33020 = ( n19781 & n33018 ) | ( n19781 & ~n33019 ) | ( n33018 & ~n33019 ) ;
  assign n33021 = n8399 ^ n6271 ^ 1'b0 ;
  assign n33022 = n33020 & ~n33021 ;
  assign n33023 = n7229 | n12588 ;
  assign n33024 = n33023 ^ n5812 ^ 1'b0 ;
  assign n33025 = n21622 & n33024 ;
  assign n33026 = n4275 & n33025 ;
  assign n33027 = n14035 ^ n3985 ^ 1'b0 ;
  assign n33028 = n33027 ^ n5022 ^ 1'b0 ;
  assign n33029 = n3704 & ~n31889 ;
  assign n33030 = x130 | n2202 ;
  assign n33031 = n5847 | n23273 ;
  assign n33032 = n33031 ^ n18571 ^ 1'b0 ;
  assign n33033 = n24127 ^ n14740 ^ 1'b0 ;
  assign n33034 = n16255 | n33033 ;
  assign n33035 = n33034 ^ n2120 ^ 1'b0 ;
  assign n33036 = ~n21901 & n33035 ;
  assign n33037 = ~n3444 & n20547 ;
  assign n33038 = n8048 | n33037 ;
  assign n33039 = n16072 & ~n16911 ;
  assign n33040 = ~n33038 & n33039 ;
  assign n33041 = n13399 | n22116 ;
  assign n33042 = n28698 | n33041 ;
  assign n33043 = ~n10177 & n33042 ;
  assign n33044 = n33043 ^ n21712 ^ 1'b0 ;
  assign n33045 = n25866 ^ n21856 ^ 1'b0 ;
  assign n33046 = n20145 & ~n33045 ;
  assign n33047 = n7141 | n32614 ;
  assign n33048 = ~n7046 & n10628 ;
  assign n33049 = n19348 ^ n3981 ^ 1'b0 ;
  assign n33050 = n33049 ^ n23297 ^ 1'b0 ;
  assign n33051 = n6602 | n14281 ;
  assign n33052 = n33051 ^ n9504 ^ 1'b0 ;
  assign n33053 = n3039 | n33052 ;
  assign n33054 = n33053 ^ n10610 ^ 1'b0 ;
  assign n33055 = n15770 & ~n24570 ;
  assign n33056 = n15575 | n33055 ;
  assign n33057 = n6592 ^ n5659 ^ n3509 ;
  assign n33058 = n31761 & ~n33057 ;
  assign n33059 = n4974 & ~n30698 ;
  assign n33060 = ~n4635 & n33059 ;
  assign n33061 = n466 | n4511 ;
  assign n33062 = n2431 | n6202 ;
  assign n33063 = n10043 | n33062 ;
  assign n33064 = n10397 & n15311 ;
  assign n33065 = n33064 ^ n15098 ^ 1'b0 ;
  assign n33066 = ~n10356 & n33065 ;
  assign n33067 = n5759 | n6999 ;
  assign n33068 = n29439 ^ n14902 ^ 1'b0 ;
  assign n33069 = n33067 & ~n33068 ;
  assign n33070 = n33069 ^ n5282 ^ 1'b0 ;
  assign n33071 = n14501 | n16178 ;
  assign n33072 = n16535 | n33071 ;
  assign n33073 = n7888 | n9803 ;
  assign n33074 = n29049 ^ n13693 ^ n10637 ;
  assign n33075 = n33074 ^ n1830 ^ 1'b0 ;
  assign n33076 = ~n33073 & n33075 ;
  assign n33077 = n11522 ^ n4764 ^ n2622 ;
  assign n33078 = n10310 | n32039 ;
  assign n33080 = n20629 ^ n6978 ^ 1'b0 ;
  assign n33081 = ~n3744 & n33080 ;
  assign n33079 = ( n9466 & n21893 ) | ( n9466 & n25200 ) | ( n21893 & n25200 ) ;
  assign n33082 = n33081 ^ n33079 ^ 1'b0 ;
  assign n33083 = n16864 | n33082 ;
  assign n33084 = ~n7617 & n16228 ;
  assign n33085 = ~n705 & n8947 ;
  assign n33086 = n33085 ^ n4838 ^ 1'b0 ;
  assign n33087 = n32018 ^ n2122 ^ 1'b0 ;
  assign n33088 = ~n12394 & n33087 ;
  assign n33089 = n4638 | n9531 ;
  assign n33090 = n3977 & ~n33089 ;
  assign n33091 = n5509 & ~n33090 ;
  assign n33092 = ~n22658 & n33091 ;
  assign n33093 = n33092 ^ n1603 ^ 1'b0 ;
  assign n33094 = n781 & n23094 ;
  assign n33095 = n33094 ^ n6642 ^ 1'b0 ;
  assign n33096 = n20799 ^ n6378 ^ 1'b0 ;
  assign n33097 = n3668 | n33096 ;
  assign n33098 = n6642 & ~n11138 ;
  assign n33099 = ~n16903 & n33098 ;
  assign n33100 = n11923 & ~n27667 ;
  assign n33101 = n17548 ^ n9674 ^ n6817 ;
  assign n33102 = ( ~n8897 & n9967 ) | ( ~n8897 & n25600 ) | ( n9967 & n25600 ) ;
  assign n33103 = n2178 & ~n33102 ;
  assign n33104 = n17970 | n24941 ;
  assign n33105 = n33104 ^ n31645 ^ 1'b0 ;
  assign n33106 = ~n2944 & n15461 ;
  assign n33107 = n33106 ^ n7222 ^ 1'b0 ;
  assign n33108 = n10629 | n33107 ;
  assign n33109 = ~n12066 & n24524 ;
  assign n33110 = n25495 ^ n13776 ^ 1'b0 ;
  assign n33111 = n33109 & ~n33110 ;
  assign n33112 = n33111 ^ n25511 ^ 1'b0 ;
  assign n33113 = n8940 & n29319 ;
  assign n33114 = ~n3396 & n33113 ;
  assign n33115 = n33114 ^ n16663 ^ 1'b0 ;
  assign n33118 = n7972 ^ n2883 ^ 1'b0 ;
  assign n33119 = n14437 | n33118 ;
  assign n33116 = n5700 ^ n1707 ^ 1'b0 ;
  assign n33117 = n25906 & n33116 ;
  assign n33120 = n33119 ^ n33117 ^ 1'b0 ;
  assign n33121 = n18104 ^ n6120 ^ 1'b0 ;
  assign n33122 = n25236 & n33121 ;
  assign n33123 = ~n796 & n33122 ;
  assign n33124 = n33123 ^ n19966 ^ 1'b0 ;
  assign n33125 = n30977 ^ n8066 ^ n3092 ;
  assign n33126 = n33125 ^ n8627 ^ 1'b0 ;
  assign n33127 = n3705 & n14363 ;
  assign n33128 = n3867 | n23904 ;
  assign n33129 = n12817 | n13330 ;
  assign n33130 = n33129 ^ n4643 ^ 1'b0 ;
  assign n33131 = n33130 ^ n14459 ^ 1'b0 ;
  assign n33132 = n31399 & n33131 ;
  assign n33133 = n20536 ^ n7838 ^ 1'b0 ;
  assign n33134 = n33133 ^ n20450 ^ 1'b0 ;
  assign n33135 = n22680 & ~n26534 ;
  assign n33136 = n33135 ^ n20797 ^ 1'b0 ;
  assign n33137 = n9640 & n29524 ;
  assign n33138 = n12887 & n33137 ;
  assign n33139 = n28829 & ~n33138 ;
  assign n33140 = n13653 & n25750 ;
  assign n33141 = n3163 & n28837 ;
  assign n33142 = x251 & n26892 ;
  assign n33143 = ~n4157 & n33142 ;
  assign n33145 = n21048 ^ n4832 ^ n2122 ;
  assign n33144 = n6939 & ~n30287 ;
  assign n33146 = n33145 ^ n33144 ^ 1'b0 ;
  assign n33147 = n33114 ^ n11625 ^ 1'b0 ;
  assign n33148 = ( n6059 & ~n9041 ) | ( n6059 & n33147 ) | ( ~n9041 & n33147 ) ;
  assign n33149 = ( n6451 & n19285 ) | ( n6451 & n19823 ) | ( n19285 & n19823 ) ;
  assign n33150 = n27402 ^ n6307 ^ 1'b0 ;
  assign n33151 = n31559 & ~n33150 ;
  assign n33152 = n15456 ^ n542 ^ 1'b0 ;
  assign n33153 = n33152 ^ n3117 ^ 1'b0 ;
  assign n33154 = n2155 & ~n33153 ;
  assign n33155 = n25018 ^ n2961 ^ 1'b0 ;
  assign n33156 = ~n15131 & n31197 ;
  assign n33157 = n33156 ^ n9210 ^ 1'b0 ;
  assign n33158 = n14725 ^ n9815 ^ 1'b0 ;
  assign n33159 = n32930 ^ n14136 ^ 1'b0 ;
  assign n33160 = n13121 | n32682 ;
  assign n33161 = n9560 | n33160 ;
  assign n33162 = n24514 ^ n3908 ^ 1'b0 ;
  assign n33163 = n9407 ^ n6862 ^ 1'b0 ;
  assign n33164 = n30537 & n33163 ;
  assign n33165 = n8098 & ~n13689 ;
  assign n33166 = n10555 & n33165 ;
  assign n33167 = n33166 ^ n8404 ^ 1'b0 ;
  assign n33168 = n9928 & n31052 ;
  assign n33169 = n906 & n8150 ;
  assign n33170 = x30 & n25671 ;
  assign n33171 = n33169 & n33170 ;
  assign n33172 = n13720 | n24595 ;
  assign n33173 = n5754 ^ n5522 ^ 1'b0 ;
  assign n33174 = n33173 ^ n22363 ^ 1'b0 ;
  assign n33175 = ~n3529 & n33174 ;
  assign n33176 = n30681 ^ n23123 ^ 1'b0 ;
  assign n33177 = n1653 & n33176 ;
  assign n33178 = n17330 & n29299 ;
  assign n33179 = n5091 & ~n11722 ;
  assign n33180 = ~n5091 & n33179 ;
  assign n33181 = n4934 & ~n19639 ;
  assign n33182 = x244 | n8618 ;
  assign n33183 = n33182 ^ n25128 ^ 1'b0 ;
  assign n33184 = n10225 | n11041 ;
  assign n33185 = n9533 | n18948 ;
  assign n33186 = n11199 & n14138 ;
  assign n33187 = n17901 | n33186 ;
  assign n33188 = n458 & n15711 ;
  assign n33189 = n33188 ^ n20107 ^ 1'b0 ;
  assign n33190 = n30873 ^ n11056 ^ n5665 ;
  assign n33191 = ~n29464 & n33190 ;
  assign n33192 = n5652 & ~n7398 ;
  assign n33193 = ( n10416 & ~n27206 ) | ( n10416 & n33192 ) | ( ~n27206 & n33192 ) ;
  assign n33194 = x143 & n882 ;
  assign n33195 = n33194 ^ n9310 ^ n8133 ;
  assign n33196 = n2789 & ~n33195 ;
  assign n33197 = n29215 ^ n16525 ^ 1'b0 ;
  assign n33198 = ~n5380 & n24443 ;
  assign n33199 = n17220 & ~n33198 ;
  assign n33200 = ~n3000 & n19126 ;
  assign n33201 = n11583 ^ n1148 ^ 1'b0 ;
  assign n33202 = ( n14739 & n22867 ) | ( n14739 & ~n33201 ) | ( n22867 & ~n33201 ) ;
  assign n33203 = n765 | n32709 ;
  assign n33204 = n2040 | n33203 ;
  assign n33205 = n32130 & ~n33204 ;
  assign n33206 = n33205 ^ n4453 ^ 1'b0 ;
  assign n33207 = n33206 ^ n29031 ^ n20447 ;
  assign n33208 = n2940 & ~n28507 ;
  assign n33209 = ~n10860 & n33208 ;
  assign n33210 = ( ~n4377 & n14087 ) | ( ~n4377 & n15977 ) | ( n14087 & n15977 ) ;
  assign n33211 = n33210 ^ n26535 ^ 1'b0 ;
  assign n33212 = ~n25057 & n33211 ;
  assign n33213 = n20739 | n22913 ;
  assign n33214 = n2226 & ~n2375 ;
  assign n33215 = n4706 & n33214 ;
  assign n33216 = n5100 | n33215 ;
  assign n33217 = n33216 ^ n12848 ^ n1835 ;
  assign n33218 = ~n15565 & n18361 ;
  assign n33219 = n33218 ^ n25240 ^ 1'b0 ;
  assign n33220 = n11857 & n15453 ;
  assign n33221 = n1443 | n9072 ;
  assign n33222 = n258 & ~n33221 ;
  assign n33223 = n361 & ~n496 ;
  assign n33224 = n33222 | n33223 ;
  assign n33225 = n1547 | n33224 ;
  assign n33226 = n3087 & ~n21259 ;
  assign n33227 = n1048 & n33226 ;
  assign n33228 = ~n33225 & n33227 ;
  assign n33229 = n12503 & n32892 ;
  assign n33230 = n3385 & ~n5362 ;
  assign n33231 = ( n5177 & ~n31174 ) | ( n5177 & n33230 ) | ( ~n31174 & n33230 ) ;
  assign n33232 = x164 & n11623 ;
  assign n33233 = n3215 & n33232 ;
  assign n33234 = n21109 | n33233 ;
  assign n33235 = n2366 & ~n3954 ;
  assign n33236 = x56 & n28862 ;
  assign n33237 = n22829 ^ n8406 ^ 1'b0 ;
  assign n33238 = n817 & n14263 ;
  assign n33239 = n18758 ^ n11182 ^ n3879 ;
  assign n33240 = n25230 & ~n33239 ;
  assign n33241 = n7895 ^ n6429 ^ 1'b0 ;
  assign n33242 = n6114 & n33241 ;
  assign n33243 = n10376 ^ n7472 ^ 1'b0 ;
  assign n33244 = n8751 & ~n24062 ;
  assign n33245 = n33244 ^ n12699 ^ 1'b0 ;
  assign n33246 = n4918 & ~n11995 ;
  assign n33247 = n16340 & n33246 ;
  assign n33248 = n10079 | n19361 ;
  assign n33249 = n15065 ^ n7025 ^ x223 ;
  assign n33250 = n22461 & n33249 ;
  assign n33251 = n33250 ^ n23996 ^ 1'b0 ;
  assign n33252 = n6297 & ~n24941 ;
  assign n33253 = n8375 ^ n6525 ^ 1'b0 ;
  assign n33254 = ~n31783 & n33253 ;
  assign n33255 = n1048 & n30475 ;
  assign n33256 = n21871 & n33255 ;
  assign n33257 = n7350 & ~n18161 ;
  assign n33259 = n30587 ^ n12696 ^ 1'b0 ;
  assign n33260 = n4875 | n33259 ;
  assign n33258 = n11852 & n29936 ;
  assign n33261 = n33260 ^ n33258 ^ 1'b0 ;
  assign n33262 = ~n5261 & n27103 ;
  assign n33263 = ~n17176 & n33262 ;
  assign n33264 = n8280 ^ n2182 ^ 1'b0 ;
  assign n33265 = ~n25023 & n33264 ;
  assign n33266 = n6359 ^ n317 ^ 1'b0 ;
  assign n33267 = n24717 & ~n33266 ;
  assign n33268 = n8322 & n13511 ;
  assign n33269 = n11433 & n33268 ;
  assign n33270 = n13097 & ~n29686 ;
  assign n33271 = n10849 & n33270 ;
  assign n33272 = n4122 & ~n29408 ;
  assign n33273 = n10336 ^ n5163 ^ 1'b0 ;
  assign n33274 = n16859 & n19524 ;
  assign n33275 = ~n24739 & n33274 ;
  assign n33276 = n19215 ^ n3505 ^ 1'b0 ;
  assign n33277 = n28748 ^ n15145 ^ 1'b0 ;
  assign n33278 = n33276 & ~n33277 ;
  assign n33279 = n5619 & n9816 ;
  assign n33280 = n7974 | n9545 ;
  assign n33281 = n9706 & ~n33280 ;
  assign n33282 = ( x2 & n15574 ) | ( x2 & n33281 ) | ( n15574 & n33281 ) ;
  assign n33283 = ~n10985 & n33282 ;
  assign n33284 = n17352 | n21700 ;
  assign n33285 = n13231 & ~n33284 ;
  assign n33286 = n4598 | n12328 ;
  assign n33287 = n27347 ^ n21720 ^ 1'b0 ;
  assign n33288 = n1439 | n33287 ;
  assign n33290 = n7743 & n9864 ;
  assign n33289 = ~n24778 & n30779 ;
  assign n33291 = n33290 ^ n33289 ^ 1'b0 ;
  assign n33292 = n12669 | n18485 ;
  assign n33293 = n4284 | n21233 ;
  assign n33294 = ~n739 & n1971 ;
  assign n33295 = n4003 ^ n3213 ^ 1'b0 ;
  assign n33296 = n20252 & ~n33295 ;
  assign n33297 = n9863 & n33296 ;
  assign n33298 = n7450 ^ n1579 ^ 1'b0 ;
  assign n33299 = n8406 & ~n33298 ;
  assign n33300 = n20449 ^ n12699 ^ 1'b0 ;
  assign n33301 = n17041 ^ x20 ^ 1'b0 ;
  assign n33302 = n11162 ^ x141 ^ 1'b0 ;
  assign n33303 = n10807 | n33302 ;
  assign n33304 = n23382 ^ n15666 ^ 1'b0 ;
  assign n33305 = n20550 & ~n33304 ;
  assign n33306 = ( n451 & n28033 ) | ( n451 & ~n33305 ) | ( n28033 & ~n33305 ) ;
  assign n33307 = n12963 & n28347 ;
  assign n33308 = n2725 | n12142 ;
  assign n33309 = ~n24376 & n33308 ;
  assign n33310 = n13580 & ~n23599 ;
  assign n33311 = ( n943 & ~n4375 ) | ( n943 & n15252 ) | ( ~n4375 & n15252 ) ;
  assign n33312 = n31039 & ~n33311 ;
  assign n33313 = n14971 & n33312 ;
  assign n33314 = n18502 ^ n6741 ^ 1'b0 ;
  assign n33315 = n12381 & n33314 ;
  assign n33316 = n5980 | n33315 ;
  assign n33317 = n33316 ^ n31431 ^ 1'b0 ;
  assign n33321 = n12831 ^ n3855 ^ 1'b0 ;
  assign n33322 = ~n9813 & n33321 ;
  assign n33318 = n10299 & ~n17338 ;
  assign n33319 = n5932 & n33318 ;
  assign n33320 = n10498 | n33319 ;
  assign n33323 = n33322 ^ n33320 ^ n12499 ;
  assign n33324 = n21843 ^ n13584 ^ 1'b0 ;
  assign n33325 = n2150 ^ n1382 ^ 1'b0 ;
  assign n33326 = n5094 | n33325 ;
  assign n33327 = ~n10006 & n21164 ;
  assign n33328 = n33326 | n33327 ;
  assign n33329 = n8674 & ~n10061 ;
  assign n33330 = ~n794 & n33329 ;
  assign n33331 = n33330 ^ n30495 ^ n13856 ;
  assign n33332 = n33331 ^ n12256 ^ 1'b0 ;
  assign n33333 = n1791 | n33332 ;
  assign n33334 = x61 & ~n33333 ;
  assign n33335 = n19746 ^ n9992 ^ 1'b0 ;
  assign n33336 = n31174 ^ n3420 ^ 1'b0 ;
  assign n33337 = ( n8907 & n12679 ) | ( n8907 & n33336 ) | ( n12679 & n33336 ) ;
  assign n33338 = n31378 ^ n7519 ^ 1'b0 ;
  assign n33339 = n25114 | n33338 ;
  assign n33340 = n3052 & ~n4643 ;
  assign n33341 = n33340 ^ n4302 ^ 1'b0 ;
  assign n33342 = ~n15575 & n33341 ;
  assign n33343 = n25415 & n33342 ;
  assign n33344 = n33343 ^ n26930 ^ 1'b0 ;
  assign n33347 = n8994 ^ n3707 ^ 1'b0 ;
  assign n33345 = n15473 ^ n5975 ^ 1'b0 ;
  assign n33346 = n19677 & ~n33345 ;
  assign n33348 = n33347 ^ n33346 ^ n11567 ;
  assign n33350 = n7573 | n7967 ;
  assign n33349 = n3195 & ~n10062 ;
  assign n33351 = n33350 ^ n33349 ^ 1'b0 ;
  assign n33352 = n33351 ^ n24854 ^ n22019 ;
  assign n33353 = n17126 ^ n4494 ^ n2657 ;
  assign n33354 = n9912 & ~n24266 ;
  assign n33355 = n33354 ^ n10570 ^ 1'b0 ;
  assign n33356 = n1776 & ~n11328 ;
  assign n33357 = n1025 & ~n2600 ;
  assign n33358 = n9499 & n33357 ;
  assign n33359 = ~n13976 & n14109 ;
  assign n33360 = n33359 ^ n8360 ^ 1'b0 ;
  assign n33361 = n13510 & n30555 ;
  assign n33362 = ~n18108 & n33361 ;
  assign n33363 = ~n23163 & n24992 ;
  assign n33364 = ~n5746 & n19370 ;
  assign n33365 = n33364 ^ n26463 ^ 1'b0 ;
  assign n33366 = n3385 | n16679 ;
  assign n33367 = n13612 ^ n10150 ^ 1'b0 ;
  assign n33368 = n5154 & n33367 ;
  assign n33369 = n2102 & ~n16571 ;
  assign n33370 = n25267 | n33369 ;
  assign n33371 = n1133 & ~n23271 ;
  assign n33372 = n8178 & n33371 ;
  assign n33373 = ~n3111 & n8822 ;
  assign n33374 = n3111 & n33373 ;
  assign n33375 = ~n22521 & n22928 ;
  assign n33376 = n33374 & n33375 ;
  assign n33377 = n33376 ^ n2740 ^ 1'b0 ;
  assign n33378 = n24504 & ~n33377 ;
  assign n33379 = n18729 ^ n12530 ^ 1'b0 ;
  assign n33380 = ~n776 & n19671 ;
  assign n33381 = n33379 & n33380 ;
  assign n33382 = n5617 ^ n2216 ^ 1'b0 ;
  assign n33383 = n12328 | n32822 ;
  assign n33384 = n18006 | n21096 ;
  assign n33385 = n12355 & ~n13366 ;
  assign n33386 = n33385 ^ n24551 ^ 1'b0 ;
  assign n33387 = ~n21460 & n29049 ;
  assign n33388 = n8129 & ~n30524 ;
  assign n33389 = n22584 ^ x215 ^ 1'b0 ;
  assign n33390 = n11685 & n22265 ;
  assign n33391 = ( ~n5081 & n32700 ) | ( ~n5081 & n33390 ) | ( n32700 & n33390 ) ;
  assign n33392 = n2343 & n11701 ;
  assign n33393 = n5023 | n14025 ;
  assign n33394 = n33393 ^ n1167 ^ 1'b0 ;
  assign n33395 = ~n1153 & n27081 ;
  assign n33396 = n33395 ^ n14059 ^ 1'b0 ;
  assign n33397 = n6256 & n13091 ;
  assign n33398 = n14445 & ~n16669 ;
  assign n33399 = n33398 ^ n10776 ^ 1'b0 ;
  assign n33400 = n33397 & n33399 ;
  assign n33401 = n33400 ^ n2164 ^ 1'b0 ;
  assign n33402 = n1519 & n2370 ;
  assign n33403 = ( n5481 & n6886 ) | ( n5481 & ~n33402 ) | ( n6886 & ~n33402 ) ;
  assign n33404 = n13184 & ~n22632 ;
  assign n33405 = n13502 & n13774 ;
  assign n33406 = ~n9006 & n33405 ;
  assign n33407 = n12653 & ~n16838 ;
  assign n33408 = n33407 ^ n9007 ^ 1'b0 ;
  assign n33409 = n4368 & n33408 ;
  assign n33410 = n27569 & n33409 ;
  assign n33411 = n33410 ^ n4241 ^ 1'b0 ;
  assign n33412 = ~n440 & n16068 ;
  assign n33413 = ~n22554 & n33412 ;
  assign n33414 = n2684 & n7258 ;
  assign n33415 = n33414 ^ n5619 ^ 1'b0 ;
  assign n33416 = n23951 ^ n4979 ^ 1'b0 ;
  assign n33417 = n20453 ^ n15137 ^ 1'b0 ;
  assign n33418 = n6358 ^ n1876 ^ 1'b0 ;
  assign n33419 = n4815 ^ n3010 ^ 1'b0 ;
  assign n33420 = ~n25273 & n33419 ;
  assign n33421 = n9970 & ~n32563 ;
  assign n33422 = ~n33420 & n33421 ;
  assign n33423 = n16012 ^ n13538 ^ n11253 ;
  assign n33424 = n33423 ^ n25088 ^ x182 ;
  assign n33425 = ( n395 & n4861 ) | ( n395 & ~n27214 ) | ( n4861 & ~n27214 ) ;
  assign n33427 = n10554 | n20125 ;
  assign n33428 = n33427 ^ n4711 ^ 1'b0 ;
  assign n33426 = n15348 & n17010 ;
  assign n33429 = n33428 ^ n33426 ^ 1'b0 ;
  assign n33430 = n15255 ^ n4438 ^ 1'b0 ;
  assign n33431 = n18277 | n27094 ;
  assign n33432 = n21758 & ~n33431 ;
  assign n33433 = ~n23504 & n28373 ;
  assign n33434 = ~n1482 & n30242 ;
  assign n33435 = n33434 ^ n27146 ^ 1'b0 ;
  assign n33436 = n8587 | n31889 ;
  assign n33437 = n33436 ^ n13809 ^ 1'b0 ;
  assign n33438 = n5884 & n6696 ;
  assign n33439 = ( n5963 & ~n17190 ) | ( n5963 & n33438 ) | ( ~n17190 & n33438 ) ;
  assign n33440 = n12996 & n18959 ;
  assign n33441 = ~n20578 & n33440 ;
  assign n33442 = n5657 & ~n31957 ;
  assign n33443 = ~n10676 & n17127 ;
  assign n33444 = n7922 | n33443 ;
  assign n33445 = ~n24581 & n33444 ;
  assign n33446 = n2953 & n33445 ;
  assign n33447 = n21726 ^ n9377 ^ n1032 ;
  assign n33448 = n5983 & n23765 ;
  assign n33449 = n10112 ^ n9976 ^ 1'b0 ;
  assign n33450 = n19830 ^ n13606 ^ 1'b0 ;
  assign n33451 = ~n25188 & n25696 ;
  assign n33452 = n6161 & n33451 ;
  assign n33453 = n33450 & ~n33452 ;
  assign n33454 = n19815 ^ n19303 ^ 1'b0 ;
  assign n33455 = ~n5353 & n33454 ;
  assign n33456 = ~x89 & n5418 ;
  assign n33457 = n31819 & n33456 ;
  assign n33458 = ~n8520 & n31089 ;
  assign n33459 = ~n19671 & n33458 ;
  assign n33460 = n2211 & n16720 ;
  assign n33461 = ~n376 & n7219 ;
  assign n33462 = n10991 & n33461 ;
  assign n33463 = n11496 ^ n705 ^ 1'b0 ;
  assign n33464 = n30331 ^ n13126 ^ n11911 ;
  assign n33465 = n28581 ^ n10805 ^ 1'b0 ;
  assign n33466 = ~n8991 & n12446 ;
  assign n33467 = ~n12446 & n33466 ;
  assign n33468 = n9905 & ~n33467 ;
  assign n33469 = n33468 ^ n1730 ^ 1'b0 ;
  assign n33470 = n33469 ^ n1103 ^ 1'b0 ;
  assign n33471 = ( n4465 & n8321 ) | ( n4465 & n16149 ) | ( n8321 & n16149 ) ;
  assign n33472 = n33471 ^ n11816 ^ 1'b0 ;
  assign n33473 = n28362 ^ n16932 ^ n14236 ;
  assign n33474 = n27718 | n33473 ;
  assign n33475 = ( n4496 & ~n22656 ) | ( n4496 & n26833 ) | ( ~n22656 & n26833 ) ;
  assign n33476 = n9117 ^ n3396 ^ 1'b0 ;
  assign n33477 = n8682 & n33476 ;
  assign n33478 = n11270 ^ x45 ^ 1'b0 ;
  assign n33479 = n1899 & n6714 ;
  assign n33480 = n33478 & n33479 ;
  assign n33484 = n20354 & ~n30234 ;
  assign n33481 = ~n1575 & n28672 ;
  assign n33482 = n30015 & n33481 ;
  assign n33483 = n24676 | n33482 ;
  assign n33485 = n33484 ^ n33483 ^ 1'b0 ;
  assign n33486 = n17287 & n33485 ;
  assign n33487 = n21863 & n33486 ;
  assign n33488 = x202 & n374 ;
  assign n33489 = n33488 ^ n15131 ^ 1'b0 ;
  assign n33490 = n33489 ^ n7629 ^ 1'b0 ;
  assign n33491 = n4520 & n33490 ;
  assign n33492 = n12036 ^ n10876 ^ 1'b0 ;
  assign n33493 = ( n5392 & ~n25205 ) | ( n5392 & n32123 ) | ( ~n25205 & n32123 ) ;
  assign n33494 = n613 & n33062 ;
  assign n33495 = n24977 & n33494 ;
  assign n33496 = n2178 | n4755 ;
  assign n33497 = n6203 & ~n33496 ;
  assign n33498 = n33495 & n33497 ;
  assign n33500 = n4899 ^ n4157 ^ 1'b0 ;
  assign n33501 = ~n6144 & n33500 ;
  assign n33499 = n6315 | n29919 ;
  assign n33502 = n33501 ^ n33499 ^ 1'b0 ;
  assign n33503 = n20918 ^ n15653 ^ 1'b0 ;
  assign n33504 = ~n4491 & n33503 ;
  assign n33506 = ~n8676 & n13947 ;
  assign n33505 = n9824 & n10650 ;
  assign n33507 = n33506 ^ n33505 ^ 1'b0 ;
  assign n33508 = n20386 | n21990 ;
  assign n33509 = n33507 & ~n33508 ;
  assign n33510 = n31515 & ~n33509 ;
  assign n33511 = n7666 ^ n3835 ^ 1'b0 ;
  assign n33512 = n15392 & n33511 ;
  assign n33513 = n1596 & n33512 ;
  assign n33514 = n33513 ^ n14930 ^ 1'b0 ;
  assign n33515 = n13259 ^ n3243 ^ 1'b0 ;
  assign n33516 = ~n26906 & n33515 ;
  assign n33517 = n33516 ^ n3640 ^ 1'b0 ;
  assign n33518 = n23131 ^ n2055 ^ 1'b0 ;
  assign n33519 = ~n19726 & n24449 ;
  assign n33520 = n31351 | n33519 ;
  assign n33521 = n5355 & n23270 ;
  assign n33522 = n33521 ^ n16467 ^ 1'b0 ;
  assign n33524 = n27119 ^ x173 ^ 1'b0 ;
  assign n33523 = n23150 ^ n8141 ^ 1'b0 ;
  assign n33525 = n33524 ^ n33523 ^ n29004 ;
  assign n33526 = n13095 & n26283 ;
  assign n33527 = n19435 ^ n786 ^ 1'b0 ;
  assign n33528 = n33526 & ~n33527 ;
  assign n33529 = n13546 & n15131 ;
  assign n33530 = ~n711 & n33529 ;
  assign n33531 = n19502 | n33530 ;
  assign n33532 = x84 & ~n27415 ;
  assign n33533 = n21873 & n33532 ;
  assign n33534 = ~n6881 & n23423 ;
  assign n33535 = n33534 ^ n9594 ^ n378 ;
  assign n33536 = n33533 | n33535 ;
  assign n33537 = n33536 ^ n13505 ^ 1'b0 ;
  assign n33538 = n9496 | n32582 ;
  assign n33539 = n33538 ^ n25872 ^ 1'b0 ;
  assign n33540 = n7384 & n9569 ;
  assign n33541 = n33540 ^ n15181 ^ 1'b0 ;
  assign n33542 = n5811 ^ x22 ^ 1'b0 ;
  assign n33543 = x207 & ~n33542 ;
  assign n33544 = n33543 ^ n3389 ^ 1'b0 ;
  assign n33545 = ~n30751 & n33544 ;
  assign n33546 = n14620 ^ n12226 ^ n595 ;
  assign n33547 = n1092 & n5983 ;
  assign n33548 = n33547 ^ n8082 ^ 1'b0 ;
  assign n33549 = n28206 ^ n17763 ^ 1'b0 ;
  assign n33550 = ~n33548 & n33549 ;
  assign n33551 = n12719 ^ n4458 ^ 1'b0 ;
  assign n33552 = n1272 & ~n33551 ;
  assign n33553 = n7085 ^ x192 ^ 1'b0 ;
  assign n33554 = n27244 & ~n33553 ;
  assign n33555 = n17009 ^ n13582 ^ 1'b0 ;
  assign n33556 = n33555 ^ n13991 ^ 1'b0 ;
  assign n33557 = n10480 ^ n4443 ^ n2170 ;
  assign n33558 = ~n9686 & n18394 ;
  assign n33559 = n12275 ^ n10808 ^ 1'b0 ;
  assign n33560 = ~n5089 & n33559 ;
  assign n33561 = n7255 & n10259 ;
  assign n33562 = ~n33560 & n33561 ;
  assign n33563 = n12700 ^ x20 ^ 1'b0 ;
  assign n33564 = n8304 | n33563 ;
  assign n33565 = n27003 & ~n33564 ;
  assign n33566 = x231 & ~n3134 ;
  assign n33567 = n33566 ^ n18164 ^ 1'b0 ;
  assign n33568 = n27864 ^ n8273 ^ 1'b0 ;
  assign n33570 = n799 | n2661 ;
  assign n33571 = n2661 & ~n33570 ;
  assign n33572 = x169 | n7124 ;
  assign n33573 = n7124 & ~n33572 ;
  assign n33574 = n33573 ^ n1997 ^ 1'b0 ;
  assign n33575 = n33574 ^ n3030 ^ 1'b0 ;
  assign n33576 = n33571 | n33575 ;
  assign n33569 = n2274 & ~n4818 ;
  assign n33577 = n33576 ^ n33569 ^ 1'b0 ;
  assign n33581 = ( ~x163 & n16594 ) | ( ~x163 & n23405 ) | ( n16594 & n23405 ) ;
  assign n33578 = n9794 | n23044 ;
  assign n33579 = x247 ^ x129 ^ 1'b0 ;
  assign n33580 = ~n33578 & n33579 ;
  assign n33582 = n33581 ^ n33580 ^ 1'b0 ;
  assign n33583 = n18924 ^ n14694 ^ 1'b0 ;
  assign n33584 = n12730 | n20916 ;
  assign n33585 = n11372 ^ n5737 ^ 1'b0 ;
  assign n33586 = n5209 & ~n33585 ;
  assign n33587 = n4555 & n33586 ;
  assign n33588 = ~n25396 & n33587 ;
  assign n33589 = ~n19243 & n26139 ;
  assign n33590 = n1133 & n9202 ;
  assign n33591 = n1977 & n4547 ;
  assign n33592 = ~n33590 & n33591 ;
  assign n33593 = n28802 ^ n15319 ^ 1'b0 ;
  assign n33594 = n7173 | n24426 ;
  assign n33595 = n33594 ^ n27710 ^ 1'b0 ;
  assign n33596 = ( n18331 & n32620 ) | ( n18331 & ~n33595 ) | ( n32620 & ~n33595 ) ;
  assign n33597 = n1373 | n5893 ;
  assign n33598 = ~n3385 & n4919 ;
  assign n33599 = ~n23662 & n33598 ;
  assign n33600 = ~n14676 & n18428 ;
  assign n33601 = n33600 ^ n10911 ^ 1'b0 ;
  assign n33602 = n33601 ^ n3750 ^ 1'b0 ;
  assign n33603 = n6633 & n33114 ;
  assign n33604 = n3755 & ~n27244 ;
  assign n33607 = n372 & n22122 ;
  assign n33605 = n9738 & ~n17185 ;
  assign n33606 = n33605 ^ n2912 ^ 1'b0 ;
  assign n33608 = n33607 ^ n33606 ^ n622 ;
  assign n33609 = n8351 & ~n13737 ;
  assign n33610 = n33609 ^ n5058 ^ x143 ;
  assign n33611 = n863 & n20099 ;
  assign n33612 = n12565 ^ n9429 ^ 1'b0 ;
  assign n33613 = n5276 & n33612 ;
  assign n33614 = n25923 & n33613 ;
  assign n33615 = n33614 ^ n28190 ^ 1'b0 ;
  assign n33616 = n3880 | n25733 ;
  assign n33617 = ~n6551 & n8978 ;
  assign n33618 = n33617 ^ n22837 ^ 1'b0 ;
  assign n33619 = n25481 ^ n16964 ^ 1'b0 ;
  assign n33620 = n29846 & ~n33619 ;
  assign n33621 = n22117 ^ n1303 ^ 1'b0 ;
  assign n33622 = n26663 & n33621 ;
  assign n33623 = n33622 ^ n29002 ^ 1'b0 ;
  assign n33624 = n18568 ^ n16177 ^ 1'b0 ;
  assign n33625 = ( n1336 & ~n11458 ) | ( n1336 & n33624 ) | ( ~n11458 & n33624 ) ;
  assign n33626 = n21486 ^ n296 ^ 1'b0 ;
  assign n33627 = n11498 & n33626 ;
  assign n33628 = n33625 & n33627 ;
  assign n33629 = n4092 | n24290 ;
  assign n33630 = n22910 ^ n15445 ^ n13011 ;
  assign n33631 = n826 & n18136 ;
  assign n33632 = n12335 | n16665 ;
  assign n33633 = n18825 & ~n33632 ;
  assign n33634 = n19292 & ~n33633 ;
  assign n33635 = n11854 & n20648 ;
  assign n33636 = ~n7732 & n33635 ;
  assign n33637 = ~n6246 & n32517 ;
  assign n33638 = n33636 & n33637 ;
  assign n33639 = n1361 & ~n33638 ;
  assign n33640 = n33639 ^ n9852 ^ 1'b0 ;
  assign n33641 = n10174 & n21980 ;
  assign n33642 = n17889 ^ n1508 ^ 1'b0 ;
  assign n33643 = n5565 ^ n3843 ^ 1'b0 ;
  assign n33644 = n15985 & n33643 ;
  assign n33645 = n13716 ^ n622 ^ 1'b0 ;
  assign n33646 = ~n5367 & n33645 ;
  assign n33647 = n31743 ^ n25652 ^ 1'b0 ;
  assign n33648 = n29552 | n33647 ;
  assign n33649 = n11796 | n33648 ;
  assign n33650 = n2724 | n33649 ;
  assign n33651 = n6276 ^ n3546 ^ 1'b0 ;
  assign n33652 = n6276 | n33651 ;
  assign n33653 = n4801 | n10889 ;
  assign n33654 = n16408 ^ n1051 ^ 1'b0 ;
  assign n33655 = n33653 | n33654 ;
  assign n33666 = n15983 ^ n13151 ^ 1'b0 ;
  assign n33667 = n7866 & n33666 ;
  assign n33656 = n6700 & ~n27336 ;
  assign n33657 = n33656 ^ n10731 ^ 1'b0 ;
  assign n33658 = n2535 & ~n15699 ;
  assign n33659 = n9039 & n33658 ;
  assign n33660 = n33659 ^ n15795 ^ 1'b0 ;
  assign n33661 = n8814 ^ n1247 ^ 1'b0 ;
  assign n33662 = n33661 ^ n23907 ^ 1'b0 ;
  assign n33663 = n33660 & ~n33662 ;
  assign n33664 = ~n22451 & n33663 ;
  assign n33665 = ~n33657 & n33664 ;
  assign n33668 = n33667 ^ n33665 ^ 1'b0 ;
  assign n33669 = ~n33655 & n33668 ;
  assign n33670 = n494 | n14546 ;
  assign n33671 = n33669 | n33670 ;
  assign n33672 = n32669 ^ n28514 ^ 1'b0 ;
  assign n33673 = n14637 ^ n349 ^ 1'b0 ;
  assign n33674 = n5542 & n8112 ;
  assign n33675 = n17590 & n33674 ;
  assign n33676 = n32107 | n33675 ;
  assign n33677 = n7173 ^ n3216 ^ 1'b0 ;
  assign n33678 = n3393 | n33677 ;
  assign n33679 = n10449 & n10577 ;
  assign n33680 = n33679 ^ n1419 ^ 1'b0 ;
  assign n33681 = n10373 & n30444 ;
  assign n33682 = ~n25440 & n32957 ;
  assign n33683 = ~n3755 & n33682 ;
  assign n33684 = n27507 ^ n19810 ^ 1'b0 ;
  assign n33685 = n6992 & n17839 ;
  assign n33686 = n6612 & n33685 ;
  assign n33688 = n27444 ^ n22556 ^ 1'b0 ;
  assign n33689 = n33688 ^ n12235 ^ 1'b0 ;
  assign n33687 = n22556 & ~n30820 ;
  assign n33690 = n33689 ^ n33687 ^ 1'b0 ;
  assign n33691 = n12218 ^ n10884 ^ 1'b0 ;
  assign n33692 = ~n2661 & n33691 ;
  assign n33693 = n11287 & ~n16471 ;
  assign n33694 = ~n17923 & n18700 ;
  assign n33695 = n6700 & n10510 ;
  assign n33696 = n33695 ^ n15022 ^ 1'b0 ;
  assign n33697 = n18548 ^ n11265 ^ 1'b0 ;
  assign n33698 = n33696 & n33697 ;
  assign n33699 = n33698 ^ n8566 ^ 1'b0 ;
  assign n33700 = n5997 & n7788 ;
  assign n33701 = n25305 & ~n33111 ;
  assign n33702 = n21868 ^ n17717 ^ 1'b0 ;
  assign n33703 = ~n13407 & n33702 ;
  assign n33704 = n1148 & ~n6612 ;
  assign n33705 = ~n6122 & n33704 ;
  assign n33706 = ~n3934 & n33705 ;
  assign n33707 = ( n11799 & n17987 ) | ( n11799 & n21516 ) | ( n17987 & n21516 ) ;
  assign n33712 = ~n9683 & n19813 ;
  assign n33713 = n3386 & n33712 ;
  assign n33708 = n1588 & n7301 ;
  assign n33709 = ~n4964 & n33708 ;
  assign n33710 = n33709 ^ n21843 ^ 1'b0 ;
  assign n33711 = n11155 & ~n33710 ;
  assign n33714 = n33713 ^ n33711 ^ n711 ;
  assign n33715 = n5720 & n17488 ;
  assign n33716 = n33714 & n33715 ;
  assign n33717 = n13084 & ~n33716 ;
  assign n33718 = n2170 ^ x181 ^ 1'b0 ;
  assign n33719 = n11204 & ~n33718 ;
  assign n33720 = n14740 | n31870 ;
  assign n33721 = n24640 & ~n28125 ;
  assign n33722 = ~n17308 & n20702 ;
  assign n33723 = n26553 & ~n33722 ;
  assign n33724 = ~n1382 & n3929 ;
  assign n33725 = n33724 ^ n19719 ^ 1'b0 ;
  assign n33726 = n14617 & n33725 ;
  assign n33727 = n6436 & n33726 ;
  assign n33728 = n1919 & ~n5665 ;
  assign n33729 = ~n1919 & n33728 ;
  assign n33730 = x112 & ~n10564 ;
  assign n33731 = n33730 ^ n12708 ^ 1'b0 ;
  assign n33732 = ~n7550 & n33731 ;
  assign n33733 = n29926 ^ n14640 ^ 1'b0 ;
  assign n33734 = ~n1876 & n33733 ;
  assign n33735 = n31643 ^ n17278 ^ 1'b0 ;
  assign n33736 = n530 & ~n33735 ;
  assign n33737 = n16398 ^ n4426 ^ 1'b0 ;
  assign n33739 = n14529 | n29403 ;
  assign n33738 = n12169 | n29855 ;
  assign n33740 = n33739 ^ n33738 ^ 1'b0 ;
  assign n33741 = n27187 ^ n18358 ^ 1'b0 ;
  assign n33742 = n25229 ^ n11903 ^ 1'b0 ;
  assign n33743 = n23020 | n33742 ;
  assign n33744 = ~n5145 & n20160 ;
  assign n33745 = n33260 ^ n28953 ^ n20891 ;
  assign n33746 = n11091 ^ n5725 ^ 1'b0 ;
  assign n33747 = n5690 ^ n954 ^ 1'b0 ;
  assign n33748 = n16267 ^ n876 ^ 1'b0 ;
  assign n33749 = n33747 & n33748 ;
  assign n33750 = ( n24498 & n33746 ) | ( n24498 & n33749 ) | ( n33746 & n33749 ) ;
  assign n33751 = n33750 ^ n5315 ^ 1'b0 ;
  assign n33758 = n30537 ^ n18362 ^ 1'b0 ;
  assign n33752 = n6769 & ~n6798 ;
  assign n33753 = n5554 ^ n938 ^ 1'b0 ;
  assign n33754 = n33752 & n33753 ;
  assign n33755 = ~n22607 & n33754 ;
  assign n33756 = ~n12326 & n33755 ;
  assign n33757 = n20794 | n33756 ;
  assign n33759 = n33758 ^ n33757 ^ 1'b0 ;
  assign n33760 = x188 & ~n33158 ;
  assign n33761 = n33760 ^ n29904 ^ 1'b0 ;
  assign n33762 = n33761 ^ x203 ^ 1'b0 ;
  assign n33763 = n3335 | n11819 ;
  assign n33764 = ( n5043 & n11430 ) | ( n5043 & n33501 ) | ( n11430 & n33501 ) ;
  assign n33765 = n33764 ^ n29397 ^ 1'b0 ;
  assign n33766 = ~n6951 & n33765 ;
  assign n33767 = n1954 | n8250 ;
  assign n33768 = n33767 ^ n3536 ^ 1'b0 ;
  assign n33769 = n14857 & n22053 ;
  assign n33770 = ~n8231 & n13158 ;
  assign n33771 = n7310 & n33770 ;
  assign n33772 = n33769 & ~n33771 ;
  assign n33773 = n22909 & n33772 ;
  assign n33774 = n11600 | n15449 ;
  assign n33775 = n1718 | n20413 ;
  assign n33776 = n3082 & ~n33775 ;
  assign n33777 = n13650 | n33776 ;
  assign n33778 = n393 & ~n33777 ;
  assign n33779 = ~n5511 & n9959 ;
  assign n33780 = n2458 & n33779 ;
  assign n33781 = n33780 ^ n13444 ^ 1'b0 ;
  assign n33782 = n24977 ^ n9495 ^ 1'b0 ;
  assign n33783 = n4325 & n33782 ;
  assign n33784 = n663 & ~n24936 ;
  assign n33785 = n3805 & ~n33784 ;
  assign n33786 = n33785 ^ n3351 ^ 1'b0 ;
  assign n33787 = n16697 ^ n16231 ^ 1'b0 ;
  assign n33788 = ( ~n2228 & n5732 ) | ( ~n2228 & n26341 ) | ( n5732 & n26341 ) ;
  assign n33789 = ~n6008 & n33788 ;
  assign n33790 = n33789 ^ n15594 ^ 1'b0 ;
  assign n33791 = n2580 & n23280 ;
  assign n33792 = n28687 ^ n27353 ^ 1'b0 ;
  assign n33793 = n10170 | n23755 ;
  assign n33794 = n17695 & ~n33793 ;
  assign n33797 = n11880 ^ n6734 ^ 1'b0 ;
  assign n33795 = ~n11705 & n15259 ;
  assign n33796 = n26939 & n33795 ;
  assign n33798 = n33797 ^ n33796 ^ 1'b0 ;
  assign n33799 = n1217 & ~n27494 ;
  assign n33800 = ~n1049 & n9499 ;
  assign n33801 = n33152 ^ n2580 ^ 1'b0 ;
  assign n33802 = n33801 ^ n17452 ^ 1'b0 ;
  assign n33803 = n33800 & n33802 ;
  assign n33804 = ~n33626 & n33803 ;
  assign n33805 = n3412 ^ n2982 ^ 1'b0 ;
  assign n33806 = n33805 ^ n14239 ^ n13061 ;
  assign n33807 = ( x57 & n19328 ) | ( x57 & ~n33806 ) | ( n19328 & ~n33806 ) ;
  assign n33808 = n16608 ^ x207 ^ 1'b0 ;
  assign n33809 = n5474 & n33808 ;
  assign n33810 = n33809 ^ n3370 ^ 1'b0 ;
  assign n33811 = n6259 & ~n11353 ;
  assign n33812 = n13409 & ~n29686 ;
  assign n33813 = n33812 ^ n21304 ^ 1'b0 ;
  assign n33814 = n24858 ^ n10860 ^ 1'b0 ;
  assign n33815 = n1850 & ~n7118 ;
  assign n33816 = ~n27689 & n33815 ;
  assign n33817 = n9534 | n13849 ;
  assign n33818 = n17889 & ~n26272 ;
  assign n33819 = n33817 & n33818 ;
  assign n33821 = n24376 ^ n13183 ^ 1'b0 ;
  assign n33820 = n20997 & n31308 ;
  assign n33822 = n33821 ^ n33820 ^ 1'b0 ;
  assign n33823 = n4256 & ~n10852 ;
  assign n33824 = n33823 ^ n7328 ^ 1'b0 ;
  assign n33825 = n33824 ^ n30984 ^ 1'b0 ;
  assign n33826 = n9175 & n11503 ;
  assign n33827 = n10353 & n11458 ;
  assign n33828 = ~n16710 & n33827 ;
  assign n33829 = n6361 | n33828 ;
  assign n33831 = x248 & ~n913 ;
  assign n33832 = n913 & n33831 ;
  assign n33833 = n15308 | n33832 ;
  assign n33834 = ~n3986 & n33833 ;
  assign n33835 = n33834 ^ x105 ^ 1'b0 ;
  assign n33830 = n24290 ^ n22156 ^ n6383 ;
  assign n33836 = n33835 ^ n33830 ^ 1'b0 ;
  assign n33837 = n16627 ^ n8249 ^ 1'b0 ;
  assign n33838 = ( n6025 & n9157 ) | ( n6025 & ~n29602 ) | ( n9157 & ~n29602 ) ;
  assign n33842 = n8547 ^ n7579 ^ 1'b0 ;
  assign n33843 = n5418 | n33842 ;
  assign n33839 = n27482 ^ n16719 ^ 1'b0 ;
  assign n33840 = n8571 | n33839 ;
  assign n33841 = n33190 | n33840 ;
  assign n33844 = n33843 ^ n33841 ^ 1'b0 ;
  assign n33845 = n13472 | n19032 ;
  assign n33846 = n33845 ^ n18008 ^ 1'b0 ;
  assign n33847 = n30301 & n33846 ;
  assign n33848 = ~n14679 & n33847 ;
  assign n33849 = n7220 ^ x112 ^ 1'b0 ;
  assign n33850 = n7899 & ~n33849 ;
  assign n33851 = n33850 ^ n13127 ^ 1'b0 ;
  assign n33852 = n13443 ^ n4522 ^ 1'b0 ;
  assign n33853 = n4708 & n33852 ;
  assign n33854 = n12230 & ~n33853 ;
  assign n33855 = n19528 ^ n14695 ^ 1'b0 ;
  assign n33856 = n6300 & n33204 ;
  assign n33857 = ~n33855 & n33856 ;
  assign n33858 = n7315 & n15975 ;
  assign n33859 = n24625 & n33858 ;
  assign n33860 = n15269 & ~n33859 ;
  assign n33861 = n33860 ^ n9714 ^ 1'b0 ;
  assign n33862 = ~n4608 & n25499 ;
  assign n33863 = n4027 | n5354 ;
  assign n33864 = ~n2155 & n33863 ;
  assign n33865 = ~n10682 & n28838 ;
  assign n33866 = ( n794 & n1219 ) | ( n794 & n11762 ) | ( n1219 & n11762 ) ;
  assign n33867 = ~n6431 & n9027 ;
  assign n33868 = n1786 & n5975 ;
  assign n33869 = n33867 | n33868 ;
  assign n33870 = n33866 | n33869 ;
  assign n33871 = n33454 ^ n27600 ^ 1'b0 ;
  assign n33872 = n33870 & n33871 ;
  assign n33873 = n4259 & n4465 ;
  assign n33874 = ~n33872 & n33873 ;
  assign n33876 = n26656 ^ x166 ^ 1'b0 ;
  assign n33875 = n6524 & n19533 ;
  assign n33877 = n33876 ^ n33875 ^ 1'b0 ;
  assign n33878 = n17370 ^ n9876 ^ 1'b0 ;
  assign n33879 = n5810 | n33878 ;
  assign n33880 = n33879 ^ n5296 ^ n886 ;
  assign n33881 = n7141 & n26905 ;
  assign n33882 = n25134 & n33881 ;
  assign n33883 = n33414 ^ n26780 ^ 1'b0 ;
  assign n33884 = n18164 | n32730 ;
  assign n33885 = n33884 ^ n20708 ^ 1'b0 ;
  assign n33886 = n26118 & ~n33885 ;
  assign n33887 = n2177 | n4864 ;
  assign n33888 = n33887 ^ n14429 ^ 1'b0 ;
  assign n33889 = n12676 ^ n8277 ^ n4714 ;
  assign n33890 = n17341 ^ n5984 ^ n4290 ;
  assign n33891 = n7183 | n17336 ;
  assign n33892 = n2252 & ~n33891 ;
  assign n33893 = n22043 ^ n13757 ^ 1'b0 ;
  assign n33894 = n33892 | n33893 ;
  assign n33895 = n13737 & n33894 ;
  assign n33896 = n4711 & n8745 ;
  assign n33897 = ~n5769 & n33896 ;
  assign n33898 = ~n9560 & n33897 ;
  assign n33899 = n14240 & n33898 ;
  assign n33900 = n11879 ^ n2960 ^ n2004 ;
  assign n33901 = ~n9694 & n33900 ;
  assign n33902 = ~n11669 & n33901 ;
  assign n33903 = x160 & ~n1254 ;
  assign n33904 = n1254 & n33903 ;
  assign n33905 = n21347 | n33904 ;
  assign n33906 = n7651 | n33905 ;
  assign n33907 = n4282 & ~n33906 ;
  assign n33908 = n13571 | n13776 ;
  assign n33909 = n15191 & ~n33908 ;
  assign n33910 = n33909 ^ n20816 ^ 1'b0 ;
  assign n33911 = n33907 | n33910 ;
  assign n33912 = n15366 & ~n21694 ;
  assign n33913 = n33912 ^ n14777 ^ 1'b0 ;
  assign n33914 = n15515 & ~n33913 ;
  assign n33915 = ( ~n5235 & n27698 ) | ( ~n5235 & n32331 ) | ( n27698 & n32331 ) ;
  assign n33916 = n4366 & ~n8365 ;
  assign n33917 = n15617 & ~n23068 ;
  assign n33918 = n33917 ^ n24602 ^ 1'b0 ;
  assign n33919 = n5988 & n33918 ;
  assign n33920 = n25762 & ~n27509 ;
  assign n33921 = ~n8785 & n33804 ;
  assign n33922 = n2055 | n6400 ;
  assign n33923 = n33922 ^ n11819 ^ 1'b0 ;
  assign n33924 = ~n3900 & n33923 ;
  assign n33925 = n26601 & n33924 ;
  assign n33927 = n17052 & n23780 ;
  assign n33926 = ~n6269 & n24695 ;
  assign n33928 = n33927 ^ n33926 ^ 1'b0 ;
  assign n33929 = n33731 ^ n26612 ^ 1'b0 ;
  assign n33930 = n3805 & ~n12224 ;
  assign n33931 = n33930 ^ n862 ^ 1'b0 ;
  assign n33932 = ( ~n4237 & n8566 ) | ( ~n4237 & n33931 ) | ( n8566 & n33931 ) ;
  assign n33933 = n29511 ^ n26930 ^ 1'b0 ;
  assign n33934 = ~n520 & n11747 ;
  assign n33935 = n15973 & ~n33934 ;
  assign n33936 = ~n3496 & n33935 ;
  assign n33937 = n6966 ^ n4809 ^ 1'b0 ;
  assign n33938 = n23110 | n33937 ;
  assign n33939 = n378 & ~n33938 ;
  assign n33940 = n13047 ^ n7689 ^ n975 ;
  assign n33941 = ~n2098 & n2606 ;
  assign n33942 = n33940 & n33941 ;
  assign n33943 = n28604 ^ n2193 ^ 1'b0 ;
  assign n33944 = n9099 & ~n33943 ;
  assign n33945 = n33944 ^ n6627 ^ 1'b0 ;
  assign n33946 = n3265 & ~n7119 ;
  assign n33947 = n15840 & n33946 ;
  assign n33948 = ~x82 & n33947 ;
  assign n33949 = n1758 | n8233 ;
  assign n33950 = n1487 & ~n33949 ;
  assign n33951 = n738 | n33950 ;
  assign n33952 = ~n21046 & n21164 ;
  assign n33953 = n33952 ^ n28544 ^ n2120 ;
  assign n33954 = n15889 ^ n3342 ^ 1'b0 ;
  assign n33955 = n5913 ^ n501 ^ 1'b0 ;
  assign n33956 = n23174 ^ n7130 ^ 1'b0 ;
  assign n33957 = n33955 & ~n33956 ;
  assign n33958 = ~n11142 & n23396 ;
  assign n33959 = ~n33957 & n33958 ;
  assign n33960 = n24286 | n28795 ;
  assign n33961 = n17676 & ~n33960 ;
  assign n33962 = n33961 ^ n11650 ^ 1'b0 ;
  assign n33963 = ~n675 & n33962 ;
  assign n33964 = n17805 & ~n28830 ;
  assign n33965 = n33964 ^ n624 ^ 1'b0 ;
  assign n33966 = n1383 & n33965 ;
  assign n33967 = ~n15263 & n33966 ;
  assign n33968 = ~n16045 & n33967 ;
  assign n33969 = n25551 & n33968 ;
  assign n33971 = n16204 ^ n5116 ^ 1'b0 ;
  assign n33972 = x200 & ~n33971 ;
  assign n33970 = n9674 | n22095 ;
  assign n33973 = n33972 ^ n33970 ^ 1'b0 ;
  assign n33974 = x80 & n794 ;
  assign n33975 = n4962 & n33974 ;
  assign n33976 = n27434 ^ n9603 ^ 1'b0 ;
  assign n33977 = n33975 | n33976 ;
  assign n33978 = n14440 ^ n11201 ^ 1'b0 ;
  assign n33979 = n30129 & n33978 ;
  assign n33980 = n33979 ^ n12650 ^ 1'b0 ;
  assign n33981 = n8325 ^ n6429 ^ 1'b0 ;
  assign n33982 = n1151 & n33981 ;
  assign n33983 = n15930 & n29003 ;
  assign n33984 = n1784 & n33983 ;
  assign n33985 = n7387 & n33984 ;
  assign n33986 = n7734 & n18673 ;
  assign n33987 = n33986 ^ n2369 ^ 1'b0 ;
  assign n33988 = n33987 ^ n4589 ^ 1'b0 ;
  assign n33989 = n7629 & ~n24073 ;
  assign n33990 = n33989 ^ n21045 ^ 1'b0 ;
  assign n33991 = n33990 ^ x112 ^ 1'b0 ;
  assign n33992 = n10586 | n17040 ;
  assign n33993 = ~n9886 & n12418 ;
  assign n33994 = ~n12551 & n33993 ;
  assign n33995 = ( ~n1028 & n3861 ) | ( ~n1028 & n5438 ) | ( n3861 & n5438 ) ;
  assign n33996 = n3329 | n18163 ;
  assign n33997 = n33995 & ~n33996 ;
  assign n33998 = ~n30781 & n33997 ;
  assign n33999 = ~n10483 & n10508 ;
  assign n34000 = ~n5478 & n33999 ;
  assign n34001 = n33769 ^ n6640 ^ 1'b0 ;
  assign n34002 = ~n34000 & n34001 ;
  assign n34003 = n14240 ^ n10731 ^ 1'b0 ;
  assign n34004 = n5720 & n34003 ;
  assign n34005 = n25307 & n34004 ;
  assign n34006 = n15230 & n34005 ;
  assign n34007 = ( n4150 & n4927 ) | ( n4150 & ~n5911 ) | ( n4927 & ~n5911 ) ;
  assign n34008 = n11807 & ~n34007 ;
  assign n34009 = n7495 & ~n31754 ;
  assign n34010 = n34009 ^ n17251 ^ 1'b0 ;
  assign n34011 = n23572 ^ n14229 ^ 1'b0 ;
  assign n34012 = n13392 & ~n34011 ;
  assign n34013 = n34012 ^ n17827 ^ 1'b0 ;
  assign n34014 = n34010 & n34013 ;
  assign n34015 = ~n305 & n1020 ;
  assign n34016 = ~n15010 & n28586 ;
  assign n34017 = ~n1956 & n3323 ;
  assign n34018 = n32793 ^ n10382 ^ 1'b0 ;
  assign n34019 = n14471 & ~n34018 ;
  assign n34020 = n4652 & ~n32876 ;
  assign n34021 = n27852 & n30581 ;
  assign n34026 = n21100 ^ n6053 ^ 1'b0 ;
  assign n34027 = n2715 | n19310 ;
  assign n34028 = ( n9741 & ~n34026 ) | ( n9741 & n34027 ) | ( ~n34026 & n34027 ) ;
  assign n34022 = n3408 | n25319 ;
  assign n34023 = n34022 ^ n7522 ^ 1'b0 ;
  assign n34024 = n34023 ^ n12439 ^ 1'b0 ;
  assign n34025 = n17859 | n34024 ;
  assign n34029 = n34028 ^ n34025 ^ 1'b0 ;
  assign n34030 = n5398 | n16813 ;
  assign n34031 = n26087 ^ n25359 ^ 1'b0 ;
  assign n34032 = n13026 & n34031 ;
  assign n34033 = ~n4553 & n8336 ;
  assign n34034 = n34033 ^ n7727 ^ n2375 ;
  assign n34035 = n3412 & ~n34034 ;
  assign n34036 = x184 & n34035 ;
  assign n34037 = n13624 & ~n15338 ;
  assign n34038 = n19195 ^ n2439 ^ n1595 ;
  assign n34039 = n9974 & ~n21520 ;
  assign n34040 = ~n26950 & n34039 ;
  assign n34041 = n11963 & ~n20529 ;
  assign n34042 = n34041 ^ n14723 ^ 1'b0 ;
  assign n34043 = n8520 | n30400 ;
  assign n34044 = n18482 & ~n29627 ;
  assign n34045 = n34043 & n34044 ;
  assign n34046 = n29267 ^ n7907 ^ 1'b0 ;
  assign n34047 = ~n21135 & n22660 ;
  assign n34048 = n29061 & n34047 ;
  assign n34049 = n5163 & n12632 ;
  assign n34050 = ( ~n4555 & n31264 ) | ( ~n4555 & n34049 ) | ( n31264 & n34049 ) ;
  assign n34051 = ( x3 & ~x191 ) | ( x3 & n4242 ) | ( ~x191 & n4242 ) ;
  assign n34052 = n34051 ^ n12471 ^ 1'b0 ;
  assign n34053 = n34052 ^ n2752 ^ 1'b0 ;
  assign n34055 = n28586 ^ n15479 ^ 1'b0 ;
  assign n34056 = ~n21114 & n34055 ;
  assign n34054 = n21201 ^ x116 ^ 1'b0 ;
  assign n34057 = n34056 ^ n34054 ^ 1'b0 ;
  assign n34058 = ~n4662 & n34057 ;
  assign n34059 = n34058 ^ n17406 ^ 1'b0 ;
  assign n34060 = ~n1473 & n15490 ;
  assign n34061 = ~n638 & n16481 ;
  assign n34062 = ~n19986 & n34061 ;
  assign n34063 = n7530 ^ n4835 ^ 1'b0 ;
  assign n34064 = n13171 & ~n17183 ;
  assign n34065 = n34064 ^ n1550 ^ 1'b0 ;
  assign n34066 = n26179 ^ n25151 ^ 1'b0 ;
  assign n34067 = n25029 | n34066 ;
  assign n34068 = n21695 ^ n18889 ^ 1'b0 ;
  assign n34069 = n26056 & ~n34068 ;
  assign n34070 = n29364 ^ n21090 ^ 1'b0 ;
  assign n34071 = n34069 | n34070 ;
  assign n34072 = n34071 ^ n3806 ^ 1'b0 ;
  assign n34073 = ~n3753 & n3796 ;
  assign n34074 = n34072 & n34073 ;
  assign n34075 = ~n296 & n11146 ;
  assign n34076 = n34075 ^ n9578 ^ 1'b0 ;
  assign n34077 = ~n31686 & n34076 ;
  assign n34078 = n4567 & n30475 ;
  assign n34079 = n19545 | n20853 ;
  assign n34080 = n2247 | n34079 ;
  assign n34081 = n9865 | n10689 ;
  assign n34082 = n29650 & n34081 ;
  assign n34083 = n11333 ^ n10851 ^ 1'b0 ;
  assign n34084 = ~n31070 & n34083 ;
  assign n34085 = ~n4622 & n8287 ;
  assign n34086 = n34085 ^ n14488 ^ 1'b0 ;
  assign n34087 = n2356 & ~n5876 ;
  assign n34088 = n11874 | n28740 ;
  assign n34089 = ~n4565 & n34088 ;
  assign n34090 = n23672 ^ n5613 ^ 1'b0 ;
  assign n34091 = n23055 | n34090 ;
  assign n34092 = n5959 ^ n4222 ^ 1'b0 ;
  assign n34093 = ~n3078 & n22053 ;
  assign n34094 = n34092 & n34093 ;
  assign n34095 = n34094 ^ n25640 ^ 1'b0 ;
  assign n34096 = n20772 & n22879 ;
  assign n34097 = n22173 & n34096 ;
  assign n34098 = n5598 & ~n34097 ;
  assign n34099 = n21434 | n31093 ;
  assign n34100 = n31580 ^ n7850 ^ 1'b0 ;
  assign n34101 = n34099 & n34100 ;
  assign n34102 = n33651 ^ n31551 ^ 1'b0 ;
  assign n34103 = n8353 & ~n34102 ;
  assign n34104 = n10835 | n12195 ;
  assign n34105 = n2487 & ~n33496 ;
  assign n34106 = n17093 ^ n14507 ^ 1'b0 ;
  assign n34107 = n34105 | n34106 ;
  assign n34108 = n6731 & ~n34107 ;
  assign n34109 = n19064 & n22615 ;
  assign n34110 = ( ~n2406 & n15037 ) | ( ~n2406 & n15854 ) | ( n15037 & n15854 ) ;
  assign n34111 = n5576 & ~n25492 ;
  assign n34112 = n3704 | n8892 ;
  assign n34113 = n4239 & n34112 ;
  assign n34114 = n708 & n11211 ;
  assign n34115 = ~n5382 & n19752 ;
  assign n34116 = ( n8684 & ~n18513 ) | ( n8684 & n19038 ) | ( ~n18513 & n19038 ) ;
  assign n34117 = n24941 ^ n22998 ^ n6868 ;
  assign n34118 = n34116 & n34117 ;
  assign n34119 = n34115 & n34118 ;
  assign n34120 = n15282 ^ n9788 ^ n2180 ;
  assign n34121 = n19336 & ~n34120 ;
  assign n34122 = ( n906 & n17388 ) | ( n906 & n33769 ) | ( n17388 & n33769 ) ;
  assign n34123 = n31984 ^ n19016 ^ 1'b0 ;
  assign n34124 = n8764 & ~n34123 ;
  assign n34125 = n23872 ^ n14912 ^ 1'b0 ;
  assign n34126 = n518 | n14595 ;
  assign n34127 = n34126 ^ n2420 ^ 1'b0 ;
  assign n34128 = n4838 & n34127 ;
  assign n34129 = ~n32671 & n34128 ;
  assign n34130 = n3944 ^ n2484 ^ 1'b0 ;
  assign n34131 = n6476 & n34130 ;
  assign n34132 = n34131 ^ n6406 ^ 1'b0 ;
  assign n34133 = n34129 | n34132 ;
  assign n34134 = n1353 | n20315 ;
  assign n34135 = n34134 ^ n23902 ^ n17141 ;
  assign n34137 = n2877 | n12513 ;
  assign n34136 = n10867 & ~n18688 ;
  assign n34138 = n34137 ^ n34136 ^ 1'b0 ;
  assign n34139 = n2564 & ~n19244 ;
  assign n34140 = n21129 & n34139 ;
  assign n34141 = ( n11571 & n34138 ) | ( n11571 & n34140 ) | ( n34138 & n34140 ) ;
  assign n34142 = n4932 | n15275 ;
  assign n34144 = n17536 | n21808 ;
  assign n34145 = n10187 & ~n34144 ;
  assign n34143 = n1973 & ~n9180 ;
  assign n34146 = n34145 ^ n34143 ^ 1'b0 ;
  assign n34147 = n2647 & ~n27433 ;
  assign n34148 = n5650 & n34147 ;
  assign n34149 = n34148 ^ x241 ^ 1'b0 ;
  assign n34150 = ~n34146 & n34149 ;
  assign n34151 = n6629 & n8308 ;
  assign n34152 = n13433 & ~n34151 ;
  assign n34153 = n8762 & n32150 ;
  assign n34154 = n34153 ^ n17047 ^ 1'b0 ;
  assign n34155 = ~n10797 & n15614 ;
  assign n34156 = ~n32028 & n34155 ;
  assign n34157 = ~n11034 & n33946 ;
  assign n34158 = n1069 & n34157 ;
  assign n34159 = n2319 & ~n26488 ;
  assign n34162 = x27 & n29938 ;
  assign n34160 = ~n8164 & n11472 ;
  assign n34161 = ~n18715 & n34160 ;
  assign n34163 = n34162 ^ n34161 ^ 1'b0 ;
  assign n34164 = n12197 | n31920 ;
  assign n34165 = n27029 | n34164 ;
  assign n34166 = n19536 | n20598 ;
  assign n34167 = n12338 & ~n34166 ;
  assign n34168 = n34167 ^ x6 ^ 1'b0 ;
  assign n34169 = n15026 & ~n19946 ;
  assign n34170 = n34168 & n34169 ;
  assign n34172 = n14516 & n23602 ;
  assign n34171 = n24612 & ~n34046 ;
  assign n34173 = n34172 ^ n34171 ^ 1'b0 ;
  assign n34174 = n5422 & ~n21824 ;
  assign n34176 = n12621 & n26521 ;
  assign n34175 = n6719 & n8301 ;
  assign n34177 = n34176 ^ n34175 ^ n29587 ;
  assign n34178 = x31 & n1833 ;
  assign n34179 = x207 | n2144 ;
  assign n34180 = n12564 & ~n26369 ;
  assign n34181 = n33555 ^ n25450 ^ 1'b0 ;
  assign n34182 = ~n5328 & n34181 ;
  assign n34183 = n34182 ^ n6404 ^ 1'b0 ;
  assign n34184 = ~n3935 & n20653 ;
  assign n34185 = n34184 ^ n15992 ^ n3985 ;
  assign n34186 = ~n20614 & n34185 ;
  assign n34187 = ~n3594 & n34186 ;
  assign n34188 = n5422 | n17910 ;
  assign n34189 = n34188 ^ n27035 ^ 1'b0 ;
  assign n34190 = n7783 & ~n15652 ;
  assign n34191 = n34190 ^ n9720 ^ 1'b0 ;
  assign n34192 = n34191 ^ n16693 ^ 1'b0 ;
  assign n34193 = ( n5569 & ~n8725 ) | ( n5569 & n34192 ) | ( ~n8725 & n34192 ) ;
  assign n34194 = n14742 & n20644 ;
  assign n34195 = n4169 & n34194 ;
  assign n34196 = n34195 ^ n2615 ^ 1'b0 ;
  assign n34197 = ~n13122 & n34196 ;
  assign n34198 = n34197 ^ n19002 ^ 1'b0 ;
  assign n34199 = n4934 & ~n5862 ;
  assign n34200 = n34199 ^ n26125 ^ 1'b0 ;
  assign n34201 = n20214 ^ n5573 ^ 1'b0 ;
  assign n34202 = ~n3267 & n32793 ;
  assign n34203 = n10003 & ~n29065 ;
  assign n34204 = ~x181 & n34203 ;
  assign n34205 = n28627 & ~n34204 ;
  assign n34206 = n15680 & n21249 ;
  assign n34207 = n4824 & n14755 ;
  assign n34208 = n34207 ^ n20348 ^ n13981 ;
  assign n34209 = ~n1757 & n17889 ;
  assign n34210 = ~n6441 & n18168 ;
  assign n34213 = n15089 & ~n29480 ;
  assign n34211 = n31063 ^ n4725 ^ 1'b0 ;
  assign n34212 = ~n32541 & n34211 ;
  assign n34214 = n34213 ^ n34212 ^ 1'b0 ;
  assign n34215 = n24751 ^ n8728 ^ n1573 ;
  assign n34216 = ~n4821 & n34215 ;
  assign n34217 = n34216 ^ n3683 ^ 1'b0 ;
  assign n34218 = n4788 & ~n30493 ;
  assign n34219 = ~n5292 & n34218 ;
  assign n34222 = ~n15510 & n16872 ;
  assign n34223 = n19562 & n34222 ;
  assign n34220 = n5509 & n8863 ;
  assign n34221 = ~n14435 & n34220 ;
  assign n34224 = n34223 ^ n34221 ^ n19172 ;
  assign n34225 = ( n8900 & ~n10455 ) | ( n8900 & n30328 ) | ( ~n10455 & n30328 ) ;
  assign n34230 = ~n2178 & n5616 ;
  assign n34231 = n34230 ^ n4423 ^ 1'b0 ;
  assign n34232 = n7093 | n34231 ;
  assign n34233 = n1333 & ~n34232 ;
  assign n34226 = n3946 | n18420 ;
  assign n34227 = n16061 ^ n1950 ^ 1'b0 ;
  assign n34228 = n34226 & n34227 ;
  assign n34229 = ~n8816 & n34228 ;
  assign n34234 = n34233 ^ n34229 ^ 1'b0 ;
  assign n34235 = n6985 ^ n3286 ^ 1'b0 ;
  assign n34236 = n4363 & ~n34235 ;
  assign n34237 = n34236 ^ n12488 ^ 1'b0 ;
  assign n34238 = n34237 ^ n12029 ^ 1'b0 ;
  assign n34239 = n9703 & ~n16145 ;
  assign n34240 = n34239 ^ n6144 ^ 1'b0 ;
  assign n34241 = n17717 ^ n10992 ^ 1'b0 ;
  assign n34242 = n34240 & n34241 ;
  assign n34243 = n25467 & ~n30283 ;
  assign n34244 = n3884 & n34243 ;
  assign n34245 = ~n13585 & n13691 ;
  assign n34246 = ~x123 & n28442 ;
  assign n34247 = n34245 & n34246 ;
  assign n34248 = n7414 | n18281 ;
  assign n34249 = n29002 ^ n26606 ^ n25272 ;
  assign n34250 = x0 & n18265 ;
  assign n34251 = n34250 ^ n5610 ^ 1'b0 ;
  assign n34252 = n4417 & ~n16428 ;
  assign n34253 = n4880 & ~n9114 ;
  assign n34254 = n6565 ^ n4502 ^ 1'b0 ;
  assign n34255 = ( n1185 & n9628 ) | ( n1185 & n12792 ) | ( n9628 & n12792 ) ;
  assign n34256 = n7948 | n16466 ;
  assign n34257 = n34256 ^ n15950 ^ 1'b0 ;
  assign n34258 = n15785 ^ n558 ^ 1'b0 ;
  assign n34259 = n34257 & ~n34258 ;
  assign n34260 = n16818 ^ n7908 ^ 1'b0 ;
  assign n34261 = n3279 | n34260 ;
  assign n34262 = n5051 ^ n3272 ^ 1'b0 ;
  assign n34263 = n3440 & n34262 ;
  assign n34264 = ~n34261 & n34263 ;
  assign n34265 = n31152 ^ n16675 ^ 1'b0 ;
  assign n34266 = n22641 & n34265 ;
  assign n34267 = n34266 ^ n18221 ^ n3124 ;
  assign n34268 = n680 & n8191 ;
  assign n34269 = n31603 & n34268 ;
  assign n34270 = n5961 & n34269 ;
  assign n34271 = ( x128 & n27604 ) | ( x128 & n34270 ) | ( n27604 & n34270 ) ;
  assign n34272 = ~n20033 & n28305 ;
  assign n34273 = n453 & n29439 ;
  assign n34274 = ~n34272 & n34273 ;
  assign n34275 = n8103 ^ n4788 ^ 1'b0 ;
  assign n34276 = n20998 & n34275 ;
  assign n34277 = n8225 | n28265 ;
  assign n34278 = n34007 & ~n34277 ;
  assign n34279 = n8375 ^ n1569 ^ 1'b0 ;
  assign n34280 = ~n34278 & n34279 ;
  assign n34281 = x56 & ~n5445 ;
  assign n34282 = n34281 ^ n1805 ^ 1'b0 ;
  assign n34283 = ~n11416 & n34282 ;
  assign n34284 = ~n2638 & n6989 ;
  assign n34285 = n11024 & n34284 ;
  assign n34286 = n31294 & ~n34285 ;
  assign n34287 = ~n3000 & n4983 ;
  assign n34288 = ~n25659 & n34287 ;
  assign n34291 = ~n9889 & n17202 ;
  assign n34292 = n1204 & n34291 ;
  assign n34289 = ( ~n11908 & n23904 ) | ( ~n11908 & n24627 ) | ( n23904 & n24627 ) ;
  assign n34290 = n19812 & ~n34289 ;
  assign n34293 = n34292 ^ n34290 ^ 1'b0 ;
  assign n34294 = ~n15385 & n26302 ;
  assign n34295 = n15637 ^ n6603 ^ 1'b0 ;
  assign n34296 = ~n1220 & n3216 ;
  assign n34297 = n34296 ^ n1185 ^ 1'b0 ;
  assign n34298 = n2297 | n28258 ;
  assign n34299 = n34297 | n34298 ;
  assign n34300 = n34299 ^ n18221 ^ n17155 ;
  assign n34301 = n25715 ^ n14510 ^ 1'b0 ;
  assign n34302 = n5782 ^ n1435 ^ 1'b0 ;
  assign n34303 = n9540 | n34302 ;
  assign n34304 = n34303 ^ n17929 ^ n2055 ;
  assign n34305 = n3579 | n4338 ;
  assign n34306 = n10926 & ~n34305 ;
  assign n34307 = n34306 ^ n23313 ^ 1'b0 ;
  assign n34308 = n34307 ^ n18791 ^ n3951 ;
  assign n34309 = n17932 ^ n963 ^ 1'b0 ;
  assign n34310 = n13631 ^ n8578 ^ 1'b0 ;
  assign n34311 = n3316 | n23726 ;
  assign n34312 = n30756 & ~n34311 ;
  assign n34313 = n33965 ^ n13339 ^ n1503 ;
  assign n34314 = n34313 ^ n877 ^ 1'b0 ;
  assign n34315 = n2535 & ~n34314 ;
  assign n34316 = ~n7464 & n18096 ;
  assign n34317 = n34316 ^ n13028 ^ 1'b0 ;
  assign n34318 = n14845 & n34317 ;
  assign n34319 = n11237 | n25334 ;
  assign n34320 = n34318 | n34319 ;
  assign n34321 = n30101 ^ n23017 ^ n1495 ;
  assign n34322 = ~n9267 & n12113 ;
  assign n34323 = n34322 ^ n17842 ^ 1'b0 ;
  assign n34324 = n5838 ^ n2577 ^ 1'b0 ;
  assign n34325 = n3845 & ~n34324 ;
  assign n34326 = n34325 ^ n23130 ^ 1'b0 ;
  assign n34327 = n7884 & ~n13487 ;
  assign n34328 = n34327 ^ n9507 ^ 1'b0 ;
  assign n34329 = ~n14829 & n34328 ;
  assign n34330 = ( n3440 & ~n4775 ) | ( n3440 & n15750 ) | ( ~n4775 & n15750 ) ;
  assign n34331 = n8523 & ~n34330 ;
  assign n34334 = n19255 ^ n18658 ^ 1'b0 ;
  assign n34335 = n8707 & n34334 ;
  assign n34336 = ~n28030 & n34335 ;
  assign n34332 = n21819 ^ n20450 ^ 1'b0 ;
  assign n34333 = x207 & n34332 ;
  assign n34337 = n34336 ^ n34333 ^ n5635 ;
  assign n34338 = n22667 | n26245 ;
  assign n34339 = n9275 ^ n3680 ^ 1'b0 ;
  assign n34340 = n17012 | n34339 ;
  assign n34341 = n4794 & ~n34340 ;
  assign n34342 = ~n23907 & n34341 ;
  assign n34343 = ( ~n6657 & n16642 ) | ( ~n6657 & n19923 ) | ( n16642 & n19923 ) ;
  assign n34344 = n12158 ^ n6479 ^ 1'b0 ;
  assign n34345 = ( n6524 & n20743 ) | ( n6524 & n34344 ) | ( n20743 & n34344 ) ;
  assign n34346 = n14935 & n23686 ;
  assign n34347 = n14714 & n27392 ;
  assign n34348 = n28168 & n34347 ;
  assign n34349 = n3655 & n8087 ;
  assign n34350 = ~n19972 & n20390 ;
  assign n34358 = n15375 ^ n8520 ^ 1'b0 ;
  assign n34359 = ~n12738 & n34358 ;
  assign n34352 = ~n1714 & n8087 ;
  assign n34353 = ~n3174 & n34352 ;
  assign n34354 = n7433 | n34353 ;
  assign n34355 = n5385 | n34354 ;
  assign n34351 = n1748 & n11685 ;
  assign n34356 = n34355 ^ n34351 ^ 1'b0 ;
  assign n34357 = n14518 | n34356 ;
  assign n34360 = n34359 ^ n34357 ^ 1'b0 ;
  assign n34361 = ~n2587 & n24541 ;
  assign n34362 = n34361 ^ n9402 ^ 1'b0 ;
  assign n34363 = ~x221 & n4608 ;
  assign n34364 = n3468 & ~n34363 ;
  assign n34365 = ~n1279 & n8884 ;
  assign n34366 = n33850 & ~n34365 ;
  assign n34367 = n18658 & ~n25459 ;
  assign n34368 = n9520 & n30825 ;
  assign n34369 = ~n9956 & n34368 ;
  assign n34370 = n22410 & n33538 ;
  assign n34371 = n5209 ^ n5075 ^ n826 ;
  assign n34372 = n10732 ^ n2615 ^ 1'b0 ;
  assign n34373 = n25674 | n34372 ;
  assign n34374 = n34373 ^ n30605 ^ 1'b0 ;
  assign n34375 = ~n3344 & n15398 ;
  assign n34376 = n34375 ^ n17854 ^ 1'b0 ;
  assign n34377 = n34376 ^ n28873 ^ n4905 ;
  assign n34378 = n14916 ^ n4923 ^ 1'b0 ;
  assign n34379 = n18285 & ~n34378 ;
  assign n34380 = n15082 ^ n3110 ^ 1'b0 ;
  assign n34381 = ~n15137 & n34380 ;
  assign n34382 = n30723 ^ n11929 ^ 1'b0 ;
  assign n34383 = n15026 & ~n19984 ;
  assign n34384 = n34382 | n34383 ;
  assign n34385 = n23178 ^ n20047 ^ 1'b0 ;
  assign n34386 = n22721 ^ n8927 ^ 1'b0 ;
  assign n34387 = n2747 & ~n14553 ;
  assign n34388 = n11963 & n34387 ;
  assign n34389 = ~n7185 & n31879 ;
  assign n34390 = ~n21600 & n34389 ;
  assign n34391 = n11999 ^ n9883 ^ n6842 ;
  assign n34392 = ( ~n5210 & n13149 ) | ( ~n5210 & n31337 ) | ( n13149 & n31337 ) ;
  assign n34393 = ~n13014 & n13239 ;
  assign n34394 = ~n16674 & n34393 ;
  assign n34395 = n10297 & ~n34394 ;
  assign n34396 = n12209 & n34395 ;
  assign n34397 = n320 & ~n31188 ;
  assign n34398 = n17482 & n18196 ;
  assign n34399 = n34398 ^ n22754 ^ 1'b0 ;
  assign n34400 = n24247 ^ n5488 ^ 1'b0 ;
  assign n34401 = n6322 ^ n6043 ^ 1'b0 ;
  assign n34402 = n7409 & n27082 ;
  assign n34403 = ~n10637 & n11237 ;
  assign n34404 = n7224 & ~n34403 ;
  assign n34405 = n26185 ^ n4381 ^ 1'b0 ;
  assign n34406 = n18888 & n27271 ;
  assign n34407 = ( n16101 & n17900 ) | ( n16101 & ~n34406 ) | ( n17900 & ~n34406 ) ;
  assign n34408 = n8816 & ~n17676 ;
  assign n34409 = ~n8816 & n34408 ;
  assign n34410 = n34409 ^ n28101 ^ n10501 ;
  assign n34411 = n12269 ^ n3959 ^ 1'b0 ;
  assign n34412 = n3529 | n5074 ;
  assign n34413 = n34411 | n34412 ;
  assign n34414 = n21492 ^ n5183 ^ 1'b0 ;
  assign n34415 = n17688 | n18875 ;
  assign n34416 = n34415 ^ n4327 ^ 1'b0 ;
  assign n34417 = ( n12787 & ~n22665 ) | ( n12787 & n34416 ) | ( ~n22665 & n34416 ) ;
  assign n34418 = n18455 & n34417 ;
  assign n34419 = n15056 | n34418 ;
  assign n34420 = n13954 & ~n34419 ;
  assign n34421 = n34420 ^ n13563 ^ 1'b0 ;
  assign n34422 = n14175 & ~n19579 ;
  assign n34423 = n31595 ^ n25462 ^ 1'b0 ;
  assign n34424 = n33190 ^ n10042 ^ 1'b0 ;
  assign n34425 = n10858 | n34424 ;
  assign n34427 = ~n5054 & n18117 ;
  assign n34428 = ~n9518 & n34427 ;
  assign n34426 = n21402 ^ n2246 ^ n1259 ;
  assign n34429 = n34428 ^ n34426 ^ n16087 ;
  assign n34430 = n4169 & n8891 ;
  assign n34431 = n34429 & n34430 ;
  assign n34432 = ~n6895 & n12555 ;
  assign n34433 = n883 & n34432 ;
  assign n34434 = n1754 | n14729 ;
  assign n34435 = n34433 & ~n34434 ;
  assign n34436 = n12068 ^ n5291 ^ 1'b0 ;
  assign n34437 = ~n9213 & n24798 ;
  assign n34438 = ~n34436 & n34437 ;
  assign n34439 = n21748 ^ n18774 ^ n983 ;
  assign n34440 = n34439 ^ n34246 ^ 1'b0 ;
  assign n34441 = n13628 | n21345 ;
  assign n34442 = ( n26865 & ~n27545 ) | ( n26865 & n32952 ) | ( ~n27545 & n32952 ) ;
  assign n34443 = n34442 ^ n23495 ^ 1'b0 ;
  assign n34444 = n13985 ^ n7899 ^ 1'b0 ;
  assign n34445 = n34444 ^ n5386 ^ 1'b0 ;
  assign n34446 = n13370 & n34445 ;
  assign n34447 = ~n4359 & n33815 ;
  assign n34448 = ~n3465 & n5595 ;
  assign n34449 = n34448 ^ n4260 ^ 1'b0 ;
  assign n34450 = ~n8312 & n21438 ;
  assign n34451 = n34450 ^ n7407 ^ 1'b0 ;
  assign n34452 = n12032 | n14470 ;
  assign n34453 = n34451 & ~n34452 ;
  assign n34454 = n20075 ^ n5946 ^ 1'b0 ;
  assign n34455 = n829 | n2443 ;
  assign n34456 = n7654 & n34455 ;
  assign n34457 = n19393 & n34456 ;
  assign n34458 = n23473 & ~n34457 ;
  assign n34459 = n18756 & n34458 ;
  assign n34460 = n3158 & n5871 ;
  assign n34461 = ( ~n8581 & n30802 ) | ( ~n8581 & n34460 ) | ( n30802 & n34460 ) ;
  assign n34462 = n34461 ^ n5284 ^ x74 ;
  assign n34463 = n18102 ^ n16589 ^ 1'b0 ;
  assign n34464 = ~n3820 & n20696 ;
  assign n34465 = n34464 ^ n13961 ^ 1'b0 ;
  assign n34466 = n11963 | n34465 ;
  assign n34467 = n32496 & ~n34466 ;
  assign n34468 = n6374 | n34467 ;
  assign n34469 = n34468 ^ n33489 ^ 1'b0 ;
  assign n34470 = n5484 & ~n19828 ;
  assign n34471 = n34470 ^ n5089 ^ 1'b0 ;
  assign n34472 = n34469 & n34471 ;
  assign n34473 = n27673 | n30299 ;
  assign n34474 = n4934 & ~n12479 ;
  assign n34475 = n34474 ^ n4327 ^ 1'b0 ;
  assign n34476 = n34475 ^ n5168 ^ 1'b0 ;
  assign n34477 = n30840 ^ n6374 ^ 1'b0 ;
  assign n34478 = n4794 & ~n34477 ;
  assign n34479 = n15324 ^ n3572 ^ 1'b0 ;
  assign n34480 = n14572 & ~n34479 ;
  assign n34481 = n5565 ^ n1667 ^ 1'b0 ;
  assign n34482 = n16661 ^ n7766 ^ 1'b0 ;
  assign n34483 = n34481 & ~n34482 ;
  assign n34484 = ~n1047 & n5987 ;
  assign n34485 = n34484 ^ n5082 ^ 1'b0 ;
  assign n34486 = n19385 & ~n34485 ;
  assign n34487 = ( n25192 & ~n34483 ) | ( n25192 & n34486 ) | ( ~n34483 & n34486 ) ;
  assign n34488 = ( n2924 & ~n9479 ) | ( n2924 & n34487 ) | ( ~n9479 & n34487 ) ;
  assign n34489 = n32791 ^ n6555 ^ 1'b0 ;
  assign n34490 = n4494 & ~n21683 ;
  assign n34491 = ~n6893 & n34490 ;
  assign n34492 = n33771 & n34491 ;
  assign n34493 = n18532 ^ n710 ^ 1'b0 ;
  assign n34494 = x250 & ~n30022 ;
  assign n34495 = n33739 ^ n17788 ^ 1'b0 ;
  assign n34496 = ~n18563 & n34495 ;
  assign n34497 = n30610 & n34496 ;
  assign n34498 = ~n34494 & n34497 ;
  assign n34499 = ~n1200 & n1490 ;
  assign n34500 = ~n21191 & n34499 ;
  assign n34501 = n34500 ^ x69 ^ 1'b0 ;
  assign n34502 = n13954 & ~n34501 ;
  assign n34503 = n15197 & n34502 ;
  assign n34504 = ~n18617 & n34503 ;
  assign n34505 = n34504 ^ n12480 ^ 1'b0 ;
  assign n34506 = n3417 & ~n14487 ;
  assign n34507 = ~n9502 & n34506 ;
  assign n34508 = n1021 & n34507 ;
  assign n34509 = n5402 & n11152 ;
  assign n34510 = ~n21670 & n34509 ;
  assign n34511 = ( ~n3712 & n19408 ) | ( ~n3712 & n23155 ) | ( n19408 & n23155 ) ;
  assign n34512 = ( n1961 & n34510 ) | ( n1961 & n34511 ) | ( n34510 & n34511 ) ;
  assign n34513 = n11964 & n26046 ;
  assign n34514 = ( n1575 & ~n2316 ) | ( n1575 & n34513 ) | ( ~n2316 & n34513 ) ;
  assign n34515 = n24165 | n34514 ;
  assign n34516 = ( n957 & n28489 ) | ( n957 & n34515 ) | ( n28489 & n34515 ) ;
  assign n34517 = n16228 | n23104 ;
  assign n34518 = n34517 ^ n8425 ^ 1'b0 ;
  assign n34519 = ~n8347 & n34518 ;
  assign n34520 = n14584 | n30357 ;
  assign n34521 = n34520 ^ n8936 ^ 1'b0 ;
  assign n34523 = n7568 | n21428 ;
  assign n34522 = x226 & n23388 ;
  assign n34524 = n34523 ^ n34522 ^ 1'b0 ;
  assign n34525 = n19649 ^ n2048 ^ 1'b0 ;
  assign n34526 = n17160 | n34525 ;
  assign n34527 = n19961 & ~n25699 ;
  assign n34528 = n34527 ^ n6582 ^ 1'b0 ;
  assign n34529 = n26516 & ~n27744 ;
  assign n34530 = n28866 ^ n14723 ^ 1'b0 ;
  assign n34531 = n11545 ^ n992 ^ 1'b0 ;
  assign n34532 = n13901 ^ n11020 ^ 1'b0 ;
  assign n34533 = n34531 & ~n34532 ;
  assign n34534 = ~n10690 & n22177 ;
  assign n34535 = n3400 & ~n6336 ;
  assign n34536 = ~n9628 & n34535 ;
  assign n34537 = n11730 ^ n9170 ^ 1'b0 ;
  assign n34538 = n26322 ^ n17113 ^ 1'b0 ;
  assign n34539 = n7608 & ~n9589 ;
  assign n34540 = n29748 ^ n13077 ^ 1'b0 ;
  assign n34541 = n2755 | n12287 ;
  assign n34542 = n276 & ~n34541 ;
  assign n34543 = n9147 ^ n5749 ^ 1'b0 ;
  assign n34544 = ~n3059 & n34543 ;
  assign n34545 = n30393 ^ n5118 ^ 1'b0 ;
  assign n34546 = n535 & ~n34545 ;
  assign n34547 = n16932 & n25104 ;
  assign n34548 = n34547 ^ n23846 ^ 1'b0 ;
  assign n34549 = ~n22547 & n34548 ;
  assign n34550 = n34549 ^ n14915 ^ 1'b0 ;
  assign n34551 = ~n9578 & n34550 ;
  assign n34552 = n2023 & n5869 ;
  assign n34553 = ~n5774 & n34552 ;
  assign n34554 = n946 | n20282 ;
  assign n34555 = ~n34553 & n34554 ;
  assign n34556 = n9870 & n24401 ;
  assign n34557 = n34556 ^ n2514 ^ 1'b0 ;
  assign n34558 = n2110 & ~n34557 ;
  assign n34559 = n10242 & n11189 ;
  assign n34560 = n12308 & ~n34559 ;
  assign n34561 = n19199 | n26582 ;
  assign n34562 = n14147 ^ n9400 ^ 1'b0 ;
  assign n34563 = n34561 | n34562 ;
  assign n34564 = n26742 ^ n17859 ^ 1'b0 ;
  assign n34565 = n11612 | n25024 ;
  assign n34566 = n34565 ^ n3267 ^ 1'b0 ;
  assign n34567 = ~n8993 & n34566 ;
  assign n34568 = n14732 ^ x150 ^ 1'b0 ;
  assign n34569 = n12361 & ~n34568 ;
  assign n34570 = n2380 | n8377 ;
  assign n34571 = ~n4202 & n4389 ;
  assign n34572 = n34571 ^ n1153 ^ 1'b0 ;
  assign n34573 = n2545 & n2936 ;
  assign n34574 = n34573 ^ n22182 ^ 1'b0 ;
  assign n34575 = n4027 & n34574 ;
  assign n34576 = n28140 & n34575 ;
  assign n34577 = n34576 ^ n12123 ^ 1'b0 ;
  assign n34578 = x152 | n14025 ;
  assign n34579 = n1129 & n17478 ;
  assign n34580 = ~n943 & n34579 ;
  assign n34581 = n34580 ^ n11514 ^ 1'b0 ;
  assign n34582 = n4670 | n6506 ;
  assign n34583 = ( n498 & n34581 ) | ( n498 & n34582 ) | ( n34581 & n34582 ) ;
  assign n34585 = n5080 | n10090 ;
  assign n34586 = n34585 ^ x107 ^ 1'b0 ;
  assign n34584 = n7699 ^ n4372 ^ 1'b0 ;
  assign n34587 = n34586 ^ n34584 ^ n20375 ;
  assign n34588 = n27960 ^ n23654 ^ 1'b0 ;
  assign n34589 = n4296 & ~n4611 ;
  assign n34590 = n12725 | n13452 ;
  assign n34591 = n34590 ^ n29414 ^ 1'b0 ;
  assign n34593 = n701 & n17970 ;
  assign n34592 = n12923 & ~n16591 ;
  assign n34594 = n34593 ^ n34592 ^ 1'b0 ;
  assign n34595 = n3328 & ~n24269 ;
  assign n34596 = n9049 ^ n3666 ^ 1'b0 ;
  assign n34598 = ~n6497 & n12072 ;
  assign n34599 = n34598 ^ n1620 ^ 1'b0 ;
  assign n34597 = ~n17149 & n21196 ;
  assign n34600 = n34599 ^ n34597 ^ 1'b0 ;
  assign n34601 = n4953 & ~n28343 ;
  assign n34602 = n2155 & n4309 ;
  assign n34603 = n25779 ^ n22934 ^ 1'b0 ;
  assign n34604 = ~n7893 & n18682 ;
  assign n34605 = n34604 ^ n1462 ^ 1'b0 ;
  assign n34606 = n25665 ^ n10231 ^ 1'b0 ;
  assign n34607 = n12713 & ~n34606 ;
  assign n34608 = n6447 & ~n21849 ;
  assign n34609 = n8493 & ~n27719 ;
  assign n34610 = n4745 & n13562 ;
  assign n34611 = n8874 ^ n1552 ^ 1'b0 ;
  assign n34612 = ~n1648 & n34611 ;
  assign n34614 = ~n765 & n15575 ;
  assign n34613 = n27494 ^ n9175 ^ 1'b0 ;
  assign n34615 = n34614 ^ n34613 ^ 1'b0 ;
  assign n34616 = n34612 & ~n34615 ;
  assign n34617 = n11379 | n26339 ;
  assign n34618 = n3845 ^ n3379 ^ 1'b0 ;
  assign n34619 = ~n595 & n2466 ;
  assign n34620 = ~n5280 & n5937 ;
  assign n34621 = n4585 | n31969 ;
  assign n34622 = n10938 | n34621 ;
  assign n34623 = ~n3685 & n34622 ;
  assign n34624 = n18804 ^ n17499 ^ 1'b0 ;
  assign n34625 = n7157 ^ n6621 ^ 1'b0 ;
  assign n34626 = n997 | n1997 ;
  assign n34627 = n34626 ^ n24233 ^ 1'b0 ;
  assign n34628 = ~n19025 & n19046 ;
  assign n34629 = ~n34627 & n34628 ;
  assign n34630 = n20280 ^ n18781 ^ n13023 ;
  assign n34631 = ~n2743 & n19634 ;
  assign n34632 = n1116 ^ n335 ^ 1'b0 ;
  assign n34633 = n7632 | n10978 ;
  assign n34634 = ~n1225 & n8745 ;
  assign n34635 = ~n34633 & n34634 ;
  assign n34636 = n21369 ^ n17455 ^ 1'b0 ;
  assign n34637 = ~n9262 & n9636 ;
  assign n34638 = n16623 ^ n4368 ^ 1'b0 ;
  assign n34639 = ~n34637 & n34638 ;
  assign n34640 = ~n9982 & n24189 ;
  assign n34641 = n15239 & n34640 ;
  assign n34642 = n34641 ^ n8172 ^ 1'b0 ;
  assign n34643 = n30022 ^ n10374 ^ 1'b0 ;
  assign n34644 = n32311 & ~n34643 ;
  assign n34645 = n15553 & ~n32269 ;
  assign n34646 = n29181 & n34645 ;
  assign n34647 = n30577 ^ n24428 ^ x43 ;
  assign n34648 = n17642 ^ n8671 ^ 1'b0 ;
  assign n34649 = n28099 | n34648 ;
  assign n34650 = n25990 | n28286 ;
  assign n34651 = x146 | n34650 ;
  assign n34652 = n3171 & n3939 ;
  assign n34653 = n8830 | n34652 ;
  assign n34654 = n9053 & n19985 ;
  assign n34655 = n34654 ^ n8839 ^ 1'b0 ;
  assign n34656 = n13606 & n23065 ;
  assign n34657 = n6248 & n8745 ;
  assign n34658 = n34657 ^ n20954 ^ 1'b0 ;
  assign n34659 = ~n19344 & n34658 ;
  assign n34660 = n6137 | n14312 ;
  assign n34661 = n34660 ^ n29996 ^ 1'b0 ;
  assign n34662 = ~n13263 & n14769 ;
  assign n34663 = n18514 ^ n488 ^ 1'b0 ;
  assign n34664 = n34662 & ~n34663 ;
  assign n34665 = n3234 & ~n6615 ;
  assign n34666 = n34665 ^ n18033 ^ 1'b0 ;
  assign n34668 = n2901 & n13404 ;
  assign n34669 = n34668 ^ n8955 ^ 1'b0 ;
  assign n34667 = n7379 & n23511 ;
  assign n34670 = n34669 ^ n34667 ^ 1'b0 ;
  assign n34671 = ~n10870 & n16403 ;
  assign n34672 = ~n17178 & n34671 ;
  assign n34673 = n34670 & ~n34672 ;
  assign n34674 = n11482 | n12133 ;
  assign n34675 = n4275 & ~n34674 ;
  assign n34676 = n6567 | n12840 ;
  assign n34677 = n34676 ^ x143 ^ 1'b0 ;
  assign n34678 = n8326 | n34677 ;
  assign n34679 = ( n13856 & n24713 ) | ( n13856 & n34678 ) | ( n24713 & n34678 ) ;
  assign n34680 = n9353 & ~n32249 ;
  assign n34681 = n5756 ^ n1487 ^ 1'b0 ;
  assign n34682 = n4733 & ~n34681 ;
  assign n34683 = n34682 ^ n16815 ^ 1'b0 ;
  assign n34684 = n22740 & ~n34683 ;
  assign n34685 = n19941 | n26524 ;
  assign n34686 = n34684 & ~n34685 ;
  assign n34687 = n21899 ^ n14384 ^ 1'b0 ;
  assign n34688 = n23128 & ~n34687 ;
  assign n34689 = x14 & n16085 ;
  assign n34690 = ~n16085 & n34689 ;
  assign n34692 = n14398 & ~n19955 ;
  assign n34691 = n12653 & n15243 ;
  assign n34693 = n34692 ^ n34691 ^ n8414 ;
  assign n34694 = ( n18567 & n21979 ) | ( n18567 & n26342 ) | ( n21979 & n26342 ) ;
  assign n34695 = n6387 & ~n19417 ;
  assign n34696 = n32339 ^ n26532 ^ n10637 ;
  assign n34697 = ( n5118 & ~n12426 ) | ( n5118 & n25109 ) | ( ~n12426 & n25109 ) ;
  assign n34698 = n34696 & ~n34697 ;
  assign n34700 = n3142 | n12812 ;
  assign n34699 = ~n5637 & n6152 ;
  assign n34701 = n34700 ^ n34699 ^ 1'b0 ;
  assign n34702 = n17029 ^ n8814 ^ 1'b0 ;
  assign n34703 = ~n31721 & n34702 ;
  assign n34704 = n24699 ^ n15405 ^ 1'b0 ;
  assign n34705 = n24365 ^ n10451 ^ 1'b0 ;
  assign n34706 = n4222 | n17067 ;
  assign n34707 = n24907 | n34706 ;
  assign n34708 = ~n1689 & n14620 ;
  assign n34709 = n34708 ^ n29823 ^ 1'b0 ;
  assign n34710 = n28002 ^ n16947 ^ 1'b0 ;
  assign n34711 = n2367 | n8713 ;
  assign n34712 = n34711 ^ n8845 ^ 1'b0 ;
  assign n34713 = ~n4387 & n34712 ;
  assign n34714 = n34713 ^ n10291 ^ 1'b0 ;
  assign n34715 = n14929 & ~n23694 ;
  assign n34716 = n18750 | n31017 ;
  assign n34717 = n9095 & ~n23054 ;
  assign n34718 = ~n10657 & n34717 ;
  assign n34719 = n30810 ^ n7806 ^ n2663 ;
  assign n34720 = ( n17763 & n34718 ) | ( n17763 & n34719 ) | ( n34718 & n34719 ) ;
  assign n34721 = ~n310 & n4635 ;
  assign n34722 = n34721 ^ n34564 ^ 1'b0 ;
  assign n34723 = ~n18256 & n34722 ;
  assign n34724 = n9505 & n32853 ;
  assign n34725 = n33805 ^ n27475 ^ 1'b0 ;
  assign n34726 = ~n3050 & n12969 ;
  assign n34727 = ( n4216 & n4953 ) | ( n4216 & ~n5735 ) | ( n4953 & ~n5735 ) ;
  assign n34728 = n1589 & n34727 ;
  assign n34729 = n34728 ^ n2246 ^ 1'b0 ;
  assign n34730 = n34726 & ~n34729 ;
  assign n34732 = n8702 ^ n3411 ^ 1'b0 ;
  assign n34731 = ~n3129 & n13938 ;
  assign n34733 = n34732 ^ n34731 ^ n16396 ;
  assign n34734 = n17123 ^ n9974 ^ 1'b0 ;
  assign n34735 = n34734 ^ n3928 ^ 1'b0 ;
  assign n34736 = n17258 & n34735 ;
  assign n34737 = n30444 ^ n4964 ^ 1'b0 ;
  assign n34740 = x6 & x25 ;
  assign n34741 = n1990 & n34740 ;
  assign n34738 = n9484 & n11416 ;
  assign n34739 = n34738 ^ n2993 ^ 1'b0 ;
  assign n34742 = n34741 ^ n34739 ^ n3823 ;
  assign n34743 = n1262 & n5206 ;
  assign n34744 = n34743 ^ n27816 ^ 1'b0 ;
  assign n34745 = n23333 ^ n2719 ^ 1'b0 ;
  assign n34746 = n2502 ^ n334 ^ 1'b0 ;
  assign n34747 = n12413 & n34746 ;
  assign n34748 = n34747 ^ n16435 ^ 1'b0 ;
  assign n34749 = n24319 & n34748 ;
  assign n34750 = n34749 ^ n22520 ^ 1'b0 ;
  assign n34751 = n25937 ^ n14690 ^ 1'b0 ;
  assign n34752 = ~n21716 & n34751 ;
  assign n34753 = n7601 & n11923 ;
  assign n34754 = n33133 ^ n15252 ^ n6370 ;
  assign n34755 = n27606 ^ n25084 ^ 1'b0 ;
  assign n34756 = n30041 | n34755 ;
  assign n34757 = n34756 ^ n11369 ^ 1'b0 ;
  assign n34758 = n2540 & ~n34757 ;
  assign n34759 = ( n15594 & n22378 ) | ( n15594 & n25017 ) | ( n22378 & n25017 ) ;
  assign n34760 = n16137 ^ n1766 ^ 1'b0 ;
  assign n34761 = n34759 & n34760 ;
  assign n34762 = n20914 & ~n34761 ;
  assign n34763 = n12754 ^ n7350 ^ 1'b0 ;
  assign n34764 = n24247 ^ n7858 ^ 1'b0 ;
  assign n34765 = n10652 & ~n34764 ;
  assign n34766 = n11232 ^ n1653 ^ 1'b0 ;
  assign n34767 = n8424 & n34766 ;
  assign n34768 = n11354 & n34767 ;
  assign n34769 = n9958 ^ n9856 ^ 1'b0 ;
  assign n34770 = ~n5328 & n22249 ;
  assign n34771 = ~n3106 & n34770 ;
  assign n34772 = n13458 | n34771 ;
  assign n34773 = n34772 ^ n5846 ^ 1'b0 ;
  assign n34774 = ~n10929 & n21590 ;
  assign n34775 = n4090 ^ n3134 ^ 1'b0 ;
  assign n34776 = n4426 | n34775 ;
  assign n34777 = ( n7574 & n17682 ) | ( n7574 & n34776 ) | ( n17682 & n34776 ) ;
  assign n34778 = n2602 & n12418 ;
  assign n34779 = ~n7523 & n34778 ;
  assign n34780 = ~n34777 & n34779 ;
  assign n34781 = ( ~n858 & n11986 ) | ( ~n858 & n17741 ) | ( n11986 & n17741 ) ;
  assign n34782 = n21137 ^ n2062 ^ 1'b0 ;
  assign n34783 = n34782 ^ n17509 ^ 1'b0 ;
  assign n34784 = n21413 ^ n7255 ^ 1'b0 ;
  assign n34785 = n34783 & n34784 ;
  assign n34786 = n34781 & n34785 ;
  assign n34787 = n3106 | n14952 ;
  assign n34788 = n34787 ^ n5586 ^ 1'b0 ;
  assign n34789 = ( ~n1251 & n5511 ) | ( ~n1251 & n28516 ) | ( n5511 & n28516 ) ;
  assign n34790 = n15867 & n34789 ;
  assign n34791 = n9533 & ~n23281 ;
  assign n34792 = ( ~n19011 & n27005 ) | ( ~n19011 & n27490 ) | ( n27005 & n27490 ) ;
  assign n34793 = n8642 ^ n6881 ^ 1'b0 ;
  assign n34794 = n21990 ^ n20265 ^ 1'b0 ;
  assign n34795 = n34793 & ~n34794 ;
  assign n34796 = n16146 & n18526 ;
  assign n34797 = n34796 ^ n18235 ^ 1'b0 ;
  assign n34798 = ~n2701 & n15574 ;
  assign n34799 = n34798 ^ n15138 ^ 1'b0 ;
  assign n34800 = n9993 ^ n6506 ^ 1'b0 ;
  assign n34801 = n509 | n7691 ;
  assign n34802 = ( n3951 & n14010 ) | ( n3951 & ~n34801 ) | ( n14010 & ~n34801 ) ;
  assign n34804 = ( n1997 & n8117 ) | ( n1997 & ~n9892 ) | ( n8117 & ~n9892 ) ;
  assign n34803 = n9391 & n17896 ;
  assign n34805 = n34804 ^ n34803 ^ 1'b0 ;
  assign n34806 = n19712 & ~n34805 ;
  assign n34807 = n1283 & n34806 ;
  assign n34808 = n34807 ^ n21262 ^ n16374 ;
  assign n34809 = ~n7382 & n30303 ;
  assign n34810 = n608 | n26102 ;
  assign n34811 = n34809 & ~n34810 ;
  assign n34812 = n34811 ^ n29555 ^ 1'b0 ;
  assign n34813 = ~n2957 & n34812 ;
  assign n34814 = n25517 ^ n1710 ^ 1'b0 ;
  assign n34815 = ~n12909 & n16594 ;
  assign n34816 = n34814 & n34815 ;
  assign n34817 = n10899 | n34051 ;
  assign n34818 = ~n14222 & n34817 ;
  assign n34821 = n30671 ^ n10177 ^ 1'b0 ;
  assign n34819 = n16708 & n23475 ;
  assign n34820 = ~n19712 & n34819 ;
  assign n34822 = n34821 ^ n34820 ^ 1'b0 ;
  assign n34823 = n6067 | n27072 ;
  assign n34824 = n18475 & ~n31479 ;
  assign n34825 = n26827 & n34824 ;
  assign n34826 = n22559 ^ n18320 ^ 1'b0 ;
  assign n34827 = x145 | n13268 ;
  assign n34828 = n19372 ^ n3014 ^ 1'b0 ;
  assign n34829 = ( ~n11572 & n33152 ) | ( ~n11572 & n34828 ) | ( n33152 & n34828 ) ;
  assign n34830 = n20939 ^ n3439 ^ 1'b0 ;
  assign n34831 = n34829 & ~n34830 ;
  assign n34832 = n7506 & n15669 ;
  assign n34833 = ~n12253 & n34832 ;
  assign n34834 = ( ~n3886 & n24371 ) | ( ~n3886 & n34833 ) | ( n24371 & n34833 ) ;
  assign n34835 = n34834 ^ n23494 ^ n17305 ;
  assign n34836 = n26752 ^ n23751 ^ n1148 ;
  assign n34837 = ~n1695 & n2164 ;
  assign n34838 = ~n2409 & n34837 ;
  assign n34839 = n34838 ^ n15277 ^ n12247 ;
  assign n34840 = n7987 & ~n34839 ;
  assign n34841 = n26816 & n34840 ;
  assign n34842 = n10190 ^ n3258 ^ 1'b0 ;
  assign n34843 = n34842 ^ n3139 ^ 1'b0 ;
  assign n34844 = n10046 | n34843 ;
  assign n34845 = n25802 ^ n3962 ^ n3237 ;
  assign n34846 = ~n2362 & n34845 ;
  assign n34847 = n714 | n34846 ;
  assign n34848 = n2884 | n34847 ;
  assign n34849 = n1420 | n3465 ;
  assign n34850 = n4931 & ~n34849 ;
  assign n34851 = n11365 & n34850 ;
  assign n34852 = ( n2846 & ~n31298 ) | ( n2846 & n33764 ) | ( ~n31298 & n33764 ) ;
  assign n34853 = n6782 | n27955 ;
  assign n34854 = n21580 ^ n558 ^ 1'b0 ;
  assign n34855 = ~n9540 & n34854 ;
  assign n34856 = n8535 & n23485 ;
  assign n34857 = n34856 ^ n8499 ^ 1'b0 ;
  assign n34858 = n34857 ^ n13221 ^ 1'b0 ;
  assign n34859 = n33713 ^ n1814 ^ 1'b0 ;
  assign n34860 = n24181 ^ n14768 ^ n10287 ;
  assign n34861 = n34860 ^ n15070 ^ 1'b0 ;
  assign n34862 = n2158 ^ n1681 ^ 1'b0 ;
  assign n34863 = n34861 & ~n34862 ;
  assign n34864 = n22603 ^ n14167 ^ 1'b0 ;
  assign n34865 = n9270 ^ n9104 ^ 1'b0 ;
  assign n34866 = ( n2353 & n24669 ) | ( n2353 & ~n26982 ) | ( n24669 & ~n26982 ) ;
  assign n34867 = n2493 & n13626 ;
  assign n34868 = ~n32336 & n34867 ;
  assign n34869 = n33896 & n34124 ;
  assign n34870 = n34869 ^ n18938 ^ 1'b0 ;
  assign n34871 = ( ~n2047 & n3801 ) | ( ~n2047 & n5496 ) | ( n3801 & n5496 ) ;
  assign n34872 = n5253 & ~n34871 ;
  assign n34873 = n34872 ^ n28544 ^ 1'b0 ;
  assign n34874 = n1129 & n18104 ;
  assign n34875 = n34874 ^ n16878 ^ 1'b0 ;
  assign n34876 = n34875 ^ n2915 ^ 1'b0 ;
  assign n34877 = n4622 | n34876 ;
  assign n34879 = n680 | n23957 ;
  assign n34878 = ~n11891 & n14760 ;
  assign n34880 = n34879 ^ n34878 ^ 1'b0 ;
  assign n34881 = x137 & n34880 ;
  assign n34882 = n9330 & n34881 ;
  assign n34883 = n4840 & ~n34882 ;
  assign n34884 = n34883 ^ x192 ^ 1'b0 ;
  assign n34885 = x143 & ~n11963 ;
  assign n34886 = n7310 & n34885 ;
  assign n34887 = n34886 ^ n18472 ^ n2291 ;
  assign n34888 = n19283 & n34887 ;
  assign n34889 = n32733 ^ n20349 ^ 1'b0 ;
  assign n34890 = n33090 | n34889 ;
  assign n34891 = n5368 | n8463 ;
  assign n34892 = n14310 & n25685 ;
  assign n34893 = n19608 & n34892 ;
  assign n34894 = ~n24172 & n24214 ;
  assign n34895 = n7966 & n34894 ;
  assign n34896 = n15626 & n19435 ;
  assign n34897 = n34896 ^ n4436 ^ 1'b0 ;
  assign n34898 = ( n10523 & ~n14307 ) | ( n10523 & n20724 ) | ( ~n14307 & n20724 ) ;
  assign n34899 = n32178 & n34898 ;
  assign n34900 = ~n34897 & n34899 ;
  assign n34901 = ~n5418 & n17654 ;
  assign n34902 = ~n4348 & n15615 ;
  assign n34903 = ~n4153 & n34902 ;
  assign n34904 = n34903 ^ n19622 ^ 1'b0 ;
  assign n34905 = n882 & n13952 ;
  assign n34906 = n20817 | n34905 ;
  assign n34907 = ( n5237 & n34904 ) | ( n5237 & n34906 ) | ( n34904 & n34906 ) ;
  assign n34908 = n30330 ^ n28780 ^ 1'b0 ;
  assign n34909 = n3272 | n4682 ;
  assign n34910 = n2128 | n34909 ;
  assign n34911 = n34910 ^ n34518 ^ 1'b0 ;
  assign n34912 = n5016 & n8077 ;
  assign n34913 = n34912 ^ n17519 ^ 1'b0 ;
  assign n34914 = n18930 & n27332 ;
  assign n34915 = n34914 ^ n27791 ^ 1'b0 ;
  assign n34916 = n15385 & ~n23254 ;
  assign n34917 = n34916 ^ n14805 ^ 1'b0 ;
  assign n34918 = ~n9708 & n24776 ;
  assign n34919 = n12553 & n14536 ;
  assign n34920 = n34919 ^ n27301 ^ 1'b0 ;
  assign n34921 = n34681 ^ n18364 ^ n10333 ;
  assign n34922 = n4691 & ~n33435 ;
  assign n34923 = x215 & n6639 ;
  assign n34924 = ~n8742 & n34923 ;
  assign n34925 = ~n724 & n17843 ;
  assign n34926 = n34925 ^ n9377 ^ 1'b0 ;
  assign n34927 = n19639 ^ n2641 ^ n491 ;
  assign n34928 = ( n13670 & n34926 ) | ( n13670 & ~n34927 ) | ( n34926 & ~n34927 ) ;
  assign n34929 = n9173 ^ n2307 ^ 1'b0 ;
  assign n34930 = x13 & n34929 ;
  assign n34931 = n8023 & ~n34930 ;
  assign n34932 = n4888 & ~n4965 ;
  assign n34933 = n34932 ^ n4752 ^ 1'b0 ;
  assign n34934 = n2211 & n34933 ;
  assign n34935 = ~n4821 & n22522 ;
  assign n34936 = n9755 & n23818 ;
  assign n34937 = n34936 ^ n15490 ^ 1'b0 ;
  assign n34938 = n1219 | n29926 ;
  assign n34939 = n14739 | n34938 ;
  assign n34940 = n28323 | n34939 ;
  assign n34941 = ~n34937 & n34940 ;
  assign n34942 = n5488 & n9365 ;
  assign n34943 = n34942 ^ n18298 ^ 1'b0 ;
  assign n34944 = ~n11371 & n34943 ;
  assign n34945 = n34941 | n34944 ;
  assign n34946 = n6875 & n34945 ;
  assign n34947 = ~n28616 & n34946 ;
  assign n34948 = n17176 ^ n15137 ^ 1'b0 ;
  assign n34949 = ~n1899 & n9982 ;
  assign n34950 = n5355 & n34949 ;
  assign n34951 = n34950 ^ n3855 ^ 1'b0 ;
  assign n34952 = n34951 ^ n26273 ^ n23953 ;
  assign n34953 = n34948 & n34952 ;
  assign n34954 = ~n11462 & n34953 ;
  assign n34955 = ~x153 & n1611 ;
  assign n34956 = n6116 ^ n686 ^ 1'b0 ;
  assign n34957 = n4298 ^ n716 ^ 1'b0 ;
  assign n34958 = n20772 & ~n34957 ;
  assign n34959 = n12556 ^ n1487 ^ 1'b0 ;
  assign n34960 = ~n27165 & n34959 ;
  assign n34961 = n34960 ^ n4637 ^ 1'b0 ;
  assign n34962 = n6688 & ~n28424 ;
  assign n34963 = ~n34961 & n34962 ;
  assign n34964 = n33553 ^ n10652 ^ 1'b0 ;
  assign n34965 = x140 & ~n34964 ;
  assign n34966 = n13954 & n34965 ;
  assign n34967 = n12696 & n34966 ;
  assign n34968 = ~n16037 & n33830 ;
  assign n34969 = ( ~n367 & n13633 ) | ( ~n367 & n15520 ) | ( n13633 & n15520 ) ;
  assign n34970 = n34969 ^ n8351 ^ n4957 ;
  assign n34971 = n34970 ^ n15683 ^ 1'b0 ;
  assign n34972 = n3793 | n32496 ;
  assign n34973 = n34972 ^ n2968 ^ 1'b0 ;
  assign n34974 = n27832 ^ n3003 ^ 1'b0 ;
  assign n34975 = n18133 | n18873 ;
  assign n34976 = n20201 & ~n34975 ;
  assign n34977 = n17911 ^ n8368 ^ 1'b0 ;
  assign n34978 = n12633 & n16654 ;
  assign n34979 = ( n3016 & n10085 ) | ( n3016 & n22312 ) | ( n10085 & n22312 ) ;
  assign n34980 = n25066 ^ n8421 ^ 1'b0 ;
  assign n34981 = n1242 & n34980 ;
  assign n34982 = n21109 ^ n17041 ^ 1'b0 ;
  assign n34983 = n5963 | n34982 ;
  assign n34984 = n3716 & ~n15733 ;
  assign n34985 = n7484 & n34984 ;
  assign n34986 = n34985 ^ n4522 ^ 1'b0 ;
  assign n34987 = n9833 & n34986 ;
  assign n34988 = n18972 ^ n10299 ^ n2368 ;
  assign n34989 = n5003 & n22039 ;
  assign n34990 = n34989 ^ n2370 ^ 1'b0 ;
  assign n34991 = n1032 & n6781 ;
  assign n34992 = n5446 & n34991 ;
  assign n34993 = n19333 ^ n8344 ^ 1'b0 ;
  assign n34994 = n34992 | n34993 ;
  assign n34995 = n18726 ^ n2426 ^ 1'b0 ;
  assign n34996 = ~n21901 & n34995 ;
  assign n34997 = n34996 ^ n11696 ^ 1'b0 ;
  assign n34998 = ~n19297 & n34997 ;
  assign n34999 = n16193 & n34998 ;
  assign n35000 = n34999 ^ n529 ^ 1'b0 ;
  assign n35001 = n24573 ^ n21164 ^ 1'b0 ;
  assign n35002 = n3704 & n35001 ;
  assign n35003 = n11166 ^ n2999 ^ 1'b0 ;
  assign n35004 = ~n5195 & n8428 ;
  assign n35005 = ~n2404 & n35004 ;
  assign n35006 = ( x61 & n784 ) | ( x61 & n34166 ) | ( n784 & n34166 ) ;
  assign n35007 = n19955 ^ n14296 ^ n5001 ;
  assign n35008 = n35006 & n35007 ;
  assign n35009 = n26868 ^ n16723 ^ 1'b0 ;
  assign n35010 = n12855 & n35009 ;
  assign n35011 = n24139 ^ n5173 ^ n1684 ;
  assign n35012 = n34613 ^ n7596 ^ 1'b0 ;
  assign n35013 = n33607 | n35012 ;
  assign n35014 = x208 & ~n5534 ;
  assign n35015 = n7474 & n35014 ;
  assign n35016 = n3576 & ~n35015 ;
  assign n35017 = n28636 ^ n20372 ^ 1'b0 ;
  assign n35018 = n35016 & n35017 ;
  assign n35019 = n34335 ^ n25070 ^ 1'b0 ;
  assign n35020 = n21949 | n35019 ;
  assign n35021 = n35020 ^ n22471 ^ 1'b0 ;
  assign n35022 = n274 & n25694 ;
  assign n35023 = n31047 ^ n14641 ^ 1'b0 ;
  assign n35024 = n35022 & ~n35023 ;
  assign n35025 = n21491 & ~n27162 ;
  assign n35026 = n35025 ^ n13883 ^ 1'b0 ;
  assign n35027 = n16571 ^ n3646 ^ 1'b0 ;
  assign n35028 = ( ~n984 & n22014 ) | ( ~n984 & n35027 ) | ( n22014 & n35027 ) ;
  assign n35029 = n20313 ^ n14317 ^ 1'b0 ;
  assign n35030 = ~x62 & n35029 ;
  assign n35031 = ~n17780 & n35030 ;
  assign n35032 = n35031 ^ n33184 ^ 1'b0 ;
  assign n35033 = n30168 ^ n8700 ^ 1'b0 ;
  assign n35034 = ~n26461 & n35033 ;
  assign n35035 = n5421 ^ n4616 ^ x113 ;
  assign n35036 = n35035 ^ n6256 ^ 1'b0 ;
  assign n35037 = n830 & n33725 ;
  assign n35038 = n21917 | n35037 ;
  assign n35041 = n20257 ^ n14114 ^ 1'b0 ;
  assign n35042 = n28135 | n35041 ;
  assign n35039 = n26225 & n32823 ;
  assign n35040 = ~n19292 & n35039 ;
  assign n35043 = n35042 ^ n35040 ^ 1'b0 ;
  assign n35044 = n12569 ^ n1384 ^ 1'b0 ;
  assign n35045 = n20505 & n35044 ;
  assign n35046 = n16989 ^ n8505 ^ 1'b0 ;
  assign n35047 = n13343 & n35046 ;
  assign n35048 = n5767 | n22661 ;
  assign n35049 = n19546 | n35048 ;
  assign n35050 = n11767 & n35049 ;
  assign n35051 = n17089 & n35050 ;
  assign n35052 = n6184 & n21995 ;
  assign n35053 = n35052 ^ n27043 ^ 1'b0 ;
  assign n35054 = n25977 ^ n9072 ^ 1'b0 ;
  assign n35055 = n15553 & ~n35054 ;
  assign n35056 = n11628 & ~n12532 ;
  assign n35057 = ~n12231 & n28295 ;
  assign n35058 = ~n6583 & n28625 ;
  assign n35059 = n10942 | n23386 ;
  assign n35060 = n35058 | n35059 ;
  assign n35062 = n10006 ^ n2782 ^ 1'b0 ;
  assign n35063 = ~n16066 & n35062 ;
  assign n35061 = n18477 ^ n17447 ^ 1'b0 ;
  assign n35064 = n35063 ^ n35061 ^ n18548 ;
  assign n35065 = n4794 & n35064 ;
  assign n35066 = ~n7015 & n10794 ;
  assign n35067 = n35066 ^ n21563 ^ n20805 ;
  assign n35068 = n4122 | n5485 ;
  assign n35069 = n35068 ^ n22141 ^ 1'b0 ;
  assign n35070 = n27509 ^ n6269 ^ 1'b0 ;
  assign n35071 = n35070 ^ n21879 ^ 1'b0 ;
  assign n35072 = n5594 & ~n6456 ;
  assign n35073 = n9452 | n35072 ;
  assign n35074 = n5134 & n21306 ;
  assign n35075 = n4330 & n35074 ;
  assign n35076 = n28008 | n35075 ;
  assign n35077 = n34444 ^ n16395 ^ 1'b0 ;
  assign n35078 = n8087 & ~n8630 ;
  assign n35079 = n27126 ^ n9611 ^ 1'b0 ;
  assign n35080 = n19931 ^ n5458 ^ 1'b0 ;
  assign n35081 = n12778 & ~n30799 ;
  assign n35082 = n10150 | n19200 ;
  assign n35083 = n9773 ^ x11 ^ 1'b0 ;
  assign n35084 = n35082 & ~n35083 ;
  assign n35085 = n7581 & n8192 ;
  assign n35086 = n35085 ^ n16640 ^ 1'b0 ;
  assign n35087 = ~n2216 & n35086 ;
  assign n35088 = n35087 ^ n13890 ^ 1'b0 ;
  assign n35089 = n8077 ^ n7486 ^ n5428 ;
  assign n35090 = n35089 ^ n33111 ^ n9009 ;
  assign n35091 = n35090 ^ n2988 ^ 1'b0 ;
  assign n35092 = ( n869 & n3082 ) | ( n869 & ~n35091 ) | ( n3082 & ~n35091 ) ;
  assign n35093 = n35092 ^ n6499 ^ 1'b0 ;
  assign n35094 = ~n6253 & n35093 ;
  assign n35095 = n7814 & n31320 ;
  assign n35096 = n3607 & n16885 ;
  assign n35097 = ~n9288 & n35096 ;
  assign n35098 = n1343 & n5720 ;
  assign n35099 = n35097 & ~n35098 ;
  assign n35100 = n8125 & n35099 ;
  assign n35101 = n12896 ^ n5617 ^ 1'b0 ;
  assign n35102 = ~n26964 & n35101 ;
  assign n35103 = ~n4241 & n14183 ;
  assign n35104 = n22905 ^ n707 ^ 1'b0 ;
  assign n35105 = n24773 & ~n35104 ;
  assign n35106 = n35105 ^ n11255 ^ 1'b0 ;
  assign n35107 = n16956 ^ n9708 ^ 1'b0 ;
  assign n35108 = n33750 & ~n35107 ;
  assign n35109 = n24004 ^ n7620 ^ 1'b0 ;
  assign n35110 = n35108 & n35109 ;
  assign n35111 = n11410 ^ n4375 ^ 1'b0 ;
  assign n35112 = ~x99 & n25125 ;
  assign n35113 = n32585 | n35112 ;
  assign n35115 = x105 & n20153 ;
  assign n35114 = ~n7035 & n11134 ;
  assign n35116 = n35115 ^ n35114 ^ 1'b0 ;
  assign n35117 = n27716 | n35116 ;
  assign n35118 = n5187 ^ n4428 ^ 1'b0 ;
  assign n35119 = ( n9513 & n13292 ) | ( n9513 & n35118 ) | ( n13292 & n35118 ) ;
  assign n35120 = n29703 ^ n4124 ^ 1'b0 ;
  assign n35121 = n6864 | n20495 ;
  assign n35122 = ~n3812 & n35121 ;
  assign n35123 = n31507 & ~n35122 ;
  assign n35124 = n8198 | n32746 ;
  assign n35125 = n2385 & ~n28158 ;
  assign n35126 = ~n2706 & n25495 ;
  assign n35127 = n18361 ^ n16906 ^ 1'b0 ;
  assign n35128 = n35127 ^ n34662 ^ 1'b0 ;
  assign n35129 = n30865 ^ n19626 ^ 1'b0 ;
  assign n35130 = x205 & ~n3966 ;
  assign n35131 = n16026 & n35130 ;
  assign n35132 = n35131 ^ n17143 ^ n6733 ;
  assign n35133 = n35129 & ~n35132 ;
  assign n35134 = n20103 & n35133 ;
  assign n35135 = n35134 ^ n10944 ^ 1'b0 ;
  assign n35136 = n18067 & n20181 ;
  assign n35137 = n14188 ^ n11770 ^ n1112 ;
  assign n35138 = n23364 & n35137 ;
  assign n35139 = ~n35136 & n35138 ;
  assign n35140 = ~n4896 & n28649 ;
  assign n35141 = n35140 ^ n22114 ^ 1'b0 ;
  assign n35142 = n8011 & n35141 ;
  assign n35143 = n9019 ^ n6112 ^ 1'b0 ;
  assign n35144 = n26626 ^ n20152 ^ 1'b0 ;
  assign n35145 = n18123 | n35144 ;
  assign n35146 = n12225 | n35145 ;
  assign n35147 = n35146 ^ n31805 ^ 1'b0 ;
  assign n35148 = ( n19290 & n35143 ) | ( n19290 & n35147 ) | ( n35143 & n35147 ) ;
  assign n35149 = ~n15347 & n26663 ;
  assign n35150 = n35149 ^ n14584 ^ 1'b0 ;
  assign n35151 = x202 & ~n801 ;
  assign n35152 = ~x202 & n35151 ;
  assign n35153 = n1500 | n35152 ;
  assign n35154 = n4095 & n35153 ;
  assign n35155 = n35154 ^ n15353 ^ 1'b0 ;
  assign n35156 = n12608 & ~n15725 ;
  assign n35157 = n35156 ^ n2951 ^ 1'b0 ;
  assign n35158 = n35157 ^ n31871 ^ 1'b0 ;
  assign n35159 = n25132 ^ n12650 ^ 1'b0 ;
  assign n35160 = n11659 & n15875 ;
  assign n35161 = ~n20547 & n35160 ;
  assign n35162 = n16364 ^ n16122 ^ 1'b0 ;
  assign n35163 = n33530 & n35162 ;
  assign n35165 = n13176 ^ n3483 ^ 1'b0 ;
  assign n35164 = ~n5151 & n10501 ;
  assign n35166 = n35165 ^ n35164 ^ 1'b0 ;
  assign n35167 = n6024 & ~n35166 ;
  assign n35168 = n35167 ^ n20786 ^ 1'b0 ;
  assign n35169 = n4762 | n29285 ;
  assign n35170 = n2192 & n11055 ;
  assign n35171 = n35170 ^ n28795 ^ 1'b0 ;
  assign n35172 = ~n35169 & n35171 ;
  assign n35173 = n29623 & n35172 ;
  assign n35174 = n10915 ^ n3234 ^ 1'b0 ;
  assign n35175 = n35174 ^ n8188 ^ n772 ;
  assign n35176 = n28383 ^ n16591 ^ n2528 ;
  assign n35177 = n6257 & ~n12734 ;
  assign n35178 = n35177 ^ n13249 ^ 1'b0 ;
  assign n35181 = n9856 | n11355 ;
  assign n35182 = n11764 & ~n35181 ;
  assign n35180 = n5356 & ~n11017 ;
  assign n35183 = n35182 ^ n35180 ^ n10767 ;
  assign n35179 = ~n1095 & n15224 ;
  assign n35184 = n35183 ^ n35179 ^ 1'b0 ;
  assign n35185 = n3823 ^ x61 ^ 1'b0 ;
  assign n35186 = n19792 & n35185 ;
  assign n35187 = n35186 ^ n25524 ^ 1'b0 ;
  assign n35188 = ~n10134 & n11685 ;
  assign n35189 = ~n25070 & n35188 ;
  assign n35190 = n22655 & ~n35189 ;
  assign n35191 = n5705 ^ n4563 ^ 1'b0 ;
  assign n35192 = n8722 | n35191 ;
  assign n35193 = n4044 & ~n17550 ;
  assign n35194 = n25257 & n30802 ;
  assign n35195 = n35194 ^ n3920 ^ 1'b0 ;
  assign n35196 = ~n12944 & n31765 ;
  assign n35197 = ~n35195 & n35196 ;
  assign n35198 = n24592 ^ n16763 ^ 1'b0 ;
  assign n35199 = n23335 ^ n13313 ^ 1'b0 ;
  assign n35200 = n25628 ^ n3206 ^ 1'b0 ;
  assign n35201 = n22295 & ~n35200 ;
  assign n35202 = n15240 & n15446 ;
  assign n35203 = ( ~n710 & n9362 ) | ( ~n710 & n21474 ) | ( n9362 & n21474 ) ;
  assign n35204 = n19462 ^ n19185 ^ 1'b0 ;
  assign n35205 = n14575 ^ n4208 ^ 1'b0 ;
  assign n35206 = n33018 & n35205 ;
  assign n35207 = n2678 ^ x185 ^ 1'b0 ;
  assign n35208 = n2643 & n35207 ;
  assign n35209 = n21252 ^ n19865 ^ 1'b0 ;
  assign n35210 = n35208 & n35209 ;
  assign n35211 = ~n1051 & n35210 ;
  assign n35212 = n27164 & n35211 ;
  assign n35213 = ~n8236 & n23065 ;
  assign n35214 = n10480 & n35213 ;
  assign n35215 = ~n8468 & n35214 ;
  assign n35216 = n35215 ^ n5315 ^ 1'b0 ;
  assign n35217 = n4035 & n23629 ;
  assign n35218 = n2097 ^ x208 ^ 1'b0 ;
  assign n35219 = n2415 & n35218 ;
  assign n35220 = n35219 ^ n6297 ^ 1'b0 ;
  assign n35221 = n15137 | n19373 ;
  assign n35222 = n35220 | n35221 ;
  assign n35223 = ( n29318 & n35217 ) | ( n29318 & n35222 ) | ( n35217 & n35222 ) ;
  assign n35224 = n3525 & n19369 ;
  assign n35225 = ~n17392 & n35224 ;
  assign n35226 = n12972 ^ n11253 ^ 1'b0 ;
  assign n35227 = ~n12450 & n35226 ;
  assign n35228 = n10737 & n12542 ;
  assign n35229 = n8547 ^ n3837 ^ 1'b0 ;
  assign n35230 = ~n35228 & n35229 ;
  assign n35232 = n13515 ^ n11097 ^ n5391 ;
  assign n35231 = n20450 & ~n26322 ;
  assign n35233 = n35232 ^ n35231 ^ 1'b0 ;
  assign n35234 = ~n858 & n26595 ;
  assign n35235 = ~n5619 & n18180 ;
  assign n35236 = n13465 & n35235 ;
  assign n35237 = ~n14553 & n35236 ;
  assign n35238 = ~n3537 & n16608 ;
  assign n35239 = ( n1154 & n20813 ) | ( n1154 & ~n35238 ) | ( n20813 & ~n35238 ) ;
  assign n35240 = n14298 & n15466 ;
  assign n35241 = n1989 & ~n32819 ;
  assign n35242 = n18083 | n21601 ;
  assign n35243 = n35242 ^ n14470 ^ 1'b0 ;
  assign n35244 = n15113 ^ n6500 ^ 1'b0 ;
  assign n35245 = ~n4226 & n35244 ;
  assign n35247 = n4152 & n7149 ;
  assign n35248 = ~n2827 & n35247 ;
  assign n35246 = n3795 & ~n12576 ;
  assign n35249 = n35248 ^ n35246 ^ 1'b0 ;
  assign n35250 = ~n5252 & n22527 ;
  assign n35251 = n35250 ^ n8165 ^ 1'b0 ;
  assign n35252 = n4472 & n8646 ;
  assign n35253 = ~n35251 & n35252 ;
  assign n35254 = n31051 ^ n29162 ^ 1'b0 ;
  assign n35255 = ~n17056 & n35254 ;
  assign n35256 = ( x100 & n16620 ) | ( x100 & n17933 ) | ( n16620 & n17933 ) ;
  assign n35257 = n34223 ^ n21926 ^ 1'b0 ;
  assign n35258 = n35256 & n35257 ;
  assign n35259 = n1656 | n24005 ;
  assign n35260 = n16599 | n35259 ;
  assign n35261 = n35260 ^ n20483 ^ n3177 ;
  assign n35262 = n11330 ^ n8914 ^ 1'b0 ;
  assign n35263 = n289 & n35262 ;
  assign n35264 = n14398 & ~n34652 ;
  assign n35265 = n30769 ^ n8835 ^ 1'b0 ;
  assign n35266 = n35264 | n35265 ;
  assign n35267 = n31012 ^ n1623 ^ 1'b0 ;
  assign n35268 = n3601 & ~n35267 ;
  assign n35269 = n11114 | n22631 ;
  assign n35270 = n23885 & ~n35269 ;
  assign n35271 = n35270 ^ n23534 ^ 1'b0 ;
  assign n35272 = ~n13138 & n35271 ;
  assign n35273 = ( n19025 & ~n24640 ) | ( n19025 & n25402 ) | ( ~n24640 & n25402 ) ;
  assign n35274 = n14955 & ~n25091 ;
  assign n35275 = n35274 ^ n10161 ^ 1'b0 ;
  assign n35276 = ( ~n907 & n4840 ) | ( ~n907 & n9237 ) | ( n4840 & n9237 ) ;
  assign n35277 = n7492 & ~n15485 ;
  assign n35278 = n9784 & n35277 ;
  assign n35279 = n2889 & n17178 ;
  assign n35280 = n35278 | n35279 ;
  assign n35281 = n19178 & ~n35280 ;
  assign n35282 = n35276 & ~n35281 ;
  assign n35283 = n608 | n5163 ;
  assign n35284 = n35283 ^ n3898 ^ 1'b0 ;
  assign n35285 = n35284 ^ n11578 ^ 1'b0 ;
  assign n35286 = n12556 ^ n3066 ^ 1'b0 ;
  assign n35287 = ~n35285 & n35286 ;
  assign n35288 = ~n3007 & n14558 ;
  assign n35289 = ~n840 & n25371 ;
  assign n35290 = n2067 & n4152 ;
  assign n35291 = n5252 & n35290 ;
  assign n35292 = n17602 & ~n35291 ;
  assign n35293 = n35292 ^ n4088 ^ 1'b0 ;
  assign n35294 = n30294 ^ n17473 ^ 1'b0 ;
  assign n35295 = n16154 ^ n12749 ^ 1'b0 ;
  assign n35296 = n23700 | n35295 ;
  assign n35297 = n13198 ^ n7558 ^ 1'b0 ;
  assign n35298 = n34211 ^ n12992 ^ 1'b0 ;
  assign n35299 = n7226 ^ x14 ^ 1'b0 ;
  assign n35300 = n29999 | n35299 ;
  assign n35301 = n3360 | n7028 ;
  assign n35302 = n1111 | n35301 ;
  assign n35303 = n5794 & n35302 ;
  assign n35304 = n35303 ^ n22113 ^ n21395 ;
  assign n35311 = ~n1151 & n13012 ;
  assign n35306 = n11371 & ~n11415 ;
  assign n35307 = n35306 ^ n17019 ^ 1'b0 ;
  assign n35308 = n18142 & n35307 ;
  assign n35305 = n8219 | n16519 ;
  assign n35309 = n35308 ^ n35305 ^ 1'b0 ;
  assign n35310 = n10004 | n35309 ;
  assign n35312 = n35311 ^ n35310 ^ 1'b0 ;
  assign n35313 = ( n4450 & ~n30840 ) | ( n4450 & n33894 ) | ( ~n30840 & n33894 ) ;
  assign n35314 = n31819 ^ n20573 ^ 1'b0 ;
  assign n35315 = n23586 ^ n3110 ^ 1'b0 ;
  assign n35316 = n2959 & ~n35315 ;
  assign n35317 = ~n26300 & n35316 ;
  assign n35318 = n35317 ^ n30952 ^ 1'b0 ;
  assign n35319 = n3225 & n18526 ;
  assign n35320 = n11450 ^ n1522 ^ 1'b0 ;
  assign n35321 = n4925 | n12670 ;
  assign n35322 = ~n26185 & n35321 ;
  assign n35323 = n2372 & ~n6581 ;
  assign n35324 = ~n35322 & n35323 ;
  assign n35325 = n17566 ^ n10239 ^ 1'b0 ;
  assign n35326 = n2624 & n9459 ;
  assign n35327 = n12278 & n35326 ;
  assign n35328 = n9958 | n31679 ;
  assign n35329 = n35328 ^ n1671 ^ 1'b0 ;
  assign n35330 = n35327 & n35329 ;
  assign n35331 = n28933 ^ n10010 ^ 1'b0 ;
  assign n35333 = n32582 ^ n7431 ^ n2317 ;
  assign n35332 = ~n5063 & n13392 ;
  assign n35334 = n35333 ^ n35332 ^ 1'b0 ;
  assign n35335 = n20826 | n35334 ;
  assign n35336 = n26413 | n35335 ;
  assign n35337 = n7359 & n35183 ;
  assign n35338 = n14811 ^ n14555 ^ 1'b0 ;
  assign n35339 = n24626 | n35338 ;
  assign n35340 = n35339 ^ n5994 ^ n2738 ;
  assign n35341 = n2516 & ~n20611 ;
  assign n35342 = n21187 ^ n18092 ^ 1'b0 ;
  assign n35343 = ~n6497 & n35342 ;
  assign n35344 = n982 & ~n26597 ;
  assign n35345 = ~n35343 & n35344 ;
  assign n35346 = n7707 | n29363 ;
  assign n35347 = n29734 ^ n7646 ^ 1'b0 ;
  assign n35348 = n35346 | n35347 ;
  assign n35349 = n6981 & n30592 ;
  assign n35350 = n7839 & ~n14067 ;
  assign n35351 = n16932 | n29214 ;
  assign n35352 = n7586 ^ n675 ^ 1'b0 ;
  assign n35353 = n35352 ^ n8340 ^ x154 ;
  assign n35354 = n31744 | n35353 ;
  assign n35355 = n19594 ^ n5456 ^ 1'b0 ;
  assign n35356 = n24273 | n35355 ;
  assign n35357 = n3081 | n34614 ;
  assign n35358 = n28454 & ~n35357 ;
  assign n35359 = ~n12273 & n35358 ;
  assign n35360 = n4210 ^ n2950 ^ 1'b0 ;
  assign n35361 = n35360 ^ n26161 ^ 1'b0 ;
  assign n35362 = n790 | n8504 ;
  assign n35363 = n3275 | n35362 ;
  assign n35364 = n8337 & ~n25632 ;
  assign n35365 = n21146 & n35364 ;
  assign n35366 = n35365 ^ n8298 ^ 1'b0 ;
  assign n35367 = n30059 ^ n277 ^ 1'b0 ;
  assign n35368 = n26560 ^ n11699 ^ 1'b0 ;
  assign n35369 = n4153 & n35368 ;
  assign n35370 = ~n12734 & n27126 ;
  assign n35371 = ~n35369 & n35370 ;
  assign n35372 = n21092 & n29232 ;
  assign n35373 = n35372 ^ n26069 ^ 1'b0 ;
  assign n35374 = n8130 ^ n3989 ^ 1'b0 ;
  assign n35375 = ~n3007 & n9034 ;
  assign n35376 = n13466 & n35375 ;
  assign n35377 = ~n30372 & n35376 ;
  assign n35378 = n6974 & ~n13472 ;
  assign n35379 = n17525 | n21448 ;
  assign n35380 = n22272 ^ n1223 ^ 1'b0 ;
  assign n35381 = n29533 & ~n35380 ;
  assign n35382 = ( ~n6119 & n25652 ) | ( ~n6119 & n34635 ) | ( n25652 & n34635 ) ;
  assign n35383 = n27331 ^ n5792 ^ 1'b0 ;
  assign n35384 = n6510 | n25365 ;
  assign n35385 = n29607 ^ n5835 ^ 1'b0 ;
  assign n35386 = n1839 & ~n9617 ;
  assign n35387 = n35386 ^ n9526 ^ 1'b0 ;
  assign n35388 = n7934 & n22235 ;
  assign n35389 = n9993 & n35388 ;
  assign n35390 = n1815 | n19688 ;
  assign n35391 = n35390 ^ n7094 ^ 1'b0 ;
  assign n35392 = ( n14236 & n14364 ) | ( n14236 & ~n15958 ) | ( n14364 & ~n15958 ) ;
  assign n35393 = n17430 | n35392 ;
  assign n35394 = n5589 ^ n1710 ^ 1'b0 ;
  assign n35395 = n4219 | n35394 ;
  assign n35396 = n10637 | n20902 ;
  assign n35397 = ~n20724 & n35396 ;
  assign n35398 = n14716 & ~n35397 ;
  assign n35399 = n1392 | n12013 ;
  assign n35400 = n35399 ^ n15564 ^ n2143 ;
  assign n35401 = n35400 ^ n17905 ^ 1'b0 ;
  assign n35402 = n24526 & n35401 ;
  assign n35403 = n6735 & ~n9578 ;
  assign n35404 = n35403 ^ n18262 ^ 1'b0 ;
  assign n35405 = n35404 ^ n13481 ^ n1528 ;
  assign n35406 = n35405 ^ n7219 ^ 1'b0 ;
  assign n35407 = ~n21592 & n35406 ;
  assign n35408 = n35407 ^ n15509 ^ 1'b0 ;
  assign n35409 = n15321 ^ n3362 ^ 1'b0 ;
  assign n35410 = n10247 | n17503 ;
  assign n35411 = n2242 & ~n35410 ;
  assign n35412 = n21371 & n35411 ;
  assign n35413 = n35409 & n35412 ;
  assign n35414 = ~n7166 & n18298 ;
  assign n35415 = n7166 & n35414 ;
  assign n35416 = n15644 | n35415 ;
  assign n35417 = n34177 ^ n4919 ^ 1'b0 ;
  assign n35418 = n3016 ^ n1554 ^ 1'b0 ;
  assign n35419 = n16150 ^ n10678 ^ 1'b0 ;
  assign n35420 = n2316 & ~n35419 ;
  assign n35421 = n35418 & n35420 ;
  assign n35422 = n2098 | n8627 ;
  assign n35423 = n10085 | n35422 ;
  assign n35424 = ~n9116 & n19719 ;
  assign n35425 = n5831 & ~n17648 ;
  assign n35426 = ~n18540 & n32334 ;
  assign n35427 = ~n30010 & n35426 ;
  assign n35428 = n24695 | n25763 ;
  assign n35429 = n35427 & ~n35428 ;
  assign n35430 = n8038 ^ n4131 ^ n3634 ;
  assign n35431 = ~n18703 & n35430 ;
  assign n35432 = ( n14042 & n20224 ) | ( n14042 & n32948 ) | ( n20224 & n32948 ) ;
  assign n35434 = n8157 & n20761 ;
  assign n35435 = n35434 ^ x249 ^ 1'b0 ;
  assign n35433 = n2226 | n18862 ;
  assign n35436 = n35435 ^ n35433 ^ 1'b0 ;
  assign n35437 = ~n11659 & n25066 ;
  assign n35438 = n35437 ^ n5650 ^ 1'b0 ;
  assign n35439 = n27256 ^ n22881 ^ 1'b0 ;
  assign n35440 = n9652 | n35439 ;
  assign n35441 = n2623 & ~n21628 ;
  assign n35442 = n35440 & n35441 ;
  assign n35443 = n10270 ^ n2944 ^ 1'b0 ;
  assign n35444 = ~n13671 & n35443 ;
  assign n35445 = n12148 & n35444 ;
  assign n35446 = n11585 & n35445 ;
  assign n35447 = n35446 ^ n672 ^ 1'b0 ;
  assign n35448 = n18120 ^ n2394 ^ 1'b0 ;
  assign n35449 = ~n8425 & n15273 ;
  assign n35450 = ~n35448 & n35449 ;
  assign n35451 = n27602 ^ n12552 ^ 1'b0 ;
  assign n35452 = n10870 | n35451 ;
  assign n35453 = n9630 & n9890 ;
  assign n35454 = n9259 & n18008 ;
  assign n35455 = n35454 ^ n35145 ^ 1'b0 ;
  assign n35456 = ~n35453 & n35455 ;
  assign n35457 = ~n8254 & n19986 ;
  assign n35458 = n12001 ^ n1707 ^ 1'b0 ;
  assign n35459 = n35457 & n35458 ;
  assign n35460 = n23846 ^ n5082 ^ 1'b0 ;
  assign n35461 = n15743 & n28952 ;
  assign n35462 = x208 & n8048 ;
  assign n35463 = n31236 ^ n20187 ^ 1'b0 ;
  assign n35464 = ~n1336 & n2679 ;
  assign n35465 = n1318 & n35464 ;
  assign n35466 = n35465 ^ n1716 ^ 1'b0 ;
  assign n35467 = n7800 & ~n12884 ;
  assign n35468 = ~n31858 & n33801 ;
  assign n35469 = n34252 & ~n35468 ;
  assign n35470 = n35469 ^ n9271 ^ 1'b0 ;
  assign n35471 = ( ~n19069 & n22775 ) | ( ~n19069 & n31647 ) | ( n22775 & n31647 ) ;
  assign n35472 = ~n3172 & n5339 ;
  assign n35473 = n20044 ^ n9670 ^ 1'b0 ;
  assign n35474 = n2580 & n17626 ;
  assign n35475 = n5097 & n35474 ;
  assign n35476 = n2209 | n35475 ;
  assign n35477 = n35476 ^ n12699 ^ 1'b0 ;
  assign n35478 = n17361 | n17852 ;
  assign n35479 = n35477 & ~n35478 ;
  assign n35480 = n11257 ^ x55 ^ 1'b0 ;
  assign n35481 = n3010 & n35480 ;
  assign n35482 = ~n5879 & n35481 ;
  assign n35483 = n31189 & n35482 ;
  assign n35484 = n11371 ^ n1447 ^ 1'b0 ;
  assign n35485 = n4575 & n35484 ;
  assign n35486 = n3260 & n35485 ;
  assign n35490 = n3508 | n27690 ;
  assign n35487 = n8704 ^ n1402 ^ 1'b0 ;
  assign n35488 = n8109 | n35487 ;
  assign n35489 = n18295 & ~n35488 ;
  assign n35491 = n35490 ^ n35489 ^ 1'b0 ;
  assign n35492 = n17968 ^ n1879 ^ 1'b0 ;
  assign n35493 = n35491 | n35492 ;
  assign n35494 = n35493 ^ n1428 ^ 1'b0 ;
  assign n35495 = n35486 & n35494 ;
  assign n35496 = ~n24024 & n35495 ;
  assign n35497 = n35496 ^ n31237 ^ 1'b0 ;
  assign n35498 = n8993 ^ n7447 ^ 1'b0 ;
  assign n35499 = n26527 ^ n21057 ^ n3685 ;
  assign n35500 = n35499 ^ n18213 ^ n4818 ;
  assign n35501 = n315 & ~n2065 ;
  assign n35502 = ( n5173 & n16393 ) | ( n5173 & n35501 ) | ( n16393 & n35501 ) ;
  assign n35503 = ~n2374 & n4824 ;
  assign n35504 = n35503 ^ n12978 ^ 1'b0 ;
  assign n35505 = ( n8728 & n11943 ) | ( n8728 & ~n30843 ) | ( n11943 & ~n30843 ) ;
  assign n35506 = n29851 ^ n29332 ^ n1671 ;
  assign n35507 = ( n4972 & ~n8808 ) | ( n4972 & n35506 ) | ( ~n8808 & n35506 ) ;
  assign n35509 = ~n6062 & n8781 ;
  assign n35510 = n30837 | n35509 ;
  assign n35508 = n1843 & ~n15783 ;
  assign n35511 = n35510 ^ n35508 ^ 1'b0 ;
  assign n35512 = n8666 & n10831 ;
  assign n35513 = n580 & n5508 ;
  assign n35514 = n14252 & n35513 ;
  assign n35515 = n35512 | n35514 ;
  assign n35516 = n13060 ^ n6311 ^ 1'b0 ;
  assign n35517 = n5463 ^ n1523 ^ 1'b0 ;
  assign n35518 = ~n17448 & n35517 ;
  assign n35519 = n7160 & ~n11612 ;
  assign n35520 = n17765 & n35519 ;
  assign n35521 = n35518 & ~n35520 ;
  assign n35522 = ~n17297 & n35521 ;
  assign n35523 = ~n14124 & n31044 ;
  assign n35524 = n35523 ^ n7605 ^ 1'b0 ;
  assign n35525 = ( n19235 & n31975 ) | ( n19235 & ~n35524 ) | ( n31975 & ~n35524 ) ;
  assign n35526 = ~n13541 & n18094 ;
  assign n35527 = n3041 & n35526 ;
  assign n35528 = n4818 ^ n2062 ^ 1'b0 ;
  assign n35529 = n16723 & ~n31174 ;
  assign n35530 = ~n628 & n35529 ;
  assign n35531 = ~n7538 & n16112 ;
  assign n35532 = n35531 ^ n3467 ^ 1'b0 ;
  assign n35533 = n13574 & ~n35532 ;
  assign n35534 = n1534 & n2736 ;
  assign n35535 = n35534 ^ n18948 ^ 1'b0 ;
  assign n35538 = ~n2491 & n6385 ;
  assign n35536 = n10614 & ~n14172 ;
  assign n35537 = ~n15774 & n35536 ;
  assign n35539 = n35538 ^ n35537 ^ 1'b0 ;
  assign n35540 = n29874 ^ n2741 ^ 1'b0 ;
  assign n35541 = n27599 ^ n15189 ^ 1'b0 ;
  assign n35542 = n24184 & ~n35541 ;
  assign n35543 = n6114 ^ n4815 ^ 1'b0 ;
  assign n35544 = n8325 & n34906 ;
  assign n35545 = n16920 | n21704 ;
  assign n35546 = n35545 ^ n4543 ^ 1'b0 ;
  assign n35547 = n30465 ^ n26539 ^ n5954 ;
  assign n35548 = n7796 & n12943 ;
  assign n35549 = n35547 & n35548 ;
  assign n35550 = ~n15492 & n35549 ;
  assign n35553 = n12778 & n19113 ;
  assign n35554 = n35553 ^ n18147 ^ 1'b0 ;
  assign n35551 = n18557 ^ n4568 ^ 1'b0 ;
  assign n35552 = n17483 | n35551 ;
  assign n35555 = n35554 ^ n35552 ^ 1'b0 ;
  assign n35556 = n6533 | n17578 ;
  assign n35557 = n935 & n16549 ;
  assign n35558 = n29538 & n35557 ;
  assign n35559 = n9252 | n26035 ;
  assign n35560 = n1492 ^ n634 ^ 1'b0 ;
  assign n35561 = n8471 & n35560 ;
  assign n35562 = n29568 ^ n17918 ^ n14674 ;
  assign n35563 = ~n3481 & n35562 ;
  assign n35564 = ~n35561 & n35563 ;
  assign n35565 = n20533 ^ n17449 ^ 1'b0 ;
  assign n35566 = ( n2312 & n12064 ) | ( n2312 & n17012 ) | ( n12064 & n17012 ) ;
  assign n35567 = n12625 ^ n1259 ^ 1'b0 ;
  assign n35568 = n14972 & ~n35567 ;
  assign n35569 = n3011 | n17701 ;
  assign n35570 = n8415 & n10356 ;
  assign n35571 = n22709 & n35570 ;
  assign n35572 = n14855 | n35571 ;
  assign n35573 = n26112 ^ n905 ^ 1'b0 ;
  assign n35574 = n35573 ^ n25512 ^ 1'b0 ;
  assign n35575 = n21612 & ~n35574 ;
  assign n35576 = n14612 | n24849 ;
  assign n35577 = n7884 & n35576 ;
  assign n35578 = n18904 ^ n18583 ^ n5154 ;
  assign n35579 = n12224 | n35578 ;
  assign n35580 = n25280 | n35579 ;
  assign n35581 = n6676 | n14565 ;
  assign n35582 = ( ~n3223 & n4903 ) | ( ~n3223 & n15509 ) | ( n4903 & n15509 ) ;
  assign n35583 = n35582 ^ n9447 ^ 1'b0 ;
  assign n35584 = n17509 | n35583 ;
  assign n35585 = ~n16073 & n18011 ;
  assign n35586 = n29586 & n35585 ;
  assign n35587 = n17621 & ~n21862 ;
  assign n35588 = n7867 | n35587 ;
  assign n35589 = n35588 ^ n1854 ^ 1'b0 ;
  assign n35590 = n4271 & n9391 ;
  assign n35591 = n35590 ^ n24226 ^ 1'b0 ;
  assign n35592 = n15488 ^ n8796 ^ 1'b0 ;
  assign n35593 = n35591 & ~n35592 ;
  assign n35594 = n6916 | n19339 ;
  assign n35595 = n35594 ^ n15278 ^ 1'b0 ;
  assign n35596 = ~n4660 & n11609 ;
  assign n35597 = n35596 ^ n14463 ^ 1'b0 ;
  assign n35598 = n25374 & n33914 ;
  assign n35599 = n35598 ^ n27539 ^ 1'b0 ;
  assign n35600 = n308 | n10726 ;
  assign n35601 = n35600 ^ n8710 ^ 1'b0 ;
  assign n35602 = n7722 & n35601 ;
  assign n35603 = n9310 & ~n29456 ;
  assign n35604 = n35603 ^ n29364 ^ 1'b0 ;
  assign n35605 = ( n3959 & n19521 ) | ( n3959 & n35604 ) | ( n19521 & n35604 ) ;
  assign n35606 = n9161 ^ n1913 ^ 1'b0 ;
  assign n35607 = n35606 ^ n3157 ^ 1'b0 ;
  assign n35608 = ~n7188 & n23097 ;
  assign n35609 = ~n8082 & n35608 ;
  assign n35610 = n5282 & n35609 ;
  assign n35611 = n14337 ^ n1151 ^ 1'b0 ;
  assign n35612 = n35611 ^ n24422 ^ 1'b0 ;
  assign n35613 = ~n19785 & n35612 ;
  assign n35614 = x77 & n16149 ;
  assign n35615 = n35614 ^ n18450 ^ 1'b0 ;
  assign n35616 = ~n10000 & n10377 ;
  assign n35617 = n35616 ^ n6789 ^ 1'b0 ;
  assign n35618 = n7597 & ~n35617 ;
  assign n35619 = ( n28804 & ~n30917 ) | ( n28804 & n35618 ) | ( ~n30917 & n35618 ) ;
  assign n35620 = n17805 ^ n1129 ^ 1'b0 ;
  assign n35621 = n23545 | n25294 ;
  assign n35622 = n35620 & ~n35621 ;
  assign n35623 = ~n14952 & n19650 ;
  assign n35624 = n4321 & n35623 ;
  assign n35625 = ~n17263 & n22901 ;
  assign n35626 = ~n15463 & n35625 ;
  assign n35627 = n35626 ^ n14032 ^ n6687 ;
  assign n35628 = n10430 | n29494 ;
  assign n35629 = n31777 ^ n8674 ^ 1'b0 ;
  assign n35630 = ( x72 & n4993 ) | ( x72 & ~n31079 ) | ( n4993 & ~n31079 ) ;
  assign n35631 = n11053 & n35630 ;
  assign n35632 = n3177 & n14075 ;
  assign n35633 = ~n638 & n20939 ;
  assign n35634 = ~n35632 & n35633 ;
  assign n35635 = n19201 ^ n7737 ^ 1'b0 ;
  assign n35636 = n29423 ^ n7387 ^ 1'b0 ;
  assign n35637 = n32194 ^ n10690 ^ n3679 ;
  assign n35638 = n16503 & ~n35637 ;
  assign n35639 = n3686 | n10900 ;
  assign n35640 = n6388 & n11010 ;
  assign n35641 = n35640 ^ n15128 ^ 1'b0 ;
  assign n35642 = n24501 ^ n867 ^ 1'b0 ;
  assign n35643 = n35641 | n35642 ;
  assign n35644 = ~n11613 & n12120 ;
  assign n35645 = n14879 ^ n4802 ^ 1'b0 ;
  assign n35646 = ( n2029 & n33385 ) | ( n2029 & n35645 ) | ( n33385 & n35645 ) ;
  assign n35647 = n8323 & ~n31664 ;
  assign n35648 = n31355 ^ n2231 ^ 1'b0 ;
  assign n35649 = n17520 & n35648 ;
  assign n35650 = n25267 ^ n8298 ^ 1'b0 ;
  assign n35651 = x82 & ~n6761 ;
  assign n35652 = n35651 ^ n11265 ^ 1'b0 ;
  assign n35653 = n9057 ^ n5105 ^ n4910 ;
  assign n35654 = n35653 ^ n7141 ^ n3640 ;
  assign n35655 = n7958 & ~n12894 ;
  assign n35656 = n35655 ^ n1896 ^ 1'b0 ;
  assign n35657 = n2016 & n10010 ;
  assign n35658 = n34926 ^ n3184 ^ 1'b0 ;
  assign n35659 = n9067 & ~n35658 ;
  assign n35660 = n4261 & n14818 ;
  assign n35661 = ~n16384 & n35660 ;
  assign n35662 = n3377 & n14634 ;
  assign n35663 = n35662 ^ n3360 ^ 1'b0 ;
  assign n35664 = x45 & ~n6970 ;
  assign n35665 = n35664 ^ n7028 ^ 1'b0 ;
  assign n35666 = ~n29487 & n35665 ;
  assign n35667 = ~n35663 & n35666 ;
  assign n35668 = n22879 ^ n7433 ^ 1'b0 ;
  assign n35669 = n30424 & ~n35668 ;
  assign n35670 = n19956 ^ n12068 ^ n10514 ;
  assign n35671 = ~n444 & n35670 ;
  assign n35672 = ( n20150 & n35669 ) | ( n20150 & ~n35671 ) | ( n35669 & ~n35671 ) ;
  assign n35673 = n35402 ^ n30725 ^ 1'b0 ;
  assign n35674 = n3420 & ~n26473 ;
  assign n35675 = n28930 & n35674 ;
  assign n35676 = n1153 & ~n8022 ;
  assign n35677 = n35676 ^ n2252 ^ 1'b0 ;
  assign n35678 = n2925 | n26888 ;
  assign n35679 = n19885 | n30372 ;
  assign n35680 = n27786 & ~n35679 ;
  assign n35681 = n32462 ^ n31331 ^ 1'b0 ;
  assign n35682 = n6046 | n35681 ;
  assign n35683 = ~n16969 & n35682 ;
  assign n35684 = n17226 ^ n2020 ^ 1'b0 ;
  assign n35685 = n22487 ^ n11982 ^ 1'b0 ;
  assign n35686 = ( n29040 & n35684 ) | ( n29040 & n35685 ) | ( n35684 & n35685 ) ;
  assign n35687 = n10244 & n29241 ;
  assign n35688 = n24416 & n35318 ;
  assign n35689 = n35688 ^ n32499 ^ 1'b0 ;
  assign n35690 = ( n5497 & n6010 ) | ( n5497 & n6632 ) | ( n6010 & n6632 ) ;
  assign n35691 = n35690 ^ n15255 ^ 1'b0 ;
  assign n35692 = ~n6646 & n21701 ;
  assign n35693 = n15492 & ~n35692 ;
  assign n35694 = ~n8867 & n35693 ;
  assign n35695 = n33147 ^ n4256 ^ 1'b0 ;
  assign n35696 = n35694 | n35695 ;
  assign n35697 = n35696 ^ n16897 ^ 1'b0 ;
  assign n35698 = n1735 & n35697 ;
  assign n35699 = n15639 & n24595 ;
  assign n35700 = x47 & ~n1591 ;
  assign n35701 = ( n12636 & n35699 ) | ( n12636 & n35700 ) | ( n35699 & n35700 ) ;
  assign n35702 = ( n9104 & ~n11627 ) | ( n9104 & n29220 ) | ( ~n11627 & n29220 ) ;
  assign n35703 = n5650 | n35702 ;
  assign n35704 = n35703 ^ n12268 ^ 1'b0 ;
  assign n35705 = n7809 & ~n13630 ;
  assign n35706 = n35705 ^ n19575 ^ 1'b0 ;
  assign n35707 = n3873 | n35706 ;
  assign n35708 = n5152 & n11913 ;
  assign n35709 = n16231 ^ n14836 ^ n1853 ;
  assign n35710 = n35709 ^ n5301 ^ 1'b0 ;
  assign n35711 = n35708 | n35710 ;
  assign n35712 = n25618 | n35711 ;
  assign n35713 = n3288 & ~n4003 ;
  assign n35714 = n5406 & n35573 ;
  assign n35715 = n35714 ^ n4033 ^ 1'b0 ;
  assign n35716 = n11755 & ~n35212 ;
  assign n35717 = n15834 & n35716 ;
  assign n35718 = n21077 | n34552 ;
  assign n35719 = ~n26076 & n26758 ;
  assign n35720 = n35719 ^ n7601 ^ 1'b0 ;
  assign n35721 = n1748 & n16257 ;
  assign n35722 = n35418 & n35721 ;
  assign n35723 = n416 & ~n13647 ;
  assign n35724 = ~n13288 & n35723 ;
  assign n35725 = n35724 ^ n18513 ^ 1'b0 ;
  assign n35726 = n35725 ^ n33130 ^ n471 ;
  assign n35727 = n17279 ^ n15564 ^ 1'b0 ;
  assign n35728 = n7819 ^ n5619 ^ 1'b0 ;
  assign n35729 = n35728 ^ n23155 ^ 1'b0 ;
  assign n35730 = ~n8331 & n12829 ;
  assign n35731 = ~n20530 & n35730 ;
  assign n35732 = n4895 & n9944 ;
  assign n35733 = n2848 & n35732 ;
  assign n35734 = n10826 & n35733 ;
  assign n35735 = n649 & ~n971 ;
  assign n35736 = n17145 ^ n17075 ^ n12281 ;
  assign n35737 = n26738 ^ n14964 ^ n2995 ;
  assign n35738 = n7113 & ~n21363 ;
  assign n35739 = ~n35737 & n35738 ;
  assign n35740 = n12400 | n35739 ;
  assign n35741 = n35740 ^ n725 ^ 1'b0 ;
  assign n35742 = n449 & n23567 ;
  assign n35743 = n5192 & ~n14296 ;
  assign n35744 = n9481 ^ n7518 ^ 1'b0 ;
  assign n35745 = ~n13242 & n35744 ;
  assign n35747 = n8018 & ~n24215 ;
  assign n35746 = n4400 & ~n20387 ;
  assign n35748 = n35747 ^ n35746 ^ 1'b0 ;
  assign n35749 = n3935 | n35748 ;
  assign n35750 = ~n335 & n28716 ;
  assign n35751 = n35750 ^ n9479 ^ 1'b0 ;
  assign n35752 = n11299 & n19213 ;
  assign n35753 = n35752 ^ n29379 ^ 1'b0 ;
  assign n35754 = n11290 & ~n11776 ;
  assign n35763 = ~n821 & n1064 ;
  assign n35762 = n2875 & n12120 ;
  assign n35764 = n35763 ^ n35762 ^ 1'b0 ;
  assign n35757 = n4138 ^ n1259 ^ 1'b0 ;
  assign n35758 = n4565 & n35757 ;
  assign n35755 = n9031 ^ n1851 ^ 1'b0 ;
  assign n35756 = n35755 ^ n5362 ^ 1'b0 ;
  assign n35759 = n35758 ^ n35756 ^ 1'b0 ;
  assign n35760 = n29377 | n35759 ;
  assign n35761 = n22552 & ~n35760 ;
  assign n35765 = n35764 ^ n35761 ^ 1'b0 ;
  assign n35766 = n14229 & ~n16068 ;
  assign n35767 = ~n16699 & n22764 ;
  assign n35768 = ~n10250 & n35767 ;
  assign n35769 = n12642 & n19668 ;
  assign n35770 = n35769 ^ n14057 ^ 1'b0 ;
  assign n35771 = n35770 ^ n19832 ^ n7985 ;
  assign n35772 = ~n24009 & n35771 ;
  assign n35773 = ~n5278 & n35772 ;
  assign n35774 = n8990 & ~n15773 ;
  assign n35775 = n35774 ^ n9200 ^ 1'b0 ;
  assign n35776 = ( n2119 & ~n10208 ) | ( n2119 & n35775 ) | ( ~n10208 & n35775 ) ;
  assign n35777 = n20838 & n35776 ;
  assign n35778 = ~n8547 & n15235 ;
  assign n35779 = n4290 & n35778 ;
  assign n35780 = n4916 & n7617 ;
  assign n35781 = n23943 & ~n35780 ;
  assign n35782 = n35779 & n35781 ;
  assign n35783 = n11365 & ~n21523 ;
  assign n35784 = n5878 | n7239 ;
  assign n35785 = n35784 ^ n5746 ^ 1'b0 ;
  assign n35786 = ( n3696 & ~n8053 ) | ( n3696 & n35785 ) | ( ~n8053 & n35785 ) ;
  assign n35787 = n2516 ^ n1867 ^ 1'b0 ;
  assign n35788 = n5396 & ~n14317 ;
  assign n35795 = n2026 & ~n5326 ;
  assign n35790 = ( ~n5611 & n15196 ) | ( ~n5611 & n30599 ) | ( n15196 & n30599 ) ;
  assign n35791 = n35790 ^ n7850 ^ 1'b0 ;
  assign n35792 = ~n9045 & n35791 ;
  assign n35789 = n14994 & ~n21426 ;
  assign n35793 = n35792 ^ n35789 ^ 1'b0 ;
  assign n35794 = n23229 & ~n35793 ;
  assign n35796 = n35795 ^ n35794 ^ 1'b0 ;
  assign n35797 = n5893 & ~n13144 ;
  assign n35798 = ~n19110 & n24292 ;
  assign n35799 = n35798 ^ n17519 ^ 1'b0 ;
  assign n35800 = n9224 & n21928 ;
  assign n35802 = n2606 & ~n2984 ;
  assign n35801 = ( n1081 & ~n7568 ) | ( n1081 & n13691 ) | ( ~n7568 & n13691 ) ;
  assign n35803 = n35802 ^ n35801 ^ 1'b0 ;
  assign n35804 = n35803 ^ n33208 ^ n2533 ;
  assign n35805 = n31549 ^ n17073 ^ n8192 ;
  assign n35808 = n3515 | n14272 ;
  assign n35806 = n8633 & ~n18343 ;
  assign n35807 = ~n6370 & n35806 ;
  assign n35809 = n35808 ^ n35807 ^ 1'b0 ;
  assign n35810 = ( ~n9207 & n18894 ) | ( ~n9207 & n20485 ) | ( n18894 & n20485 ) ;
  assign n35811 = n18935 | n21268 ;
  assign n35812 = n445 & ~n16489 ;
  assign n35813 = ~n35811 & n35812 ;
  assign n35814 = n3845 | n7056 ;
  assign n35815 = n10349 | n35814 ;
  assign n35816 = n35815 ^ n18433 ^ n9607 ;
  assign n35817 = n16615 | n23725 ;
  assign n35818 = n5692 & ~n24349 ;
  assign n35819 = n14760 & n24000 ;
  assign n35820 = ~n5442 & n20878 ;
  assign n35821 = n35820 ^ n9630 ^ 1'b0 ;
  assign n35822 = ~n19204 & n35821 ;
  assign n35823 = n35822 ^ n25684 ^ 1'b0 ;
  assign n35824 = ~n1846 & n13003 ;
  assign n35825 = n2821 & ~n9036 ;
  assign n35826 = n12967 | n29480 ;
  assign n35827 = n22334 ^ n4172 ^ 1'b0 ;
  assign n35828 = ~n24399 & n35827 ;
  assign n35829 = ( x129 & n8993 ) | ( x129 & n26418 ) | ( n8993 & n26418 ) ;
  assign n35830 = n35828 & ~n35829 ;
  assign n35831 = ~n5237 & n6952 ;
  assign n35832 = n35831 ^ n15758 ^ 1'b0 ;
  assign n35833 = n35830 & ~n35832 ;
  assign n35834 = n17091 & n30729 ;
  assign n35835 = ~x78 & n35834 ;
  assign n35836 = n9930 ^ n2301 ^ 1'b0 ;
  assign n35837 = n28362 & ~n35836 ;
  assign n35838 = n3542 & n12812 ;
  assign n35839 = n22123 | n35838 ;
  assign n35840 = n35839 ^ x88 ^ 1'b0 ;
  assign n35841 = n22336 ^ n10333 ^ 1'b0 ;
  assign n35842 = ~n17167 & n35841 ;
  assign n35843 = n7358 & n35183 ;
  assign n35844 = ~n8092 & n8915 ;
  assign n35845 = n4696 & ~n25239 ;
  assign n35846 = ~n35515 & n35845 ;
  assign n35847 = n13468 ^ n1501 ^ 1'b0 ;
  assign n35848 = ~n23681 & n35847 ;
  assign n35849 = n420 & n28840 ;
  assign n35850 = n4657 & n35849 ;
  assign n35851 = ~n1912 & n12359 ;
  assign n35852 = n35851 ^ n31760 ^ 1'b0 ;
  assign n35853 = n29546 & n35852 ;
  assign n35854 = ~n2070 & n17308 ;
  assign n35856 = n11313 | n16473 ;
  assign n35857 = n35856 ^ n5362 ^ 1'b0 ;
  assign n35855 = n10869 ^ n1161 ^ n786 ;
  assign n35858 = n35857 ^ n35855 ^ n19959 ;
  assign n35859 = ( n7266 & n12646 ) | ( n7266 & n22758 ) | ( n12646 & n22758 ) ;
  assign n35860 = n16674 & ~n34510 ;
  assign n35861 = n34964 & n35860 ;
  assign n35862 = n10158 ^ n1620 ^ 1'b0 ;
  assign n35863 = n10897 & n35862 ;
  assign n35864 = n35863 ^ n19923 ^ 1'b0 ;
  assign n35865 = n20667 & ~n20937 ;
  assign n35866 = n35865 ^ n10133 ^ 1'b0 ;
  assign n35867 = ~n823 & n17659 ;
  assign n35868 = n35867 ^ n9162 ^ 1'b0 ;
  assign n35869 = n7462 & ~n35868 ;
  assign n35870 = n22987 | n35869 ;
  assign n35871 = n28225 | n35870 ;
  assign n35872 = ~n382 & n17768 ;
  assign n35873 = n35872 ^ n17508 ^ 1'b0 ;
  assign n35874 = n35873 ^ n33460 ^ 1'b0 ;
  assign n35875 = ( ~n15125 & n29391 ) | ( ~n15125 & n35874 ) | ( n29391 & n35874 ) ;
  assign n35876 = n9532 & n35875 ;
  assign n35877 = n35876 ^ n5722 ^ 1'b0 ;
  assign n35878 = n33350 ^ n5363 ^ 1'b0 ;
  assign n35879 = n6146 & ~n10374 ;
  assign n35880 = n10374 & n35879 ;
  assign n35881 = n20211 | n35880 ;
  assign n35882 = n35880 & ~n35881 ;
  assign n35883 = ~n959 & n11091 ;
  assign n35884 = n35882 & n35883 ;
  assign n35885 = n35884 ^ n21695 ^ n11383 ;
  assign n35886 = ~n4122 & n23451 ;
  assign n35887 = ~n15874 & n17641 ;
  assign n35888 = n35887 ^ n6597 ^ 1'b0 ;
  assign n35889 = ~n35886 & n35888 ;
  assign n35890 = ~n661 & n3826 ;
  assign n35893 = ~n1570 & n14507 ;
  assign n35891 = n29805 ^ n10944 ^ 1'b0 ;
  assign n35892 = x61 & ~n35891 ;
  assign n35894 = n35893 ^ n35892 ^ n7197 ;
  assign n35895 = ~n14185 & n21320 ;
  assign n35896 = n11447 & n35895 ;
  assign n35897 = n33936 ^ n32732 ^ 1'b0 ;
  assign n35898 = n14236 ^ n3689 ^ 1'b0 ;
  assign n35899 = n18793 & n21904 ;
  assign n35901 = n8499 & ~n24519 ;
  assign n35900 = ~n18082 & n22277 ;
  assign n35902 = n35901 ^ n35900 ^ 1'b0 ;
  assign n35903 = ( n14821 & n30191 ) | ( n14821 & ~n35902 ) | ( n30191 & ~n35902 ) ;
  assign n35904 = n7491 ^ n7204 ^ n4165 ;
  assign n35905 = n35904 ^ n436 ^ 1'b0 ;
  assign n35906 = n35905 ^ n23295 ^ n13789 ;
  assign n35907 = ~n18746 & n33676 ;
  assign n35908 = n724 | n17410 ;
  assign n35909 = n7648 & ~n14206 ;
  assign n35910 = ~n8184 & n35909 ;
  assign n35911 = n19974 | n35910 ;
  assign n35912 = n35911 ^ n365 ^ 1'b0 ;
  assign n35913 = n9742 | n33997 ;
  assign n35914 = n1824 & ~n8185 ;
  assign n35915 = n33806 ^ n13738 ^ 1'b0 ;
  assign n35916 = n29911 & n35915 ;
  assign n35917 = n3619 & ~n9134 ;
  assign n35918 = ~n6849 & n35917 ;
  assign n35919 = n1742 & ~n8520 ;
  assign n35920 = n3640 & n35919 ;
  assign n35921 = n32775 ^ n15615 ^ 1'b0 ;
  assign n35922 = ~n35920 & n35921 ;
  assign n35923 = n35918 | n35922 ;
  assign n35924 = n26539 | n30792 ;
  assign n35925 = n22469 ^ n8717 ^ 1'b0 ;
  assign n35926 = n3686 | n18726 ;
  assign n35927 = n31688 ^ n29391 ^ 1'b0 ;
  assign n35928 = n1997 | n35927 ;
  assign n35930 = n4239 ^ n1632 ^ 1'b0 ;
  assign n35929 = n4386 & ~n10205 ;
  assign n35931 = n35930 ^ n35929 ^ 1'b0 ;
  assign n35932 = n32360 | n32676 ;
  assign n35933 = n23493 ^ n547 ^ 1'b0 ;
  assign n35934 = n1413 & n35933 ;
  assign n35935 = n22615 ^ x188 ^ 1'b0 ;
  assign n35936 = n4449 & ~n35935 ;
  assign n35937 = n28845 ^ n1183 ^ 1'b0 ;
  assign n35938 = n8487 | n35937 ;
  assign n35939 = n13254 & n14435 ;
  assign n35940 = n35939 ^ n22079 ^ 1'b0 ;
  assign n35941 = ~n4187 & n35940 ;
  assign n35942 = n35941 ^ n24885 ^ 1'b0 ;
  assign n35943 = n13686 ^ n637 ^ 1'b0 ;
  assign n35944 = n2533 & ~n35943 ;
  assign n35945 = n35944 ^ n3996 ^ n2343 ;
  assign n35946 = n35942 & ~n35945 ;
  assign n35947 = ( n7643 & ~n13424 ) | ( n7643 & n28638 ) | ( ~n13424 & n28638 ) ;
  assign n35948 = n11576 | n35947 ;
  assign n35949 = n35946 | n35948 ;
  assign n35950 = n711 | n17345 ;
  assign n35951 = n13466 & ~n35950 ;
  assign n35952 = n35951 ^ n11583 ^ 1'b0 ;
  assign n35953 = n4905 | n23859 ;
  assign n35954 = n12427 | n35953 ;
  assign n35955 = n35954 ^ n34043 ^ 1'b0 ;
  assign n35956 = n33200 ^ n30972 ^ 1'b0 ;
  assign n35957 = n5231 & ~n35956 ;
  assign n35958 = ~n12014 & n13834 ;
  assign n35959 = n35958 ^ n13204 ^ 1'b0 ;
  assign n35960 = n16609 & n32278 ;
  assign n35961 = n35960 ^ n15279 ^ 1'b0 ;
  assign n35962 = n5494 | n35961 ;
  assign n35963 = n13827 & ~n35962 ;
  assign n35964 = n13424 ^ n12586 ^ 1'b0 ;
  assign n35965 = n17825 | n35964 ;
  assign n35966 = n21926 | n34441 ;
  assign n35967 = n9998 ^ n4202 ^ 1'b0 ;
  assign n35968 = ~n5900 & n35967 ;
  assign n35969 = n18829 & n35968 ;
  assign n35970 = n8220 ^ x215 ^ x30 ;
  assign n35971 = n3088 & n25150 ;
  assign n35972 = n35970 | n35971 ;
  assign n35973 = n33739 | n35972 ;
  assign n35974 = n33490 ^ n23450 ^ 1'b0 ;
  assign n35975 = n9539 ^ n5229 ^ 1'b0 ;
  assign n35976 = ~n2566 & n35975 ;
  assign n35977 = n17316 ^ n8011 ^ n4269 ;
  assign n35978 = n1397 | n35977 ;
  assign n35979 = n35978 ^ n21227 ^ 1'b0 ;
  assign n35980 = n4739 & ~n35979 ;
  assign n35981 = n26738 ^ n20835 ^ n8234 ;
  assign n35982 = n8167 | n35981 ;
  assign n35983 = n34056 | n35982 ;
  assign n35984 = n20089 ^ n17025 ^ 1'b0 ;
  assign n35985 = n35983 & ~n35984 ;
  assign n35986 = n15123 ^ n779 ^ 1'b0 ;
  assign n35987 = n23386 ^ n12948 ^ 1'b0 ;
  assign n35988 = ( n1433 & n29081 ) | ( n1433 & n35987 ) | ( n29081 & n35987 ) ;
  assign n35989 = n10765 & n24385 ;
  assign n35990 = n19722 ^ n15418 ^ 1'b0 ;
  assign n35991 = n22199 & ~n35990 ;
  assign n35992 = n6207 & n32278 ;
  assign n35993 = ~x70 & n17538 ;
  assign n35994 = n35993 ^ n17748 ^ 1'b0 ;
  assign n35995 = n32744 | n35994 ;
  assign n35996 = n10472 & ~n30443 ;
  assign n35997 = ~n6847 & n12068 ;
  assign n35998 = n35997 ^ n25122 ^ n1120 ;
  assign n35999 = n20435 ^ n15042 ^ 1'b0 ;
  assign n36000 = n32703 & ~n35999 ;
  assign n36001 = n36000 ^ n1796 ^ 1'b0 ;
  assign n36002 = n34948 ^ n1525 ^ 1'b0 ;
  assign n36003 = n25570 ^ n13946 ^ 1'b0 ;
  assign n36004 = n2375 | n18352 ;
  assign n36005 = n36004 ^ n14641 ^ 1'b0 ;
  assign n36006 = n35129 ^ n7107 ^ 1'b0 ;
  assign n36007 = n36005 & ~n36006 ;
  assign n36008 = n8371 & n36007 ;
  assign n36009 = ~n12597 & n12655 ;
  assign n36010 = n36009 ^ n25290 ^ 1'b0 ;
  assign n36011 = n2476 ^ n369 ^ 1'b0 ;
  assign n36012 = n10931 & n36011 ;
  assign n36013 = n36012 ^ n15975 ^ 1'b0 ;
  assign n36014 = n34481 & n36013 ;
  assign n36015 = n2915 & ~n7318 ;
  assign n36016 = n36015 ^ n8395 ^ 1'b0 ;
  assign n36017 = n28794 | n36016 ;
  assign n36018 = n25426 ^ n19287 ^ 1'b0 ;
  assign n36019 = n36017 | n36018 ;
  assign n36020 = n5221 ^ n5181 ^ 1'b0 ;
  assign n36021 = n2396 & n36020 ;
  assign n36022 = ~n13230 & n36021 ;
  assign n36023 = n1300 & ~n12224 ;
  assign n36024 = n5799 | n20279 ;
  assign n36031 = n7285 ^ n2231 ^ 1'b0 ;
  assign n36030 = ~n12867 & n26746 ;
  assign n36032 = n36031 ^ n36030 ^ 1'b0 ;
  assign n36027 = n15437 ^ n12569 ^ 1'b0 ;
  assign n36025 = n1856 & n18528 ;
  assign n36026 = n10068 & ~n36025 ;
  assign n36028 = n36027 ^ n36026 ^ 1'b0 ;
  assign n36029 = n21651 & n36028 ;
  assign n36033 = n36032 ^ n36029 ^ n3302 ;
  assign n36034 = ~n1660 & n18629 ;
  assign n36035 = n36034 ^ n14218 ^ 1'b0 ;
  assign n36036 = n15255 & ~n22272 ;
  assign n36037 = n36036 ^ n886 ^ 1'b0 ;
  assign n36038 = n36037 ^ n35045 ^ 1'b0 ;
  assign n36039 = ~n4830 & n14900 ;
  assign n36040 = ~n581 & n36039 ;
  assign n36041 = n7373 & ~n27470 ;
  assign n36042 = n36040 & n36041 ;
  assign n36043 = ~n9452 & n13261 ;
  assign n36044 = n26236 ^ n2083 ^ 1'b0 ;
  assign n36045 = n36043 | n36044 ;
  assign n36046 = n36045 ^ n29996 ^ 1'b0 ;
  assign n36047 = n19822 ^ n5611 ^ n1977 ;
  assign n36048 = n11569 ^ n9803 ^ 1'b0 ;
  assign n36049 = n15020 | n36048 ;
  assign n36050 = ( n9806 & ~n36047 ) | ( n9806 & n36049 ) | ( ~n36047 & n36049 ) ;
  assign n36051 = n2199 | n29602 ;
  assign n36052 = n618 | n27200 ;
  assign n36053 = n36052 ^ n22485 ^ 1'b0 ;
  assign n36054 = ~n2225 & n25863 ;
  assign n36055 = n365 | n8832 ;
  assign n36056 = n16467 | n36055 ;
  assign n36057 = n9841 & n36056 ;
  assign n36058 = n9393 & n36057 ;
  assign n36059 = n10709 & n13778 ;
  assign n36060 = n36059 ^ n33578 ^ 1'b0 ;
  assign n36061 = n3634 & ~n12987 ;
  assign n36062 = n31768 ^ n5100 ^ 1'b0 ;
  assign n36063 = n4799 & ~n36062 ;
  assign n36064 = n8580 & n13068 ;
  assign n36065 = n10389 & ~n17981 ;
  assign n36066 = n36065 ^ n23994 ^ 1'b0 ;
  assign n36067 = n6151 & ~n25593 ;
  assign n36068 = n35907 ^ n33073 ^ 1'b0 ;
  assign n36069 = ~n7855 & n36068 ;
  assign n36070 = n24909 ^ n3014 ^ 1'b0 ;
  assign n36071 = x144 & n36070 ;
  assign n36072 = n14405 ^ n6992 ^ 1'b0 ;
  assign n36073 = n36071 & n36072 ;
  assign n36074 = n9930 ^ n2443 ^ 1'b0 ;
  assign n36075 = ~n4055 & n36074 ;
  assign n36076 = ~n9416 & n36075 ;
  assign n36077 = ~n6187 & n26814 ;
  assign n36078 = x57 & n914 ;
  assign n36079 = n1682 & ~n36078 ;
  assign n36080 = n9336 & n36079 ;
  assign n36082 = n9504 ^ n2369 ^ n1103 ;
  assign n36081 = n6974 | n20603 ;
  assign n36083 = n36082 ^ n36081 ^ 1'b0 ;
  assign n36084 = n36083 ^ n7384 ^ 1'b0 ;
  assign n36085 = ~n3007 & n16252 ;
  assign n36086 = n12605 ^ n4657 ^ x156 ;
  assign n36087 = n36086 ^ n26633 ^ n19411 ;
  assign n36088 = n36087 ^ n28101 ^ 1'b0 ;
  assign n36089 = n2098 ^ n1960 ^ 1'b0 ;
  assign n36090 = n9144 & n18847 ;
  assign n36091 = ~n17471 & n29757 ;
  assign n36092 = n19439 ^ n7666 ^ 1'b0 ;
  assign n36093 = n15057 | n36092 ;
  assign n36094 = n2362 | n9995 ;
  assign n36095 = n11386 ^ n5432 ^ 1'b0 ;
  assign n36096 = n36094 & n36095 ;
  assign n36097 = n34460 ^ n1290 ^ 1'b0 ;
  assign n36098 = n36096 & n36097 ;
  assign n36099 = ( n4331 & n9967 ) | ( n4331 & n11147 ) | ( n9967 & n11147 ) ;
  assign n36101 = n1795 & ~n8236 ;
  assign n36100 = ~n12902 & n20776 ;
  assign n36102 = n36101 ^ n36100 ^ n20407 ;
  assign n36103 = n9501 & n36102 ;
  assign n36104 = n13401 & n19916 ;
  assign n36105 = n36104 ^ n3851 ^ 1'b0 ;
  assign n36106 = n24628 ^ n20081 ^ 1'b0 ;
  assign n36107 = n26742 ^ n24484 ^ 1'b0 ;
  assign n36108 = n5105 & ~n36107 ;
  assign n36109 = n7799 & n36108 ;
  assign n36110 = n16137 ^ n8893 ^ 1'b0 ;
  assign n36111 = n29036 ^ n12935 ^ 1'b0 ;
  assign n36112 = n36110 & ~n36111 ;
  assign n36113 = n13635 & ~n29631 ;
  assign n36114 = n23567 | n35829 ;
  assign n36115 = n12471 & n19139 ;
  assign n36116 = n36115 ^ n32813 ^ 1'b0 ;
  assign n36117 = n18784 & ~n20079 ;
  assign n36118 = n3868 | n14557 ;
  assign n36119 = n36118 ^ n23328 ^ 1'b0 ;
  assign n36120 = ~n22532 & n36119 ;
  assign n36121 = n9638 & ~n30292 ;
  assign n36122 = n36121 ^ n23463 ^ 1'b0 ;
  assign n36123 = n22338 ^ n20916 ^ 1'b0 ;
  assign n36124 = n22537 ^ n15065 ^ 1'b0 ;
  assign n36125 = n30756 ^ n15577 ^ 1'b0 ;
  assign n36126 = ~n357 & n25990 ;
  assign n36127 = n36126 ^ n17566 ^ n13469 ;
  assign n36128 = n14998 ^ n6341 ^ n3508 ;
  assign n36129 = ~n8493 & n36128 ;
  assign n36130 = n36127 & n36129 ;
  assign n36131 = n4491 & ~n15097 ;
  assign n36132 = n2959 & n9552 ;
  assign n36133 = n36132 ^ n8131 ^ 1'b0 ;
  assign n36134 = ~n1048 & n20838 ;
  assign n36135 = n36134 ^ n6037 ^ 1'b0 ;
  assign n36136 = n30825 & n36135 ;
  assign n36137 = n3588 & n36136 ;
  assign n36138 = n29553 & ~n30078 ;
  assign n36139 = n4216 & ~n30846 ;
  assign n36140 = n8904 & n9266 ;
  assign n36141 = n5900 | n7293 ;
  assign n36142 = n36141 ^ n27230 ^ n7382 ;
  assign n36143 = ~n2041 & n36142 ;
  assign n36144 = n5675 | n18144 ;
  assign n36145 = n36144 ^ n18061 ^ 1'b0 ;
  assign n36149 = ~n13167 & n21882 ;
  assign n36150 = n18240 & n36149 ;
  assign n36146 = n4908 | n30056 ;
  assign n36147 = n36146 ^ n3197 ^ 1'b0 ;
  assign n36148 = ~n5731 & n36147 ;
  assign n36151 = n36150 ^ n36148 ^ 1'b0 ;
  assign n36152 = ~n15119 & n23557 ;
  assign n36153 = n21103 ^ n4001 ^ 1'b0 ;
  assign n36154 = n9377 | n36153 ;
  assign n36155 = ~n2900 & n21683 ;
  assign n36156 = n36155 ^ n10299 ^ 1'b0 ;
  assign n36157 = n36156 ^ n9649 ^ 1'b0 ;
  assign n36158 = n9792 & n36157 ;
  assign n36159 = n17172 ^ n10649 ^ n1820 ;
  assign n36160 = n7135 ^ n3416 ^ 1'b0 ;
  assign n36161 = ~n12095 & n36160 ;
  assign n36162 = n36161 ^ n8015 ^ 1'b0 ;
  assign n36163 = n36162 ^ n9496 ^ 1'b0 ;
  assign n36164 = n20921 | n35577 ;
  assign n36165 = n36164 ^ n24311 ^ 1'b0 ;
  assign n36166 = n8595 ^ n874 ^ 1'b0 ;
  assign n36167 = n3457 | n36166 ;
  assign n36168 = n36167 ^ n25315 ^ 1'b0 ;
  assign n36169 = n27069 ^ n2942 ^ 1'b0 ;
  assign n36170 = n3323 & n36169 ;
  assign n36171 = n23140 ^ n22035 ^ 1'b0 ;
  assign n36172 = n33655 | n36171 ;
  assign n36173 = ~n2845 & n36172 ;
  assign n36174 = n4830 | n5560 ;
  assign n36175 = n36174 ^ n30864 ^ n1456 ;
  assign n36176 = n2508 & n26719 ;
  assign n36177 = n36176 ^ n12704 ^ 1'b0 ;
  assign n36178 = ~n1048 & n36177 ;
  assign n36180 = n6261 & n18764 ;
  assign n36181 = n36180 ^ n26995 ^ 1'b0 ;
  assign n36179 = n35538 ^ n22425 ^ 1'b0 ;
  assign n36182 = n36181 ^ n36179 ^ n20095 ;
  assign n36183 = n9099 & ~n36182 ;
  assign n36184 = x172 | n5206 ;
  assign n36185 = ~n4341 & n36184 ;
  assign n36186 = n36185 ^ n31236 ^ 1'b0 ;
  assign n36187 = n564 | n36186 ;
  assign n36188 = n19654 ^ n13899 ^ 1'b0 ;
  assign n36190 = n16370 ^ n5685 ^ n4797 ;
  assign n36191 = ~n7716 & n36190 ;
  assign n36189 = n5504 & n6540 ;
  assign n36192 = n36191 ^ n36189 ^ n20208 ;
  assign n36193 = x192 | n28606 ;
  assign n36194 = n4723 & ~n36193 ;
  assign n36195 = n36194 ^ n34197 ^ 1'b0 ;
  assign n36196 = n14017 & ~n21802 ;
  assign n36197 = ( n3901 & ~n7162 ) | ( n3901 & n36196 ) | ( ~n7162 & n36196 ) ;
  assign n36198 = n36197 ^ n26873 ^ 1'b0 ;
  assign n36199 = n16368 & n36198 ;
  assign n36200 = n36199 ^ n1458 ^ 1'b0 ;
  assign n36201 = n4117 | n9066 ;
  assign n36202 = n3619 | n36201 ;
  assign n36203 = n27438 ^ n9758 ^ 1'b0 ;
  assign n36204 = n36202 & ~n36203 ;
  assign n36205 = n31520 ^ n28292 ^ 1'b0 ;
  assign n36206 = n20648 & n36205 ;
  assign n36207 = n1989 & ~n14886 ;
  assign n36208 = n23027 ^ n2443 ^ 1'b0 ;
  assign n36209 = n5921 | n36208 ;
  assign n36210 = n6886 ^ n537 ^ 1'b0 ;
  assign n36211 = n30836 & ~n36210 ;
  assign n36212 = n11265 | n16926 ;
  assign n36213 = n12952 & ~n36212 ;
  assign n36214 = n36213 ^ n11333 ^ 1'b0 ;
  assign n36215 = ( ~n6703 & n9061 ) | ( ~n6703 & n36214 ) | ( n9061 & n36214 ) ;
  assign n36216 = n10746 ^ n5187 ^ 1'b0 ;
  assign n36217 = n9026 & ~n36216 ;
  assign n36218 = ~n6010 & n36217 ;
  assign n36219 = n18296 & n19166 ;
  assign n36221 = n12426 ^ n1885 ^ 1'b0 ;
  assign n36220 = ~n14120 & n26647 ;
  assign n36222 = n36221 ^ n36220 ^ 1'b0 ;
  assign n36223 = ~n2735 & n7773 ;
  assign n36224 = n6896 & n9681 ;
  assign n36225 = n36224 ^ n5676 ^ 1'b0 ;
  assign n36226 = n23557 & ~n36225 ;
  assign n36227 = n20638 ^ n14078 ^ 1'b0 ;
  assign n36228 = x143 & n30171 ;
  assign n36229 = x249 | n13676 ;
  assign n36230 = n35593 & ~n36229 ;
  assign n36231 = n5387 & n12354 ;
  assign n36232 = n25583 ^ n5734 ^ 1'b0 ;
  assign n36233 = n15814 ^ n4585 ^ 1'b0 ;
  assign n36234 = ~n7738 & n36233 ;
  assign n36235 = ~n4065 & n12647 ;
  assign n36237 = n1805 | n12030 ;
  assign n36238 = n36237 ^ n7805 ^ 1'b0 ;
  assign n36236 = n4568 | n20332 ;
  assign n36239 = n36238 ^ n36236 ^ 1'b0 ;
  assign n36240 = n2932 & ~n36239 ;
  assign n36241 = n10738 ^ n10499 ^ 1'b0 ;
  assign n36242 = n2790 | n36241 ;
  assign n36243 = n983 | n5038 ;
  assign n36244 = n36242 & ~n36243 ;
  assign n36245 = n18356 & ~n36244 ;
  assign n36246 = n36245 ^ n22711 ^ 1'b0 ;
  assign n36247 = n7316 | n29256 ;
  assign n36248 = n18954 ^ n5531 ^ 1'b0 ;
  assign n36249 = n26896 & ~n36248 ;
  assign n36250 = n13083 ^ n1980 ^ 1'b0 ;
  assign n36251 = n3218 & ~n36250 ;
  assign n36252 = n36251 ^ n11187 ^ 1'b0 ;
  assign n36253 = n4576 & n12549 ;
  assign n36254 = n36253 ^ n6545 ^ 1'b0 ;
  assign n36255 = n26562 | n36254 ;
  assign n36256 = n36255 ^ n1575 ^ 1'b0 ;
  assign n36257 = ~n14425 & n33276 ;
  assign n36258 = n9289 & ~n34718 ;
  assign n36259 = n17376 & n36258 ;
  assign n36260 = n3378 & ~n21513 ;
  assign n36261 = n25512 & n36260 ;
  assign n36262 = n4038 ^ n589 ^ 1'b0 ;
  assign n36263 = n8276 | n36262 ;
  assign n36264 = n5728 | n22683 ;
  assign n36265 = n5130 & ~n8728 ;
  assign n36266 = n20735 & n36265 ;
  assign n36267 = n12287 ^ n2319 ^ 1'b0 ;
  assign n36268 = n10475 & ~n36267 ;
  assign n36269 = n36268 ^ n22275 ^ 1'b0 ;
  assign n36270 = n22702 ^ n871 ^ 1'b0 ;
  assign n36271 = n9676 & ~n22860 ;
  assign n36272 = n36271 ^ n29182 ^ 1'b0 ;
  assign n36273 = n2881 | n3513 ;
  assign n36274 = n3371 | n36273 ;
  assign n36275 = n36274 ^ n25747 ^ n7035 ;
  assign n36276 = n8000 & ~n36275 ;
  assign n36277 = n36276 ^ n31081 ^ 1'b0 ;
  assign n36278 = n7902 & ~n8983 ;
  assign n36279 = n36278 ^ n14576 ^ 1'b0 ;
  assign n36280 = n20177 | n29539 ;
  assign n36281 = n36279 | n36280 ;
  assign n36282 = n22941 ^ n12022 ^ 1'b0 ;
  assign n36283 = n10158 & ~n36282 ;
  assign n36284 = n9669 & n19708 ;
  assign n36285 = n4144 & n32813 ;
  assign n36286 = ( n29566 & n36284 ) | ( n29566 & ~n36285 ) | ( n36284 & ~n36285 ) ;
  assign n36287 = n18315 & ~n21856 ;
  assign n36288 = ~x165 & n36287 ;
  assign n36289 = n15338 ^ n8980 ^ n1828 ;
  assign n36290 = ~n36288 & n36289 ;
  assign n36291 = n12699 | n36290 ;
  assign n36292 = n3199 & n16419 ;
  assign n36293 = n12714 ^ n11731 ^ 1'b0 ;
  assign n36294 = n36292 & ~n36293 ;
  assign n36295 = n5563 ^ n3064 ^ 1'b0 ;
  assign n36296 = n36295 ^ n34501 ^ 1'b0 ;
  assign n36297 = n17417 & n36296 ;
  assign n36298 = ~n3290 & n36297 ;
  assign n36299 = n611 | n2701 ;
  assign n36300 = n4827 | n36299 ;
  assign n36301 = n36300 ^ n22135 ^ 1'b0 ;
  assign n36302 = ~n20094 & n36301 ;
  assign n36303 = ~n21315 & n36302 ;
  assign n36304 = n23945 ^ n15643 ^ 1'b0 ;
  assign n36305 = n28316 ^ n977 ^ 1'b0 ;
  assign n36306 = ~n36304 & n36305 ;
  assign n36307 = n18055 ^ n14612 ^ 1'b0 ;
  assign n36311 = ~n1879 & n9200 ;
  assign n36308 = ~n13419 & n14887 ;
  assign n36309 = ~n20709 & n36308 ;
  assign n36310 = n11186 | n36309 ;
  assign n36312 = n36311 ^ n36310 ^ 1'b0 ;
  assign n36313 = n7467 & ~n20030 ;
  assign n36314 = n9496 & ~n22351 ;
  assign n36315 = n36314 ^ n4753 ^ 1'b0 ;
  assign n36316 = n5507 & n36315 ;
  assign n36317 = ~n9202 & n36316 ;
  assign n36318 = n9864 & n12083 ;
  assign n36319 = n8236 & n12642 ;
  assign n36320 = n10356 & n36319 ;
  assign n36321 = n7184 & ~n18499 ;
  assign n36322 = ~n36320 & n36321 ;
  assign n36323 = n18019 ^ n4723 ^ 1'b0 ;
  assign n36324 = n13582 & n18466 ;
  assign n36325 = n16038 | n27469 ;
  assign n36326 = n36324 & ~n36325 ;
  assign n36327 = n31662 ^ n30531 ^ 1'b0 ;
  assign n36328 = n26297 | n36327 ;
  assign n36329 = ( ~n2491 & n36326 ) | ( ~n2491 & n36328 ) | ( n36326 & n36328 ) ;
  assign n36330 = n8607 ^ n8096 ^ 1'b0 ;
  assign n36331 = n36330 ^ n9562 ^ 1'b0 ;
  assign n36332 = n36331 ^ n4562 ^ 1'b0 ;
  assign n36333 = ~n2103 & n7877 ;
  assign n36334 = n36332 & n36333 ;
  assign n36335 = n9360 & ~n26153 ;
  assign n36336 = n27230 ^ n26822 ^ 1'b0 ;
  assign n36337 = n36335 & ~n36336 ;
  assign n36338 = n2301 | n8545 ;
  assign n36339 = n9340 & ~n36338 ;
  assign n36340 = n6549 | n8941 ;
  assign n36341 = n13452 | n36340 ;
  assign n36343 = n29745 ^ n25348 ^ 1'b0 ;
  assign n36342 = n5393 & ~n29756 ;
  assign n36344 = n36343 ^ n36342 ^ 1'b0 ;
  assign n36345 = n13193 & n21515 ;
  assign n36346 = n3197 & n13938 ;
  assign n36347 = n36346 ^ n6485 ^ 1'b0 ;
  assign n36348 = n7066 & ~n10682 ;
  assign n36349 = n36347 & n36348 ;
  assign n36350 = n4539 | n36349 ;
  assign n36351 = x94 | n36350 ;
  assign n36352 = ~n1364 & n36351 ;
  assign n36353 = n36352 ^ n8347 ^ 1'b0 ;
  assign n36354 = ~n471 & n8064 ;
  assign n36355 = ~n17858 & n36354 ;
  assign n36356 = ( n15255 & n31686 ) | ( n15255 & n36355 ) | ( n31686 & n36355 ) ;
  assign n36357 = n3903 ^ n448 ^ 1'b0 ;
  assign n36358 = n36357 ^ n33384 ^ 1'b0 ;
  assign n36359 = n12266 & ~n12466 ;
  assign n36360 = n33815 & n36359 ;
  assign n36361 = n5659 ^ n4712 ^ 1'b0 ;
  assign n36362 = n5400 & ~n12136 ;
  assign n36363 = n19624 & ~n22758 ;
  assign n36364 = ~n2493 & n36363 ;
  assign n36365 = n36364 ^ n25012 ^ n1343 ;
  assign n36366 = n921 & ~n5103 ;
  assign n36367 = n1294 & ~n7808 ;
  assign n36368 = n34927 | n36367 ;
  assign n36369 = n36368 ^ n18707 ^ 1'b0 ;
  assign n36370 = ~n9788 & n36369 ;
  assign n36371 = ~n9252 & n26260 ;
  assign n36372 = n34483 ^ n19971 ^ 1'b0 ;
  assign n36373 = n36371 | n36372 ;
  assign n36374 = n16845 ^ n1011 ^ n514 ;
  assign n36375 = ~n2045 & n28842 ;
  assign n36376 = ~n34228 & n36375 ;
  assign n36377 = n9317 & n22276 ;
  assign n36378 = n19538 ^ n3838 ^ 1'b0 ;
  assign n36379 = n36377 & n36378 ;
  assign n36380 = n12330 ^ n8025 ^ 1'b0 ;
  assign n36381 = n19948 ^ n1309 ^ 1'b0 ;
  assign n36382 = x88 & ~n36381 ;
  assign n36383 = n3478 ^ n2542 ^ 1'b0 ;
  assign n36384 = n8216 & ~n15343 ;
  assign n36385 = n28296 ^ x53 ^ 1'b0 ;
  assign n36386 = ~n36178 & n36385 ;
  assign n36387 = n5659 ^ n3604 ^ 1'b0 ;
  assign n36388 = n6518 | n36387 ;
  assign n36389 = n4514 | n36388 ;
  assign n36390 = ~n15931 & n36389 ;
  assign n36391 = n32562 ^ n264 ^ 1'b0 ;
  assign n36392 = n36390 & n36391 ;
  assign n36393 = n19932 ^ n14444 ^ 1'b0 ;
  assign n36394 = n5442 ^ n3368 ^ 1'b0 ;
  assign n36395 = n36394 ^ n10407 ^ n9072 ;
  assign n36396 = n10071 ^ n1374 ^ 1'b0 ;
  assign n36397 = n18906 ^ n12260 ^ 1'b0 ;
  assign n36398 = ~n17642 & n36397 ;
  assign n36399 = ~n12167 & n16737 ;
  assign n36400 = n36399 ^ n13306 ^ 1'b0 ;
  assign n36401 = ~n10639 & n15704 ;
  assign n36402 = n36401 ^ n20659 ^ 1'b0 ;
  assign n36403 = n20833 & n36402 ;
  assign n36404 = ~n638 & n3195 ;
  assign n36405 = ~n12409 & n36404 ;
  assign n36406 = n1796 & n36405 ;
  assign n36407 = n10321 ^ n8935 ^ 1'b0 ;
  assign n36408 = ~n33223 & n36407 ;
  assign n36409 = n15314 ^ n394 ^ 1'b0 ;
  assign n36410 = n36408 & n36409 ;
  assign n36411 = n36410 ^ n16298 ^ 1'b0 ;
  assign n36412 = n13607 ^ n10733 ^ n4997 ;
  assign n36413 = ~n14947 & n36412 ;
  assign n36414 = n36413 ^ n29001 ^ n17274 ;
  assign n36415 = n2050 & n12845 ;
  assign n36416 = n5946 & n36415 ;
  assign n36417 = n13170 & ~n22452 ;
  assign n36418 = n20388 & n36417 ;
  assign n36419 = n8937 ^ n629 ^ 1'b0 ;
  assign n36420 = n1217 & n36419 ;
  assign n36421 = n5649 & n36420 ;
  assign n36423 = n5949 & n16407 ;
  assign n36424 = n36423 ^ n4551 ^ 1'b0 ;
  assign n36422 = n28084 ^ n26925 ^ n8676 ;
  assign n36425 = n36424 ^ n36422 ^ 1'b0 ;
  assign n36426 = n6707 & n36425 ;
  assign n36427 = n342 & n36426 ;
  assign n36428 = n13781 | n33102 ;
  assign n36429 = n24246 ^ n6582 ^ 1'b0 ;
  assign n36430 = n36429 ^ n7606 ^ n2112 ;
  assign n36431 = n16008 | n20153 ;
  assign n36432 = n25297 | n36431 ;
  assign n36433 = n2213 & ~n20608 ;
  assign n36434 = n22951 | n36433 ;
  assign n36435 = n16379 & ~n36434 ;
  assign n36436 = ~n13152 & n14586 ;
  assign n36437 = n4305 & n36436 ;
  assign n36438 = x245 & ~n4767 ;
  assign n36439 = n1342 | n36438 ;
  assign n36440 = ~n310 & n3710 ;
  assign n36441 = ( n4009 & n27041 ) | ( n4009 & n36440 ) | ( n27041 & n36440 ) ;
  assign n36442 = ( ~n372 & n11776 ) | ( ~n372 & n36441 ) | ( n11776 & n36441 ) ;
  assign n36443 = ( n19312 & n28761 ) | ( n19312 & n36442 ) | ( n28761 & n36442 ) ;
  assign n36444 = n2549 | n12696 ;
  assign n36445 = n36444 ^ n12078 ^ 1'b0 ;
  assign n36446 = ~n1159 & n36445 ;
  assign n36447 = ~n9919 & n36446 ;
  assign n36448 = ~n9990 & n16236 ;
  assign n36449 = ~n21382 & n36448 ;
  assign n36450 = n11660 ^ n938 ^ 1'b0 ;
  assign n36451 = ( n7935 & n25338 ) | ( n7935 & ~n36450 ) | ( n25338 & ~n36450 ) ;
  assign n36452 = n35758 | n36451 ;
  assign n36453 = n5763 & n36452 ;
  assign n36454 = x221 & n31734 ;
  assign n36455 = n13154 & n36454 ;
  assign n36456 = n8390 & ~n14272 ;
  assign n36457 = ~n20742 & n36456 ;
  assign n36458 = n36457 ^ n35180 ^ 1'b0 ;
  assign n36459 = n11701 ^ n8607 ^ 1'b0 ;
  assign n36460 = n1577 ^ n935 ^ 1'b0 ;
  assign n36461 = n10648 | n36460 ;
  assign n36462 = n2466 & n18142 ;
  assign n36463 = ( x86 & n30360 ) | ( x86 & n36462 ) | ( n30360 & n36462 ) ;
  assign n36464 = n23257 ^ n3802 ^ 1'b0 ;
  assign n36465 = n36463 & n36464 ;
  assign n36466 = n24194 ^ n14801 ^ n1478 ;
  assign n36467 = ~n1376 & n36466 ;
  assign n36468 = n15275 & n18399 ;
  assign n36469 = ~n6753 & n36468 ;
  assign n36470 = ~n928 & n6288 ;
  assign n36471 = n36470 ^ n7868 ^ 1'b0 ;
  assign n36472 = ( n8030 & n20628 ) | ( n8030 & n36471 ) | ( n20628 & n36471 ) ;
  assign n36473 = n36472 ^ n20673 ^ 1'b0 ;
  assign n36474 = n36469 & n36473 ;
  assign n36475 = n31790 ^ n10256 ^ 1'b0 ;
  assign n36476 = n1424 & ~n9660 ;
  assign n36477 = ~n9365 & n17566 ;
  assign n36478 = x215 & ~n17113 ;
  assign n36479 = ( ~n6529 & n8123 ) | ( ~n6529 & n14055 ) | ( n8123 & n14055 ) ;
  assign n36480 = n27730 ^ n22897 ^ 1'b0 ;
  assign n36481 = n7298 | n36480 ;
  assign n36482 = n4754 ^ n3152 ^ 1'b0 ;
  assign n36483 = ~n10781 & n36482 ;
  assign n36484 = n36483 ^ n33346 ^ n6678 ;
  assign n36485 = n1492 & n36484 ;
  assign n36486 = n32220 ^ n19961 ^ 1'b0 ;
  assign n36487 = ~n28073 & n36486 ;
  assign n36492 = n19700 ^ n9481 ^ 1'b0 ;
  assign n36488 = ( n423 & n1219 ) | ( n423 & ~n16353 ) | ( n1219 & ~n16353 ) ;
  assign n36489 = n11078 | n36488 ;
  assign n36490 = n36489 ^ n3663 ^ 1'b0 ;
  assign n36491 = n23715 | n36490 ;
  assign n36493 = n36492 ^ n36491 ^ n24965 ;
  assign n36494 = n10517 ^ n4997 ^ 1'b0 ;
  assign n36495 = ~n29025 & n36494 ;
  assign n36496 = ~n13207 & n36495 ;
  assign n36497 = n813 & n36496 ;
  assign n36498 = n15252 ^ n3265 ^ 1'b0 ;
  assign n36499 = n3769 & n9973 ;
  assign n36500 = ~n31154 & n36499 ;
  assign n36501 = ~n36498 & n36500 ;
  assign n36502 = n32553 ^ n22572 ^ 1'b0 ;
  assign n36503 = n26920 & ~n36502 ;
  assign n36504 = ~n7646 & n20840 ;
  assign n36505 = n9481 | n19602 ;
  assign n36506 = n36504 & ~n36505 ;
  assign n36507 = n31757 | n36506 ;
  assign n36508 = n27336 & ~n36507 ;
  assign n36509 = n36508 ^ n29318 ^ x186 ;
  assign n36510 = ~n10448 & n34937 ;
  assign n36511 = n36510 ^ n7648 ^ 1'b0 ;
  assign n36513 = ( n293 & n7807 ) | ( n293 & ~n8639 ) | ( n7807 & ~n8639 ) ;
  assign n36512 = n16977 & ~n19356 ;
  assign n36514 = n36513 ^ n36512 ^ 1'b0 ;
  assign n36515 = n799 | n6861 ;
  assign n36516 = n36515 ^ n2389 ^ 1'b0 ;
  assign n36517 = n10776 | n36516 ;
  assign n36518 = n36517 ^ n28573 ^ 1'b0 ;
  assign n36519 = n36514 & ~n36518 ;
  assign n36520 = n9515 & n26539 ;
  assign n36521 = x228 & n34937 ;
  assign n36522 = n26185 ^ n16599 ^ 1'b0 ;
  assign n36523 = n15483 & ~n19685 ;
  assign n36524 = n6352 & n36523 ;
  assign n36525 = n18551 | n36524 ;
  assign n36526 = n11044 ^ n7209 ^ n2953 ;
  assign n36527 = n4047 & n36526 ;
  assign n36528 = ( n5189 & ~n9934 ) | ( n5189 & n12350 ) | ( ~n9934 & n12350 ) ;
  assign n36529 = n36528 ^ n9627 ^ 1'b0 ;
  assign n36530 = n3240 & n4708 ;
  assign n36531 = ~n36529 & n36530 ;
  assign n36532 = n15423 ^ n3704 ^ 1'b0 ;
  assign n36533 = n3506 & ~n36532 ;
  assign n36534 = n1937 & n34439 ;
  assign n36535 = n35112 ^ n1010 ^ 1'b0 ;
  assign n36536 = n17372 ^ n13048 ^ 1'b0 ;
  assign n36537 = n10610 & n36536 ;
  assign n36538 = n36537 ^ n29238 ^ 1'b0 ;
  assign n36539 = n3721 | n36156 ;
  assign n36540 = n36539 ^ n18298 ^ 1'b0 ;
  assign n36541 = n28121 | n33194 ;
  assign n36542 = n10317 | n36541 ;
  assign n36543 = n34168 & ~n36542 ;
  assign n36544 = n5804 ^ n5446 ^ 1'b0 ;
  assign n36545 = n4009 & ~n6514 ;
  assign n36546 = n36545 ^ n17406 ^ n5650 ;
  assign n36547 = n5725 | n17678 ;
  assign n36548 = n2158 & ~n36547 ;
  assign n36549 = ( ~n389 & n11204 ) | ( ~n389 & n36548 ) | ( n11204 & n36548 ) ;
  assign n36550 = n18734 | n35011 ;
  assign n36551 = n5238 ^ n4807 ^ 1'b0 ;
  assign n36552 = ~n4876 & n36551 ;
  assign n36553 = n15391 & n36552 ;
  assign n36554 = ~n5003 & n36553 ;
  assign n36555 = n25166 ^ n5373 ^ 1'b0 ;
  assign n36556 = ~n21741 & n30657 ;
  assign n36557 = n28395 ^ n4773 ^ x156 ;
  assign n36558 = n22069 ^ n11651 ^ 1'b0 ;
  assign n36559 = n10271 | n36558 ;
  assign n36560 = n27363 & n36559 ;
  assign n36561 = n23724 | n30947 ;
  assign n36562 = n36561 ^ n21942 ^ 1'b0 ;
  assign n36563 = n33106 | n36562 ;
  assign n36564 = n20629 ^ n11102 ^ n2771 ;
  assign n36565 = n20995 | n36564 ;
  assign n36566 = n18948 & ~n24375 ;
  assign n36567 = n17588 | n35133 ;
  assign n36568 = n7386 | n30252 ;
  assign n36569 = x158 & n5192 ;
  assign n36570 = n36569 ^ n8693 ^ 1'b0 ;
  assign n36571 = n6726 | n36570 ;
  assign n36572 = n13942 & n33133 ;
  assign n36573 = n36572 ^ x51 ^ 1'b0 ;
  assign n36574 = n31467 ^ n25975 ^ 1'b0 ;
  assign n36575 = n5205 & n11863 ;
  assign n36576 = n14167 ^ n6992 ^ 1'b0 ;
  assign n36577 = n382 & n2326 ;
  assign n36578 = n4685 | n21841 ;
  assign n36579 = n2678 | n36578 ;
  assign n36580 = n36579 ^ n23746 ^ 1'b0 ;
  assign n36581 = n36580 ^ n35528 ^ 1'b0 ;
  assign n36582 = n23440 ^ n11285 ^ 1'b0 ;
  assign n36583 = ~n14514 & n18194 ;
  assign n36584 = n13198 & n24157 ;
  assign n36585 = n36583 & n36584 ;
  assign n36586 = n18910 | n24290 ;
  assign n36587 = n1606 & ~n7536 ;
  assign n36588 = n2653 & n36587 ;
  assign n36589 = ( ~n16307 & n16786 ) | ( ~n16307 & n16799 ) | ( n16786 & n16799 ) ;
  assign n36590 = n36588 | n36589 ;
  assign n36594 = n24657 & ~n25402 ;
  assign n36591 = n24514 | n28917 ;
  assign n36592 = n8557 | n36591 ;
  assign n36593 = n12571 & n36592 ;
  assign n36595 = n36594 ^ n36593 ^ 1'b0 ;
  assign n36596 = n36128 ^ n7631 ^ 1'b0 ;
  assign n36597 = ~n22357 & n36596 ;
  assign n36598 = n5140 ^ n1730 ^ 1'b0 ;
  assign n36599 = n36597 & n36598 ;
  assign n36600 = ~n21213 & n26610 ;
  assign n36601 = n36600 ^ n25361 ^ 1'b0 ;
  assign n36602 = ~n13802 & n36601 ;
  assign n36603 = n36602 ^ n6524 ^ 1'b0 ;
  assign n36604 = n21734 & n35829 ;
  assign n36605 = n8734 & n11002 ;
  assign n36606 = n1232 & n18935 ;
  assign n36607 = n420 | n25517 ;
  assign n36608 = n18300 ^ n9520 ^ n1203 ;
  assign n36609 = n10106 | n31949 ;
  assign n36610 = n36609 ^ n22243 ^ 1'b0 ;
  assign n36611 = n3707 & n4773 ;
  assign n36612 = ~n23539 & n36611 ;
  assign n36613 = n10071 | n19741 ;
  assign n36614 = n3138 & ~n36613 ;
  assign n36615 = n12224 ^ n2487 ^ 1'b0 ;
  assign n36616 = n14256 & ~n36615 ;
  assign n36617 = ~n23980 & n36616 ;
  assign n36618 = n29309 ^ n28135 ^ 1'b0 ;
  assign n36619 = n12709 | n36618 ;
  assign n36620 = n36619 ^ n35609 ^ 1'b0 ;
  assign n36621 = n36620 ^ n33814 ^ 1'b0 ;
  assign n36622 = n9586 ^ n6748 ^ 1'b0 ;
  assign n36623 = n2897 | n36622 ;
  assign n36624 = n36623 ^ n32253 ^ 1'b0 ;
  assign n36625 = n30464 & ~n32381 ;
  assign n36626 = ~n31181 & n32124 ;
  assign n36627 = n36626 ^ n7732 ^ 1'b0 ;
  assign n36628 = ~n16768 & n20769 ;
  assign n36629 = n31724 ^ n8844 ^ n3668 ;
  assign n36630 = n34586 ^ n6550 ^ 1'b0 ;
  assign n36631 = n5403 | n15977 ;
  assign n36632 = n36631 ^ n15889 ^ 1'b0 ;
  assign n36633 = n8674 | n12123 ;
  assign n36634 = n26822 ^ n16135 ^ 1'b0 ;
  assign n36635 = n14008 & ~n27347 ;
  assign n36636 = n21436 ^ n10941 ^ n1441 ;
  assign n36637 = n9999 ^ n2242 ^ 1'b0 ;
  assign n36638 = n29447 & n36637 ;
  assign n36639 = ~n4111 & n36638 ;
  assign n36640 = n12006 & ~n15678 ;
  assign n36641 = n36639 & n36640 ;
  assign n36642 = n34465 ^ n30483 ^ 1'b0 ;
  assign n36643 = ~n10489 & n10606 ;
  assign n36644 = n36643 ^ n19592 ^ 1'b0 ;
  assign n36645 = ~n18970 & n36644 ;
  assign n36646 = n29740 ^ n4161 ^ 1'b0 ;
  assign n36647 = ~n36645 & n36646 ;
  assign n36648 = n7766 & n18948 ;
  assign n36649 = n36648 ^ n18291 ^ 1'b0 ;
  assign n36650 = n3751 | n9334 ;
  assign n36651 = n8278 | n36650 ;
  assign n36652 = n11657 | n36651 ;
  assign n36653 = n31081 ^ n3271 ^ 1'b0 ;
  assign n36654 = n708 & ~n21798 ;
  assign n36655 = n4364 ^ n619 ^ 1'b0 ;
  assign n36656 = n4728 & ~n36655 ;
  assign n36657 = n36656 ^ n18781 ^ 1'b0 ;
  assign n36659 = n11529 & n27648 ;
  assign n36658 = ~n24731 & n31129 ;
  assign n36660 = n36659 ^ n36658 ^ 1'b0 ;
  assign n36661 = n1813 & n32029 ;
  assign n36662 = n9866 | n20637 ;
  assign n36664 = n24745 & ~n24870 ;
  assign n36663 = n20243 & ~n26688 ;
  assign n36665 = n36664 ^ n36663 ^ 1'b0 ;
  assign n36666 = n36665 ^ n19491 ^ n9253 ;
  assign n36667 = n34369 ^ n1912 ^ 1'b0 ;
  assign n36668 = n453 & n36651 ;
  assign n36669 = ~n1694 & n7019 ;
  assign n36670 = n36669 ^ n28138 ^ 1'b0 ;
  assign n36671 = ~n20831 & n20989 ;
  assign n36672 = n3054 & ~n5234 ;
  assign n36673 = ( n2589 & n15733 ) | ( n2589 & ~n36672 ) | ( n15733 & ~n36672 ) ;
  assign n36674 = n23419 ^ n3490 ^ 1'b0 ;
  assign n36675 = n7349 & n36674 ;
  assign n36676 = n4629 & n6810 ;
  assign n36677 = n36676 ^ n13678 ^ n9994 ;
  assign n36678 = n18966 | n36677 ;
  assign n36679 = n35333 ^ n5291 ^ 1'b0 ;
  assign n36680 = n11071 | n36679 ;
  assign n36681 = n11191 & ~n23070 ;
  assign n36682 = ~n36680 & n36681 ;
  assign n36683 = ~n18943 & n36682 ;
  assign n36684 = n21187 ^ n1645 ^ 1'b0 ;
  assign n36685 = ~n19443 & n36684 ;
  assign n36686 = n18819 & ~n24228 ;
  assign n36687 = n8375 & n36686 ;
  assign n36688 = n7873 | n36687 ;
  assign n36689 = n36685 | n36688 ;
  assign n36691 = n9693 ^ n767 ^ x95 ;
  assign n36692 = n36691 ^ n21006 ^ 1'b0 ;
  assign n36693 = n6291 | n36692 ;
  assign n36690 = n8174 & n23324 ;
  assign n36694 = n36693 ^ n36690 ^ 1'b0 ;
  assign n36695 = ~n2799 & n8632 ;
  assign n36696 = n4851 & n5890 ;
  assign n36697 = n24881 & n36696 ;
  assign n36698 = n18233 | n34670 ;
  assign n36699 = x55 & n28674 ;
  assign n36700 = n36699 ^ n4434 ^ 1'b0 ;
  assign n36702 = ~n5067 & n9836 ;
  assign n36703 = ~n9781 & n36702 ;
  assign n36701 = n4062 & n16026 ;
  assign n36704 = n36703 ^ n36701 ^ 1'b0 ;
  assign n36705 = n30018 & n36704 ;
  assign n36706 = n7909 & ~n34808 ;
  assign n36707 = n36706 ^ x119 ^ 1'b0 ;
  assign n36708 = n16502 ^ n12340 ^ n8524 ;
  assign n36709 = n36708 ^ n15146 ^ n10041 ;
  assign n36710 = n7150 & ~n23284 ;
  assign n36711 = ( n31833 & n36709 ) | ( n31833 & ~n36710 ) | ( n36709 & ~n36710 ) ;
  assign n36712 = n9967 ^ n6147 ^ 1'b0 ;
  assign n36713 = n15238 ^ n14090 ^ n6177 ;
  assign n36717 = n30766 ^ n17919 ^ n17330 ;
  assign n36714 = n6607 & n20974 ;
  assign n36715 = n1778 & n36714 ;
  assign n36716 = ~n1059 & n36715 ;
  assign n36718 = n36717 ^ n36716 ^ 1'b0 ;
  assign n36719 = n13586 ^ n6284 ^ 1'b0 ;
  assign n36720 = n21237 & ~n29360 ;
  assign n36721 = n36720 ^ n5456 ^ 1'b0 ;
  assign n36722 = n1077 & ~n36721 ;
  assign n36723 = n36722 ^ n15779 ^ n15472 ;
  assign n36724 = n2123 & n12944 ;
  assign n36725 = n22786 ^ n18290 ^ 1'b0 ;
  assign n36726 = n4621 | n21092 ;
  assign n36727 = n20772 ^ x205 ^ 1'b0 ;
  assign n36728 = ~n14282 & n20372 ;
  assign n36729 = n19360 ^ n12733 ^ 1'b0 ;
  assign n36730 = n27291 ^ n5182 ^ 1'b0 ;
  assign n36731 = ~n36729 & n36730 ;
  assign n36732 = ~n14246 & n16475 ;
  assign n36733 = n4534 | n10664 ;
  assign n36734 = n13420 & n22316 ;
  assign n36735 = ~n13420 & n36734 ;
  assign n36736 = n8479 ^ n4794 ^ 1'b0 ;
  assign n36737 = n36735 | n36736 ;
  assign n36738 = n36737 ^ n28412 ^ 1'b0 ;
  assign n36739 = n36733 & n36738 ;
  assign n36740 = n15315 & n29285 ;
  assign n36741 = n36740 ^ n2569 ^ 1'b0 ;
  assign n36742 = n19640 & n36741 ;
  assign n36743 = ( n26546 & ~n35322 ) | ( n26546 & n36742 ) | ( ~n35322 & n36742 ) ;
  assign n36744 = ~n485 & n27535 ;
  assign n36745 = n36744 ^ n19986 ^ 1'b0 ;
  assign n36746 = n9009 ^ n2710 ^ 1'b0 ;
  assign n36747 = ~n1566 & n8366 ;
  assign n36748 = n36747 ^ n17118 ^ n11493 ;
  assign n36749 = n36746 & ~n36748 ;
  assign n36750 = n6711 | n25269 ;
  assign n36751 = n21908 & ~n36750 ;
  assign n36752 = ~n5596 & n22477 ;
  assign n36753 = n9260 & ~n9846 ;
  assign n36754 = ~n36752 & n36753 ;
  assign n36755 = ~n3571 & n25500 ;
  assign n36756 = ~n34842 & n36755 ;
  assign n36757 = n14569 & ~n19983 ;
  assign n36758 = n36757 ^ n3377 ^ 1'b0 ;
  assign n36759 = n3243 & ~n14007 ;
  assign n36760 = n36759 ^ n21026 ^ n6688 ;
  assign n36766 = n15230 ^ n4121 ^ 1'b0 ;
  assign n36767 = n5481 | n36766 ;
  assign n36768 = n4368 & n9224 ;
  assign n36769 = n36767 & n36768 ;
  assign n36761 = n11061 & n15078 ;
  assign n36762 = ~n28953 & n36761 ;
  assign n36763 = n10608 ^ n9832 ^ 1'b0 ;
  assign n36764 = n36762 | n36763 ;
  assign n36765 = n16183 & ~n36764 ;
  assign n36770 = n36769 ^ n36765 ^ 1'b0 ;
  assign n36771 = n7807 | n9959 ;
  assign n36772 = n36771 ^ n36453 ^ 1'b0 ;
  assign n36773 = n12980 & ~n14775 ;
  assign n36774 = n5796 & n36773 ;
  assign n36775 = ~n490 & n6064 ;
  assign n36776 = n36775 ^ n11749 ^ 1'b0 ;
  assign n36777 = ( n1664 & ~n5347 ) | ( n1664 & n36776 ) | ( ~n5347 & n36776 ) ;
  assign n36778 = n5359 & ~n6868 ;
  assign n36779 = n7763 ^ n5987 ^ 1'b0 ;
  assign n36780 = n36779 ^ n26067 ^ 1'b0 ;
  assign n36781 = n10800 | n36780 ;
  assign n36782 = ~n18150 & n20281 ;
  assign n36783 = n21289 | n23465 ;
  assign n36784 = n24726 ^ n11955 ^ n5984 ;
  assign n36785 = n12812 | n29212 ;
  assign n36786 = n36785 ^ n23911 ^ 1'b0 ;
  assign n36787 = ~n36784 & n36786 ;
  assign n36788 = n1734 | n20012 ;
  assign n36790 = n5998 | n9267 ;
  assign n36789 = ~n4512 & n6148 ;
  assign n36791 = n36790 ^ n36789 ^ 1'b0 ;
  assign n36792 = n4783 & n16594 ;
  assign n36793 = n20297 & n36792 ;
  assign n36794 = n5138 & n17896 ;
  assign n36795 = n36794 ^ n11116 ^ 1'b0 ;
  assign n36796 = n4424 | n22442 ;
  assign n36797 = n5111 & n8252 ;
  assign n36798 = n36797 ^ n4602 ^ 1'b0 ;
  assign n36799 = n3408 | n22253 ;
  assign n36800 = n36798 & ~n36799 ;
  assign n36801 = n1627 & n26539 ;
  assign n36802 = n36801 ^ n25915 ^ 1'b0 ;
  assign n36803 = n7648 & ~n36802 ;
  assign n36804 = ( n8442 & n36800 ) | ( n8442 & ~n36803 ) | ( n36800 & ~n36803 ) ;
  assign n36805 = ( ~n5115 & n8822 ) | ( ~n5115 & n14190 ) | ( n8822 & n14190 ) ;
  assign n36806 = n6099 | n7989 ;
  assign n36807 = ~n22198 & n36806 ;
  assign n36808 = n4299 & n36807 ;
  assign n36809 = n13354 & ~n33159 ;
  assign n36810 = n11365 & n13486 ;
  assign n36811 = n349 | n7185 ;
  assign n36812 = n7392 & ~n36811 ;
  assign n36813 = n20829 & n36812 ;
  assign n36814 = ( ~n4126 & n16947 ) | ( ~n4126 & n36813 ) | ( n16947 & n36813 ) ;
  assign n36815 = ( ~n16508 & n16751 ) | ( ~n16508 & n36814 ) | ( n16751 & n36814 ) ;
  assign n36816 = n12967 ^ n3502 ^ 1'b0 ;
  assign n36817 = n28036 & n36816 ;
  assign n36818 = n17007 ^ n11296 ^ 1'b0 ;
  assign n36819 = n36817 & ~n36818 ;
  assign n36820 = n36813 ^ n33828 ^ n21594 ;
  assign n36821 = n9693 & n36820 ;
  assign n36822 = n34550 ^ n5335 ^ 1'b0 ;
  assign n36823 = n3506 & ~n36822 ;
  assign n36824 = n17666 ^ n6080 ^ n5827 ;
  assign n36825 = ~n18486 & n36824 ;
  assign n36826 = x107 & ~n30489 ;
  assign n36827 = n36826 ^ n11148 ^ 1'b0 ;
  assign n36828 = n29686 ^ n19309 ^ n18733 ;
  assign n36829 = n36828 ^ n26639 ^ 1'b0 ;
  assign n36830 = n31994 ^ n14794 ^ n7216 ;
  assign n36831 = n666 & ~n26397 ;
  assign n36832 = n19430 & n36831 ;
  assign n36833 = n18410 | n32935 ;
  assign n36834 = n17688 ^ n1021 ^ 1'b0 ;
  assign n36836 = ~n3704 & n9695 ;
  assign n36835 = n2922 & ~n18188 ;
  assign n36837 = n36836 ^ n36835 ^ 1'b0 ;
  assign n36838 = n35302 ^ n1664 ^ 1'b0 ;
  assign n36839 = n24418 & n36838 ;
  assign n36840 = ~n23180 & n31378 ;
  assign n36841 = n20006 | n23574 ;
  assign n36842 = n33953 ^ n26520 ^ 1'b0 ;
  assign n36843 = n1324 | n3793 ;
  assign n36844 = n36843 ^ n11809 ^ n10026 ;
  assign n36845 = ~n11017 & n23688 ;
  assign n36846 = n14898 & n16191 ;
  assign n36847 = ~n5162 & n36846 ;
  assign n36848 = n11449 ^ n3100 ^ 1'b0 ;
  assign n36849 = ~n2988 & n36848 ;
  assign n36850 = n2140 & n16168 ;
  assign n36851 = ( n8442 & n18569 ) | ( n8442 & ~n24735 ) | ( n18569 & ~n24735 ) ;
  assign n36852 = ~n2075 & n36782 ;
  assign n36853 = ~n21057 & n36324 ;
  assign n36854 = n9076 & n36853 ;
  assign n36855 = ~n5792 & n36854 ;
  assign n36856 = n7590 & n31779 ;
  assign n36857 = ~x128 & n36856 ;
  assign n36861 = n8936 ^ n5490 ^ 1'b0 ;
  assign n36862 = ~n10236 & n36861 ;
  assign n36863 = n492 & n36862 ;
  assign n36864 = n19064 & n36863 ;
  assign n36865 = n36864 ^ n5292 ^ 1'b0 ;
  assign n36858 = x229 & n18841 ;
  assign n36859 = n20739 | n36858 ;
  assign n36860 = n36859 ^ n26824 ^ 1'b0 ;
  assign n36866 = n36865 ^ n36860 ^ n24311 ;
  assign n36867 = n23077 ^ n10846 ^ 1'b0 ;
  assign n36868 = n6629 & n29920 ;
  assign n36869 = n4341 | n19427 ;
  assign n36870 = n36869 ^ n32732 ^ 1'b0 ;
  assign n36873 = n13735 | n18628 ;
  assign n36871 = n10606 ^ n6053 ^ n5849 ;
  assign n36872 = n36871 ^ n7242 ^ 1'b0 ;
  assign n36874 = n36873 ^ n36872 ^ n4804 ;
  assign n36875 = n36874 ^ n1971 ^ 1'b0 ;
  assign n36876 = ( ~n6632 & n14663 ) | ( ~n6632 & n28690 ) | ( n14663 & n28690 ) ;
  assign n36877 = n29529 ^ n19722 ^ 1'b0 ;
  assign n36878 = n18129 & ~n31046 ;
  assign n36879 = ~n14015 & n27580 ;
  assign n36880 = ( n2576 & n9496 ) | ( n2576 & ~n10215 ) | ( n9496 & ~n10215 ) ;
  assign n36881 = ~n36879 & n36880 ;
  assign n36882 = n36881 ^ n5574 ^ 1'b0 ;
  assign n36883 = n21213 ^ n15863 ^ 1'b0 ;
  assign n36884 = x177 & ~n36883 ;
  assign n36885 = n30418 | n36697 ;
  assign n36886 = n4638 & ~n24981 ;
  assign n36887 = ( n2047 & n28362 ) | ( n2047 & ~n36886 ) | ( n28362 & ~n36886 ) ;
  assign n36888 = n32954 ^ n30046 ^ n20456 ;
  assign n36889 = n28046 & n30048 ;
  assign n36890 = n36651 ^ n3088 ^ 1'b0 ;
  assign n36891 = ~n1065 & n36890 ;
  assign n36892 = n36891 ^ n6155 ^ 1'b0 ;
  assign n36893 = n28793 ^ n3668 ^ 1'b0 ;
  assign n36894 = n22995 ^ n12818 ^ 1'b0 ;
  assign n36895 = ~n4150 & n36894 ;
  assign n36896 = n36895 ^ n7493 ^ 1'b0 ;
  assign n36897 = ~n36893 & n36896 ;
  assign n36898 = n28833 & n31514 ;
  assign n36899 = n7648 & ~n9041 ;
  assign n36900 = n36899 ^ n23996 ^ n6950 ;
  assign n36901 = n11031 & n19873 ;
  assign n36902 = n13534 | n33222 ;
  assign n36903 = n36901 & ~n36902 ;
  assign n36904 = n34851 ^ n5025 ^ 1'b0 ;
  assign n36905 = n13942 ^ n9113 ^ 1'b0 ;
  assign n36906 = n17858 & n36905 ;
  assign n36907 = n36906 ^ n8151 ^ 1'b0 ;
  assign n36908 = n21503 ^ n4428 ^ 1'b0 ;
  assign n36909 = n36907 & n36908 ;
  assign n36910 = n20524 & n29827 ;
  assign n36911 = n36910 ^ n19195 ^ 1'b0 ;
  assign n36912 = n30186 ^ n17642 ^ n3290 ;
  assign n36913 = n8925 | n31634 ;
  assign n36914 = n36913 ^ n21515 ^ 1'b0 ;
  assign n36915 = n5156 | n19200 ;
  assign n36916 = n5156 & ~n36915 ;
  assign n36917 = ( n10074 & n20464 ) | ( n10074 & n36916 ) | ( n20464 & n36916 ) ;
  assign n36918 = n10483 ^ n2915 ^ 1'b0 ;
  assign n36919 = n13054 | n36918 ;
  assign n36920 = n1471 | n20896 ;
  assign n36921 = n36920 ^ n397 ^ 1'b0 ;
  assign n36924 = n12646 ^ n7784 ^ 1'b0 ;
  assign n36925 = ~n18404 & n36924 ;
  assign n36922 = ~n12714 & n20506 ;
  assign n36923 = n21310 | n36922 ;
  assign n36926 = n36925 ^ n36923 ^ 1'b0 ;
  assign n36927 = n23862 ^ n21873 ^ 1'b0 ;
  assign n36928 = n24960 ^ n9686 ^ 1'b0 ;
  assign n36929 = ( n3574 & n6062 ) | ( n3574 & n36592 ) | ( n6062 & n36592 ) ;
  assign n36932 = ~n7516 & n16095 ;
  assign n36930 = n23378 ^ n18260 ^ 1'b0 ;
  assign n36931 = ~n9830 & n36930 ;
  assign n36933 = n36932 ^ n36931 ^ 1'b0 ;
  assign n36934 = n1389 & ~n13862 ;
  assign n36935 = n36934 ^ n24258 ^ 1'b0 ;
  assign n36939 = ( n4009 & n10311 ) | ( n4009 & n11816 ) | ( n10311 & n11816 ) ;
  assign n36940 = n15040 & ~n36939 ;
  assign n36941 = ~n7407 & n36940 ;
  assign n36942 = n14981 | n26049 ;
  assign n36943 = n36941 & ~n36942 ;
  assign n36936 = n20904 ^ n14062 ^ 1'b0 ;
  assign n36937 = n4991 & n36936 ;
  assign n36938 = n28109 & n36937 ;
  assign n36944 = n36943 ^ n36938 ^ 1'b0 ;
  assign n36945 = n18308 ^ n6305 ^ 1'b0 ;
  assign n36946 = n14929 ^ n6525 ^ 1'b0 ;
  assign n36947 = n4113 | n24214 ;
  assign n36948 = n36947 ^ n24672 ^ 1'b0 ;
  assign n36949 = ( n21625 & n36946 ) | ( n21625 & n36948 ) | ( n36946 & n36948 ) ;
  assign n36950 = n24218 ^ n10176 ^ 1'b0 ;
  assign n36951 = n2763 | n14651 ;
  assign n36952 = n36951 ^ n464 ^ 1'b0 ;
  assign n36953 = n7703 & n24317 ;
  assign n36954 = n1129 & n4898 ;
  assign n36955 = n36954 ^ n14193 ^ 1'b0 ;
  assign n36956 = n7875 | n25618 ;
  assign n36957 = n21973 ^ n3160 ^ 1'b0 ;
  assign n36958 = x158 & n36957 ;
  assign n36959 = n36958 ^ n28761 ^ 1'b0 ;
  assign n36960 = n3832 & n36959 ;
  assign n36961 = ~n25231 & n36960 ;
  assign n36962 = n36961 ^ n25598 ^ 1'b0 ;
  assign n36963 = n5188 & n36962 ;
  assign n36964 = n27031 ^ n5371 ^ 1'b0 ;
  assign n36965 = n36384 ^ n12882 ^ 1'b0 ;
  assign n36966 = n22375 & n36965 ;
  assign n36967 = n6941 & n32626 ;
  assign n36968 = n7308 ^ n6107 ^ 1'b0 ;
  assign n36969 = n7957 | n13045 ;
  assign n36970 = n36969 ^ n1820 ^ 1'b0 ;
  assign n36971 = ( n24194 & ~n36968 ) | ( n24194 & n36970 ) | ( ~n36968 & n36970 ) ;
  assign n36972 = ( n2922 & ~n15059 ) | ( n2922 & n31479 ) | ( ~n15059 & n31479 ) ;
  assign n36973 = n25731 ^ n6985 ^ 1'b0 ;
  assign n36974 = n29332 ^ n15551 ^ 1'b0 ;
  assign n36975 = n36973 | n36974 ;
  assign n36976 = n24906 ^ n8414 ^ 1'b0 ;
  assign n36977 = n24418 & ~n36976 ;
  assign n36978 = n13018 & n16903 ;
  assign n36979 = ~n6896 & n36978 ;
  assign n36980 = n19575 & ~n36979 ;
  assign n36981 = n10807 & n36980 ;
  assign n36982 = n12439 & ~n17229 ;
  assign n36983 = n36982 ^ n28975 ^ n8117 ;
  assign n36984 = n916 & n4598 ;
  assign n36985 = ~n4669 & n36984 ;
  assign n36986 = n10443 & ~n36985 ;
  assign n36987 = n36986 ^ n363 ^ 1'b0 ;
  assign n36988 = n3205 | n28694 ;
  assign n36989 = ~n15340 & n18900 ;
  assign n36990 = n8583 & ~n15941 ;
  assign n36991 = n36990 ^ n7096 ^ 1'b0 ;
  assign n36992 = ~n10443 & n36991 ;
  assign n36993 = n2528 | n9199 ;
  assign n36994 = n17178 ^ n15038 ^ 1'b0 ;
  assign n36995 = n29637 ^ n9505 ^ 1'b0 ;
  assign n36996 = n4338 & ~n17337 ;
  assign n36997 = n28655 & ~n36996 ;
  assign n36998 = n36997 ^ n5402 ^ 1'b0 ;
  assign n36999 = n21289 & ~n30863 ;
  assign n37000 = n36998 & n36999 ;
  assign n37001 = n22964 ^ n592 ^ 1'b0 ;
  assign n37002 = n27455 & n37001 ;
  assign n37003 = ~n30744 & n32776 ;
  assign n37004 = n37003 ^ n29605 ^ 1'b0 ;
  assign n37005 = n29490 ^ n10690 ^ 1'b0 ;
  assign n37006 = n29649 & n37005 ;
  assign n37007 = n37006 ^ n14843 ^ 1'b0 ;
  assign n37008 = n31125 ^ n18275 ^ n3795 ;
  assign n37009 = ~n4023 & n37008 ;
  assign n37010 = n37009 ^ n8658 ^ 1'b0 ;
  assign n37011 = n15926 | n22500 ;
  assign n37012 = n19439 ^ x168 ^ 1'b0 ;
  assign n37014 = n8085 ^ n5146 ^ 1'b0 ;
  assign n37013 = ~n2622 & n31044 ;
  assign n37015 = n37014 ^ n37013 ^ 1'b0 ;
  assign n37016 = ~n6057 & n18209 ;
  assign n37017 = n22490 & ~n33237 ;
  assign n37018 = n37017 ^ x181 ^ 1'b0 ;
  assign n37019 = n789 & ~n28512 ;
  assign n37020 = n37019 ^ n13773 ^ 1'b0 ;
  assign n37021 = ~n7737 & n10243 ;
  assign n37022 = n6817 & ~n37021 ;
  assign n37025 = n17131 ^ n17089 ^ n5333 ;
  assign n37026 = ~n23540 & n37025 ;
  assign n37023 = n12235 ^ n1048 ^ 1'b0 ;
  assign n37024 = n1378 | n37023 ;
  assign n37027 = n37026 ^ n37024 ^ 1'b0 ;
  assign n37028 = n14030 & ~n28784 ;
  assign n37029 = ~n16562 & n37028 ;
  assign n37030 = n4386 | n37029 ;
  assign n37031 = n33525 ^ n14981 ^ 1'b0 ;
  assign n37032 = n21563 ^ n19331 ^ 1'b0 ;
  assign n37033 = n30455 & n37032 ;
  assign n37034 = ~n6991 & n7944 ;
  assign n37035 = ~n28794 & n37034 ;
  assign n37036 = ~n2255 & n7124 ;
  assign n37037 = n274 & ~n12962 ;
  assign n37038 = n13961 & n37037 ;
  assign n37039 = ~n7128 & n37038 ;
  assign n37040 = n16198 & ~n37039 ;
  assign n37041 = ( ~n32530 & n33119 ) | ( ~n32530 & n37040 ) | ( n33119 & n37040 ) ;
  assign n37042 = n867 & ~n6928 ;
  assign n37043 = n37042 ^ n2887 ^ 1'b0 ;
  assign n37044 = n20915 ^ n8766 ^ 1'b0 ;
  assign n37045 = n21126 | n37044 ;
  assign n37046 = n8988 ^ n6920 ^ 1'b0 ;
  assign n37047 = ( n37043 & ~n37045 ) | ( n37043 & n37046 ) | ( ~n37045 & n37046 ) ;
  assign n37048 = n20971 ^ n3010 ^ 1'b0 ;
  assign n37049 = n13710 | n37048 ;
  assign n37050 = n4380 ^ n3496 ^ 1'b0 ;
  assign n37051 = n5047 | n37050 ;
  assign n37052 = n37051 ^ n30790 ^ 1'b0 ;
  assign n37056 = n26770 ^ n15845 ^ 1'b0 ;
  assign n37057 = n16421 | n37056 ;
  assign n37054 = n2044 & n10609 ;
  assign n37055 = ~n21755 & n37054 ;
  assign n37058 = n37057 ^ n37055 ^ 1'b0 ;
  assign n37053 = n6381 & ~n11247 ;
  assign n37059 = n37058 ^ n37053 ^ 1'b0 ;
  assign n37060 = n13256 & n31320 ;
  assign n37061 = n15446 & ~n31933 ;
  assign n37062 = n16646 & n37061 ;
  assign n37063 = n1557 | n37062 ;
  assign n37064 = n15446 ^ n13047 ^ 1'b0 ;
  assign n37065 = ~n4795 & n28459 ;
  assign n37066 = n19006 ^ n7263 ^ 1'b0 ;
  assign n37067 = n35127 ^ n14749 ^ 1'b0 ;
  assign n37068 = ~n2472 & n37067 ;
  assign n37069 = n4470 & n23182 ;
  assign n37070 = n30018 ^ n1926 ^ 1'b0 ;
  assign n37071 = n37069 & n37070 ;
  assign n37072 = ( n23672 & ~n37068 ) | ( n23672 & n37071 ) | ( ~n37068 & n37071 ) ;
  assign n37073 = ~n9659 & n20899 ;
  assign n37074 = n19107 | n19888 ;
  assign n37075 = n12231 & n25648 ;
  assign n37076 = n18287 & n37075 ;
  assign n37077 = n32123 ^ x56 ^ 1'b0 ;
  assign n37078 = ~n37076 & n37077 ;
  assign n37079 = n10765 ^ n10149 ^ 1'b0 ;
  assign n37080 = ~x207 & n1867 ;
  assign n37081 = n26247 ^ n10847 ^ 1'b0 ;
  assign n37082 = n37080 & ~n37081 ;
  assign n37083 = n35677 ^ n34486 ^ n27197 ;
  assign n37084 = n37082 & ~n37083 ;
  assign n37085 = n12225 & n29311 ;
  assign n37086 = n1441 | n6581 ;
  assign n37087 = n970 & n32162 ;
  assign n37088 = n37087 ^ n4752 ^ 1'b0 ;
  assign n37089 = n4797 | n20735 ;
  assign n37090 = n8510 | n37089 ;
  assign n37091 = n37088 & ~n37090 ;
  assign n37092 = n6851 & ~n20916 ;
  assign n37093 = n7247 & n37092 ;
  assign n37094 = ( x107 & n12861 ) | ( x107 & n37093 ) | ( n12861 & n37093 ) ;
  assign n37095 = ~n37091 & n37094 ;
  assign n37096 = n4689 & ~n21537 ;
  assign n37097 = n10907 | n20593 ;
  assign n37098 = n37096 & ~n37097 ;
  assign n37099 = n37098 ^ n28891 ^ n19702 ;
  assign n37100 = n27968 ^ n14752 ^ 1'b0 ;
  assign n37101 = n16059 & n37100 ;
  assign n37102 = n26515 ^ n23044 ^ 1'b0 ;
  assign n37103 = n37101 & n37102 ;
  assign n37104 = ~n765 & n11732 ;
  assign n37105 = n14492 & n37104 ;
  assign n37106 = n25637 ^ n5749 ^ 1'b0 ;
  assign n37107 = n29796 | n37106 ;
  assign n37108 = n37107 ^ n22979 ^ 1'b0 ;
  assign n37109 = n15025 & ~n16080 ;
  assign n37110 = n1775 | n23133 ;
  assign n37111 = n37110 ^ n34353 ^ n5708 ;
  assign n37112 = ~n23152 & n23473 ;
  assign n37113 = n37112 ^ n18296 ^ 1'b0 ;
  assign n37114 = n10208 & n37113 ;
  assign n37115 = n2409 ^ n772 ^ 1'b0 ;
  assign n37116 = n37115 ^ n9813 ^ 1'b0 ;
  assign n37117 = n3455 | n37116 ;
  assign n37118 = n17949 ^ n13306 ^ n2507 ;
  assign n37119 = n485 | n4234 ;
  assign n37120 = n6722 ^ n1999 ^ 1'b0 ;
  assign n37121 = ~n3634 & n10636 ;
  assign n37122 = n37121 ^ n20940 ^ 1'b0 ;
  assign n37123 = n37120 & n37122 ;
  assign n37124 = n4292 & n37123 ;
  assign n37125 = n26956 & ~n37124 ;
  assign n37126 = n37125 ^ n17903 ^ 1'b0 ;
  assign n37127 = n34275 ^ n20499 ^ 1'b0 ;
  assign n37128 = n14797 & n37127 ;
  assign n37129 = n24927 & ~n37128 ;
  assign n37130 = ~n20739 & n21535 ;
  assign n37131 = ~n20794 & n29716 ;
  assign n37132 = n15745 ^ n4551 ^ 1'b0 ;
  assign n37133 = n4222 ^ n740 ^ 1'b0 ;
  assign n37134 = n35780 ^ n23891 ^ n8395 ;
  assign n37135 = n2547 | n32567 ;
  assign n37136 = n17490 ^ n5933 ^ 1'b0 ;
  assign n37137 = ~x225 & n12369 ;
  assign n37138 = n37137 ^ n3385 ^ 1'b0 ;
  assign n37139 = ~n606 & n37138 ;
  assign n37140 = n37139 ^ n6968 ^ 1'b0 ;
  assign n37141 = n3805 & n12176 ;
  assign n37142 = n37141 ^ n26155 ^ 1'b0 ;
  assign n37143 = n37071 & ~n37142 ;
  assign n37144 = n37143 ^ n3059 ^ 1'b0 ;
  assign n37145 = n17522 ^ n11762 ^ 1'b0 ;
  assign n37146 = ~n1023 & n37145 ;
  assign n37147 = ~n15895 & n37146 ;
  assign n37148 = n11681 ^ n10657 ^ 1'b0 ;
  assign n37149 = n27735 & ~n37148 ;
  assign n37150 = n10832 & n13468 ;
  assign n37151 = n37150 ^ n3594 ^ 1'b0 ;
  assign n37152 = n37151 ^ n23133 ^ 1'b0 ;
  assign n37153 = n37152 ^ n16379 ^ 1'b0 ;
  assign n37154 = n932 & n37153 ;
  assign n37155 = n14080 | n27974 ;
  assign n37156 = n18530 & ~n37155 ;
  assign n37157 = n35705 & ~n37156 ;
  assign n37158 = n2674 & n6120 ;
  assign n37159 = n37158 ^ n21990 ^ 1'b0 ;
  assign n37160 = ~n8888 & n37159 ;
  assign n37161 = n37160 ^ n891 ^ 1'b0 ;
  assign n37163 = n1160 & ~n9943 ;
  assign n37162 = n3249 & n29734 ;
  assign n37164 = n37163 ^ n37162 ^ 1'b0 ;
  assign n37165 = n37164 ^ n24938 ^ 1'b0 ;
  assign n37166 = ~n16436 & n37165 ;
  assign n37167 = ( n1527 & n20838 ) | ( n1527 & ~n30256 ) | ( n20838 & ~n30256 ) ;
  assign n37168 = n24079 ^ n2267 ^ 1'b0 ;
  assign n37169 = n37168 ^ n30281 ^ n26275 ;
  assign n37170 = n26185 & ~n30200 ;
  assign n37171 = n36332 & n37170 ;
  assign n37172 = n9798 ^ n8406 ^ 1'b0 ;
  assign n37173 = n22417 | n37172 ;
  assign n37174 = n13688 | n37173 ;
  assign n37175 = n37174 ^ n6994 ^ 1'b0 ;
  assign n37176 = n15770 & ~n27380 ;
  assign n37177 = ~n15046 & n37176 ;
  assign n37178 = n25802 ^ n3930 ^ 1'b0 ;
  assign n37179 = ~n32170 & n33877 ;
  assign n37180 = ~n1929 & n37179 ;
  assign n37181 = n28925 ^ n24961 ^ 1'b0 ;
  assign n37182 = n13429 & n37181 ;
  assign n37183 = n13672 ^ n8216 ^ 1'b0 ;
  assign n37184 = n15911 | n37183 ;
  assign n37185 = n1442 & n26843 ;
  assign n37186 = n3416 & n24691 ;
  assign n37187 = n12722 & n37186 ;
  assign n37188 = n37187 ^ n12123 ^ 1'b0 ;
  assign n37189 = n22118 ^ n5639 ^ 1'b0 ;
  assign n37190 = n9628 & ~n26303 ;
  assign n37191 = n37190 ^ n8978 ^ 1'b0 ;
  assign n37192 = n7020 | n10433 ;
  assign n37193 = n4415 & ~n29267 ;
  assign n37194 = n37193 ^ n15998 ^ 1'b0 ;
  assign n37195 = n30824 & ~n37194 ;
  assign n37196 = n37195 ^ n6270 ^ 1'b0 ;
  assign n37197 = n7035 ^ n6303 ^ 1'b0 ;
  assign n37198 = n2370 | n32219 ;
  assign n37199 = n31065 | n37198 ;
  assign n37200 = n9378 | n13541 ;
  assign n37201 = n13482 & ~n37200 ;
  assign n37202 = x112 | n29894 ;
  assign n37203 = n16313 ^ n3190 ^ 1'b0 ;
  assign n37204 = n22739 | n24960 ;
  assign n37205 = ~n27818 & n37204 ;
  assign n37206 = ~n29653 & n30500 ;
  assign n37207 = n28826 ^ n274 ^ 1'b0 ;
  assign n37208 = ~n15707 & n36465 ;
  assign n37209 = n37208 ^ n3590 ^ 1'b0 ;
  assign n37210 = n7860 & ~n13966 ;
  assign n37211 = n25187 & n30423 ;
  assign n37212 = n29082 & n37211 ;
  assign n37213 = n15707 ^ n13037 ^ 1'b0 ;
  assign n37214 = ~n37212 & n37213 ;
  assign n37215 = n920 & ~n7605 ;
  assign n37216 = n37215 ^ n24455 ^ 1'b0 ;
  assign n37217 = n19885 ^ x172 ^ 1'b0 ;
  assign n37218 = n16500 ^ n2499 ^ 1'b0 ;
  assign n37219 = n1395 & n35785 ;
  assign n37220 = ~x29 & n23504 ;
  assign n37221 = n22147 ^ n16233 ^ n3036 ;
  assign n37222 = n22301 | n37221 ;
  assign n37223 = n37220 & ~n37222 ;
  assign n37224 = n15503 ^ n3412 ^ n1185 ;
  assign n37226 = n31336 ^ n17152 ^ n8734 ;
  assign n37225 = ~n12688 & n19453 ;
  assign n37227 = n37226 ^ n37225 ^ 1'b0 ;
  assign n37228 = ( n12830 & ~n37224 ) | ( n12830 & n37227 ) | ( ~n37224 & n37227 ) ;
  assign n37229 = n37228 ^ n26896 ^ n12564 ;
  assign n37230 = n1553 & n4404 ;
  assign n37231 = n37230 ^ n18415 ^ 1'b0 ;
  assign n37232 = ~n14941 & n25305 ;
  assign n37233 = n9202 & n37232 ;
  assign n37234 = n37233 ^ n13240 ^ 1'b0 ;
  assign n37235 = n14236 | n15025 ;
  assign n37236 = n9321 | n10273 ;
  assign n37237 = n35944 | n37236 ;
  assign n37238 = x115 & ~n15887 ;
  assign n37239 = ~n37237 & n37238 ;
  assign n37240 = ( n359 & ~n6731 ) | ( n359 & n12854 ) | ( ~n6731 & n12854 ) ;
  assign n37241 = n7085 ^ n2797 ^ 1'b0 ;
  assign n37242 = n18478 ^ n5510 ^ 1'b0 ;
  assign n37243 = n14121 & ~n37242 ;
  assign n37244 = n4608 ^ n2121 ^ 1'b0 ;
  assign n37245 = ~n5676 & n37244 ;
  assign n37246 = ( ~n16003 & n37243 ) | ( ~n16003 & n37245 ) | ( n37243 & n37245 ) ;
  assign n37247 = n10982 & ~n36642 ;
  assign n37248 = ~n37246 & n37247 ;
  assign n37249 = n29043 ^ n22787 ^ 1'b0 ;
  assign n37250 = n4849 & ~n26245 ;
  assign n37251 = n37250 ^ n1249 ^ 1'b0 ;
  assign n37252 = n9494 & ~n37251 ;
  assign n37253 = n1944 & ~n4253 ;
  assign n37254 = ~n3714 & n37253 ;
  assign n37255 = n37254 ^ n11982 ^ 1'b0 ;
  assign n37256 = ~n15427 & n37255 ;
  assign n37257 = ( n18543 & ~n23073 ) | ( n18543 & n37256 ) | ( ~n23073 & n37256 ) ;
  assign n37258 = n25459 ^ n17914 ^ 1'b0 ;
  assign n37259 = n35435 & n37258 ;
  assign n37260 = n22220 ^ n10932 ^ 1'b0 ;
  assign n37262 = ~n5958 & n7480 ;
  assign n37263 = n3712 & n37262 ;
  assign n37264 = n37263 ^ n27464 ^ 1'b0 ;
  assign n37261 = n29292 | n29902 ;
  assign n37265 = n37264 ^ n37261 ^ 1'b0 ;
  assign n37266 = n15353 | n17594 ;
  assign n37267 = n37266 ^ n6644 ^ n1945 ;
  assign n37269 = n16909 & n34662 ;
  assign n37268 = n5056 & ~n32990 ;
  assign n37270 = n37269 ^ n37268 ^ n2493 ;
  assign n37271 = n1636 | n20783 ;
  assign n37272 = n37271 ^ x180 ^ 1'b0 ;
  assign n37273 = n5622 & ~n19169 ;
  assign n37274 = n12460 | n16576 ;
  assign n37275 = n28030 | n37274 ;
  assign n37276 = n12787 & ~n37275 ;
  assign n37277 = n37133 ^ n15785 ^ 1'b0 ;
  assign n37278 = n2831 | n17369 ;
  assign n37279 = n27480 ^ n17950 ^ 1'b0 ;
  assign n37280 = ~n7022 & n37279 ;
  assign n37281 = n20337 & n37280 ;
  assign n37282 = ~n37278 & n37281 ;
  assign n37284 = n13500 ^ n10022 ^ n7714 ;
  assign n37283 = n7399 | n11071 ;
  assign n37285 = n37284 ^ n37283 ^ 1'b0 ;
  assign n37286 = n12140 & n37285 ;
  assign n37287 = n16803 & n18046 ;
  assign n37288 = n31694 & ~n37287 ;
  assign n37289 = n32147 ^ n13513 ^ 1'b0 ;
  assign n37290 = ( ~x100 & n677 ) | ( ~x100 & n25697 ) | ( n677 & n25697 ) ;
  assign n37291 = n37290 ^ n30626 ^ n4190 ;
  assign n37292 = n37291 ^ n3400 ^ 1'b0 ;
  assign n37293 = n15534 & ~n33188 ;
  assign n37294 = n1864 & n37293 ;
  assign n37295 = n6182 | n13737 ;
  assign n37296 = ~n4338 & n10439 ;
  assign n37297 = n37296 ^ n29575 ^ 1'b0 ;
  assign n37298 = n37295 & ~n37297 ;
  assign n37299 = n17488 & n37298 ;
  assign n37300 = n23150 ^ n5986 ^ 1'b0 ;
  assign n37301 = n37300 ^ n30024 ^ n2746 ;
  assign n37305 = ~n1147 & n2623 ;
  assign n37306 = ~n2623 & n37305 ;
  assign n37307 = ~n3555 & n5722 ;
  assign n37308 = n3555 & n37307 ;
  assign n37309 = ~n3178 & n37308 ;
  assign n37310 = n8210 & ~n37309 ;
  assign n37311 = ( n1963 & n37306 ) | ( n1963 & n37310 ) | ( n37306 & n37310 ) ;
  assign n37312 = n812 | n7781 ;
  assign n37313 = n812 & ~n37312 ;
  assign n37314 = n4130 | n37313 ;
  assign n37315 = n4130 & ~n37314 ;
  assign n37316 = n763 & n37315 ;
  assign n37317 = n37316 ^ n12041 ^ 1'b0 ;
  assign n37318 = n37311 & ~n37317 ;
  assign n37302 = n7043 | n13541 ;
  assign n37303 = n37302 ^ n4323 ^ 1'b0 ;
  assign n37304 = n29220 | n37303 ;
  assign n37319 = n37318 ^ n37304 ^ 1'b0 ;
  assign n37320 = n6619 & n15941 ;
  assign n37321 = n22941 & n37320 ;
  assign n37322 = n28567 ^ n10744 ^ 1'b0 ;
  assign n37323 = ~n3319 & n37322 ;
  assign n37324 = n37323 ^ n3672 ^ 1'b0 ;
  assign n37325 = n10928 & ~n32135 ;
  assign n37326 = n37325 ^ n24769 ^ n17229 ;
  assign n37327 = n6159 & ~n37212 ;
  assign n37329 = ~n6606 & n12720 ;
  assign n37328 = ~n5368 & n15469 ;
  assign n37330 = n37329 ^ n37328 ^ 1'b0 ;
  assign n37331 = ~n17069 & n37330 ;
  assign n37332 = n12745 | n17835 ;
  assign n37333 = n23493 ^ n14440 ^ 1'b0 ;
  assign n37334 = n2120 & n37333 ;
  assign n37335 = n23156 ^ n4718 ^ 1'b0 ;
  assign n37336 = ~n30729 & n37335 ;
  assign n37337 = n7749 ^ n3701 ^ 1'b0 ;
  assign n37338 = n17543 ^ n10074 ^ 1'b0 ;
  assign n37339 = ~n5709 & n37338 ;
  assign n37340 = n37339 ^ n17190 ^ 1'b0 ;
  assign n37341 = x31 & ~n37340 ;
  assign n37342 = n37341 ^ n18701 ^ n3768 ;
  assign n37343 = n4124 & n8632 ;
  assign n37344 = n34523 ^ n22618 ^ 1'b0 ;
  assign n37345 = n37343 & n37344 ;
  assign n37346 = n1742 & ~n12297 ;
  assign n37347 = n12459 ^ n7879 ^ 1'b0 ;
  assign n37348 = n12383 | n37347 ;
  assign n37349 = n37346 | n37348 ;
  assign n37350 = n14768 ^ n4139 ^ 1'b0 ;
  assign n37352 = n9540 ^ x187 ^ 1'b0 ;
  assign n37351 = n14470 | n16014 ;
  assign n37353 = n37352 ^ n37351 ^ 1'b0 ;
  assign n37354 = n37353 ^ n11204 ^ 1'b0 ;
  assign n37355 = n24343 ^ n3195 ^ 1'b0 ;
  assign n37356 = n21990 | n37355 ;
  assign n37357 = n2272 & ~n37356 ;
  assign n37358 = n17619 ^ n675 ^ 1'b0 ;
  assign n37359 = n22054 ^ n4458 ^ 1'b0 ;
  assign n37360 = ~n4055 & n37359 ;
  assign n37361 = ~n10790 & n37360 ;
  assign n37362 = n20667 ^ n17012 ^ n2681 ;
  assign n37363 = n37361 & n37362 ;
  assign n37365 = n24946 ^ n2011 ^ 1'b0 ;
  assign n37366 = ~n5119 & n37365 ;
  assign n37367 = n13805 & n37366 ;
  assign n37368 = n37367 ^ n4834 ^ 1'b0 ;
  assign n37369 = n37368 ^ n826 ^ 1'b0 ;
  assign n37364 = n1966 & n35214 ;
  assign n37370 = n37369 ^ n37364 ^ 1'b0 ;
  assign n37371 = n7455 & n8307 ;
  assign n37372 = n37371 ^ n13518 ^ 1'b0 ;
  assign n37373 = ~n5076 & n20684 ;
  assign n37374 = n8295 & n37373 ;
  assign n37375 = ( ~n5790 & n37372 ) | ( ~n5790 & n37374 ) | ( n37372 & n37374 ) ;
  assign n37378 = ~n4193 & n27388 ;
  assign n37379 = n277 & n37378 ;
  assign n37376 = n19523 & n33074 ;
  assign n37377 = n37376 ^ n33586 ^ 1'b0 ;
  assign n37380 = n37379 ^ n37377 ^ n11181 ;
  assign n37381 = n3403 | n9742 ;
  assign n37385 = n31621 ^ n23779 ^ 1'b0 ;
  assign n37386 = n8939 | n37385 ;
  assign n37387 = n30313 ^ n11522 ^ 1'b0 ;
  assign n37388 = n37386 | n37387 ;
  assign n37382 = n5885 | n24203 ;
  assign n37383 = n5987 & ~n37382 ;
  assign n37384 = n2258 & ~n37383 ;
  assign n37389 = n37388 ^ n37384 ^ 1'b0 ;
  assign n37390 = n8978 & ~n31754 ;
  assign n37391 = n37390 ^ n4559 ^ 1'b0 ;
  assign n37392 = n37391 ^ n24283 ^ 1'b0 ;
  assign n37393 = ~n6548 & n17201 ;
  assign n37394 = n37393 ^ n15998 ^ 1'b0 ;
  assign n37395 = n4327 & ~n37394 ;
  assign n37396 = n540 & ~n9853 ;
  assign n37397 = n37396 ^ n16341 ^ 1'b0 ;
  assign n37398 = ~n9754 & n15838 ;
  assign n37399 = n37398 ^ n12627 ^ 1'b0 ;
  assign n37400 = n6934 & n37399 ;
  assign n37401 = n31236 & n37400 ;
  assign n37402 = n3772 & n19650 ;
  assign n37403 = n1853 | n23087 ;
  assign n37404 = n37403 ^ n24770 ^ 1'b0 ;
  assign n37405 = ~n1744 & n30756 ;
  assign n37406 = n20064 & n37405 ;
  assign n37407 = n37406 ^ n34112 ^ 1'b0 ;
  assign n37408 = n1866 & ~n22982 ;
  assign n37409 = ~n6920 & n10898 ;
  assign n37411 = n547 & n13934 ;
  assign n37412 = n29393 & n37411 ;
  assign n37410 = n8042 | n13576 ;
  assign n37413 = n37412 ^ n37410 ^ 1'b0 ;
  assign n37414 = n31070 & ~n33756 ;
  assign n37417 = n8319 | n9515 ;
  assign n37415 = n4970 ^ n3698 ^ 1'b0 ;
  assign n37416 = n9705 & n37415 ;
  assign n37418 = n37417 ^ n37416 ^ 1'b0 ;
  assign n37419 = ~n15438 & n37418 ;
  assign n37420 = n453 & n10196 ;
  assign n37421 = n6226 | n15003 ;
  assign n37422 = n2564 | n37421 ;
  assign n37423 = n37422 ^ n37400 ^ n11159 ;
  assign n37424 = n9855 | n15303 ;
  assign n37425 = n7729 & n12789 ;
  assign n37426 = n37425 ^ n14754 ^ 1'b0 ;
  assign n37427 = n23152 & ~n32194 ;
  assign n37428 = n37426 & n37427 ;
  assign n37429 = n883 | n5425 ;
  assign n37430 = n883 & ~n37429 ;
  assign n37431 = n10437 & ~n37430 ;
  assign n37432 = ~n10437 & n37431 ;
  assign n37433 = n1778 & ~n37432 ;
  assign n37434 = ~n8684 & n37433 ;
  assign n37435 = ( n6188 & n19336 ) | ( n6188 & ~n37434 ) | ( n19336 & ~n37434 ) ;
  assign n37436 = n30989 ^ n2023 ^ 1'b0 ;
  assign n37437 = n37435 & n37436 ;
  assign n37438 = n34071 ^ n30181 ^ n26089 ;
  assign n37439 = ~n3513 & n9708 ;
  assign n37440 = n14372 ^ n6566 ^ n3725 ;
  assign n37441 = n5604 | n37440 ;
  assign n37442 = n8994 & ~n31125 ;
  assign n37443 = n1896 & ~n24172 ;
  assign n37444 = n29299 ^ n6864 ^ 1'b0 ;
  assign n37445 = ~x92 & n4691 ;
  assign n37446 = n32021 ^ n15437 ^ 1'b0 ;
  assign n37447 = n17728 ^ n11473 ^ 1'b0 ;
  assign n37448 = n26300 ^ n21819 ^ 1'b0 ;
  assign n37449 = n37447 & ~n37448 ;
  assign n37450 = n37449 ^ n16385 ^ 1'b0 ;
  assign n37451 = n17412 & ~n37450 ;
  assign n37452 = x163 & ~n34355 ;
  assign n37453 = n9209 ^ n4473 ^ n3440 ;
  assign n37458 = ~n317 & n7207 ;
  assign n37459 = n317 & n37458 ;
  assign n37460 = ~n3996 & n37459 ;
  assign n37461 = ~n709 & n2211 ;
  assign n37462 = ~n2211 & n37461 ;
  assign n37463 = n37460 & ~n37462 ;
  assign n37464 = ~n37460 & n37463 ;
  assign n37465 = n1708 & n37464 ;
  assign n37454 = n747 & n2757 ;
  assign n37455 = ~n747 & n37454 ;
  assign n37456 = n2272 & ~n37455 ;
  assign n37457 = n19507 & ~n37456 ;
  assign n37466 = n37465 ^ n37457 ^ 1'b0 ;
  assign n37467 = n14590 | n18356 ;
  assign n37468 = n14845 ^ n14770 ^ 1'b0 ;
  assign n37469 = n3917 | n9207 ;
  assign n37470 = n2922 | n37469 ;
  assign n37471 = n22238 & n37470 ;
  assign n37472 = n37471 ^ n30361 ^ 1'b0 ;
  assign n37473 = n361 & n11386 ;
  assign n37474 = ~n37115 & n37473 ;
  assign n37475 = n10492 ^ n5519 ^ n613 ;
  assign n37476 = n37475 ^ n25537 ^ 1'b0 ;
  assign n37477 = n12536 ^ n10499 ^ 1'b0 ;
  assign n37478 = n14715 ^ n6516 ^ 1'b0 ;
  assign n37479 = n9024 & ~n37478 ;
  assign n37480 = n37479 ^ n5580 ^ 1'b0 ;
  assign n37481 = n37480 ^ n20337 ^ n19319 ;
  assign n37482 = n12262 | n37481 ;
  assign n37483 = n7183 & ~n37482 ;
  assign n37484 = n6260 ^ n2644 ^ 1'b0 ;
  assign n37485 = n20645 ^ n815 ^ 1'b0 ;
  assign n37486 = n37484 & n37485 ;
  assign n37487 = n28869 & ~n29724 ;
  assign n37488 = n37487 ^ n7555 ^ 1'b0 ;
  assign n37489 = n24987 ^ n11981 ^ 1'b0 ;
  assign n37490 = ~n7752 & n14652 ;
  assign n37491 = ~n37489 & n37490 ;
  assign n37492 = n11784 ^ n8195 ^ 1'b0 ;
  assign n37493 = n4906 ^ n2142 ^ n553 ;
  assign n37494 = ( n17619 & n37492 ) | ( n17619 & ~n37493 ) | ( n37492 & ~n37493 ) ;
  assign n37495 = n13960 & n27192 ;
  assign n37496 = n33438 & n34990 ;
  assign n37497 = n37496 ^ n16307 ^ 1'b0 ;
  assign n37500 = n2041 & n2269 ;
  assign n37501 = ~n4642 & n37500 ;
  assign n37498 = n25467 ^ n20041 ^ 1'b0 ;
  assign n37499 = ~n19693 & n37498 ;
  assign n37502 = n37501 ^ n37499 ^ 1'b0 ;
  assign n37503 = n15910 ^ n7229 ^ 1'b0 ;
  assign n37504 = ~n18023 & n37503 ;
  assign n37505 = n37504 ^ n10234 ^ 1'b0 ;
  assign n37506 = n25963 ^ n8349 ^ 1'b0 ;
  assign n37507 = ~n28104 & n31271 ;
  assign n37508 = n14487 & n27929 ;
  assign n37509 = n37508 ^ n4910 ^ 1'b0 ;
  assign n37510 = n37509 ^ n18385 ^ 1'b0 ;
  assign n37511 = n32751 & ~n37510 ;
  assign n37512 = n809 & n7721 ;
  assign n37513 = n5879 & n37512 ;
  assign n37514 = n7195 & n11431 ;
  assign n37515 = n37514 ^ n17609 ^ 1'b0 ;
  assign n37516 = n7191 ^ x17 ^ 1'b0 ;
  assign n37517 = ~n30116 & n37516 ;
  assign n37518 = n23164 ^ n5119 ^ 1'b0 ;
  assign n37519 = n37517 & n37518 ;
  assign n37520 = ( n4431 & n12373 ) | ( n4431 & ~n32024 ) | ( n12373 & ~n32024 ) ;
  assign n37521 = n22532 ^ n13347 ^ 1'b0 ;
  assign n37522 = n19016 ^ n12052 ^ 1'b0 ;
  assign n37523 = n4934 ^ n635 ^ 1'b0 ;
  assign n37524 = n33347 | n37523 ;
  assign n37525 = n11206 ^ n4619 ^ 1'b0 ;
  assign n37526 = x180 & ~n33602 ;
  assign n37527 = n37526 ^ n8835 ^ 1'b0 ;
  assign n37528 = n37383 ^ n7050 ^ 1'b0 ;
  assign n37530 = ( n613 & n11978 ) | ( n613 & ~n20772 ) | ( n11978 & ~n20772 ) ;
  assign n37529 = ( ~n6187 & n7716 ) | ( ~n6187 & n30810 ) | ( n7716 & n30810 ) ;
  assign n37531 = n37530 ^ n37529 ^ 1'b0 ;
  assign n37532 = n9829 & ~n26505 ;
  assign n37533 = n35000 ^ n22490 ^ 1'b0 ;
  assign n37534 = n28745 & n37533 ;
  assign n37535 = ~n922 & n17326 ;
  assign n37536 = n3728 ^ n679 ^ 1'b0 ;
  assign n37537 = n25682 & ~n37536 ;
  assign n37538 = n37537 ^ n911 ^ 1'b0 ;
  assign n37539 = ~n3362 & n21475 ;
  assign n37540 = n16102 ^ n5051 ^ 1'b0 ;
  assign n37541 = n6414 | n37540 ;
  assign n37542 = n37541 ^ n34814 ^ 1'b0 ;
  assign n37543 = n7775 | n30698 ;
  assign n37544 = n19690 & ~n37543 ;
  assign n37545 = n4222 & ~n37544 ;
  assign n37546 = n37545 ^ n6190 ^ 1'b0 ;
  assign n37547 = n2912 ^ n2537 ^ 1'b0 ;
  assign n37548 = n37546 & n37547 ;
  assign n37549 = n1521 & ~n28848 ;
  assign n37550 = ~n16058 & n37549 ;
  assign n37551 = ( n8873 & n24449 ) | ( n8873 & n25978 ) | ( n24449 & n25978 ) ;
  assign n37552 = ~n3996 & n33484 ;
  assign n37553 = n21434 & n37552 ;
  assign n37554 = n12728 | n23910 ;
  assign n37555 = ~n9965 & n18670 ;
  assign n37556 = n11253 & ~n15008 ;
  assign n37557 = n6274 | n18785 ;
  assign n37558 = n37557 ^ n7972 ^ 1'b0 ;
  assign n37559 = n3458 & ~n37558 ;
  assign n37560 = n3894 ^ n2848 ^ 1'b0 ;
  assign n37561 = n8467 ^ n4268 ^ 1'b0 ;
  assign n37562 = ( n30855 & ~n37560 ) | ( n30855 & n37561 ) | ( ~n37560 & n37561 ) ;
  assign n37563 = n36751 ^ n15961 ^ n7859 ;
  assign n37564 = ~n2653 & n37563 ;
  assign n37565 = n8690 ^ x3 ^ 1'b0 ;
  assign n37566 = n30371 ^ n10066 ^ 1'b0 ;
  assign n37567 = ~n11659 & n19501 ;
  assign n37568 = n1545 & n16430 ;
  assign n37569 = n16663 ^ n12124 ^ 1'b0 ;
  assign n37570 = ( n17426 & ~n37568 ) | ( n17426 & n37569 ) | ( ~n37568 & n37569 ) ;
  assign n37571 = n7113 & n36790 ;
  assign n37572 = ~n37570 & n37571 ;
  assign n37573 = n10695 & ~n27522 ;
  assign n37574 = n37573 ^ n21497 ^ 1'b0 ;
  assign n37575 = n11127 & ~n37574 ;
  assign n37576 = n11965 | n37575 ;
  assign n37577 = n27834 | n37576 ;
  assign n37578 = n33791 ^ n5025 ^ 1'b0 ;
  assign n37579 = n37577 & ~n37578 ;
  assign n37580 = n3420 & n11728 ;
  assign n37581 = n24468 | n37580 ;
  assign n37582 = n31564 & ~n37581 ;
  assign n37583 = n25305 ^ n1369 ^ 1'b0 ;
  assign n37584 = n37058 ^ n7961 ^ n4830 ;
  assign n37585 = n7019 | n34081 ;
  assign n37586 = n31994 ^ n27122 ^ 1'b0 ;
  assign n37587 = n5918 | n37586 ;
  assign n37588 = n7797 & n12928 ;
  assign n37590 = n7462 & n23810 ;
  assign n37589 = ~n364 & n3734 ;
  assign n37591 = n37590 ^ n37589 ^ 1'b0 ;
  assign n37592 = n37591 ^ n4254 ^ 1'b0 ;
  assign n37593 = ~n34681 & n37592 ;
  assign n37594 = n30042 ^ n14946 ^ 1'b0 ;
  assign n37595 = n26716 ^ n17279 ^ 1'b0 ;
  assign n37596 = n37594 & ~n37595 ;
  assign n37597 = n9010 ^ n8116 ^ n3812 ;
  assign n37598 = ( n8536 & n18518 ) | ( n8536 & n37597 ) | ( n18518 & n37597 ) ;
  assign n37599 = n22702 ^ n6289 ^ 1'b0 ;
  assign n37600 = n4547 & n7643 ;
  assign n37601 = n37600 ^ n7629 ^ 1'b0 ;
  assign n37602 = n10277 & n32617 ;
  assign n37603 = n37601 & n37602 ;
  assign n37604 = n12430 & n16395 ;
  assign n37605 = n37604 ^ n2549 ^ 1'b0 ;
  assign n37606 = n12138 | n13155 ;
  assign n37607 = n37606 ^ n23907 ^ n14218 ;
  assign n37608 = ~n14989 & n37607 ;
  assign n37609 = n7586 & n37608 ;
  assign n37610 = ~n9957 & n15259 ;
  assign n37611 = ( n3223 & ~n4646 ) | ( n3223 & n24311 ) | ( ~n4646 & n24311 ) ;
  assign n37612 = n3546 & n20361 ;
  assign n37613 = ( x40 & ~n22222 ) | ( x40 & n37612 ) | ( ~n22222 & n37612 ) ;
  assign n37614 = n7013 ^ n4867 ^ 1'b0 ;
  assign n37615 = n15412 ^ n9009 ^ n5590 ;
  assign n37616 = ~n37614 & n37615 ;
  assign n37617 = n34231 ^ n1107 ^ 1'b0 ;
  assign n37618 = n31805 & ~n37617 ;
  assign n37619 = n30572 & n37618 ;
  assign n37620 = ~n1648 & n19974 ;
  assign n37621 = n27787 ^ n9425 ^ 1'b0 ;
  assign n37622 = ~n18034 & n37621 ;
  assign n37623 = n4078 ^ x50 ^ 1'b0 ;
  assign n37624 = n37623 ^ n15894 ^ 1'b0 ;
  assign n37627 = n8024 ^ n300 ^ 1'b0 ;
  assign n37628 = n7579 & n37627 ;
  assign n37625 = ~n12295 & n31273 ;
  assign n37626 = n18290 & n37625 ;
  assign n37629 = n37628 ^ n37626 ^ 1'b0 ;
  assign n37634 = n9142 & ~n13924 ;
  assign n37633 = ~n3307 & n16928 ;
  assign n37635 = n37634 ^ n37633 ^ 1'b0 ;
  assign n37630 = n37615 ^ n24655 ^ 1'b0 ;
  assign n37631 = n18149 & n37630 ;
  assign n37632 = n36492 & ~n37631 ;
  assign n37636 = n37635 ^ n37632 ^ n2678 ;
  assign n37637 = n18277 ^ n16069 ^ 1'b0 ;
  assign n37638 = ~n18463 & n37637 ;
  assign n37639 = n33822 ^ n5785 ^ 1'b0 ;
  assign n37642 = ~n2789 & n4431 ;
  assign n37640 = n2396 & n2988 ;
  assign n37641 = ~n21952 & n37640 ;
  assign n37643 = n37642 ^ n37641 ^ 1'b0 ;
  assign n37644 = n4596 ^ n1748 ^ 1'b0 ;
  assign n37645 = ~n37643 & n37644 ;
  assign n37646 = n1802 & ~n12575 ;
  assign n37649 = n13780 ^ n2037 ^ 1'b0 ;
  assign n37647 = n10208 & n22490 ;
  assign n37648 = ~n2525 & n37647 ;
  assign n37650 = n37649 ^ n37648 ^ n9276 ;
  assign n37651 = n37646 & ~n37650 ;
  assign n37652 = n32626 | n32709 ;
  assign n37653 = n37652 ^ n33281 ^ 1'b0 ;
  assign n37654 = n4790 & n14742 ;
  assign n37655 = n6177 & n37654 ;
  assign n37656 = n16114 & ~n37655 ;
  assign n37657 = n34069 ^ n30571 ^ 1'b0 ;
  assign n37658 = n4244 & n12359 ;
  assign n37659 = ~n7972 & n37658 ;
  assign n37660 = n26607 ^ n26605 ^ 1'b0 ;
  assign n37661 = n29817 | n37660 ;
  assign n37662 = n2625 & n37661 ;
  assign n37663 = ~n19990 & n35589 ;
  assign n37664 = ~n21475 & n28648 ;
  assign n37665 = n21743 ^ n12860 ^ 1'b0 ;
  assign n37666 = ~n37664 & n37665 ;
  assign n37668 = n32878 & n33420 ;
  assign n37667 = ~n4877 & n7623 ;
  assign n37669 = n37668 ^ n37667 ^ 1'b0 ;
  assign n37670 = n12176 ^ n4244 ^ 1'b0 ;
  assign n37671 = ( n10632 & n12864 ) | ( n10632 & ~n37670 ) | ( n12864 & ~n37670 ) ;
  assign n37672 = n37671 ^ n26251 ^ 1'b0 ;
  assign n37673 = n4248 ^ n1232 ^ n831 ;
  assign n37674 = n14752 | n18500 ;
  assign n37675 = n37674 ^ n3558 ^ 1'b0 ;
  assign n37676 = n37675 ^ n29770 ^ n28458 ;
  assign n37677 = n6618 ^ n6166 ^ 1'b0 ;
  assign n37678 = n30832 | n37677 ;
  assign n37679 = n2264 & ~n27211 ;
  assign n37680 = n11805 & ~n14593 ;
  assign n37681 = n37680 ^ n12754 ^ 1'b0 ;
  assign n37682 = n8861 & ~n37681 ;
  assign n37683 = ~n12952 & n28791 ;
  assign n37684 = n20748 & n37683 ;
  assign n37685 = n16422 ^ n879 ^ 1'b0 ;
  assign n37686 = ~n37684 & n37685 ;
  assign n37687 = n12748 ^ n3037 ^ 1'b0 ;
  assign n37688 = n30285 & ~n37687 ;
  assign n37689 = n28627 & ~n37688 ;
  assign n37690 = n15733 & ~n26597 ;
  assign n37691 = ~n10529 & n29187 ;
  assign n37692 = n2749 ^ x8 ^ 1'b0 ;
  assign n37693 = n5009 & ~n37692 ;
  assign n37694 = n1596 & ~n7898 ;
  assign n37695 = n37694 ^ n5197 ^ 1'b0 ;
  assign n37696 = n4496 & ~n31544 ;
  assign n37697 = n22649 & ~n35189 ;
  assign n37698 = n37696 & n37697 ;
  assign n37699 = n7791 | n30661 ;
  assign n37700 = ( n13306 & n32610 ) | ( n13306 & ~n33010 ) | ( n32610 & ~n33010 ) ;
  assign n37701 = n14494 ^ n4994 ^ 1'b0 ;
  assign n37702 = n23587 ^ n18841 ^ 1'b0 ;
  assign n37703 = ~n6612 & n37702 ;
  assign n37704 = n28916 ^ n1596 ^ 1'b0 ;
  assign n37705 = n8976 & ~n29713 ;
  assign n37706 = n37705 ^ n34233 ^ 1'b0 ;
  assign n37707 = n10240 ^ n4420 ^ 1'b0 ;
  assign n37708 = n24043 ^ n22542 ^ 1'b0 ;
  assign n37709 = ~n12028 & n37708 ;
  assign n37710 = n30769 & n37709 ;
  assign n37711 = n37710 ^ n12850 ^ 1'b0 ;
  assign n37712 = n37707 & ~n37711 ;
  assign n37713 = ~n3938 & n31332 ;
  assign n37714 = n37137 ^ n16271 ^ 1'b0 ;
  assign n37715 = ( n13154 & n14900 ) | ( n13154 & n31005 ) | ( n14900 & n31005 ) ;
  assign n37716 = n9246 & ~n37715 ;
  assign n37717 = n11786 & n37716 ;
  assign n37718 = ( n12732 & n35440 ) | ( n12732 & ~n37097 ) | ( n35440 & ~n37097 ) ;
  assign n37719 = n37718 ^ n8878 ^ 1'b0 ;
  assign n37720 = n16416 & n18953 ;
  assign n37721 = ~n25569 & n37720 ;
  assign n37722 = ~n2413 & n37721 ;
  assign n37723 = x66 & ~n5363 ;
  assign n37724 = n37723 ^ n27408 ^ 1'b0 ;
  assign n37725 = n4295 ^ n2759 ^ 1'b0 ;
  assign n37726 = n22629 | n37725 ;
  assign n37727 = n657 & ~n37726 ;
  assign n37728 = ~n1801 & n37727 ;
  assign n37729 = n35027 ^ n22751 ^ 1'b0 ;
  assign n37730 = n8607 & n37729 ;
  assign n37731 = n4423 & ~n37730 ;
  assign n37732 = ( n25277 & n33194 ) | ( n25277 & n37731 ) | ( n33194 & n37731 ) ;
  assign n37734 = n14580 ^ n11402 ^ 1'b0 ;
  assign n37735 = n10819 | n37734 ;
  assign n37733 = ~n5539 & n27188 ;
  assign n37736 = n37735 ^ n37733 ^ n11571 ;
  assign n37737 = n26917 ^ n10105 ^ 1'b0 ;
  assign n37738 = n37737 ^ n25554 ^ 1'b0 ;
  assign n37739 = n30134 ^ n3191 ^ 1'b0 ;
  assign n37740 = n971 & ~n6051 ;
  assign n37741 = n6574 & n11381 ;
  assign n37742 = ~n5203 & n37741 ;
  assign n37743 = n16290 & n37742 ;
  assign n37744 = n25002 ^ n8330 ^ 1'b0 ;
  assign n37745 = n37743 | n37744 ;
  assign n37746 = n14369 | n16227 ;
  assign n37747 = ( n2743 & n32184 ) | ( n2743 & ~n37746 ) | ( n32184 & ~n37746 ) ;
  assign n37748 = n36128 ^ n18557 ^ n10888 ;
  assign n37749 = n37748 ^ n33067 ^ n3546 ;
  assign n37750 = n7679 & n17895 ;
  assign n37751 = n19333 ^ n7258 ^ 1'b0 ;
  assign n37752 = n16610 & n37751 ;
  assign n37753 = n2004 & n25326 ;
  assign n37754 = n37753 ^ n6412 ^ 1'b0 ;
  assign n37755 = n2172 & ~n37754 ;
  assign n37756 = n37755 ^ n29098 ^ 1'b0 ;
  assign n37757 = n14032 ^ n6001 ^ 1'b0 ;
  assign n37758 = n562 & n30285 ;
  assign n37759 = n37758 ^ n13554 ^ 1'b0 ;
  assign n37760 = ~n17453 & n37759 ;
  assign n37761 = n37760 ^ n19390 ^ 1'b0 ;
  assign n37762 = n10971 ^ n9336 ^ 1'b0 ;
  assign n37763 = n26488 ^ n19349 ^ 1'b0 ;
  assign n37764 = n12841 | n20369 ;
  assign n37765 = ~n2192 & n3828 ;
  assign n37766 = ~n9532 & n37765 ;
  assign n37767 = n6639 & ~n20949 ;
  assign n37775 = n23830 ^ n8421 ^ n1458 ;
  assign n37768 = n26024 ^ n9067 ^ 1'b0 ;
  assign n37769 = n10569 & ~n37768 ;
  assign n37770 = n37769 ^ n1028 ^ 1'b0 ;
  assign n37771 = ~n10075 & n37770 ;
  assign n37772 = ~n29479 & n37771 ;
  assign n37773 = n1657 & n37772 ;
  assign n37774 = n20675 & ~n37773 ;
  assign n37776 = n37775 ^ n37774 ^ 1'b0 ;
  assign n37777 = n22084 | n30524 ;
  assign n37778 = ~n11601 & n13787 ;
  assign n37779 = n37121 ^ n7584 ^ 1'b0 ;
  assign n37780 = n37778 & ~n37779 ;
  assign n37781 = n7271 | n7859 ;
  assign n37782 = n20144 | n30215 ;
  assign n37783 = n32020 | n37501 ;
  assign n37784 = n8081 ^ n3172 ^ 1'b0 ;
  assign n37785 = n1435 & n2584 ;
  assign n37786 = n37785 ^ n24024 ^ n10111 ;
  assign n37787 = n35385 & ~n37786 ;
  assign n37788 = ~n25470 & n37787 ;
  assign n37789 = n22066 ^ n7464 ^ 1'b0 ;
  assign n37790 = ~n4082 & n29450 ;
  assign n37791 = n29952 ^ n17295 ^ 1'b0 ;
  assign n37792 = n28160 ^ n3513 ^ 1'b0 ;
  assign n37793 = ( ~n4387 & n11147 ) | ( ~n4387 & n37792 ) | ( n11147 & n37792 ) ;
  assign n37794 = n37793 ^ n12488 ^ 1'b0 ;
  assign n37795 = n25142 & ~n37794 ;
  assign n37797 = ~n7658 & n14622 ;
  assign n37798 = n37797 ^ n19488 ^ 1'b0 ;
  assign n37796 = n14526 | n16593 ;
  assign n37799 = n37798 ^ n37796 ^ 1'b0 ;
  assign n37800 = n36031 | n37799 ;
  assign n37801 = n37795 | n37800 ;
  assign n37802 = ~n28626 & n33399 ;
  assign n37803 = ~n35157 & n37802 ;
  assign n37804 = n5374 ^ n2988 ^ 1'b0 ;
  assign n37805 = n12638 ^ n2570 ^ 1'b0 ;
  assign n37806 = n37804 & n37805 ;
  assign n37807 = ~n20619 & n27239 ;
  assign n37808 = n7407 & ~n35905 ;
  assign n37809 = n9657 | n12139 ;
  assign n37810 = n37809 ^ n24573 ^ 1'b0 ;
  assign n37811 = n17791 & n37810 ;
  assign n37812 = n37811 ^ n2331 ^ n1832 ;
  assign n37813 = n13710 ^ n10231 ^ 1'b0 ;
  assign n37814 = n1328 & n9119 ;
  assign n37815 = n34129 & n37814 ;
  assign n37816 = n5461 ^ n2501 ^ 1'b0 ;
  assign n37817 = ~n3036 & n32059 ;
  assign n37818 = ~n3568 & n37817 ;
  assign n37819 = ~n11400 & n37818 ;
  assign n37820 = n13620 & ~n32360 ;
  assign n37821 = ~n7676 & n8730 ;
  assign n37822 = ~n31586 & n37821 ;
  assign n37825 = n11976 & ~n12074 ;
  assign n37823 = n28148 ^ n23806 ^ 1'b0 ;
  assign n37824 = n17926 & n37823 ;
  assign n37826 = n37825 ^ n37824 ^ 1'b0 ;
  assign n37827 = n425 & n3036 ;
  assign n37828 = n8520 | n19823 ;
  assign n37829 = n37827 & ~n37828 ;
  assign n37830 = n21831 & n32147 ;
  assign n37831 = n37830 ^ n24920 ^ 1'b0 ;
  assign n37832 = n31275 & ~n37572 ;
  assign n37833 = n7583 & n37832 ;
  assign n37834 = n2516 & ~n29972 ;
  assign n37835 = ( n11485 & ~n20081 ) | ( n11485 & n28499 ) | ( ~n20081 & n28499 ) ;
  assign n37836 = n1053 & ~n16119 ;
  assign n37837 = n16348 ^ n6709 ^ 1'b0 ;
  assign n37838 = n6531 & ~n14597 ;
  assign n37839 = n3613 & ~n8282 ;
  assign n37840 = n37839 ^ n26322 ^ 1'b0 ;
  assign n37841 = n5792 ^ n317 ^ 1'b0 ;
  assign n37842 = n18003 | n37841 ;
  assign n37843 = n4039 & ~n16473 ;
  assign n37844 = n37843 ^ n9836 ^ 1'b0 ;
  assign n37845 = n6833 & ~n37844 ;
  assign n37846 = n6881 ^ n3820 ^ 1'b0 ;
  assign n37847 = n285 | n17801 ;
  assign n37848 = n8984 | n37847 ;
  assign n37849 = n37848 ^ n36088 ^ 1'b0 ;
  assign n37850 = n17488 ^ x29 ^ 1'b0 ;
  assign n37851 = n2912 | n37850 ;
  assign n37852 = n10481 | n28472 ;
  assign n37853 = n9956 ^ n1966 ^ 1'b0 ;
  assign n37854 = ~n32937 & n37853 ;
  assign n37855 = n15464 ^ n8214 ^ n6985 ;
  assign n37856 = n37855 ^ n25775 ^ 1'b0 ;
  assign n37857 = n11262 & ~n37856 ;
  assign n37858 = n5634 ^ n1147 ^ 1'b0 ;
  assign n37859 = n5432 & ~n20254 ;
  assign n37860 = n37859 ^ n20056 ^ 1'b0 ;
  assign n37861 = n32830 ^ n6522 ^ 1'b0 ;
  assign n37866 = n3012 & n6659 ;
  assign n37867 = n37866 ^ n4132 ^ 1'b0 ;
  assign n37868 = n7474 & ~n37867 ;
  assign n37865 = n9475 | n16980 ;
  assign n37869 = n37868 ^ n37865 ^ 1'b0 ;
  assign n37870 = n5482 | n37869 ;
  assign n37862 = n2481 & n11804 ;
  assign n37863 = n37862 ^ n1267 ^ 1'b0 ;
  assign n37864 = n37863 ^ n1203 ^ 1'b0 ;
  assign n37871 = n37870 ^ n37864 ^ n22625 ;
  assign n37872 = n19873 | n24545 ;
  assign n37873 = n20358 & n37872 ;
  assign n37874 = n2967 & n37873 ;
  assign n37875 = n37874 ^ n8518 ^ n7255 ;
  assign n37879 = n7786 & ~n12469 ;
  assign n37880 = n37879 ^ n977 ^ 1'b0 ;
  assign n37881 = n8499 & n37880 ;
  assign n37877 = ~n890 & n1906 ;
  assign n37878 = n1853 & n37877 ;
  assign n37882 = n37881 ^ n37878 ^ n4410 ;
  assign n37876 = n13510 & ~n28862 ;
  assign n37883 = n37882 ^ n37876 ^ 1'b0 ;
  assign n37884 = n33934 ^ n14070 ^ 1'b0 ;
  assign n37885 = n2061 & ~n12329 ;
  assign n37886 = n16429 ^ n558 ^ 1'b0 ;
  assign n37887 = n15061 & n37886 ;
  assign n37888 = n2552 & ~n16753 ;
  assign n37889 = n37888 ^ n37089 ^ 1'b0 ;
  assign n37890 = n37889 ^ n33450 ^ n2178 ;
  assign n37891 = n9019 & n32930 ;
  assign n37892 = n37891 ^ n400 ^ 1'b0 ;
  assign n37893 = n26535 ^ n15100 ^ 1'b0 ;
  assign n37894 = n34920 ^ n23574 ^ 1'b0 ;
  assign n37895 = ~n11185 & n37894 ;
  assign n37896 = n37895 ^ n4488 ^ 1'b0 ;
  assign n37897 = n8064 & ~n37896 ;
  assign n37898 = n14900 ^ n1899 ^ 1'b0 ;
  assign n37899 = n19229 ^ n9463 ^ 1'b0 ;
  assign n37901 = n1851 ^ n1736 ^ 1'b0 ;
  assign n37902 = n6059 & n37901 ;
  assign n37903 = n33169 ^ n10176 ^ 1'b0 ;
  assign n37904 = n37902 & n37903 ;
  assign n37900 = n22334 ^ n14144 ^ 1'b0 ;
  assign n37905 = n37904 ^ n37900 ^ n26056 ;
  assign n37906 = n37905 ^ n26952 ^ n20103 ;
  assign n37907 = n7390 ^ n5300 ^ n2037 ;
  assign n37908 = n2174 | n10976 ;
  assign n37909 = n1851 & ~n37908 ;
  assign n37910 = n8936 ^ n3186 ^ 1'b0 ;
  assign n37911 = ~n3795 & n37910 ;
  assign n37912 = n29916 ^ n15348 ^ n5418 ;
  assign n37913 = n37912 ^ n21901 ^ n17641 ;
  assign n37914 = n9711 & n37913 ;
  assign n37915 = ~n19319 & n23715 ;
  assign n37916 = n37915 ^ n7537 ^ 1'b0 ;
  assign n37917 = n37916 ^ n26654 ^ 1'b0 ;
  assign n37918 = ( n2392 & n27886 ) | ( n2392 & ~n30874 ) | ( n27886 & ~n30874 ) ;
  assign n37919 = n5368 ^ n4991 ^ 1'b0 ;
  assign n37920 = n8390 & ~n37919 ;
  assign n37921 = n37920 ^ n36722 ^ n16318 ;
  assign n37922 = n36838 ^ n1606 ^ 1'b0 ;
  assign n37923 = n37922 ^ n15126 ^ 1'b0 ;
  assign n37924 = ( ~n4493 & n11379 ) | ( ~n4493 & n24640 ) | ( n11379 & n24640 ) ;
  assign n37925 = n17818 ^ n3616 ^ 1'b0 ;
  assign n37926 = ~n37924 & n37925 ;
  assign n37927 = n4984 & n8254 ;
  assign n37928 = n9442 & n37927 ;
  assign n37929 = n37928 ^ n10416 ^ 1'b0 ;
  assign n37930 = ~n24340 & n37929 ;
  assign n37931 = n1083 & n3947 ;
  assign n37932 = n37931 ^ n5578 ^ 1'b0 ;
  assign n37933 = ~n35216 & n37932 ;
  assign n37934 = ~n691 & n26277 ;
  assign n37935 = n37934 ^ n4867 ^ 1'b0 ;
  assign n37936 = n7647 & n37935 ;
  assign n37937 = n20262 & n28946 ;
  assign n37938 = n37936 & n37937 ;
  assign n37939 = n37379 ^ n12522 ^ 1'b0 ;
  assign n37940 = n9079 & ~n37939 ;
  assign n37941 = ( ~n1813 & n29637 ) | ( ~n1813 & n33062 ) | ( n29637 & n33062 ) ;
  assign n37942 = n33347 ^ n23635 ^ n22566 ;
  assign n37943 = n37942 ^ n7463 ^ 1'b0 ;
  assign n37944 = ( n5326 & n24215 ) | ( n5326 & n33788 ) | ( n24215 & n33788 ) ;
  assign n37945 = n24226 ^ n3010 ^ 1'b0 ;
  assign n37946 = n37944 | n37945 ;
  assign n37947 = n13800 ^ n2385 ^ 1'b0 ;
  assign n37948 = n13349 ^ n11072 ^ 1'b0 ;
  assign n37949 = n4135 & ~n37948 ;
  assign n37950 = n23830 & n37949 ;
  assign n37951 = n8778 | n24131 ;
  assign n37952 = n29228 | n37951 ;
  assign n37953 = n8994 ^ n2112 ^ 1'b0 ;
  assign n37954 = ~n26223 & n37953 ;
  assign n37955 = ~n9817 & n37954 ;
  assign n37956 = n29075 & n37955 ;
  assign n37957 = n9393 ^ n525 ^ 1'b0 ;
  assign n37958 = n4542 & n13291 ;
  assign n37959 = n21306 ^ n7596 ^ 1'b0 ;
  assign n37960 = n8352 | n24653 ;
  assign n37961 = n37959 | n37960 ;
  assign n37962 = ~n2693 & n3205 ;
  assign n37963 = n9578 & ~n9680 ;
  assign n37964 = n16524 & ~n37963 ;
  assign n37965 = n10436 & n37964 ;
  assign n37966 = n3520 | n6518 ;
  assign n37967 = n17858 | n37966 ;
  assign n37968 = n8568 | n37967 ;
  assign n37969 = n15154 | n16560 ;
  assign n37970 = n35202 | n37969 ;
  assign n37971 = ~n3265 & n12733 ;
  assign n37972 = n37971 ^ n24678 ^ 1'b0 ;
  assign n37973 = ~n20221 & n37972 ;
  assign n37974 = n37973 ^ n2286 ^ 1'b0 ;
  assign n37975 = ~n37970 & n37974 ;
  assign n37976 = n5292 & ~n10767 ;
  assign n37977 = n32306 & n37976 ;
  assign n37978 = n920 & ~n18190 ;
  assign n37979 = n7040 | n23284 ;
  assign n37980 = n37979 ^ n12297 ^ 1'b0 ;
  assign n37981 = ~n2889 & n37980 ;
  assign n37982 = n37981 ^ n36922 ^ 1'b0 ;
  assign n37983 = n1605 & ~n22601 ;
  assign n37984 = n7086 & ~n13487 ;
  assign n37985 = n37984 ^ n5384 ^ 1'b0 ;
  assign n37986 = n12268 & ~n31793 ;
  assign n37987 = n20788 ^ n14821 ^ 1'b0 ;
  assign n37988 = n37986 & n37987 ;
  assign n37989 = n11870 ^ n2053 ^ 1'b0 ;
  assign n37990 = n10306 | n37989 ;
  assign n37991 = n37990 ^ n20047 ^ 1'b0 ;
  assign n37992 = n22117 ^ n9436 ^ n2372 ;
  assign n37993 = n2859 & ~n24399 ;
  assign n37994 = n37993 ^ n33688 ^ 1'b0 ;
  assign n37995 = ~n34692 & n37994 ;
  assign n37996 = n37995 ^ n9017 ^ 1'b0 ;
  assign n37997 = n33023 & ~n37996 ;
  assign n37998 = n16204 & ~n17733 ;
  assign n37999 = n12188 & n37998 ;
  assign n38000 = n5714 & n10578 ;
  assign n38001 = n25004 ^ n15725 ^ 1'b0 ;
  assign n38002 = n38000 & n38001 ;
  assign n38003 = n38002 ^ n19623 ^ 1'b0 ;
  assign n38004 = n4263 | n6524 ;
  assign n38006 = n6005 & ~n9124 ;
  assign n38007 = ~n12595 & n38006 ;
  assign n38008 = n5269 | n38007 ;
  assign n38009 = n13127 & ~n38008 ;
  assign n38005 = n11369 | n28901 ;
  assign n38010 = n38009 ^ n38005 ^ 1'b0 ;
  assign n38011 = n3191 & ~n25399 ;
  assign n38012 = n38011 ^ n17759 ^ 1'b0 ;
  assign n38013 = n16928 ^ n11647 ^ 1'b0 ;
  assign n38014 = n18129 ^ n6415 ^ 1'b0 ;
  assign n38015 = n16185 & n24247 ;
  assign n38016 = ( ~n4649 & n9428 ) | ( ~n4649 & n38015 ) | ( n9428 & n38015 ) ;
  assign n38017 = n37249 & n38016 ;
  assign n38018 = n5622 ^ n3223 ^ 1'b0 ;
  assign n38019 = x3 & n38018 ;
  assign n38020 = n22297 ^ n2951 ^ 1'b0 ;
  assign n38021 = n16098 & n38020 ;
  assign n38022 = n38021 ^ n12971 ^ 1'b0 ;
  assign n38023 = n723 & n14322 ;
  assign n38024 = n16969 ^ n8862 ^ 1'b0 ;
  assign n38025 = n38023 & n38024 ;
  assign n38026 = n38025 ^ n25953 ^ 1'b0 ;
  assign n38027 = n2404 & n26835 ;
  assign n38028 = ~n1516 & n3386 ;
  assign n38029 = n38028 ^ n5291 ^ n4957 ;
  assign n38030 = ~n367 & n4059 ;
  assign n38031 = n9674 & n38030 ;
  assign n38032 = n2247 & ~n30719 ;
  assign n38033 = n38032 ^ n28793 ^ 1'b0 ;
  assign n38034 = n24844 ^ n3111 ^ 1'b0 ;
  assign n38035 = n19680 & ~n21798 ;
  assign n38036 = n38035 ^ n23662 ^ 1'b0 ;
  assign n38037 = n20172 ^ n19985 ^ 1'b0 ;
  assign n38038 = n31495 & ~n38037 ;
  assign n38039 = ~n1736 & n29168 ;
  assign n38040 = n37014 | n38039 ;
  assign n38041 = n3839 | n9383 ;
  assign n38042 = n957 | n38041 ;
  assign n38043 = n755 | n3407 ;
  assign n38044 = n19488 | n38043 ;
  assign n38045 = n11769 ^ n2053 ^ 1'b0 ;
  assign n38046 = n15124 ^ n4574 ^ 1'b0 ;
  assign n38047 = n19716 ^ n13472 ^ 1'b0 ;
  assign n38048 = n38047 ^ n3049 ^ 1'b0 ;
  assign n38049 = n19082 & n25377 ;
  assign n38050 = n6923 & n26400 ;
  assign n38051 = n38050 ^ n24921 ^ 1'b0 ;
  assign n38052 = ~n18493 & n38051 ;
  assign n38053 = ~n25004 & n38052 ;
  assign n38054 = n26422 ^ n992 ^ 1'b0 ;
  assign n38055 = n15510 | n38054 ;
  assign n38056 = n4711 & ~n38055 ;
  assign n38057 = n38056 ^ n6545 ^ 1'b0 ;
  assign n38058 = n31933 | n33240 ;
  assign n38059 = n27737 & ~n38058 ;
  assign n38060 = n5657 | n6705 ;
  assign n38061 = n37352 ^ n27906 ^ 1'b0 ;
  assign n38062 = n3850 | n14845 ;
  assign n38063 = ~n3899 & n14825 ;
  assign n38064 = n22478 & ~n31006 ;
  assign n38065 = n38064 ^ n4824 ^ 1'b0 ;
  assign n38066 = n19240 ^ n14273 ^ 1'b0 ;
  assign n38067 = n4859 & ~n38066 ;
  assign n38068 = n23703 ^ n20162 ^ 1'b0 ;
  assign n38069 = n38068 ^ n501 ^ 1'b0 ;
  assign n38070 = ~n6857 & n38069 ;
  assign n38071 = ~n3475 & n5177 ;
  assign n38072 = n3475 & n38071 ;
  assign n38073 = n17426 ^ n4874 ^ 1'b0 ;
  assign n38074 = n38072 | n38073 ;
  assign n38075 = n850 & n38074 ;
  assign n38076 = n6682 & ~n13466 ;
  assign n38077 = ~n13741 & n38076 ;
  assign n38078 = n17594 | n38077 ;
  assign n38079 = n38078 ^ n25863 ^ n22053 ;
  assign n38080 = n6406 | n21871 ;
  assign n38081 = n15014 & ~n38080 ;
  assign n38082 = n22471 ^ n14276 ^ 1'b0 ;
  assign n38083 = n11303 & n38082 ;
  assign n38084 = n4911 & n26244 ;
  assign n38085 = n38084 ^ n949 ^ 1'b0 ;
  assign n38086 = n35350 | n38085 ;
  assign n38087 = ~n699 & n17494 ;
  assign n38088 = ~n4919 & n38087 ;
  assign n38089 = n5895 | n20856 ;
  assign n38090 = n38089 ^ n3242 ^ 1'b0 ;
  assign n38091 = n22994 ^ n12700 ^ 1'b0 ;
  assign n38092 = n38090 | n38091 ;
  assign n38093 = n38092 ^ n8945 ^ 1'b0 ;
  assign n38094 = n28354 & ~n38093 ;
  assign n38095 = n20893 | n25389 ;
  assign n38096 = n19248 & n36119 ;
  assign n38097 = n1712 & n38096 ;
  assign n38098 = n3166 & n23442 ;
  assign n38099 = n5862 & n38098 ;
  assign n38100 = n38097 & ~n38099 ;
  assign n38101 = ~n7896 & n11861 ;
  assign n38102 = ~n4535 & n38101 ;
  assign n38103 = n13032 & ~n38102 ;
  assign n38104 = n38103 ^ n36027 ^ 1'b0 ;
  assign n38105 = n830 | n1279 ;
  assign n38106 = n11891 & ~n38105 ;
  assign n38107 = n27442 ^ n267 ^ 1'b0 ;
  assign n38108 = ~n24437 & n25037 ;
  assign n38109 = n8771 & n15285 ;
  assign n38110 = n38109 ^ n21609 ^ 1'b0 ;
  assign n38112 = n8912 ^ n7226 ^ 1'b0 ;
  assign n38113 = n11007 & ~n38112 ;
  assign n38111 = n595 & ~n6378 ;
  assign n38114 = n38113 ^ n38111 ^ 1'b0 ;
  assign n38116 = n9251 | n34342 ;
  assign n38117 = n38116 ^ n32993 ^ 1'b0 ;
  assign n38115 = n9095 & ~n25674 ;
  assign n38118 = n38117 ^ n38115 ^ 1'b0 ;
  assign n38119 = n25998 ^ n7722 ^ 1'b0 ;
  assign n38120 = x199 & n17312 ;
  assign n38121 = n27449 | n38120 ;
  assign n38122 = n38121 ^ n7212 ^ n6781 ;
  assign n38123 = n8889 & ~n12335 ;
  assign n38124 = n13720 | n21509 ;
  assign n38125 = ( n6253 & n38123 ) | ( n6253 & n38124 ) | ( n38123 & n38124 ) ;
  assign n38126 = n20703 ^ n13381 ^ 1'b0 ;
  assign n38127 = n10064 & n38126 ;
  assign n38128 = n3937 ^ n2314 ^ n1441 ;
  assign n38129 = ~n927 & n38128 ;
  assign n38130 = ~n2761 & n38129 ;
  assign n38131 = n26816 | n38130 ;
  assign n38132 = n16169 & ~n38131 ;
  assign n38133 = n19336 ^ n6490 ^ 1'b0 ;
  assign n38134 = ~n22217 & n38133 ;
  assign n38135 = n36858 & n38134 ;
  assign n38136 = n9701 | n26833 ;
  assign n38137 = ~n5987 & n25898 ;
  assign n38138 = n38137 ^ n16545 ^ 1'b0 ;
  assign n38139 = ( n9200 & n29061 ) | ( n9200 & n29551 ) | ( n29061 & n29551 ) ;
  assign n38140 = n937 & n31101 ;
  assign n38141 = n1570 | n30147 ;
  assign n38142 = n943 & n4691 ;
  assign n38143 = n17413 & n38142 ;
  assign n38144 = n31297 ^ n18479 ^ 1'b0 ;
  assign n38145 = n5404 | n20716 ;
  assign n38146 = n38145 ^ n29696 ^ 1'b0 ;
  assign n38147 = n19185 ^ n705 ^ 1'b0 ;
  assign n38148 = n17934 & ~n38147 ;
  assign n38152 = n9686 & n25539 ;
  assign n38149 = n31382 ^ n668 ^ 1'b0 ;
  assign n38150 = n2306 & n38149 ;
  assign n38151 = n38150 ^ n18273 ^ 1'b0 ;
  assign n38153 = n38152 ^ n38151 ^ 1'b0 ;
  assign n38154 = n2911 & ~n11412 ;
  assign n38155 = ~n420 & n5448 ;
  assign n38156 = n38155 ^ x228 ^ 1'b0 ;
  assign n38157 = n38156 ^ n9109 ^ 1'b0 ;
  assign n38158 = ~n2950 & n38157 ;
  assign n38159 = n35222 & n38158 ;
  assign n38160 = n33732 ^ n9747 ^ 1'b0 ;
  assign n38161 = n28377 | n38160 ;
  assign n38162 = n27030 ^ n13960 ^ 1'b0 ;
  assign n38163 = n25685 & ~n38162 ;
  assign n38164 = x149 & ~n6529 ;
  assign n38165 = n9928 & n38164 ;
  assign n38166 = n19210 ^ n9248 ^ 1'b0 ;
  assign n38167 = n8424 & ~n9495 ;
  assign n38168 = n24683 & n38167 ;
  assign n38169 = n32395 & n38168 ;
  assign n38173 = n8381 ^ n2311 ^ 1'b0 ;
  assign n38170 = n32916 ^ n31015 ^ 1'b0 ;
  assign n38171 = n1750 | n38170 ;
  assign n38172 = n25659 | n38171 ;
  assign n38174 = n38173 ^ n38172 ^ 1'b0 ;
  assign n38175 = n10937 & n15937 ;
  assign n38176 = n10237 & n38175 ;
  assign n38177 = n38176 ^ n17662 ^ n5012 ;
  assign n38178 = n18595 ^ n5398 ^ 1'b0 ;
  assign n38179 = n8609 ^ n4085 ^ 1'b0 ;
  assign n38180 = n12696 & ~n34087 ;
  assign n38181 = n38180 ^ n9981 ^ 1'b0 ;
  assign n38182 = n6644 & ~n34765 ;
  assign n38185 = n4742 & n7276 ;
  assign n38183 = n7672 | n24682 ;
  assign n38184 = n38183 ^ n3874 ^ 1'b0 ;
  assign n38186 = n38185 ^ n38184 ^ 1'b0 ;
  assign n38187 = n14883 & ~n18248 ;
  assign n38188 = ~n27048 & n38187 ;
  assign n38189 = n13478 ^ x44 ^ 1'b0 ;
  assign n38190 = n5280 & ~n29182 ;
  assign n38191 = n18067 & n30611 ;
  assign n38192 = ~n6618 & n15636 ;
  assign n38193 = n38192 ^ n15711 ^ 1'b0 ;
  assign n38194 = n911 & n4241 ;
  assign n38195 = ~n338 & n38194 ;
  assign n38196 = n38195 ^ n22984 ^ 1'b0 ;
  assign n38197 = n26035 ^ n25287 ^ 1'b0 ;
  assign n38198 = n36270 ^ n4714 ^ 1'b0 ;
  assign n38199 = n3052 & n6282 ;
  assign n38200 = ~n6322 & n38199 ;
  assign n38201 = n38200 ^ n36135 ^ 1'b0 ;
  assign n38202 = n3214 & n38201 ;
  assign n38203 = n15452 & n27472 ;
  assign n38204 = n10377 | n38203 ;
  assign n38205 = n27971 | n38204 ;
  assign n38206 = n38205 ^ n38061 ^ 1'b0 ;
  assign n38207 = n9974 & n38206 ;
  assign n38208 = n22527 ^ n11891 ^ 1'b0 ;
  assign n38209 = n26803 & n38208 ;
  assign n38210 = n9006 ^ n5243 ^ 1'b0 ;
  assign n38211 = n38209 & n38210 ;
  assign n38212 = ( ~n8671 & n18356 ) | ( ~n8671 & n38211 ) | ( n18356 & n38211 ) ;
  assign n38213 = n18966 & n24632 ;
  assign n38217 = n385 & n1371 ;
  assign n38218 = ~n1371 & n38217 ;
  assign n38219 = x43 & ~n765 ;
  assign n38220 = n765 & n38219 ;
  assign n38221 = n38218 | n38220 ;
  assign n38222 = n38218 & ~n38221 ;
  assign n38214 = n1707 | n2394 ;
  assign n38215 = n2394 & ~n38214 ;
  assign n38216 = n30900 | n38215 ;
  assign n38223 = n38222 ^ n38216 ^ 1'b0 ;
  assign n38224 = n38223 ^ n19399 ^ 1'b0 ;
  assign n38225 = n10071 | n38224 ;
  assign n38226 = n6978 & ~n31782 ;
  assign n38227 = n38226 ^ n20442 ^ 1'b0 ;
  assign n38228 = n4470 & n36291 ;
  assign n38229 = ~n33734 & n38228 ;
  assign n38230 = n20977 ^ n20527 ^ n11879 ;
  assign n38231 = ~n2919 & n4421 ;
  assign n38232 = ~n10250 & n23518 ;
  assign n38233 = n6765 ^ n1249 ^ 1'b0 ;
  assign n38234 = n1249 & ~n5987 ;
  assign n38235 = ~n15945 & n38234 ;
  assign n38236 = n15109 & ~n38235 ;
  assign n38237 = n5913 & ~n8847 ;
  assign n38238 = n15680 & ~n28265 ;
  assign n38239 = ~x139 & n38238 ;
  assign n38240 = n28443 & n38239 ;
  assign n38241 = n38240 ^ n17250 ^ n7914 ;
  assign n38242 = ( n1051 & ~n3900 ) | ( n1051 & n38241 ) | ( ~n3900 & n38241 ) ;
  assign n38243 = n17759 ^ n15574 ^ 1'b0 ;
  assign n38244 = n33734 ^ n30240 ^ n7664 ;
  assign n38245 = ~n7742 & n12889 ;
  assign n38246 = n8839 ^ n6912 ^ 1'b0 ;
  assign n38247 = ~n11433 & n38246 ;
  assign n38248 = ~n13346 & n17410 ;
  assign n38249 = n16725 | n38248 ;
  assign n38250 = n9670 & n22306 ;
  assign n38251 = n31874 | n31935 ;
  assign n38252 = n11348 | n38251 ;
  assign n38253 = n7242 | n26923 ;
  assign n38254 = n2182 & n22644 ;
  assign n38255 = n38254 ^ n5613 ^ 1'b0 ;
  assign n38256 = n9525 & n36472 ;
  assign n38257 = n38256 ^ n5197 ^ 1'b0 ;
  assign n38258 = n15228 & n36992 ;
  assign n38259 = n2414 & ~n11853 ;
  assign n38260 = n2067 & ~n13349 ;
  assign n38261 = n38259 & n38260 ;
  assign n38262 = n7817 | n11766 ;
  assign n38263 = ( n28842 & n38261 ) | ( n28842 & ~n38262 ) | ( n38261 & ~n38262 ) ;
  assign n38264 = ( ~n860 & n21965 ) | ( ~n860 & n25137 ) | ( n21965 & n25137 ) ;
  assign n38265 = n38264 ^ n26279 ^ 1'b0 ;
  assign n38266 = ~n38263 & n38265 ;
  assign n38267 = ( ~n2040 & n26726 ) | ( ~n2040 & n31524 ) | ( n26726 & n31524 ) ;
  assign n38268 = n4943 & ~n22961 ;
  assign n38269 = n31939 ^ n6057 ^ n3677 ;
  assign n38270 = n34455 & ~n38269 ;
  assign n38271 = n13680 | n38270 ;
  assign n38272 = n9296 ^ n5696 ^ 1'b0 ;
  assign n38273 = n38272 ^ n7601 ^ 1'b0 ;
  assign n38274 = n11911 | n12297 ;
  assign n38275 = ~n37221 & n38274 ;
  assign n38276 = ~n6516 & n37925 ;
  assign n38277 = n38276 ^ n4867 ^ 1'b0 ;
  assign n38278 = ~n2644 & n38277 ;
  assign n38279 = n4552 & n38278 ;
  assign n38280 = n35137 ^ n29115 ^ 1'b0 ;
  assign n38281 = n12792 & n15981 ;
  assign n38282 = n3458 & ~n11655 ;
  assign n38283 = n38281 & n38282 ;
  assign n38284 = ~n11143 & n14984 ;
  assign n38285 = n38284 ^ n3855 ^ 1'b0 ;
  assign n38286 = n23280 & ~n36941 ;
  assign n38287 = n37043 ^ n26342 ^ n12593 ;
  assign n38288 = n38287 ^ n23725 ^ 1'b0 ;
  assign n38289 = n38286 | n38288 ;
  assign n38290 = n22346 & n28035 ;
  assign n38291 = ~n6112 & n38290 ;
  assign n38292 = n15937 & n38291 ;
  assign n38293 = n22326 & ~n38292 ;
  assign n38294 = n33106 & n38293 ;
  assign n38295 = n10773 ^ n2441 ^ 1'b0 ;
  assign n38296 = n36881 & ~n38295 ;
  assign n38297 = n9696 ^ n3042 ^ n331 ;
  assign n38298 = n22959 | n30774 ;
  assign n38299 = n38297 | n38298 ;
  assign n38300 = n36413 & n37025 ;
  assign n38301 = n4500 | n7836 ;
  assign n38302 = n3423 | n38301 ;
  assign n38303 = n16257 ^ n10527 ^ 1'b0 ;
  assign n38305 = n6624 ^ n6008 ^ 1'b0 ;
  assign n38306 = n416 | n38305 ;
  assign n38304 = n2464 | n15381 ;
  assign n38307 = n38306 ^ n38304 ^ 1'b0 ;
  assign n38308 = n36508 ^ n25730 ^ 1'b0 ;
  assign n38309 = n2730 | n24695 ;
  assign n38310 = n21249 ^ n14658 ^ 1'b0 ;
  assign n38311 = n12306 & ~n33226 ;
  assign n38312 = n22800 ^ n8931 ^ n1439 ;
  assign n38313 = n38312 ^ n1093 ^ 1'b0 ;
  assign n38314 = n19919 ^ n19514 ^ 1'b0 ;
  assign n38315 = n38313 & ~n38314 ;
  assign n38316 = n11995 ^ n9198 ^ 1'b0 ;
  assign n38317 = ~n1884 & n38316 ;
  assign n38318 = n21371 ^ n14449 ^ 1'b0 ;
  assign n38319 = n20534 | n38318 ;
  assign n38320 = ~n10516 & n17426 ;
  assign n38321 = n5798 & n38320 ;
  assign n38322 = n15404 ^ n1259 ^ 1'b0 ;
  assign n38323 = ( n2785 & n12754 ) | ( n2785 & n15091 ) | ( n12754 & n15091 ) ;
  assign n38324 = ( n1805 & n6524 ) | ( n1805 & n27926 ) | ( n6524 & n27926 ) ;
  assign n38325 = n15131 ^ n14622 ^ 1'b0 ;
  assign n38326 = n3114 | n4555 ;
  assign n38327 = n38326 ^ n29068 ^ 1'b0 ;
  assign n38328 = n930 & ~n8536 ;
  assign n38329 = n8114 & n38328 ;
  assign n38330 = n38329 ^ n8163 ^ 1'b0 ;
  assign n38331 = ~n3490 & n5213 ;
  assign n38332 = n38331 ^ n2964 ^ 1'b0 ;
  assign n38335 = n1116 | n2105 ;
  assign n38336 = n38335 ^ n2855 ^ 1'b0 ;
  assign n38337 = ( ~n3760 & n14265 ) | ( ~n3760 & n38336 ) | ( n14265 & n38336 ) ;
  assign n38333 = n5748 ^ n1803 ^ 1'b0 ;
  assign n38334 = n38333 ^ n22536 ^ 1'b0 ;
  assign n38338 = n38337 ^ n38334 ^ n5544 ;
  assign n38339 = n3022 & ~n16627 ;
  assign n38340 = ( n5838 & n12477 ) | ( n5838 & n13419 ) | ( n12477 & n13419 ) ;
  assign n38341 = n34801 ^ n6698 ^ 1'b0 ;
  assign n38342 = n8455 | n34828 ;
  assign n38343 = n9162 ^ n6406 ^ 1'b0 ;
  assign n38344 = n25103 & n38343 ;
  assign n38345 = n38342 | n38344 ;
  assign n38346 = x207 | n35252 ;
  assign n38347 = ( ~n14265 & n21269 ) | ( ~n14265 & n38346 ) | ( n21269 & n38346 ) ;
  assign n38348 = n8633 ^ n4543 ^ 1'b0 ;
  assign n38349 = n19379 ^ n11237 ^ 1'b0 ;
  assign n38350 = ~n38348 & n38349 ;
  assign n38351 = n32520 ^ n27381 ^ 1'b0 ;
  assign n38352 = n4986 & ~n38351 ;
  assign n38353 = n5118 & ~n38352 ;
  assign n38354 = ( ~n4824 & n11557 ) | ( ~n4824 & n19473 ) | ( n11557 & n19473 ) ;
  assign n38355 = n34939 ^ n23424 ^ n1330 ;
  assign n38356 = n7562 | n18649 ;
  assign n38357 = n28567 | n38356 ;
  assign n38358 = ~n5619 & n27645 ;
  assign n38359 = n38358 ^ n10270 ^ 1'b0 ;
  assign n38360 = n36402 ^ n32727 ^ n1367 ;
  assign n38361 = n21489 ^ n15434 ^ n3877 ;
  assign n38362 = n35737 ^ n13011 ^ n4856 ;
  assign n38363 = n37240 & n38362 ;
  assign n38364 = n38363 ^ n18443 ^ 1'b0 ;
  assign n38365 = ~n5105 & n6695 ;
  assign n38366 = ~n5374 & n12885 ;
  assign n38367 = ~n17417 & n38366 ;
  assign n38368 = n23553 ^ n8956 ^ 1'b0 ;
  assign n38369 = ~n38367 & n38368 ;
  assign n38370 = n2611 & ~n2810 ;
  assign n38371 = n6066 & ~n8139 ;
  assign n38372 = n38371 ^ n20534 ^ 1'b0 ;
  assign n38373 = n36524 ^ n18936 ^ 1'b0 ;
  assign n38374 = n13768 ^ n4614 ^ 1'b0 ;
  assign n38375 = n11379 ^ n4666 ^ 1'b0 ;
  assign n38376 = n1835 | n13370 ;
  assign n38377 = n12124 ^ n7407 ^ 1'b0 ;
  assign n38378 = n36021 ^ n3294 ^ 1'b0 ;
  assign n38379 = n7116 & ~n9307 ;
  assign n38380 = n10311 ^ n5664 ^ 1'b0 ;
  assign n38381 = n13102 & n24553 ;
  assign n38382 = ~n24092 & n38381 ;
  assign n38383 = n3073 & n27056 ;
  assign n38384 = n5509 & n38383 ;
  assign n38385 = n38117 ^ n3887 ^ 1'b0 ;
  assign n38386 = n31591 | n38385 ;
  assign n38387 = n11532 ^ n7431 ^ 1'b0 ;
  assign n38388 = n18852 | n38387 ;
  assign n38389 = n37214 ^ n3797 ^ 1'b0 ;
  assign n38390 = ~n23339 & n36279 ;
  assign n38391 = n4852 & n37920 ;
  assign n38392 = ( n9264 & n27010 ) | ( n9264 & n38391 ) | ( n27010 & n38391 ) ;
  assign n38393 = n38392 ^ n5091 ^ 1'b0 ;
  assign n38395 = n17288 ^ n7738 ^ 1'b0 ;
  assign n38396 = n28866 | n38395 ;
  assign n38397 = n38396 ^ n29044 ^ 1'b0 ;
  assign n38394 = ~n15573 & n35027 ;
  assign n38398 = n38397 ^ n38394 ^ 1'b0 ;
  assign n38399 = n22537 ^ n12616 ^ 1'b0 ;
  assign n38400 = ( ~n4065 & n8912 ) | ( ~n4065 & n38399 ) | ( n8912 & n38399 ) ;
  assign n38401 = n26412 ^ n3449 ^ 1'b0 ;
  assign n38402 = n13000 & ~n38401 ;
  assign n38403 = n5619 & n34004 ;
  assign n38404 = n38403 ^ n35853 ^ n31677 ;
  assign n38405 = ~n5637 & n38404 ;
  assign n38406 = n6781 ^ n6261 ^ 1'b0 ;
  assign n38407 = n3177 | n38406 ;
  assign n38408 = ( n26744 & n28058 ) | ( n26744 & ~n38407 ) | ( n28058 & ~n38407 ) ;
  assign n38409 = n33252 & ~n38408 ;
  assign n38410 = n38409 ^ n7128 ^ 1'b0 ;
  assign n38411 = ( ~n5704 & n9081 ) | ( ~n5704 & n26339 ) | ( n9081 & n26339 ) ;
  assign n38412 = n38411 ^ n26143 ^ 1'b0 ;
  assign n38413 = n38412 ^ n35873 ^ n10301 ;
  assign n38414 = ~n9742 & n12766 ;
  assign n38415 = ( n840 & ~n10992 ) | ( n840 & n38414 ) | ( ~n10992 & n38414 ) ;
  assign n38416 = ~n2082 & n26198 ;
  assign n38417 = ~n5704 & n14236 ;
  assign n38418 = n26973 ^ n15582 ^ 1'b0 ;
  assign n38419 = n38417 | n38418 ;
  assign n38420 = n38419 ^ n35032 ^ 1'b0 ;
  assign n38421 = n1028 & n38420 ;
  assign n38422 = n9814 & ~n15193 ;
  assign n38423 = n5413 ^ n838 ^ 1'b0 ;
  assign n38424 = n6576 & ~n30758 ;
  assign n38425 = ~n6903 & n7123 ;
  assign n38426 = n35409 ^ n17543 ^ 1'b0 ;
  assign n38427 = n38425 | n38426 ;
  assign n38428 = n6477 & ~n38427 ;
  assign n38429 = n21447 & n28877 ;
  assign n38430 = n38429 ^ n17883 ^ 1'b0 ;
  assign n38431 = n26341 & n38430 ;
  assign n38432 = ~n20834 & n23688 ;
  assign n38433 = n38432 ^ n1754 ^ 1'b0 ;
  assign n38434 = n20716 ^ n16422 ^ 1'b0 ;
  assign n38435 = n25990 & n38434 ;
  assign n38438 = n1371 & ~n1638 ;
  assign n38436 = n6531 & n9773 ;
  assign n38437 = n38436 ^ n6886 ^ 1'b0 ;
  assign n38439 = n38438 ^ n38437 ^ n13894 ;
  assign n38440 = n3179 & ~n11992 ;
  assign n38441 = n20047 ^ n17754 ^ 1'b0 ;
  assign n38442 = n30787 & ~n38441 ;
  assign n38443 = n28371 ^ n17388 ^ 1'b0 ;
  assign n38444 = n4463 | n12335 ;
  assign n38445 = ~n10707 & n38444 ;
  assign n38446 = n13337 & n38445 ;
  assign n38447 = n9291 ^ n2357 ^ 1'b0 ;
  assign n38448 = ~n13037 & n38447 ;
  assign n38449 = n7356 | n19093 ;
  assign n38450 = n26598 ^ n1211 ^ 1'b0 ;
  assign n38451 = n6046 ^ n1534 ^ 1'b0 ;
  assign n38452 = n8440 & n21255 ;
  assign n38453 = ~n9490 & n38452 ;
  assign n38454 = n34739 ^ n24139 ^ 1'b0 ;
  assign n38455 = n4126 & n17825 ;
  assign n38456 = n22341 ^ n6502 ^ 1'b0 ;
  assign n38457 = n23044 | n38456 ;
  assign n38458 = n34465 ^ n31966 ^ 1'b0 ;
  assign n38459 = n12983 ^ n3596 ^ 1'b0 ;
  assign n38460 = x2 & ~n14573 ;
  assign n38461 = ~n17741 & n38460 ;
  assign n38462 = n492 | n16820 ;
  assign n38463 = ~n38461 & n38462 ;
  assign n38464 = n4516 & n31845 ;
  assign n38465 = ~n15884 & n38464 ;
  assign n38468 = n22751 ^ n1057 ^ 1'b0 ;
  assign n38466 = n9782 & ~n23881 ;
  assign n38467 = n38466 ^ n1134 ^ 1'b0 ;
  assign n38469 = n38468 ^ n38467 ^ n809 ;
  assign n38470 = n5232 | n12671 ;
  assign n38471 = n7312 & n19889 ;
  assign n38472 = n38470 & n38471 ;
  assign n38473 = n17012 & ~n22935 ;
  assign n38474 = n9922 & ~n36102 ;
  assign n38475 = n6188 ^ n5867 ^ 1'b0 ;
  assign n38476 = ~n13908 & n29827 ;
  assign n38477 = ( n5970 & n11143 ) | ( n5970 & n38476 ) | ( n11143 & n38476 ) ;
  assign n38478 = n16427 | n30032 ;
  assign n38479 = n2735 & n17858 ;
  assign n38480 = n34741 & n38479 ;
  assign n38481 = n38480 ^ n25623 ^ 1'b0 ;
  assign n38482 = n7674 & ~n33413 ;
  assign n38483 = n38482 ^ n25230 ^ 1'b0 ;
  assign n38484 = n2415 & ~n38483 ;
  assign n38485 = ~n13660 & n18873 ;
  assign n38486 = n13660 & n38485 ;
  assign n38487 = n15489 & ~n27886 ;
  assign n38488 = n38487 ^ n8431 ^ 1'b0 ;
  assign n38489 = n23864 & ~n38488 ;
  assign n38490 = n3468 ^ n1023 ^ 1'b0 ;
  assign n38491 = n12969 ^ n4466 ^ 1'b0 ;
  assign n38492 = n11491 & n38491 ;
  assign n38493 = n15669 & n38492 ;
  assign n38496 = n23618 ^ x124 ^ 1'b0 ;
  assign n38497 = n21895 & ~n38496 ;
  assign n38498 = n928 | n38497 ;
  assign n38494 = n1358 & ~n12197 ;
  assign n38495 = n21416 & ~n38494 ;
  assign n38499 = n38498 ^ n38495 ^ 1'b0 ;
  assign n38500 = n27350 & ~n38499 ;
  assign n38501 = ~n8618 & n10730 ;
  assign n38502 = n38501 ^ n29007 ^ 1'b0 ;
  assign n38503 = n17303 ^ n17077 ^ 1'b0 ;
  assign n38504 = ~n38502 & n38503 ;
  assign n38505 = x54 & ~n4988 ;
  assign n38506 = n10885 | n21626 ;
  assign n38507 = n18978 ^ n8877 ^ 1'b0 ;
  assign n38508 = x194 & ~n38507 ;
  assign n38509 = n7140 & ~n38508 ;
  assign n38510 = n12367 ^ n10878 ^ n3058 ;
  assign n38511 = n38510 ^ n6485 ^ 1'b0 ;
  assign n38512 = n38511 ^ n13474 ^ 1'b0 ;
  assign n38513 = n27103 ^ n18842 ^ 1'b0 ;
  assign n38514 = ~x143 & n38513 ;
  assign n38515 = n30287 ^ n13239 ^ 1'b0 ;
  assign n38516 = n6700 & n8463 ;
  assign n38517 = n279 & n7470 ;
  assign n38518 = ~n7824 & n38517 ;
  assign n38519 = n15019 ^ n2360 ^ 1'b0 ;
  assign n38520 = n38518 | n38519 ;
  assign n38521 = n1456 & ~n25960 ;
  assign n38522 = n38521 ^ n32485 ^ 1'b0 ;
  assign n38523 = n8114 & ~n38203 ;
  assign n38524 = n38523 ^ n1522 ^ 1'b0 ;
  assign n38525 = n22109 ^ n473 ^ 1'b0 ;
  assign n38526 = n9560 & n38525 ;
  assign n38527 = n19055 ^ n2466 ^ 1'b0 ;
  assign n38528 = n5320 | n16066 ;
  assign n38529 = n38528 ^ n3359 ^ 1'b0 ;
  assign n38530 = n4104 | n17983 ;
  assign n38531 = n20529 | n30698 ;
  assign n38532 = n17919 & ~n38531 ;
  assign n38533 = n38530 | n38532 ;
  assign n38534 = ( n530 & n38529 ) | ( n530 & n38533 ) | ( n38529 & n38533 ) ;
  assign n38535 = ~n9504 & n21340 ;
  assign n38536 = n38535 ^ n21999 ^ 1'b0 ;
  assign n38537 = n25860 ^ n11692 ^ n1473 ;
  assign n38538 = n629 & ~n38537 ;
  assign n38539 = n32763 ^ n17799 ^ 1'b0 ;
  assign n38540 = n8096 ^ n2604 ^ 1'b0 ;
  assign n38541 = ~n9630 & n38540 ;
  assign n38542 = ~n7902 & n38541 ;
  assign n38543 = n31365 & n38542 ;
  assign n38544 = ( n10489 & n17815 ) | ( n10489 & ~n25150 ) | ( n17815 & ~n25150 ) ;
  assign n38545 = n24554 & ~n38544 ;
  assign n38546 = ~n30268 & n38545 ;
  assign n38547 = n8133 & ~n38546 ;
  assign n38548 = n27795 & n38547 ;
  assign n38549 = n37535 ^ n34131 ^ n10920 ;
  assign n38550 = n6716 & n11046 ;
  assign n38551 = n38550 ^ n29839 ^ 1'b0 ;
  assign n38552 = n17812 ^ x100 ^ 1'b0 ;
  assign n38553 = n24624 & n34302 ;
  assign n38554 = n38553 ^ n2993 ^ 1'b0 ;
  assign n38555 = n23466 ^ n2047 ^ 1'b0 ;
  assign n38556 = ~n38554 & n38555 ;
  assign n38557 = n6711 | n12952 ;
  assign n38558 = n2890 & ~n38557 ;
  assign n38559 = n3958 & n24506 ;
  assign n38560 = ~n17326 & n38559 ;
  assign n38561 = n35981 ^ n21658 ^ 1'b0 ;
  assign n38562 = ~n20832 & n27826 ;
  assign n38563 = n34553 & n38562 ;
  assign n38564 = n375 & ~n38198 ;
  assign n38565 = n38563 & n38564 ;
  assign n38566 = n7932 & n28592 ;
  assign n38567 = n14578 & n38566 ;
  assign n38568 = ~n15549 & n38567 ;
  assign n38569 = n10350 ^ n8664 ^ 1'b0 ;
  assign n38570 = ~n22032 & n38569 ;
  assign n38573 = n22278 & n22343 ;
  assign n38574 = ~n10529 & n38573 ;
  assign n38571 = n9973 | n21006 ;
  assign n38572 = n36130 | n38571 ;
  assign n38575 = n38574 ^ n38572 ^ 1'b0 ;
  assign n38576 = n12595 & n22201 ;
  assign n38577 = n38576 ^ n10627 ^ 1'b0 ;
  assign n38578 = n2420 & n4626 ;
  assign n38579 = ( n13631 & ~n16110 ) | ( n13631 & n27634 ) | ( ~n16110 & n27634 ) ;
  assign n38580 = n9993 | n28170 ;
  assign n38581 = n38580 ^ n25943 ^ 1'b0 ;
  assign n38582 = n9015 & ~n12854 ;
  assign n38583 = n9468 | n9573 ;
  assign n38584 = n4220 & ~n24877 ;
  assign n38585 = n24877 & n38584 ;
  assign n38586 = n27854 ^ n6516 ^ 1'b0 ;
  assign n38587 = n38585 | n38586 ;
  assign n38588 = ~n10846 & n15985 ;
  assign n38589 = ~n15985 & n38588 ;
  assign n38590 = n8772 | n38589 ;
  assign n38591 = n8772 & ~n38590 ;
  assign n38592 = n38587 | n38591 ;
  assign n38593 = n38587 & ~n38592 ;
  assign n38594 = n2107 & n33038 ;
  assign n38595 = n38594 ^ n18978 ^ 1'b0 ;
  assign n38596 = n7069 & n38595 ;
  assign n38597 = n31046 ^ n14573 ^ 1'b0 ;
  assign n38598 = n1695 | n8498 ;
  assign n38599 = n38598 ^ n12969 ^ 1'b0 ;
  assign n38600 = n38599 ^ n3617 ^ 1'b0 ;
  assign n38601 = n1125 & ~n38600 ;
  assign n38602 = ~n32383 & n35756 ;
  assign n38603 = n7973 & n24029 ;
  assign n38604 = n14497 | n18226 ;
  assign n38605 = n34416 ^ n18297 ^ n7825 ;
  assign n38606 = n6055 & ~n33482 ;
  assign n38607 = n19335 & n38606 ;
  assign n38608 = n15292 | n38607 ;
  assign n38609 = n1936 & ~n13363 ;
  assign n38610 = n310 & ~n3956 ;
  assign n38611 = n35011 ^ n8330 ^ 1'b0 ;
  assign n38612 = n30592 & n38611 ;
  assign n38613 = n11124 ^ n10995 ^ 1'b0 ;
  assign n38614 = n5909 ^ n599 ^ 1'b0 ;
  assign n38615 = n16088 | n24284 ;
  assign n38616 = n7711 | n38615 ;
  assign n38617 = n21029 ^ n8821 ^ 1'b0 ;
  assign n38618 = n38616 & n38617 ;
  assign n38619 = n35111 ^ n24871 ^ 1'b0 ;
  assign n38620 = n38474 ^ n24298 ^ 1'b0 ;
  assign n38621 = ~n20135 & n38620 ;
  assign n38622 = n10754 & ~n20259 ;
  assign n38623 = n13601 ^ n1665 ^ 1'b0 ;
  assign n38624 = n20146 & n34094 ;
  assign n38625 = n20639 | n38624 ;
  assign n38626 = n12251 | n38625 ;
  assign n38627 = n13443 ^ n1566 ^ 1'b0 ;
  assign n38628 = n2378 & ~n38627 ;
  assign n38629 = n38628 ^ n10480 ^ 1'b0 ;
  assign n38630 = ( ~n13596 & n22155 ) | ( ~n13596 & n27474 ) | ( n22155 & n27474 ) ;
  assign n38631 = ( n5513 & n16499 ) | ( n5513 & n38630 ) | ( n16499 & n38630 ) ;
  assign n38633 = n6359 & n6502 ;
  assign n38632 = ~n2615 & n14510 ;
  assign n38634 = n38633 ^ n38632 ^ 1'b0 ;
  assign n38635 = n2099 ^ n1519 ^ 1'b0 ;
  assign n38636 = n26322 | n38635 ;
  assign n38637 = n2103 | n3298 ;
  assign n38638 = n1651 & ~n38637 ;
  assign n38639 = n35886 & ~n38638 ;
  assign n38640 = n16103 ^ x74 ^ 1'b0 ;
  assign n38641 = n33516 & n38640 ;
  assign n38642 = n6255 | n10273 ;
  assign n38646 = n8237 | n9094 ;
  assign n38647 = n38646 ^ n33995 ^ 1'b0 ;
  assign n38648 = n38647 ^ n35095 ^ n21644 ;
  assign n38649 = x101 & n38648 ;
  assign n38643 = n9704 & ~n20611 ;
  assign n38644 = n38643 ^ n16108 ^ 1'b0 ;
  assign n38645 = ( n928 & n14147 ) | ( n928 & ~n38644 ) | ( n14147 & ~n38644 ) ;
  assign n38650 = n38649 ^ n38645 ^ n20413 ;
  assign n38651 = n20473 & n31181 ;
  assign n38652 = n3855 & n7311 ;
  assign n38653 = n38652 ^ n34824 ^ 1'b0 ;
  assign n38654 = n283 | n38653 ;
  assign n38655 = n8520 | n15213 ;
  assign n38656 = n38567 & ~n38655 ;
  assign n38657 = ~n18362 & n21001 ;
  assign n38658 = n32820 ^ n1152 ^ 1'b0 ;
  assign n38659 = ~n12854 & n38658 ;
  assign n38660 = n513 | n5112 ;
  assign n38661 = n705 | n38660 ;
  assign n38662 = n32455 & ~n38661 ;
  assign n38663 = n6057 | n13864 ;
  assign n38664 = n4287 & n23898 ;
  assign n38665 = n4423 & ~n11375 ;
  assign n38666 = n8591 & n38665 ;
  assign n38667 = ( n4927 & n26534 ) | ( n4927 & ~n38666 ) | ( n26534 & ~n38666 ) ;
  assign n38668 = n38667 ^ n6325 ^ 1'b0 ;
  assign n38669 = n31399 ^ n8043 ^ 1'b0 ;
  assign n38670 = ~n14065 & n17898 ;
  assign n38671 = ~n3771 & n34112 ;
  assign n38672 = ~n19680 & n38671 ;
  assign n38673 = n19975 ^ n16777 ^ 1'b0 ;
  assign n38674 = n11485 | n38673 ;
  assign n38675 = n26768 ^ n14471 ^ 1'b0 ;
  assign n38676 = ~n26366 & n38675 ;
  assign n38677 = ~n5347 & n38676 ;
  assign n38678 = n17672 ^ n12044 ^ n10768 ;
  assign n38679 = n1513 ^ n821 ^ 1'b0 ;
  assign n38680 = ~n2701 & n38679 ;
  assign n38681 = ~n10705 & n38680 ;
  assign n38682 = n38681 ^ n25289 ^ n25038 ;
  assign n38683 = n38682 ^ n14947 ^ 1'b0 ;
  assign n38685 = n21287 & n35063 ;
  assign n38684 = n943 & ~n5835 ;
  assign n38686 = n38685 ^ n38684 ^ 1'b0 ;
  assign n38687 = n28612 ^ n1069 ^ 1'b0 ;
  assign n38688 = n19474 & ~n22614 ;
  assign n38689 = ~n5135 & n38688 ;
  assign n38690 = n38689 ^ n589 ^ 1'b0 ;
  assign n38691 = n6902 | n38690 ;
  assign n38692 = n38691 ^ n12845 ^ 1'b0 ;
  assign n38693 = x99 & n1878 ;
  assign n38694 = n19162 & n38693 ;
  assign n38695 = n3530 ^ x74 ^ 1'b0 ;
  assign n38696 = n26206 ^ n25137 ^ 1'b0 ;
  assign n38697 = n38695 | n38696 ;
  assign n38698 = n32106 | n38430 ;
  assign n38699 = n10403 & n23113 ;
  assign n38700 = n20486 | n38699 ;
  assign n38701 = n32620 ^ n21590 ^ n7081 ;
  assign n38702 = n5931 ^ n1276 ^ 1'b0 ;
  assign n38703 = n38702 ^ n35005 ^ 1'b0 ;
  assign n38704 = n17839 & ~n38703 ;
  assign n38705 = n19680 ^ n9703 ^ 1'b0 ;
  assign n38706 = n11749 & n38705 ;
  assign n38707 = n6075 | n38706 ;
  assign n38708 = n5135 & n9958 ;
  assign n38709 = ~n38707 & n38708 ;
  assign n38710 = n17802 & n24191 ;
  assign n38711 = n16124 ^ n671 ^ 1'b0 ;
  assign n38712 = ~n4924 & n38711 ;
  assign n38713 = n38712 ^ n1592 ^ 1'b0 ;
  assign n38714 = ~n1894 & n25623 ;
  assign n38715 = ~n21413 & n38714 ;
  assign n38716 = x116 & n26553 ;
  assign n38717 = n38716 ^ n12517 ^ 1'b0 ;
  assign n38718 = x206 & n27198 ;
  assign n38719 = n38718 ^ n18543 ^ 1'b0 ;
  assign n38720 = n1496 & ~n30244 ;
  assign n38721 = n38720 ^ n8281 ^ 1'b0 ;
  assign n38722 = ( ~n3860 & n16732 ) | ( ~n3860 & n38721 ) | ( n16732 & n38721 ) ;
  assign n38723 = n8690 ^ n4177 ^ 1'b0 ;
  assign n38724 = ~n16810 & n38723 ;
  assign n38725 = n11643 & n38724 ;
  assign n38726 = n4153 & ~n6359 ;
  assign n38727 = n32704 & n38726 ;
  assign n38728 = n6177 & n20384 ;
  assign n38729 = ~n35520 & n38728 ;
  assign n38730 = n9619 ^ n4330 ^ 1'b0 ;
  assign n38731 = n38730 ^ n24814 ^ 1'b0 ;
  assign n38732 = n595 | n6655 ;
  assign n38733 = n38731 | n38732 ;
  assign n38734 = n21754 | n33855 ;
  assign n38735 = ~n14709 & n21804 ;
  assign n38736 = ~n31029 & n38735 ;
  assign n38737 = n38736 ^ n31982 ^ n4269 ;
  assign n38738 = n3894 | n12280 ;
  assign n38739 = n37743 & ~n38738 ;
  assign n38740 = n17949 | n27651 ;
  assign n38741 = n38740 ^ n12074 ^ 1'b0 ;
  assign n38742 = n19198 & n21702 ;
  assign n38743 = n23376 | n38742 ;
  assign n38744 = n10636 ^ n335 ^ 1'b0 ;
  assign n38745 = n38744 ^ n19005 ^ n11175 ;
  assign n38746 = ~n10287 & n29407 ;
  assign n38747 = n38746 ^ n26819 ^ 1'b0 ;
  assign n38748 = n24426 ^ n15207 ^ 1'b0 ;
  assign n38749 = n14247 & ~n27737 ;
  assign n38750 = n3829 & ~n23335 ;
  assign n38751 = ~n1624 & n38750 ;
  assign n38752 = n389 | n38751 ;
  assign n38753 = n38752 ^ n27556 ^ 1'b0 ;
  assign n38754 = n27989 | n37836 ;
  assign n38755 = n38753 | n38754 ;
  assign n38756 = ~n21349 & n30661 ;
  assign n38757 = n3696 | n26136 ;
  assign n38758 = n12300 | n38757 ;
  assign n38759 = n2554 | n8505 ;
  assign n38760 = n20718 ^ n9821 ^ 1'b0 ;
  assign n38761 = n12393 & ~n18548 ;
  assign n38762 = ( n16898 & n28047 ) | ( n16898 & ~n38761 ) | ( n28047 & ~n38761 ) ;
  assign n38763 = n25283 & ~n34681 ;
  assign n38764 = n3279 ^ n3203 ^ 1'b0 ;
  assign n38765 = n38764 ^ n27130 ^ n11331 ;
  assign n38766 = n38765 ^ n23145 ^ n1397 ;
  assign n38767 = n22821 & n38766 ;
  assign n38768 = ( n3804 & ~n24676 ) | ( n3804 & n27146 ) | ( ~n24676 & n27146 ) ;
  assign n38769 = n876 | n28213 ;
  assign n38770 = n38769 ^ n26388 ^ n10268 ;
  assign n38771 = n38770 ^ n14612 ^ 1'b0 ;
  assign n38772 = n13256 | n30270 ;
  assign n38773 = ~n27448 & n38772 ;
  assign n38774 = n38773 ^ n33692 ^ 1'b0 ;
  assign n38775 = n35920 ^ n11033 ^ n7159 ;
  assign n38776 = n29122 & n30048 ;
  assign n38777 = n38776 ^ n7111 ^ 1'b0 ;
  assign n38781 = n6965 | n10041 ;
  assign n38778 = n5454 ^ n1620 ^ 1'b0 ;
  assign n38779 = n9156 & ~n38778 ;
  assign n38780 = ~n7962 & n38779 ;
  assign n38782 = n38781 ^ n38780 ^ 1'b0 ;
  assign n38783 = n15559 | n37093 ;
  assign n38784 = n16984 & ~n38783 ;
  assign n38785 = ~n3223 & n12887 ;
  assign n38786 = n12337 & ~n22658 ;
  assign n38787 = n38371 ^ n3573 ^ 1'b0 ;
  assign n38788 = n7541 | n38787 ;
  assign n38789 = ~n3925 & n9192 ;
  assign n38790 = n34433 & n38789 ;
  assign n38791 = n22700 & ~n23574 ;
  assign n38792 = ~n9094 & n38791 ;
  assign n38793 = ~n20910 & n22798 ;
  assign n38794 = n3684 ^ n2829 ^ 1'b0 ;
  assign n38795 = n2789 & n38794 ;
  assign n38796 = n14755 & n28344 ;
  assign n38797 = n38796 ^ n3300 ^ 1'b0 ;
  assign n38798 = n7934 ^ n6785 ^ 1'b0 ;
  assign n38799 = ~n12765 & n38798 ;
  assign n38800 = n17946 & n38799 ;
  assign n38801 = n38800 ^ n5208 ^ 1'b0 ;
  assign n38802 = n38801 ^ n37335 ^ n20254 ;
  assign n38803 = ( n23683 & n29052 ) | ( n23683 & ~n38802 ) | ( n29052 & ~n38802 ) ;
  assign n38804 = n38803 ^ n17078 ^ n8822 ;
  assign n38805 = n30261 ^ n11063 ^ 1'b0 ;
  assign n38806 = n10630 & n27044 ;
  assign n38807 = n16662 | n23091 ;
  assign n38808 = n38807 ^ n13020 ^ 1'b0 ;
  assign n38810 = n6475 & ~n20799 ;
  assign n38811 = n38810 ^ n27200 ^ 1'b0 ;
  assign n38809 = n436 & n19861 ;
  assign n38812 = n38811 ^ n38809 ^ 1'b0 ;
  assign n38813 = n7806 ^ n5714 ^ 1'b0 ;
  assign n38814 = n4979 & ~n8619 ;
  assign n38815 = ~n38813 & n38814 ;
  assign n38816 = n4553 & ~n38815 ;
  assign n38817 = ~n12486 & n38816 ;
  assign n38818 = n38817 ^ n7651 ^ 1'b0 ;
  assign n38819 = ~n614 & n3154 ;
  assign n38820 = ~n1653 & n38819 ;
  assign n38822 = n2916 ^ n2047 ^ 1'b0 ;
  assign n38821 = n18763 & n30193 ;
  assign n38823 = n38822 ^ n38821 ^ 1'b0 ;
  assign n38824 = n19893 | n23378 ;
  assign n38825 = n38823 | n38824 ;
  assign n38826 = ( n4497 & ~n7964 ) | ( n4497 & n27940 ) | ( ~n7964 & n27940 ) ;
  assign n38827 = n34523 ^ n5305 ^ 1'b0 ;
  assign n38828 = n14567 & n38827 ;
  assign n38829 = n32211 & n38828 ;
  assign n38830 = n35263 | n38829 ;
  assign n38831 = n38826 & ~n38830 ;
  assign n38832 = n18563 ^ n1627 ^ 1'b0 ;
  assign n38833 = n14932 ^ n4864 ^ 1'b0 ;
  assign n38834 = n35332 ^ n26470 ^ 1'b0 ;
  assign n38835 = ~n2687 & n38834 ;
  assign n38836 = ~n13077 & n38835 ;
  assign n38837 = ~n23458 & n38836 ;
  assign n38838 = n1590 | n11274 ;
  assign n38839 = n38838 ^ n27438 ^ 1'b0 ;
  assign n38840 = n21090 ^ n9865 ^ 1'b0 ;
  assign n38841 = n38839 | n38840 ;
  assign n38842 = ~n24239 & n32823 ;
  assign n38844 = ~n23820 & n30756 ;
  assign n38845 = n38844 ^ n3455 ^ 1'b0 ;
  assign n38846 = n2615 & n38845 ;
  assign n38843 = n16062 & ~n34559 ;
  assign n38847 = n38846 ^ n38843 ^ 1'b0 ;
  assign n38848 = n12721 ^ n10443 ^ n794 ;
  assign n38849 = n3848 & n26836 ;
  assign n38850 = n2439 | n14447 ;
  assign n38851 = ~n9699 & n38850 ;
  assign n38852 = ~n4288 & n17285 ;
  assign n38853 = n38852 ^ n4730 ^ 1'b0 ;
  assign n38854 = n22530 ^ n20577 ^ n3704 ;
  assign n38855 = n20896 & ~n28948 ;
  assign n38856 = ~n2390 & n13357 ;
  assign n38857 = n5062 ^ n3821 ^ 1'b0 ;
  assign n38858 = n18761 | n38857 ;
  assign n38859 = ( n25938 & ~n27826 ) | ( n25938 & n29169 ) | ( ~n27826 & n29169 ) ;
  assign n38860 = n38858 | n38859 ;
  assign n38861 = n38860 ^ n16071 ^ 1'b0 ;
  assign n38862 = n26824 ^ n16012 ^ 1'b0 ;
  assign n38863 = ~n12856 & n38862 ;
  assign n38864 = n36758 ^ n26647 ^ 1'b0 ;
  assign n38865 = n16006 ^ n14246 ^ n8943 ;
  assign n38869 = n3601 & n20954 ;
  assign n38870 = n12812 & n38869 ;
  assign n38867 = n11572 & ~n18453 ;
  assign n38866 = n6822 & n6851 ;
  assign n38868 = n38867 ^ n38866 ^ 1'b0 ;
  assign n38871 = n38870 ^ n38868 ^ 1'b0 ;
  assign n38872 = n1352 & ~n26828 ;
  assign n38873 = n38872 ^ n20517 ^ 1'b0 ;
  assign n38874 = n22854 ^ n11802 ^ 1'b0 ;
  assign n38875 = ~n4730 & n12275 ;
  assign n38876 = n4180 ^ n1169 ^ 1'b0 ;
  assign n38877 = n9061 & ~n22607 ;
  assign n38878 = ~n13429 & n38877 ;
  assign n38879 = n38878 ^ n11927 ^ 1'b0 ;
  assign n38880 = n11235 & ~n36462 ;
  assign n38881 = ~n20517 & n38880 ;
  assign n38883 = n3123 | n21471 ;
  assign n38884 = n38883 ^ n17484 ^ n16061 ;
  assign n38885 = n3150 ^ n2701 ^ 1'b0 ;
  assign n38886 = n38884 | n38885 ;
  assign n38887 = n26671 | n38886 ;
  assign n38882 = n1001 | n29263 ;
  assign n38888 = n38887 ^ n38882 ^ 1'b0 ;
  assign n38889 = n4296 ^ n780 ^ x5 ;
  assign n38890 = n33917 & n34911 ;
  assign n38891 = n12998 & n38890 ;
  assign n38892 = n10475 | n16744 ;
  assign n38893 = n38892 ^ n27782 ^ n13650 ;
  assign n38894 = n17717 | n23864 ;
  assign n38895 = n9529 & n18454 ;
  assign n38896 = n14088 & ~n30056 ;
  assign n38897 = ~n38895 & n38896 ;
  assign n38898 = ( ~n19317 & n25660 ) | ( ~n19317 & n38897 ) | ( n25660 & n38897 ) ;
  assign n38899 = n7054 ^ n4254 ^ 1'b0 ;
  assign n38900 = n8595 ^ n8188 ^ 1'b0 ;
  assign n38901 = n6060 | n38900 ;
  assign n38902 = n13315 | n27632 ;
  assign n38903 = n34375 & ~n38902 ;
  assign n38904 = n6060 | n9013 ;
  assign n38905 = n38904 ^ n35775 ^ 1'b0 ;
  assign n38906 = n1247 & n38905 ;
  assign n38907 = n4010 & n14174 ;
  assign n38908 = n14906 | n30583 ;
  assign n38909 = n38908 ^ n7496 ^ 1'b0 ;
  assign n38910 = n14159 ^ n13240 ^ 1'b0 ;
  assign n38911 = n5246 & ~n38910 ;
  assign n38912 = n21497 | n34135 ;
  assign n38913 = n12877 ^ n8739 ^ 1'b0 ;
  assign n38914 = n29104 ^ n8241 ^ 1'b0 ;
  assign n38915 = n7071 & ~n38914 ;
  assign n38916 = n21736 ^ n18850 ^ 1'b0 ;
  assign n38917 = n38915 & ~n38916 ;
  assign n38918 = n1392 & n10880 ;
  assign n38919 = n38918 ^ n24586 ^ n8249 ;
  assign n38920 = n38663 ^ n33390 ^ 1'b0 ;
  assign n38921 = n32146 & ~n38920 ;
  assign n38922 = n16364 ^ n1638 ^ 1'b0 ;
  assign n38923 = n38922 ^ n5203 ^ 1'b0 ;
  assign n38924 = n7279 & ~n14331 ;
  assign n38925 = n27122 ^ n17556 ^ 1'b0 ;
  assign n38926 = n15661 & n38925 ;
  assign n38927 = n13381 & n38926 ;
  assign n38928 = n4343 & n8081 ;
  assign n38929 = n38928 ^ n18546 ^ 1'b0 ;
  assign n38930 = n16257 & ~n28423 ;
  assign n38931 = n38930 ^ n21185 ^ 1'b0 ;
  assign n38932 = n2728 & ~n13504 ;
  assign n38933 = n38931 & n38932 ;
  assign n38934 = n38933 ^ x108 ^ 1'b0 ;
  assign n38935 = n37014 ^ n15637 ^ 1'b0 ;
  assign n38939 = n10352 | n27712 ;
  assign n38940 = n38939 ^ n2250 ^ 1'b0 ;
  assign n38936 = n2567 | n11659 ;
  assign n38937 = n38936 ^ n11677 ^ 1'b0 ;
  assign n38938 = n2245 & n38937 ;
  assign n38941 = n38940 ^ n38938 ^ 1'b0 ;
  assign n38942 = n12798 ^ n9004 ^ 1'b0 ;
  assign n38943 = n26112 | n38942 ;
  assign n38944 = n5676 & ~n7306 ;
  assign n38945 = n8594 ^ n4249 ^ 1'b0 ;
  assign n38946 = n38944 | n38945 ;
  assign n38947 = n3271 ^ x38 ^ 1'b0 ;
  assign n38948 = ( n9114 & n15803 ) | ( n9114 & ~n38947 ) | ( n15803 & ~n38947 ) ;
  assign n38949 = n6991 | n8211 ;
  assign n38950 = n38949 ^ n5404 ^ 1'b0 ;
  assign n38951 = ( n15623 & n38948 ) | ( n15623 & n38950 ) | ( n38948 & n38950 ) ;
  assign n38952 = ( n7028 & n16484 ) | ( n7028 & n26929 ) | ( n16484 & n26929 ) ;
  assign n38954 = n4010 ^ n1125 ^ 1'b0 ;
  assign n38955 = n36552 & ~n38954 ;
  assign n38953 = ~n28512 & n29808 ;
  assign n38956 = n38955 ^ n38953 ^ 1'b0 ;
  assign n38957 = ~n2335 & n16396 ;
  assign n38958 = n38957 ^ n2817 ^ 1'b0 ;
  assign n38959 = n6981 & n15961 ;
  assign n38960 = n15845 ^ n915 ^ 1'b0 ;
  assign n38961 = n23133 & ~n38960 ;
  assign n38962 = n8330 ^ n5554 ^ 1'b0 ;
  assign n38963 = n10217 ^ n2532 ^ 1'b0 ;
  assign n38964 = n16298 ^ n5219 ^ 1'b0 ;
  assign n38965 = n26586 | n38964 ;
  assign n38966 = n38965 ^ n22825 ^ 1'b0 ;
  assign n38967 = ~n21654 & n38966 ;
  assign n38968 = n38967 ^ n25965 ^ 1'b0 ;
  assign n38969 = n13163 & n17401 ;
  assign n38970 = n12191 & ~n19373 ;
  assign n38971 = n38970 ^ n16308 ^ 1'b0 ;
  assign n38972 = ~n34145 & n38971 ;
  assign n38973 = n3845 & ~n34092 ;
  assign n38974 = n38973 ^ n35582 ^ 1'b0 ;
  assign n38975 = n38974 ^ n7569 ^ 1'b0 ;
  assign n38976 = n30821 | n38975 ;
  assign n38977 = ~n15343 & n38255 ;
  assign n38978 = n5245 | n26586 ;
  assign n38979 = n38977 | n38978 ;
  assign n38980 = ~n6856 & n26902 ;
  assign n38981 = n38980 ^ n21726 ^ 1'b0 ;
  assign n38982 = n7020 ^ n5720 ^ n1671 ;
  assign n38983 = n17722 ^ n3262 ^ 1'b0 ;
  assign n38984 = n916 & n37449 ;
  assign n38985 = n6393 | n7271 ;
  assign n38986 = n14502 | n19155 ;
  assign n38987 = n27637 & ~n38986 ;
  assign n38988 = n37993 ^ n22601 ^ 1'b0 ;
  assign n38989 = ~n6095 & n38988 ;
  assign n38991 = ~n723 & n37792 ;
  assign n38990 = n8375 | n10852 ;
  assign n38992 = n38991 ^ n38990 ^ 1'b0 ;
  assign n38993 = n17399 | n38992 ;
  assign n38994 = n8747 | n38993 ;
  assign n38995 = ~n1813 & n10064 ;
  assign n38996 = n27239 & ~n27801 ;
  assign n38997 = ~n2868 & n28856 ;
  assign n38998 = n26801 ^ n7065 ^ 1'b0 ;
  assign n38999 = n22146 ^ n6342 ^ 1'b0 ;
  assign n39000 = n24609 ^ n22016 ^ n16166 ;
  assign n39001 = n23199 & n39000 ;
  assign n39002 = n4739 & ~n31384 ;
  assign n39003 = n38644 ^ n35161 ^ 1'b0 ;
  assign n39004 = n9842 | n34071 ;
  assign n39005 = n39004 ^ n15647 ^ n15556 ;
  assign n39006 = n24073 ^ n11608 ^ 1'b0 ;
  assign n39007 = n16618 | n39006 ;
  assign n39008 = n39007 ^ n1244 ^ 1'b0 ;
  assign n39009 = n26961 ^ n16417 ^ 1'b0 ;
  assign n39010 = n25157 & ~n39009 ;
  assign n39011 = n39010 ^ x66 ^ 1'b0 ;
  assign n39013 = n11496 | n34554 ;
  assign n39012 = n32117 | n33251 ;
  assign n39014 = n39013 ^ n39012 ^ 1'b0 ;
  assign n39015 = n38179 ^ n2162 ^ 1'b0 ;
  assign n39016 = n13539 ^ n1123 ^ 1'b0 ;
  assign n39017 = ~n10909 & n39016 ;
  assign n39018 = n39017 ^ n6976 ^ 1'b0 ;
  assign n39019 = n5293 & ~n39018 ;
  assign n39020 = n9006 & n10676 ;
  assign n39021 = n39020 ^ x110 ^ 1'b0 ;
  assign n39022 = ~n21031 & n39021 ;
  assign n39023 = ~n1966 & n39022 ;
  assign n39024 = ~n5994 & n39023 ;
  assign n39025 = n16987 ^ n15236 ^ 1'b0 ;
  assign n39026 = ( n3686 & n7981 ) | ( n3686 & n39025 ) | ( n7981 & n39025 ) ;
  assign n39027 = n36184 ^ n10082 ^ n5190 ;
  assign n39028 = n17010 & ~n21766 ;
  assign n39029 = n39028 ^ n38167 ^ 1'b0 ;
  assign n39030 = ( n18557 & n39027 ) | ( n18557 & ~n39029 ) | ( n39027 & ~n39029 ) ;
  assign n39031 = ~n10251 & n25937 ;
  assign n39032 = n17507 ^ n2655 ^ 1'b0 ;
  assign n39033 = n7382 & ~n39032 ;
  assign n39034 = ( n10664 & ~n12132 ) | ( n10664 & n13691 ) | ( ~n12132 & n13691 ) ;
  assign n39035 = n39034 ^ n31943 ^ 1'b0 ;
  assign n39036 = n5257 & ~n24264 ;
  assign n39037 = n39036 ^ n32829 ^ 1'b0 ;
  assign n39038 = n4393 & ~n31600 ;
  assign n39039 = n6093 ^ n663 ^ 1'b0 ;
  assign n39040 = n5986 & n9490 ;
  assign n39041 = n26997 ^ n8759 ^ 1'b0 ;
  assign n39042 = n39040 & ~n39041 ;
  assign n39043 = x192 & n10886 ;
  assign n39044 = n9804 & ~n39043 ;
  assign n39045 = n39044 ^ n19466 ^ 1'b0 ;
  assign n39046 = n22863 & n39045 ;
  assign n39049 = n729 & n35025 ;
  assign n39047 = n11372 & n21496 ;
  assign n39048 = n39047 ^ n1450 ^ 1'b0 ;
  assign n39050 = n39049 ^ n39048 ^ n38375 ;
  assign n39051 = ~n20501 & n27744 ;
  assign n39052 = n39051 ^ n5462 ^ 1'b0 ;
  assign n39053 = n18288 | n29380 ;
  assign n39054 = n39053 ^ n6783 ^ 1'b0 ;
  assign n39055 = n8233 ^ n7560 ^ 1'b0 ;
  assign n39056 = n30444 ^ n6192 ^ n6146 ;
  assign n39057 = n2296 | n28694 ;
  assign n39058 = ~n39056 & n39057 ;
  assign n39060 = n3642 & ~n27336 ;
  assign n39061 = n39060 ^ n35157 ^ 1'b0 ;
  assign n39059 = n5308 | n5380 ;
  assign n39062 = n39061 ^ n39059 ^ 1'b0 ;
  assign n39063 = n39062 ^ n36411 ^ 1'b0 ;
  assign n39064 = n6385 & ~n21685 ;
  assign n39065 = n2944 & ~n36324 ;
  assign n39066 = n1416 | n28176 ;
  assign n39067 = n39066 ^ n10299 ^ 1'b0 ;
  assign n39068 = n34330 ^ n10111 ^ 1'b0 ;
  assign n39069 = n4845 & ~n9454 ;
  assign n39070 = n16419 & n39069 ;
  assign n39071 = n28905 ^ n25137 ^ 1'b0 ;
  assign n39072 = ~n39070 & n39071 ;
  assign n39073 = n39072 ^ x129 ^ 1'b0 ;
  assign n39074 = n2855 & ~n31384 ;
  assign n39075 = n39073 & n39074 ;
  assign n39076 = n1866 ^ n858 ^ 1'b0 ;
  assign n39077 = n2426 & ~n35708 ;
  assign n39081 = n3690 & ~n20002 ;
  assign n39082 = n39081 ^ n12497 ^ 1'b0 ;
  assign n39083 = n27184 & ~n39082 ;
  assign n39078 = n6471 | n7916 ;
  assign n39079 = n39078 ^ n38007 ^ 1'b0 ;
  assign n39080 = n26760 & n39079 ;
  assign n39084 = n39083 ^ n39080 ^ 1'b0 ;
  assign n39085 = n38642 ^ n12703 ^ 1'b0 ;
  assign n39086 = ~n19395 & n30798 ;
  assign n39087 = ~n7923 & n39086 ;
  assign n39088 = ( ~n9432 & n11523 ) | ( ~n9432 & n30275 ) | ( n11523 & n30275 ) ;
  assign n39089 = ~n39087 & n39088 ;
  assign n39090 = n9635 & ~n22335 ;
  assign n39091 = n39090 ^ n12532 ^ 1'b0 ;
  assign n39092 = n12415 ^ n10959 ^ 1'b0 ;
  assign n39093 = n39091 & n39092 ;
  assign n39095 = n8483 & ~n22933 ;
  assign n39094 = n6075 | n28567 ;
  assign n39096 = n39095 ^ n39094 ^ 1'b0 ;
  assign n39097 = ~n2625 & n21752 ;
  assign n39098 = n39097 ^ n8496 ^ 1'b0 ;
  assign n39100 = n31850 ^ n12281 ^ 1'b0 ;
  assign n39101 = n34191 & n39100 ;
  assign n39099 = ~n1109 & n7291 ;
  assign n39102 = n39101 ^ n39099 ^ 1'b0 ;
  assign n39103 = ( n1510 & n23225 ) | ( n1510 & n30272 ) | ( n23225 & n30272 ) ;
  assign n39104 = n39103 ^ n20071 ^ 1'b0 ;
  assign n39105 = ~n11632 & n28753 ;
  assign n39106 = n39105 ^ n6632 ^ 1'b0 ;
  assign n39107 = n25990 & n31041 ;
  assign n39108 = n39107 ^ n14159 ^ n6138 ;
  assign n39109 = n11339 & n18957 ;
  assign n39110 = n31768 ^ n634 ^ 1'b0 ;
  assign n39111 = ~n39109 & n39110 ;
  assign n39112 = n39111 ^ n9984 ^ 1'b0 ;
  assign n39113 = n4563 | n8827 ;
  assign n39114 = n5831 | n39113 ;
  assign n39115 = n7117 & n13114 ;
  assign n39116 = ~n39114 & n39115 ;
  assign n39117 = n3576 | n15652 ;
  assign n39118 = ~n24418 & n39117 ;
  assign n39119 = ~n14156 & n28067 ;
  assign n39120 = n39119 ^ n19656 ^ 1'b0 ;
  assign n39121 = n5802 | n9674 ;
  assign n39122 = n32115 | n39121 ;
  assign n39123 = n4248 ^ n444 ^ 1'b0 ;
  assign n39124 = n20360 & n39123 ;
  assign n39125 = n27958 ^ n1365 ^ 1'b0 ;
  assign n39126 = n25200 ^ n3479 ^ 1'b0 ;
  assign n39127 = n18181 | n31672 ;
  assign n39128 = n18454 ^ n12771 ^ 1'b0 ;
  assign n39129 = ( n6310 & n25871 ) | ( n6310 & n39128 ) | ( n25871 & n39128 ) ;
  assign n39130 = n13354 ^ n5579 ^ 1'b0 ;
  assign n39131 = n39129 & ~n39130 ;
  assign n39132 = n1864 | n3582 ;
  assign n39133 = n39132 ^ n11127 ^ 1'b0 ;
  assign n39134 = n3780 | n8646 ;
  assign n39135 = n39134 ^ n977 ^ 1'b0 ;
  assign n39136 = n19377 & n24137 ;
  assign n39137 = n31827 & n39136 ;
  assign n39138 = n19783 ^ n7880 ^ 1'b0 ;
  assign n39139 = n35353 ^ n18120 ^ n496 ;
  assign n39140 = n8341 & ~n14801 ;
  assign n39141 = n39140 ^ n4210 ^ 1'b0 ;
  assign n39142 = n11609 | n39141 ;
  assign n39143 = n294 | n27989 ;
  assign n39144 = n16005 | n39143 ;
  assign n39145 = n8024 | n12443 ;
  assign n39146 = n3251 | n5330 ;
  assign n39147 = n39145 | n39146 ;
  assign n39148 = n4296 ^ n3009 ^ 1'b0 ;
  assign n39149 = n39148 ^ n9066 ^ 1'b0 ;
  assign n39150 = n12631 ^ n7132 ^ 1'b0 ;
  assign n39151 = n10637 | n39150 ;
  assign n39152 = n26400 ^ n11665 ^ n6097 ;
  assign n39153 = n18459 ^ n1126 ^ 1'b0 ;
  assign n39154 = n39152 | n39153 ;
  assign n39155 = n18066 & ~n24098 ;
  assign n39156 = n4357 | n34653 ;
  assign n39158 = n8399 & ~n8806 ;
  assign n39157 = n5276 & ~n14010 ;
  assign n39159 = n39158 ^ n39157 ^ 1'b0 ;
  assign n39160 = n1092 & ~n11277 ;
  assign n39161 = n39160 ^ n25900 ^ 1'b0 ;
  assign n39162 = n31865 ^ n23902 ^ 1'b0 ;
  assign n39163 = ~n32991 & n39162 ;
  assign n39164 = ~n4659 & n15716 ;
  assign n39165 = n26037 ^ n4061 ^ 1'b0 ;
  assign n39166 = n4911 & ~n34162 ;
  assign n39167 = n12313 | n32795 ;
  assign n39168 = n39167 ^ n10471 ^ 1'b0 ;
  assign n39169 = n18037 & n39168 ;
  assign n39170 = ~n22334 & n39169 ;
  assign n39171 = n26965 ^ n20546 ^ 1'b0 ;
  assign n39172 = n26636 ^ n20317 ^ 1'b0 ;
  assign n39173 = n20504 | n33507 ;
  assign n39174 = n39173 ^ n31170 ^ 1'b0 ;
  assign n39175 = n8868 & ~n9808 ;
  assign n39176 = ~n7677 & n39175 ;
  assign n39177 = n15972 ^ n15472 ^ 1'b0 ;
  assign n39178 = ~n39176 & n39177 ;
  assign n39179 = n23420 ^ n2891 ^ 1'b0 ;
  assign n39180 = n946 | n39179 ;
  assign n39181 = n39180 ^ n5800 ^ n1633 ;
  assign n39182 = n7393 & n19326 ;
  assign n39183 = ~n18055 & n32940 ;
  assign n39184 = n39183 ^ n16327 ^ 1'b0 ;
  assign n39185 = n23099 & ~n39184 ;
  assign n39186 = n15056 | n36191 ;
  assign n39187 = n15662 | n39186 ;
  assign n39188 = n8041 | n14514 ;
  assign n39190 = n29949 ^ n10606 ^ 1'b0 ;
  assign n39191 = n38009 | n39190 ;
  assign n39192 = n23959 & n26640 ;
  assign n39193 = n39191 & n39192 ;
  assign n39189 = ~n13363 & n28231 ;
  assign n39194 = n39193 ^ n39189 ^ 1'b0 ;
  assign n39195 = n7290 & n14360 ;
  assign n39196 = n9904 & n24901 ;
  assign n39197 = ( ~n4182 & n7145 ) | ( ~n4182 & n39196 ) | ( n7145 & n39196 ) ;
  assign n39198 = n15598 & ~n37868 ;
  assign n39199 = n9241 ^ n2674 ^ 1'b0 ;
  assign n39200 = ( n22601 & n35684 ) | ( n22601 & n39199 ) | ( n35684 & n39199 ) ;
  assign n39201 = n16005 | n39200 ;
  assign n39202 = ~n10780 & n24452 ;
  assign n39203 = ~n3195 & n39202 ;
  assign n39204 = n39203 ^ n1961 ^ 1'b0 ;
  assign n39205 = ~n11891 & n39204 ;
  assign n39206 = n39205 ^ n6567 ^ 1'b0 ;
  assign n39207 = n5350 & ~n35928 ;
  assign n39208 = ~n10429 & n28369 ;
  assign n39209 = ( n5511 & n6606 ) | ( n5511 & ~n39208 ) | ( n6606 & ~n39208 ) ;
  assign n39210 = n13146 & ~n39209 ;
  assign n39211 = n11267 ^ n11193 ^ 1'b0 ;
  assign n39212 = n2841 | n11883 ;
  assign n39213 = n8936 & ~n12998 ;
  assign n39214 = n3393 & n39213 ;
  assign n39215 = n34570 & ~n39214 ;
  assign n39216 = n39215 ^ n15437 ^ 1'b0 ;
  assign n39217 = n16240 ^ n1750 ^ 1'b0 ;
  assign n39218 = n8471 & n39217 ;
  assign n39219 = n12833 & ~n26247 ;
  assign n39220 = n37792 ^ n7814 ^ 1'b0 ;
  assign n39221 = n3806 & ~n39220 ;
  assign n39222 = ~n5242 & n17339 ;
  assign n39223 = n25637 & n39222 ;
  assign n39224 = n5515 & ~n39223 ;
  assign n39225 = ~n39221 & n39224 ;
  assign n39226 = ~n25800 & n27757 ;
  assign n39227 = ~n21822 & n39226 ;
  assign n39228 = n14800 & n39227 ;
  assign n39229 = n4462 ^ n4008 ^ 1'b0 ;
  assign n39230 = ~n367 & n39229 ;
  assign n39231 = n39230 ^ n9848 ^ 1'b0 ;
  assign n39232 = ~n39228 & n39231 ;
  assign n39233 = ( n13668 & n15930 ) | ( n13668 & ~n31724 ) | ( n15930 & ~n31724 ) ;
  assign n39234 = n5292 & n6565 ;
  assign n39235 = n39234 ^ n37733 ^ 1'b0 ;
  assign n39236 = n8243 ^ n1192 ^ 1'b0 ;
  assign n39237 = n19347 & ~n34615 ;
  assign n39238 = ~n22566 & n39237 ;
  assign n39239 = n16690 ^ x182 ^ 1'b0 ;
  assign n39240 = ~n39238 & n39239 ;
  assign n39241 = n13759 | n22141 ;
  assign n39242 = n15282 & n32425 ;
  assign n39243 = n6518 ^ n5099 ^ 1'b0 ;
  assign n39244 = n39243 ^ n10030 ^ n2476 ;
  assign n39245 = n10193 ^ n2319 ^ 1'b0 ;
  assign n39246 = ~n6705 & n39245 ;
  assign n39247 = n39246 ^ n13862 ^ 1'b0 ;
  assign n39248 = n12617 ^ n3893 ^ 1'b0 ;
  assign n39249 = n39247 & ~n39248 ;
  assign n39251 = n23469 | n30497 ;
  assign n39250 = ~n2286 & n30962 ;
  assign n39252 = n39251 ^ n39250 ^ 1'b0 ;
  assign n39253 = n19825 ^ n18686 ^ n15695 ;
  assign n39254 = n39253 ^ n17654 ^ n8552 ;
  assign n39255 = n13680 & ~n36236 ;
  assign n39256 = ~n39254 & n39255 ;
  assign n39257 = ~n5581 & n14988 ;
  assign n39258 = n39257 ^ n23718 ^ 1'b0 ;
  assign n39259 = n9416 ^ n7714 ^ 1'b0 ;
  assign n39260 = n5933 & ~n39259 ;
  assign n39261 = n35405 ^ n14694 ^ 1'b0 ;
  assign n39262 = ~n6551 & n33580 ;
  assign n39263 = n20866 | n37217 ;
  assign n39264 = n26929 ^ n13327 ^ n7407 ;
  assign n39265 = n36485 & ~n39264 ;
  assign n39266 = n39265 ^ n1085 ^ 1'b0 ;
  assign n39267 = n13080 | n27393 ;
  assign n39268 = n12469 & ~n39267 ;
  assign n39269 = n9731 | n39268 ;
  assign n39270 = ~n5879 & n25729 ;
  assign n39271 = n11296 | n20233 ;
  assign n39273 = n6646 & n18354 ;
  assign n39274 = n39273 ^ n19994 ^ 1'b0 ;
  assign n39272 = n7778 ^ n4864 ^ 1'b0 ;
  assign n39275 = n39274 ^ n39272 ^ n5160 ;
  assign n39276 = ( n5497 & n18190 ) | ( n5497 & ~n39275 ) | ( n18190 & ~n39275 ) ;
  assign n39277 = n37748 ^ n34233 ^ n10057 ;
  assign n39278 = ~n23924 & n39277 ;
  assign n39279 = n39278 ^ n20637 ^ 1'b0 ;
  assign n39280 = n13016 ^ n7242 ^ 1'b0 ;
  assign n39281 = ~n32020 & n39280 ;
  assign n39282 = n21748 ^ n11599 ^ 1'b0 ;
  assign n39283 = n9056 | n39282 ;
  assign n39284 = n31846 & ~n39283 ;
  assign n39285 = ~n4159 & n38060 ;
  assign n39286 = ~n18836 & n39285 ;
  assign n39290 = n2903 & ~n25396 ;
  assign n39291 = n11525 & n39290 ;
  assign n39287 = n1577 | n1824 ;
  assign n39288 = n39287 ^ n12763 ^ 1'b0 ;
  assign n39289 = ~n20223 & n39288 ;
  assign n39292 = n39291 ^ n39289 ^ 1'b0 ;
  assign n39293 = n11772 & n21801 ;
  assign n39294 = n39293 ^ n36135 ^ 1'b0 ;
  assign n39295 = n27123 ^ n21034 ^ 1'b0 ;
  assign n39296 = n10529 & n10909 ;
  assign n39297 = n37246 ^ n22196 ^ 1'b0 ;
  assign n39298 = n25420 & n39297 ;
  assign n39299 = n39298 ^ n30313 ^ n2868 ;
  assign n39300 = n19269 & ~n28046 ;
  assign n39301 = n39300 ^ n6827 ^ 1'b0 ;
  assign n39302 = ~n17228 & n19026 ;
  assign n39303 = n39302 ^ n13176 ^ 1'b0 ;
  assign n39304 = ~n3357 & n5084 ;
  assign n39305 = n38269 & ~n39304 ;
  assign n39306 = n19583 ^ n9275 ^ 1'b0 ;
  assign n39307 = ( ~n1295 & n7178 ) | ( ~n1295 & n25372 ) | ( n7178 & n25372 ) ;
  assign n39308 = n39307 ^ n15366 ^ 1'b0 ;
  assign n39309 = n4380 & n39308 ;
  assign n39310 = n3920 & n39309 ;
  assign n39311 = n483 | n39310 ;
  assign n39312 = n39311 ^ n25123 ^ 1'b0 ;
  assign n39313 = n39312 ^ n18838 ^ 1'b0 ;
  assign n39314 = ~n10402 & n34076 ;
  assign n39315 = n39314 ^ n357 ^ 1'b0 ;
  assign n39316 = ~n14012 & n20077 ;
  assign n39317 = n39316 ^ n23560 ^ 1'b0 ;
  assign n39318 = n485 & ~n35410 ;
  assign n39319 = n32041 ^ n5659 ^ 1'b0 ;
  assign n39320 = n38127 & ~n39319 ;
  assign n39321 = n37039 ^ n23628 ^ n2144 ;
  assign n39323 = n18596 ^ x192 ^ 1'b0 ;
  assign n39322 = n5921 & ~n20328 ;
  assign n39324 = n39323 ^ n39322 ^ 1'b0 ;
  assign n39325 = ~n2885 & n39324 ;
  assign n39326 = n6325 & ~n9210 ;
  assign n39327 = ~n39325 & n39326 ;
  assign n39328 = n34034 ^ n13170 ^ 1'b0 ;
  assign n39329 = n18240 ^ n9612 ^ 1'b0 ;
  assign n39330 = n8943 ^ n4962 ^ 1'b0 ;
  assign n39331 = ~n13175 & n39330 ;
  assign n39332 = n39331 ^ n22539 ^ 1'b0 ;
  assign n39336 = n1589 & n3885 ;
  assign n39334 = n2320 & n7200 ;
  assign n39335 = ~n6443 & n39334 ;
  assign n39333 = ~n8275 & n12033 ;
  assign n39337 = n39336 ^ n39335 ^ n39333 ;
  assign n39338 = n32130 ^ n28991 ^ 1'b0 ;
  assign n39339 = n39338 ^ n20564 ^ 1'b0 ;
  assign n39340 = ~n26054 & n39339 ;
  assign n39341 = n3424 | n6415 ;
  assign n39342 = n8642 & ~n39341 ;
  assign n39343 = ~n3782 & n5221 ;
  assign n39344 = n18969 & ~n24201 ;
  assign n39345 = n39343 & n39344 ;
  assign n39346 = ~n19786 & n35341 ;
  assign n39347 = ~n34456 & n39346 ;
  assign n39348 = n19068 & n19408 ;
  assign n39349 = n39348 ^ n17488 ^ 1'b0 ;
  assign n39350 = n38344 ^ n617 ^ 1'b0 ;
  assign n39351 = n11313 & ~n32654 ;
  assign n39352 = n27055 ^ n5962 ^ 1'b0 ;
  assign n39353 = n28835 ^ n13101 ^ 1'b0 ;
  assign n39354 = ~n39251 & n39353 ;
  assign n39355 = n16193 ^ n2045 ^ 1'b0 ;
  assign n39356 = n23229 & n25727 ;
  assign n39357 = ~n20165 & n39356 ;
  assign n39358 = n28271 & ~n39357 ;
  assign n39359 = n39355 & n39358 ;
  assign n39360 = n12013 ^ n8627 ^ 1'b0 ;
  assign n39361 = n20332 | n39360 ;
  assign n39362 = n39361 ^ n35028 ^ n1928 ;
  assign n39363 = n26168 ^ n10668 ^ n9226 ;
  assign n39364 = n10356 ^ n1527 ^ 1'b0 ;
  assign n39365 = ( n7457 & ~n33609 ) | ( n7457 & n39364 ) | ( ~n33609 & n39364 ) ;
  assign n39366 = n26499 & n34382 ;
  assign n39367 = n39365 & n39366 ;
  assign n39368 = n28288 & ~n29728 ;
  assign n39369 = n31108 ^ n2131 ^ 1'b0 ;
  assign n39371 = n1624 & n15828 ;
  assign n39372 = n13508 & n39371 ;
  assign n39370 = ~n8963 & n35246 ;
  assign n39373 = n39372 ^ n39370 ^ 1'b0 ;
  assign n39374 = n6642 & n21371 ;
  assign n39375 = n11607 | n39374 ;
  assign n39376 = n27796 & ~n39375 ;
  assign n39377 = n2189 | n39376 ;
  assign n39378 = n15870 | n39377 ;
  assign n39379 = ~n11365 & n17708 ;
  assign n39380 = n7265 & n39379 ;
  assign n39381 = n39252 ^ n15319 ^ 1'b0 ;
  assign n39382 = n39380 | n39381 ;
  assign n39383 = ( n970 & n10696 ) | ( n970 & ~n13023 ) | ( n10696 & ~n13023 ) ;
  assign n39384 = ( n296 & n12812 ) | ( n296 & ~n39383 ) | ( n12812 & ~n39383 ) ;
  assign n39385 = n14068 & ~n39384 ;
  assign n39386 = n23169 & ~n39385 ;
  assign n39387 = n25750 & n39386 ;
  assign n39388 = n14424 & ~n39387 ;
  assign n39389 = n39388 ^ n32226 ^ 1'b0 ;
  assign n39390 = n11017 ^ n5909 ^ 1'b0 ;
  assign n39391 = n26772 | n39390 ;
  assign n39392 = n8861 & ~n19241 ;
  assign n39393 = n39392 ^ n1346 ^ 1'b0 ;
  assign n39394 = n8889 & n14787 ;
  assign n39395 = n23482 & n39394 ;
  assign n39396 = n13896 & ~n21644 ;
  assign n39397 = n39396 ^ n7201 ^ 1'b0 ;
  assign n39398 = ~n26667 & n39397 ;
  assign n39399 = n39395 & n39398 ;
  assign n39400 = n5626 & ~n8423 ;
  assign n39401 = ~n29865 & n39400 ;
  assign n39402 = n39401 ^ n19826 ^ 1'b0 ;
  assign n39403 = n20599 ^ n1257 ^ 1'b0 ;
  assign n39404 = n14360 & n39403 ;
  assign n39405 = n27816 ^ n11926 ^ 1'b0 ;
  assign n39406 = n34052 & ~n39405 ;
  assign n39407 = ~n35585 & n39406 ;
  assign n39408 = ( n26401 & n39404 ) | ( n26401 & n39407 ) | ( n39404 & n39407 ) ;
  assign n39409 = ~n9031 & n37372 ;
  assign n39410 = n39409 ^ n35520 ^ 1'b0 ;
  assign n39411 = n9729 & ~n39410 ;
  assign n39412 = n39026 ^ n4460 ^ 1'b0 ;
  assign n39413 = n1795 & ~n39412 ;
  assign n39414 = n36784 ^ n31925 ^ 1'b0 ;
  assign n39415 = n38451 ^ n18611 ^ 1'b0 ;
  assign n39416 = n33801 & ~n39415 ;
  assign n39418 = ~n4003 & n8702 ;
  assign n39419 = n39418 ^ n2110 ^ 1'b0 ;
  assign n39417 = n1547 & n14927 ;
  assign n39420 = n39419 ^ n39417 ^ n5835 ;
  assign n39421 = ~n20501 & n39420 ;
  assign n39422 = n19695 ^ n3444 ^ 1'b0 ;
  assign n39423 = ~n19562 & n20030 ;
  assign n39424 = ~n10608 & n39423 ;
  assign n39425 = n23534 ^ n18265 ^ 1'b0 ;
  assign n39426 = n18773 ^ n4874 ^ 1'b0 ;
  assign n39427 = n12877 & ~n39426 ;
  assign n39428 = n25687 & ~n29261 ;
  assign n39429 = n39428 ^ n19726 ^ 1'b0 ;
  assign n39430 = n4935 & n19269 ;
  assign n39431 = n7293 | n24781 ;
  assign n39432 = n1466 | n39431 ;
  assign n39433 = n32556 & n39432 ;
  assign n39434 = n15129 ^ n14125 ^ n9691 ;
  assign n39435 = n5692 & ~n26115 ;
  assign n39436 = n39435 ^ n7504 ^ 1'b0 ;
  assign n39437 = n12337 | n39436 ;
  assign n39438 = n39437 ^ n5453 ^ 1'b0 ;
  assign n39439 = n3012 & n39438 ;
  assign n39440 = n8847 & n39439 ;
  assign n39441 = n20449 & ~n39440 ;
  assign n39442 = ( ~n1748 & n1763 ) | ( ~n1748 & n22810 ) | ( n1763 & n22810 ) ;
  assign n39443 = n32626 & n39442 ;
  assign n39444 = ~n8724 & n36284 ;
  assign n39445 = n39444 ^ n6466 ^ 1'b0 ;
  assign n39446 = n1352 | n11456 ;
  assign n39447 = n39445 & ~n39446 ;
  assign n39448 = n2133 | n24131 ;
  assign n39449 = n7815 ^ n6415 ^ 1'b0 ;
  assign n39450 = n1034 | n35967 ;
  assign n39451 = n28437 | n29084 ;
  assign n39452 = n1417 | n39451 ;
  assign n39453 = n2748 & n4832 ;
  assign n39455 = n28648 ^ n3012 ^ 1'b0 ;
  assign n39456 = n17651 | n39455 ;
  assign n39454 = ~n13014 & n15811 ;
  assign n39457 = n39456 ^ n39454 ^ 1'b0 ;
  assign n39458 = n39457 ^ n4508 ^ 1'b0 ;
  assign n39459 = ~n5746 & n14507 ;
  assign n39460 = ( n963 & n27933 ) | ( n963 & n39459 ) | ( n27933 & n39459 ) ;
  assign n39461 = n425 & ~n3168 ;
  assign n39462 = n11700 & n36975 ;
  assign n39465 = n9862 ^ n5074 ^ 1'b0 ;
  assign n39463 = n15088 & n16805 ;
  assign n39464 = n36821 & n39463 ;
  assign n39466 = n39465 ^ n39464 ^ 1'b0 ;
  assign n39467 = x62 & ~n1454 ;
  assign n39468 = ~n30459 & n39467 ;
  assign n39469 = n19509 ^ n9673 ^ 1'b0 ;
  assign n39470 = ~n22990 & n24909 ;
  assign n39471 = ( n17100 & n29081 ) | ( n17100 & n38614 ) | ( n29081 & n38614 ) ;
  assign n39472 = n23076 | n39043 ;
  assign n39473 = n39472 ^ n20257 ^ 1'b0 ;
  assign n39474 = ~n1151 & n7495 ;
  assign n39475 = n12100 | n16943 ;
  assign n39476 = n39475 ^ n17156 ^ 1'b0 ;
  assign n39477 = n15484 & ~n39476 ;
  assign n39478 = n39474 | n39477 ;
  assign n39479 = n28880 & n39478 ;
  assign n39480 = ~n39473 & n39479 ;
  assign n39481 = n36576 ^ n20236 ^ 1'b0 ;
  assign n39482 = n32630 ^ n7289 ^ 1'b0 ;
  assign n39483 = ~n14236 & n39482 ;
  assign n39484 = n35356 ^ n30403 ^ 1'b0 ;
  assign n39485 = n19916 | n39484 ;
  assign n39486 = n10145 & ~n11665 ;
  assign n39487 = n39486 ^ n1775 ^ 1'b0 ;
  assign n39488 = n25094 & ~n39487 ;
  assign n39489 = ~n4209 & n5759 ;
  assign n39490 = ~n39488 & n39489 ;
  assign n39491 = ~n501 & n14298 ;
  assign n39492 = n13747 & ~n39491 ;
  assign n39493 = ( ~n3977 & n16267 ) | ( ~n3977 & n39492 ) | ( n16267 & n39492 ) ;
  assign n39494 = n11057 ^ x240 ^ 1'b0 ;
  assign n39495 = n8947 & ~n39494 ;
  assign n39496 = n9428 & n39495 ;
  assign n39497 = ~n14593 & n28137 ;
  assign n39498 = n39496 & n39497 ;
  assign n39499 = n18260 & ~n19215 ;
  assign n39500 = n39499 ^ n2353 ^ 1'b0 ;
  assign n39501 = n39500 ^ n8452 ^ 1'b0 ;
  assign n39502 = n14405 & ~n39501 ;
  assign n39503 = n39502 ^ n1311 ^ 1'b0 ;
  assign n39504 = n37144 ^ n26280 ^ 1'b0 ;
  assign n39505 = ~n7486 & n39504 ;
  assign n39506 = n37020 ^ n23065 ^ 1'b0 ;
  assign n39507 = ~n3613 & n39506 ;
  assign n39508 = n3676 | n37388 ;
  assign n39509 = n7887 & ~n13880 ;
  assign n39510 = n22046 & n39509 ;
  assign n39511 = ( ~n7600 & n23387 ) | ( ~n7600 & n39510 ) | ( n23387 & n39510 ) ;
  assign n39512 = n12930 & n26973 ;
  assign n39513 = n39120 ^ n23510 ^ 1'b0 ;
  assign n39514 = n17344 & ~n39513 ;
  assign n39515 = n10102 & n12845 ;
  assign n39516 = n39515 ^ n4360 ^ 1'b0 ;
  assign n39517 = n4730 & ~n17956 ;
  assign n39518 = ~n37925 & n39517 ;
  assign n39519 = n13293 & ~n14304 ;
  assign n39520 = n39519 ^ n20212 ^ 1'b0 ;
  assign n39521 = n937 & n20759 ;
  assign n39522 = n2514 & n39521 ;
  assign n39523 = ~n4377 & n5172 ;
  assign n39524 = n39523 ^ n12553 ^ 1'b0 ;
  assign n39525 = n11713 | n35205 ;
  assign n39526 = n30081 ^ n19964 ^ n17583 ;
  assign n39527 = ( n25445 & n31384 ) | ( n25445 & n39526 ) | ( n31384 & n39526 ) ;
  assign n39528 = ~n18793 & n32942 ;
  assign n39529 = n3683 & n39528 ;
  assign n39530 = n14608 ^ n7910 ^ 1'b0 ;
  assign n39531 = n39530 ^ n11730 ^ 1'b0 ;
  assign n39532 = ~n28214 & n39531 ;
  assign n39533 = x146 & n8731 ;
  assign n39534 = n2792 & n4350 ;
  assign n39535 = ~n6872 & n28833 ;
  assign n39536 = n39534 & n39535 ;
  assign n39537 = n14590 ^ n7241 ^ 1'b0 ;
  assign n39538 = n4285 & n39537 ;
  assign n39539 = ~n34809 & n39538 ;
  assign n39540 = n14551 ^ n11714 ^ 1'b0 ;
  assign n39541 = n15249 & n39540 ;
  assign n39542 = ~n10272 & n15495 ;
  assign n39543 = n39542 ^ n10329 ^ 1'b0 ;
  assign n39544 = n17922 | n39543 ;
  assign n39545 = n1204 | n13766 ;
  assign n39546 = n3488 & ~n18270 ;
  assign n39547 = n39545 & n39546 ;
  assign n39548 = n2959 & ~n34552 ;
  assign n39549 = n39547 & n39548 ;
  assign n39550 = n1311 & n39549 ;
  assign n39552 = n37601 ^ n28379 ^ 1'b0 ;
  assign n39553 = ~n5768 & n39552 ;
  assign n39554 = n32285 & n39553 ;
  assign n39555 = ~n18149 & n39554 ;
  assign n39551 = n9251 & n9377 ;
  assign n39556 = n39555 ^ n39551 ^ 1'b0 ;
  assign n39557 = n22784 ^ n5748 ^ 1'b0 ;
  assign n39558 = n32671 & ~n39557 ;
  assign n39559 = ~n2993 & n22715 ;
  assign n39560 = n39559 ^ n37569 ^ 1'b0 ;
  assign n39561 = ~n22656 & n39560 ;
  assign n39562 = n12460 & ~n20807 ;
  assign n39563 = n15955 | n39562 ;
  assign n39564 = n18329 | n39563 ;
  assign n39565 = n9151 | n22817 ;
  assign n39566 = n5049 ^ n1203 ^ 1'b0 ;
  assign n39567 = n10627 & n39566 ;
  assign n39568 = n16144 & n21417 ;
  assign n39569 = n8969 & ~n39568 ;
  assign n39570 = n39567 & n39569 ;
  assign n39571 = ~n2473 & n5729 ;
  assign n39572 = n39571 ^ n8962 ^ 1'b0 ;
  assign n39573 = n17028 ^ n1129 ^ 1'b0 ;
  assign n39574 = ~n17289 & n34821 ;
  assign n39575 = ~n39573 & n39574 ;
  assign n39576 = n15828 | n39575 ;
  assign n39577 = ~n9977 & n14994 ;
  assign n39578 = n11102 ^ n6751 ^ 1'b0 ;
  assign n39579 = n39578 ^ n27719 ^ n20058 ;
  assign n39580 = n39579 ^ n30181 ^ 1'b0 ;
  assign n39581 = n17619 | n39580 ;
  assign n39582 = n15422 ^ n11017 ^ 1'b0 ;
  assign n39583 = ~n15366 & n39582 ;
  assign n39584 = ~n12139 & n24227 ;
  assign n39585 = ~n5628 & n39584 ;
  assign n39586 = ~n4714 & n24274 ;
  assign n39587 = ~n6295 & n11414 ;
  assign n39588 = ~x143 & n13988 ;
  assign n39589 = n39139 ^ n12276 ^ 1'b0 ;
  assign n39590 = n22961 & n39589 ;
  assign n39591 = ~n8956 & n14097 ;
  assign n39592 = ~n13060 & n27249 ;
  assign n39593 = n39592 ^ n6202 ^ 1'b0 ;
  assign n39594 = ~n270 & n1505 ;
  assign n39595 = n32762 ^ n932 ^ 1'b0 ;
  assign n39596 = n39594 & n39595 ;
  assign n39597 = n2615 | n10770 ;
  assign n39598 = n20799 ^ n5242 ^ 1'b0 ;
  assign n39599 = ~n39597 & n39598 ;
  assign n39600 = n10896 ^ n10777 ^ 1'b0 ;
  assign n39601 = n39599 & n39600 ;
  assign n39602 = ~n8134 & n39601 ;
  assign n39605 = n27826 & ~n31555 ;
  assign n39603 = ~n12388 & n18842 ;
  assign n39604 = n39603 ^ n24603 ^ 1'b0 ;
  assign n39606 = n39605 ^ n39604 ^ n13275 ;
  assign n39607 = n5628 & ~n20099 ;
  assign n39608 = n2726 ^ x163 ^ 1'b0 ;
  assign n39609 = n7868 ^ n2106 ^ 1'b0 ;
  assign n39610 = n2535 & ~n39609 ;
  assign n39611 = n1585 & n39610 ;
  assign n39612 = n39611 ^ n15835 ^ 1'b0 ;
  assign n39613 = n29225 ^ n14246 ^ 1'b0 ;
  assign n39614 = ~n39612 & n39613 ;
  assign n39615 = n36911 ^ n7968 ^ 1'b0 ;
  assign n39616 = n39614 & n39615 ;
  assign n39617 = n4584 ^ n992 ^ 1'b0 ;
  assign n39618 = n5209 & ~n18444 ;
  assign n39619 = n39618 ^ n24892 ^ 1'b0 ;
  assign n39620 = n23844 ^ n6020 ^ n1172 ;
  assign n39621 = n26912 ^ n25292 ^ 1'b0 ;
  assign n39622 = n32511 & ~n39621 ;
  assign n39623 = n2657 & ~n4639 ;
  assign n39624 = n39623 ^ n1882 ^ 1'b0 ;
  assign n39627 = ~n2418 & n37737 ;
  assign n39628 = n39627 ^ n1008 ^ 1'b0 ;
  assign n39625 = x178 & ~n13719 ;
  assign n39626 = ~n26306 & n39625 ;
  assign n39629 = n39628 ^ n39626 ^ 1'b0 ;
  assign n39630 = n5536 & ~n17836 ;
  assign n39631 = n39630 ^ n29562 ^ 1'b0 ;
  assign n39632 = ~n13087 & n39631 ;
  assign n39633 = n16451 & ~n39632 ;
  assign n39634 = n2489 | n11047 ;
  assign n39635 = n39634 ^ n7798 ^ 1'b0 ;
  assign n39636 = n982 ^ n733 ^ 1'b0 ;
  assign n39637 = n39635 & ~n39636 ;
  assign n39638 = n8118 & ~n19527 ;
  assign n39639 = n19593 ^ n4642 ^ 1'b0 ;
  assign n39640 = ~n1349 & n22026 ;
  assign n39641 = n39640 ^ n9086 ^ 1'b0 ;
  assign n39642 = n12900 & ~n39641 ;
  assign n39643 = n30773 ^ n17636 ^ 1'b0 ;
  assign n39644 = n23331 ^ n1149 ^ 1'b0 ;
  assign n39645 = n39643 | n39644 ;
  assign n39646 = n38667 ^ n1672 ^ 1'b0 ;
  assign n39647 = n35029 & n39646 ;
  assign n39648 = n38628 ^ n2875 ^ 1'b0 ;
  assign n39649 = n25924 ^ n18436 ^ n9562 ;
  assign n39650 = ~n2416 & n5513 ;
  assign n39651 = ~n12962 & n26960 ;
  assign n39652 = n39650 & n39651 ;
  assign n39653 = n3140 & ~n32832 ;
  assign n39654 = n2269 | n7800 ;
  assign n39655 = n2297 | n10305 ;
  assign n39656 = n2106 & ~n11467 ;
  assign n39657 = n31923 & n39656 ;
  assign n39658 = n19002 ^ n15289 ^ 1'b0 ;
  assign n39659 = n15648 & n39658 ;
  assign n39660 = n36939 ^ n8406 ^ 1'b0 ;
  assign n39661 = n19592 ^ n3073 ^ n1001 ;
  assign n39662 = n19723 ^ n13890 ^ 1'b0 ;
  assign n39663 = n1688 & n18868 ;
  assign n39664 = n39663 ^ n35006 ^ 1'b0 ;
  assign n39665 = n39664 ^ n14701 ^ 1'b0 ;
  assign n39666 = n6424 & ~n8408 ;
  assign n39667 = n39666 ^ n5621 ^ 1'b0 ;
  assign n39670 = n27094 ^ n13740 ^ 1'b0 ;
  assign n39671 = n33824 & ~n39670 ;
  assign n39668 = n17394 ^ n7709 ^ n4033 ;
  assign n39669 = n15774 & ~n39668 ;
  assign n39672 = n39671 ^ n39669 ^ 1'b0 ;
  assign n39673 = n39672 ^ n12780 ^ 1'b0 ;
  assign n39674 = n36917 & ~n38305 ;
  assign n39675 = ~n7070 & n39674 ;
  assign n39676 = n20073 ^ n6139 ^ 1'b0 ;
  assign n39677 = ~n15689 & n39676 ;
  assign n39678 = n19901 ^ n318 ^ 1'b0 ;
  assign n39679 = n5871 & ~n24558 ;
  assign n39680 = n10655 & ~n24867 ;
  assign n39681 = n39679 & n39680 ;
  assign n39682 = ( n12539 & ~n34151 ) | ( n12539 & n39681 ) | ( ~n34151 & n39681 ) ;
  assign n39683 = n6342 & n18718 ;
  assign n39684 = ~n613 & n39683 ;
  assign n39685 = n6139 ^ n4142 ^ n3823 ;
  assign n39686 = n29578 & n39685 ;
  assign n39687 = ~n5315 & n7702 ;
  assign n39688 = n39687 ^ n38408 ^ n9911 ;
  assign n39689 = n17185 | n39688 ;
  assign n39690 = n6923 & n11645 ;
  assign n39691 = ( ~n13626 & n18018 ) | ( ~n13626 & n19581 ) | ( n18018 & n19581 ) ;
  assign n39692 = n28761 & ~n39691 ;
  assign n39693 = ~n20389 & n39692 ;
  assign n39694 = ~n39690 & n39693 ;
  assign n39695 = n18703 ^ n11695 ^ n858 ;
  assign n39696 = n24326 | n25292 ;
  assign n39697 = n32556 & ~n39696 ;
  assign n39698 = n39697 ^ n7298 ^ 1'b0 ;
  assign n39699 = ( n7212 & ~n15071 ) | ( n7212 & n19525 ) | ( ~n15071 & n19525 ) ;
  assign n39700 = n20662 ^ n970 ^ 1'b0 ;
  assign n39701 = ~n39699 & n39700 ;
  assign n39702 = n38614 ^ n14929 ^ 1'b0 ;
  assign n39703 = n1196 | n39702 ;
  assign n39704 = ( n1696 & n17262 ) | ( n1696 & n32437 ) | ( n17262 & n32437 ) ;
  assign n39705 = n25102 & n39704 ;
  assign n39706 = ~n733 & n6978 ;
  assign n39707 = n16886 & ~n24096 ;
  assign n39708 = n22567 ^ n21680 ^ 1'b0 ;
  assign n39709 = n28033 & n39708 ;
  assign n39710 = n4840 | n7321 ;
  assign n39711 = n39710 ^ x150 ^ 1'b0 ;
  assign n39712 = n23184 & ~n23482 ;
  assign n39713 = ~n39711 & n39712 ;
  assign n39714 = ~n12940 & n30807 ;
  assign n39715 = n22113 ^ n10281 ^ 1'b0 ;
  assign n39716 = n24809 | n39715 ;
  assign n39717 = n17555 ^ n14662 ^ 1'b0 ;
  assign n39718 = n34297 & ~n39717 ;
  assign n39719 = n11053 ^ n4588 ^ 1'b0 ;
  assign n39720 = n9623 ^ n8373 ^ 1'b0 ;
  assign n39721 = ~n39719 & n39720 ;
  assign n39722 = n2148 | n3483 ;
  assign n39723 = n39722 ^ n14294 ^ 1'b0 ;
  assign n39724 = n25977 & ~n39723 ;
  assign n39725 = n25565 ^ n9943 ^ 1'b0 ;
  assign n39726 = n2192 & ~n3228 ;
  assign n39727 = ( ~n16660 & n34246 ) | ( ~n16660 & n39726 ) | ( n34246 & n39726 ) ;
  assign n39728 = n39727 ^ n37366 ^ n26716 ;
  assign n39729 = n39728 ^ n13299 ^ 1'b0 ;
  assign n39730 = ( n4085 & ~n11696 ) | ( n4085 & n19893 ) | ( ~n11696 & n19893 ) ;
  assign n39731 = n13195 & n39730 ;
  assign n39732 = ~n5132 & n20129 ;
  assign n39733 = ~n18104 & n39732 ;
  assign n39734 = n8018 & ~n16372 ;
  assign n39735 = n23794 & n39734 ;
  assign n39736 = ~n1326 & n12553 ;
  assign n39737 = n39736 ^ n5830 ^ 1'b0 ;
  assign n39738 = n5418 & n12161 ;
  assign n39739 = ~n4551 & n39738 ;
  assign n39740 = n23199 ^ n5936 ^ 1'b0 ;
  assign n39741 = n17065 & ~n39740 ;
  assign n39742 = n7741 | n28281 ;
  assign n39743 = n39742 ^ n6062 ^ 1'b0 ;
  assign n39744 = n11465 & ~n16879 ;
  assign n39745 = n39744 ^ n5262 ^ 1'b0 ;
  assign n39746 = ~n2272 & n25906 ;
  assign n39747 = n39745 & n39746 ;
  assign n39748 = n4180 & ~n39088 ;
  assign n39749 = n39747 & n39748 ;
  assign n39750 = ~n6401 & n8424 ;
  assign n39751 = ~n11512 & n13101 ;
  assign n39752 = n34475 ^ n6682 ^ 1'b0 ;
  assign n39753 = ~n6561 & n14752 ;
  assign n39754 = ~n9280 & n20090 ;
  assign n39755 = n39754 ^ n34270 ^ 1'b0 ;
  assign n39756 = n14488 ^ n11863 ^ 1'b0 ;
  assign n39757 = x115 & ~n39756 ;
  assign n39758 = n2912 & ~n11349 ;
  assign n39759 = n8130 & n39758 ;
  assign n39760 = n39759 ^ n29591 ^ 1'b0 ;
  assign n39761 = n14471 & ~n39760 ;
  assign n39762 = n4245 & n22538 ;
  assign n39763 = n22558 | n39762 ;
  assign n39764 = n27787 ^ n10097 ^ 1'b0 ;
  assign n39765 = n13338 | n39764 ;
  assign n39766 = n35692 ^ n27317 ^ n287 ;
  assign n39767 = n24265 ^ n10961 ^ 1'b0 ;
  assign n39768 = n3059 | n39767 ;
  assign n39769 = n18796 & ~n19828 ;
  assign n39770 = n3785 & n39769 ;
  assign n39771 = n34442 ^ n20898 ^ 1'b0 ;
  assign n39772 = ~n39770 & n39771 ;
  assign n39773 = n13486 & n34758 ;
  assign n39774 = n3600 & ~n35853 ;
  assign n39775 = ~n13158 & n39774 ;
  assign n39776 = n18892 ^ n9121 ^ 1'b0 ;
  assign n39777 = ( n16128 & n18658 ) | ( n16128 & n39776 ) | ( n18658 & n39776 ) ;
  assign n39778 = n38746 ^ n14061 ^ n9526 ;
  assign n39779 = n2738 & ~n10225 ;
  assign n39782 = ~n19211 & n25659 ;
  assign n39783 = n39782 ^ n2794 ^ 1'b0 ;
  assign n39780 = n5773 ^ n4298 ^ 1'b0 ;
  assign n39781 = x107 & n39780 ;
  assign n39784 = n39783 ^ n39781 ^ 1'b0 ;
  assign n39785 = n13433 ^ n11061 ^ n4403 ;
  assign n39786 = n39785 ^ n28033 ^ n11371 ;
  assign n39787 = n39786 ^ n4267 ^ 1'b0 ;
  assign n39788 = n3118 & n3661 ;
  assign n39789 = n39788 ^ n25747 ^ 1'b0 ;
  assign n39790 = n8508 | n39789 ;
  assign n39791 = n16363 ^ n13261 ^ 1'b0 ;
  assign n39792 = n4869 | n39791 ;
  assign n39793 = n14774 ^ n14212 ^ 1'b0 ;
  assign n39794 = n26585 & ~n39793 ;
  assign n39795 = ~n1344 & n20407 ;
  assign n39796 = n27786 & n39795 ;
  assign n39797 = ~n6072 & n13742 ;
  assign n39798 = n35665 ^ n7887 ^ n6554 ;
  assign n39799 = n5696 | n17863 ;
  assign n39800 = n39799 ^ n14609 ^ 1'b0 ;
  assign n39801 = n12419 & ~n23513 ;
  assign n39802 = ~n11534 & n39801 ;
  assign n39803 = ~n4714 & n39802 ;
  assign n39804 = n4962 & ~n12501 ;
  assign n39805 = n1645 & ~n15874 ;
  assign n39806 = ~n12141 & n39805 ;
  assign n39807 = n11499 & n39806 ;
  assign n39808 = n11743 & ~n39807 ;
  assign n39809 = ~n9829 & n39808 ;
  assign n39810 = n8626 & ~n39809 ;
  assign n39811 = n24424 & n39810 ;
  assign n39812 = n9525 & n31052 ;
  assign n39813 = ~n6550 & n14936 ;
  assign n39814 = n39812 | n39813 ;
  assign n39815 = ( ~n11479 & n23126 ) | ( ~n11479 & n24386 ) | ( n23126 & n24386 ) ;
  assign n39816 = ~n23967 & n39815 ;
  assign n39817 = n36554 | n39816 ;
  assign n39818 = ~x196 & n9646 ;
  assign n39819 = n1990 | n10267 ;
  assign n39820 = n39819 ^ n5502 ^ 1'b0 ;
  assign n39821 = n39820 ^ n1373 ^ 1'b0 ;
  assign n39822 = ( n6097 & ~n16433 ) | ( n6097 & n27030 ) | ( ~n16433 & n27030 ) ;
  assign n39824 = n3648 ^ n1261 ^ 1'b0 ;
  assign n39825 = n24973 | n39824 ;
  assign n39823 = n2397 & n6293 ;
  assign n39826 = n39825 ^ n39823 ^ 1'b0 ;
  assign n39827 = n3957 & ~n5898 ;
  assign n39828 = n20407 | n39827 ;
  assign n39829 = n4778 | n17408 ;
  assign n39830 = n39829 ^ n1975 ^ 1'b0 ;
  assign n39831 = n5445 ^ x120 ^ 1'b0 ;
  assign n39834 = n15432 & n24066 ;
  assign n39835 = ( n20631 & n25977 ) | ( n20631 & n39834 ) | ( n25977 & n39834 ) ;
  assign n39832 = n16221 ^ n12798 ^ 1'b0 ;
  assign n39833 = ~n34512 & n39832 ;
  assign n39836 = n39835 ^ n39833 ^ 1'b0 ;
  assign n39837 = n1349 | n1499 ;
  assign n39838 = n32709 & ~n39837 ;
  assign n39843 = n1002 ^ n425 ^ 1'b0 ;
  assign n39844 = n3912 | n39843 ;
  assign n39839 = n7584 ^ n7212 ^ 1'b0 ;
  assign n39840 = n708 & n39839 ;
  assign n39841 = n2383 | n39840 ;
  assign n39842 = n13044 & n39841 ;
  assign n39845 = n39844 ^ n39842 ^ 1'b0 ;
  assign n39846 = n5881 & n9728 ;
  assign n39847 = n39846 ^ n14073 ^ 1'b0 ;
  assign n39848 = n39847 ^ n20406 ^ 1'b0 ;
  assign n39849 = ( n1905 & n4583 ) | ( n1905 & ~n9681 ) | ( n4583 & ~n9681 ) ;
  assign n39850 = n34734 ^ n13106 ^ 1'b0 ;
  assign n39851 = ~n10484 & n18434 ;
  assign n39852 = ~n3922 & n39851 ;
  assign n39853 = n3935 | n17657 ;
  assign n39854 = ( n17674 & ~n23711 ) | ( n17674 & n39853 ) | ( ~n23711 & n39853 ) ;
  assign n39855 = n3592 | n21465 ;
  assign n39856 = n39855 ^ n7781 ^ 1'b0 ;
  assign n39857 = n8123 | n14547 ;
  assign n39858 = n30353 & ~n39857 ;
  assign n39859 = n21488 ^ n8660 ^ 1'b0 ;
  assign n39860 = ~n39858 & n39859 ;
  assign n39861 = ~x26 & n16484 ;
  assign n39862 = n671 & n26335 ;
  assign n39863 = n39861 & n39862 ;
  assign n39864 = n39863 ^ n21708 ^ 1'b0 ;
  assign n39865 = n959 & n38128 ;
  assign n39866 = n4541 ^ n727 ^ 1'b0 ;
  assign n39867 = ~n39865 & n39866 ;
  assign n39873 = ~n2968 & n9447 ;
  assign n39874 = n16062 | n39873 ;
  assign n39868 = n6930 ^ n3650 ^ 1'b0 ;
  assign n39869 = n1311 & n6687 ;
  assign n39870 = ~n1600 & n39869 ;
  assign n39871 = n39870 ^ n4321 ^ 1'b0 ;
  assign n39872 = n39868 & ~n39871 ;
  assign n39875 = n39874 ^ n39872 ^ n34007 ;
  assign n39876 = n2306 & n16624 ;
  assign n39877 = n37710 ^ n25386 ^ 1'b0 ;
  assign n39878 = n38494 ^ n25368 ^ 1'b0 ;
  assign n39879 = n39062 | n39878 ;
  assign n39880 = n17642 & n30299 ;
  assign n39881 = n9970 | n29256 ;
  assign n39882 = n39881 ^ n30810 ^ 1'b0 ;
  assign n39883 = n7180 & n39882 ;
  assign n39884 = n14815 ^ n2466 ^ 1'b0 ;
  assign n39885 = n5207 | n39884 ;
  assign n39886 = ~n34170 & n39885 ;
  assign n39887 = ~n1490 & n39886 ;
  assign n39888 = n17718 | n18098 ;
  assign n39889 = n39888 ^ n13212 ^ 1'b0 ;
  assign n39890 = n31177 ^ n21220 ^ n15622 ;
  assign n39891 = n16042 & ~n39890 ;
  assign n39892 = n5959 ^ n2297 ^ 1'b0 ;
  assign n39893 = n20374 ^ n12694 ^ 1'b0 ;
  assign n39894 = n17047 | n39893 ;
  assign n39895 = ( n8632 & n39331 ) | ( n8632 & n39894 ) | ( n39331 & n39894 ) ;
  assign n39896 = ( ~n6639 & n39892 ) | ( ~n6639 & n39895 ) | ( n39892 & n39895 ) ;
  assign n39897 = ( n4685 & ~n12840 ) | ( n4685 & n22726 ) | ( ~n12840 & n22726 ) ;
  assign n39898 = n10150 & ~n39897 ;
  assign n39899 = ~n14016 & n39898 ;
  assign n39900 = ( n20902 & n22321 ) | ( n20902 & ~n39899 ) | ( n22321 & ~n39899 ) ;
  assign n39901 = n1487 | n9531 ;
  assign n39902 = n19616 | n39901 ;
  assign n39903 = n1551 & ~n3210 ;
  assign n39904 = n3913 | n20242 ;
  assign n39905 = n14172 & ~n39904 ;
  assign n39906 = n32261 ^ n12924 ^ 1'b0 ;
  assign n39907 = n13054 | n39906 ;
  assign n39908 = ( n3772 & n14845 ) | ( n3772 & n35901 ) | ( n14845 & n35901 ) ;
  assign n39909 = n18300 ^ n2678 ^ 1'b0 ;
  assign n39910 = n724 ^ x140 ^ 1'b0 ;
  assign n39911 = n5498 | n39910 ;
  assign n39912 = ~n21421 & n36733 ;
  assign n39913 = ~n26352 & n33444 ;
  assign n39914 = ( ~n5566 & n10108 ) | ( ~n5566 & n11557 ) | ( n10108 & n11557 ) ;
  assign n39915 = n1276 & ~n14890 ;
  assign n39916 = n7866 & n27385 ;
  assign n39917 = n1928 & n39916 ;
  assign n39918 = n4394 | n15423 ;
  assign n39919 = n39918 ^ n4766 ^ 1'b0 ;
  assign n39920 = n29668 & ~n39919 ;
  assign n39921 = n39917 & n39920 ;
  assign n39922 = ~n9260 & n32571 ;
  assign n39923 = n3820 | n12493 ;
  assign n39924 = ( n3646 & n23659 ) | ( n3646 & n39923 ) | ( n23659 & n39923 ) ;
  assign n39925 = n566 | n9599 ;
  assign n39926 = ~n8425 & n39925 ;
  assign n39927 = n39926 ^ n7036 ^ 1'b0 ;
  assign n39928 = n24615 ^ n6202 ^ 1'b0 ;
  assign n39929 = n39927 & n39928 ;
  assign n39930 = n39929 ^ n12584 ^ n2649 ;
  assign n39931 = n1199 & ~n6817 ;
  assign n39932 = n5811 & n39790 ;
  assign n39933 = n1738 & n23527 ;
  assign n39934 = ~n3041 & n39933 ;
  assign n39935 = n12394 & ~n39934 ;
  assign n39936 = n11153 & n39935 ;
  assign n39937 = n25570 ^ n18166 ^ 1'b0 ;
  assign n39938 = n2893 & n39937 ;
  assign n39939 = n1947 & n39938 ;
  assign n39940 = n39939 ^ n5018 ^ 1'b0 ;
  assign n39941 = n27743 & n31133 ;
  assign n39942 = n34469 ^ n8406 ^ 1'b0 ;
  assign n39943 = n16612 ^ n9739 ^ 1'b0 ;
  assign n39944 = n35831 & ~n39943 ;
  assign n39945 = n16269 | n24433 ;
  assign n39946 = n5025 | n39945 ;
  assign n39947 = n39946 ^ n15475 ^ 1'b0 ;
  assign n39948 = ~n1186 & n8063 ;
  assign n39949 = n34382 ^ n5067 ^ 1'b0 ;
  assign n39950 = n30315 | n39949 ;
  assign n39951 = n8016 & ~n13398 ;
  assign n39952 = n39950 & n39951 ;
  assign n39953 = ( n10455 & ~n14547 ) | ( n10455 & n39952 ) | ( ~n14547 & n39952 ) ;
  assign n39954 = n14369 ^ n4910 ^ 1'b0 ;
  assign n39955 = ( ~n13971 & n14476 ) | ( ~n13971 & n39954 ) | ( n14476 & n39954 ) ;
  assign n39956 = n6454 & n18352 ;
  assign n39957 = n11406 ^ n4524 ^ 1'b0 ;
  assign n39958 = n27101 & n30217 ;
  assign n39959 = n20144 ^ n7957 ^ 1'b0 ;
  assign n39960 = n8056 & ~n27480 ;
  assign n39961 = n34120 & ~n36160 ;
  assign n39962 = n11539 ^ n11175 ^ 1'b0 ;
  assign n39963 = n7411 | n39962 ;
  assign n39964 = n39963 ^ n1404 ^ 1'b0 ;
  assign n39965 = n24024 ^ n11383 ^ n4589 ;
  assign n39966 = n39965 ^ n2999 ^ 1'b0 ;
  assign n39967 = n13567 & n39966 ;
  assign n39968 = n507 & n39967 ;
  assign n39969 = n32830 ^ n12665 ^ 1'b0 ;
  assign n39970 = n31269 ^ n1021 ^ 1'b0 ;
  assign n39971 = n2037 & n39970 ;
  assign n39972 = ~n3380 & n6395 ;
  assign n39973 = ~n19545 & n36759 ;
  assign n39974 = n6415 | n17938 ;
  assign n39975 = n17602 | n39974 ;
  assign n39976 = n39975 ^ n18679 ^ 1'b0 ;
  assign n39977 = n30977 & n39976 ;
  assign n39978 = n12812 ^ n6688 ^ 1'b0 ;
  assign n39979 = n34168 ^ n4242 ^ 1'b0 ;
  assign n39980 = n28429 ^ n13100 ^ n4721 ;
  assign n39981 = n14516 | n39980 ;
  assign n39982 = n39981 ^ n4319 ^ 1'b0 ;
  assign n39983 = n14861 | n39982 ;
  assign n39984 = n8030 ^ n6367 ^ 1'b0 ;
  assign n39985 = n36457 ^ n35015 ^ 1'b0 ;
  assign n39986 = n5576 & ~n17008 ;
  assign n39987 = ~n4844 & n37094 ;
  assign n39988 = n14635 ^ n4315 ^ 1'b0 ;
  assign n39989 = n36410 ^ n35157 ^ 1'b0 ;
  assign n39990 = n9683 | n15039 ;
  assign n39991 = n39990 ^ n24541 ^ 1'b0 ;
  assign n39992 = n39991 ^ n32753 ^ n6490 ;
  assign n39993 = n6254 & ~n22652 ;
  assign n39994 = ~n30959 & n39993 ;
  assign n39995 = n39994 ^ n12998 ^ 1'b0 ;
  assign n39996 = n5130 & ~n8925 ;
  assign n39997 = ~n2382 & n39996 ;
  assign n39999 = n20166 ^ n7207 ^ 1'b0 ;
  assign n40000 = ~n5900 & n39999 ;
  assign n39998 = x76 & n4629 ;
  assign n40001 = n40000 ^ n39998 ^ 1'b0 ;
  assign n40002 = n25004 & n27281 ;
  assign n40003 = n40002 ^ n23260 ^ 1'b0 ;
  assign n40004 = n10178 & ~n33052 ;
  assign n40005 = ~n8177 & n40004 ;
  assign n40007 = n14784 ^ n6131 ^ 1'b0 ;
  assign n40008 = n14008 & n40007 ;
  assign n40009 = ~n464 & n40008 ;
  assign n40006 = n20251 & ~n22959 ;
  assign n40010 = n40009 ^ n40006 ^ 1'b0 ;
  assign n40011 = n19947 ^ n16098 ^ n5472 ;
  assign n40012 = n2014 & ~n35169 ;
  assign n40013 = n5996 & ~n13710 ;
  assign n40014 = n40013 ^ n25132 ^ 1'b0 ;
  assign n40015 = n14724 & n22249 ;
  assign n40016 = n16530 | n22931 ;
  assign n40017 = n16530 & ~n40016 ;
  assign n40018 = n1345 & n22715 ;
  assign n40019 = ~n24521 & n40018 ;
  assign n40020 = n40019 ^ n19660 ^ 1'b0 ;
  assign n40021 = n23061 & n40020 ;
  assign n40022 = n6640 & ~n34805 ;
  assign n40023 = ~n20084 & n40022 ;
  assign n40024 = n29865 ^ n9800 ^ 1'b0 ;
  assign n40025 = n26699 ^ n11665 ^ n11476 ;
  assign n40026 = n15360 ^ n4134 ^ 1'b0 ;
  assign n40027 = ~n6352 & n22537 ;
  assign n40028 = n25503 ^ n4284 ^ 1'b0 ;
  assign n40029 = ~n40027 & n40028 ;
  assign n40030 = n5442 | n40029 ;
  assign n40031 = ( n628 & ~n34127 ) | ( n628 & n36664 ) | ( ~n34127 & n36664 ) ;
  assign n40032 = n25175 | n40031 ;
  assign n40033 = n14639 & ~n35030 ;
  assign n40034 = n1096 & n5655 ;
  assign n40035 = n17113 ^ n1023 ^ 1'b0 ;
  assign n40036 = n40035 ^ n34632 ^ 1'b0 ;
  assign n40037 = n40034 & n40036 ;
  assign n40038 = n17967 ^ n13037 ^ n10322 ;
  assign n40039 = n6057 | n13362 ;
  assign n40040 = n28478 | n40039 ;
  assign n40041 = ( x185 & ~n6754 ) | ( x185 & n40040 ) | ( ~n6754 & n40040 ) ;
  assign n40042 = n15504 | n22047 ;
  assign n40043 = n40042 ^ n30751 ^ 1'b0 ;
  assign n40044 = n40043 ^ n7405 ^ 1'b0 ;
  assign n40045 = n22986 & n40044 ;
  assign n40046 = x40 & ~n4871 ;
  assign n40047 = n40046 ^ n5884 ^ 1'b0 ;
  assign n40048 = ~n8267 & n40047 ;
  assign n40049 = n40048 ^ n5748 ^ 1'b0 ;
  assign n40050 = n2081 & ~n10864 ;
  assign n40051 = n40050 ^ n5033 ^ 1'b0 ;
  assign n40052 = n20285 ^ n7830 ^ 1'b0 ;
  assign n40053 = ~n6688 & n40052 ;
  assign n40054 = n40053 ^ n15157 ^ 1'b0 ;
  assign n40055 = n7933 & n38344 ;
  assign n40056 = ~n40054 & n40055 ;
  assign n40057 = n6433 & n9348 ;
  assign n40058 = n8107 & n40057 ;
  assign n40059 = n40058 ^ n12621 ^ n4220 ;
  assign n40060 = n27594 ^ n6679 ^ 1'b0 ;
  assign n40061 = n37569 & ~n40060 ;
  assign n40062 = n26719 & n31593 ;
  assign n40063 = n40062 ^ n8276 ^ 1'b0 ;
  assign n40064 = n5165 | n39478 ;
  assign n40065 = ~n9803 & n22201 ;
  assign n40066 = n12962 & n40065 ;
  assign n40067 = n2797 & n20956 ;
  assign n40068 = n40067 ^ n26372 ^ 1'b0 ;
  assign n40069 = ~n3874 & n39610 ;
  assign n40070 = n16446 & n40069 ;
  assign n40071 = n21786 | n26656 ;
  assign n40072 = n19364 & ~n40071 ;
  assign n40073 = n26676 & n37249 ;
  assign n40074 = n18779 ^ n3018 ^ n2170 ;
  assign n40075 = n2640 | n40074 ;
  assign n40076 = n4585 ^ n3696 ^ 1'b0 ;
  assign n40077 = n40075 | n40076 ;
  assign n40078 = n34726 & n40077 ;
  assign n40079 = n5059 | n37850 ;
  assign n40080 = n40079 ^ n23357 ^ 1'b0 ;
  assign n40081 = n5231 | n18254 ;
  assign n40082 = n34197 ^ n20012 ^ 1'b0 ;
  assign n40083 = n14645 ^ n7634 ^ 1'b0 ;
  assign n40084 = n29380 ^ n13047 ^ n5357 ;
  assign n40085 = n6803 & n40084 ;
  assign n40086 = n16098 & ~n40085 ;
  assign n40087 = n40086 ^ n11703 ^ 1'b0 ;
  assign n40088 = n5949 & n21285 ;
  assign n40089 = n14036 | n40088 ;
  assign n40090 = n40089 ^ n18307 ^ 1'b0 ;
  assign n40091 = ~n2523 & n3634 ;
  assign n40092 = n40091 ^ n3066 ^ 1'b0 ;
  assign n40093 = n40092 ^ n28530 ^ 1'b0 ;
  assign n40094 = n31130 ^ n9393 ^ 1'b0 ;
  assign n40095 = n40094 ^ n11831 ^ n6767 ;
  assign n40096 = ( n11567 & ~n31586 ) | ( n11567 & n40095 ) | ( ~n31586 & n40095 ) ;
  assign n40097 = n11344 | n39128 ;
  assign n40098 = n40097 ^ n18511 ^ 1'b0 ;
  assign n40099 = n10200 | n40098 ;
  assign n40100 = n13419 | n40099 ;
  assign n40101 = n16697 ^ n6382 ^ 1'b0 ;
  assign n40102 = ~n8491 & n11825 ;
  assign n40103 = n40102 ^ n4253 ^ 1'b0 ;
  assign n40104 = n3508 & n40103 ;
  assign n40105 = n29956 & n40104 ;
  assign n40106 = n11920 | n25175 ;
  assign n40107 = n12245 & ~n40106 ;
  assign n40108 = ~n33961 & n40107 ;
  assign n40109 = ~n18777 & n29605 ;
  assign n40110 = ( n11964 & n31343 ) | ( n11964 & ~n40109 ) | ( n31343 & ~n40109 ) ;
  assign n40111 = ( n2810 & ~n12959 ) | ( n2810 & n31760 ) | ( ~n12959 & n31760 ) ;
  assign n40112 = ~n13049 & n17910 ;
  assign n40113 = n4861 & ~n25334 ;
  assign n40114 = n40112 & n40113 ;
  assign n40115 = n7140 & ~n40114 ;
  assign n40116 = n40115 ^ x63 ^ 1'b0 ;
  assign n40117 = n12330 & ~n13537 ;
  assign n40118 = n24478 & ~n35095 ;
  assign n40119 = n40118 ^ n18905 ^ 1'b0 ;
  assign n40120 = n4631 | n15987 ;
  assign n40121 = n40120 ^ n19972 ^ x46 ;
  assign n40122 = n8660 & ~n29664 ;
  assign n40123 = n40122 ^ n28321 ^ 1'b0 ;
  assign n40124 = n36630 | n40123 ;
  assign n40125 = n40124 ^ n5990 ^ 1'b0 ;
  assign n40126 = n14844 & n17085 ;
  assign n40127 = ~n27718 & n40126 ;
  assign n40128 = n28565 & n40127 ;
  assign n40129 = n5341 | n7198 ;
  assign n40130 = ~n7065 & n22440 ;
  assign n40131 = n860 & n40130 ;
  assign n40132 = n26037 | n40131 ;
  assign n40133 = ~n5367 & n22378 ;
  assign n40134 = n38454 ^ n2765 ^ 1'b0 ;
  assign n40135 = n24823 & ~n40134 ;
  assign n40136 = ( n20998 & n40133 ) | ( n20998 & ~n40135 ) | ( n40133 & ~n40135 ) ;
  assign n40138 = n12628 ^ n4341 ^ 1'b0 ;
  assign n40139 = n19778 | n40138 ;
  assign n40137 = n18195 & n29266 ;
  assign n40140 = n40139 ^ n40137 ^ 1'b0 ;
  assign n40141 = ~n8905 & n13616 ;
  assign n40142 = n40141 ^ n31685 ^ 1'b0 ;
  assign n40143 = n9692 & n40142 ;
  assign n40144 = n24336 | n27035 ;
  assign n40145 = n40144 ^ n22101 ^ 1'b0 ;
  assign n40146 = n16363 ^ n14335 ^ 1'b0 ;
  assign n40147 = n619 | n40146 ;
  assign n40148 = n31332 ^ n3740 ^ 1'b0 ;
  assign n40149 = n40147 | n40148 ;
  assign n40150 = n33231 ^ n22381 ^ 1'b0 ;
  assign n40151 = n16791 & n40150 ;
  assign n40152 = n10731 | n17426 ;
  assign n40153 = n11934 & n24897 ;
  assign n40154 = ~n40152 & n40153 ;
  assign n40155 = n40154 ^ n9056 ^ 1'b0 ;
  assign n40156 = n25231 ^ n7832 ^ 1'b0 ;
  assign n40157 = n6695 & n40156 ;
  assign n40158 = n16259 | n34808 ;
  assign n40159 = n8331 & ~n20832 ;
  assign n40160 = n10955 | n40159 ;
  assign n40161 = n9378 ^ n5311 ^ 1'b0 ;
  assign n40162 = n38387 & n40161 ;
  assign n40163 = n5461 & ~n10957 ;
  assign n40164 = ~n3329 & n18941 ;
  assign n40165 = n21612 ^ n12028 ^ 1'b0 ;
  assign n40166 = ~n1192 & n40165 ;
  assign n40167 = n40166 ^ n20267 ^ 1'b0 ;
  assign n40168 = n32755 ^ n18388 ^ 1'b0 ;
  assign n40171 = n8038 & n20047 ;
  assign n40169 = n7648 ^ n3514 ^ 1'b0 ;
  assign n40170 = n16708 & ~n40169 ;
  assign n40172 = n40171 ^ n40170 ^ 1'b0 ;
  assign n40173 = n12074 ^ n896 ^ 1'b0 ;
  assign n40174 = n16956 & ~n40173 ;
  assign n40175 = n40174 ^ n6243 ^ 1'b0 ;
  assign n40176 = n13557 | n40175 ;
  assign n40177 = n40176 ^ n946 ^ 1'b0 ;
  assign n40178 = n3367 & n40177 ;
  assign n40179 = n40178 ^ n12480 ^ 1'b0 ;
  assign n40180 = ~n4920 & n40179 ;
  assign n40181 = n2544 & ~n13807 ;
  assign n40182 = n40181 ^ n8831 ^ 1'b0 ;
  assign n40183 = n20108 & n36413 ;
  assign n40184 = n14829 ^ n9262 ^ 1'b0 ;
  assign n40185 = ~n3777 & n18326 ;
  assign n40186 = n5051 & n40185 ;
  assign n40187 = n9816 ^ n2178 ^ 1'b0 ;
  assign n40188 = n40186 | n40187 ;
  assign n40189 = n40188 ^ n21373 ^ 1'b0 ;
  assign n40190 = n34404 ^ n17107 ^ 1'b0 ;
  assign n40191 = n22973 & ~n40190 ;
  assign n40192 = n12491 ^ n2570 ^ 1'b0 ;
  assign n40193 = n15320 & ~n32028 ;
  assign n40194 = ~n40192 & n40193 ;
  assign n40195 = ~n17122 & n34392 ;
  assign n40196 = ~n13649 & n40195 ;
  assign n40197 = ~n11756 & n16953 ;
  assign n40198 = n957 | n20251 ;
  assign n40199 = n23202 ^ n16877 ^ n14840 ;
  assign n40200 = n3032 & n14017 ;
  assign n40201 = n25180 ^ n18580 ^ 1'b0 ;
  assign n40202 = n1662 & ~n10584 ;
  assign n40203 = n36275 & n40202 ;
  assign n40204 = n23236 ^ n20631 ^ 1'b0 ;
  assign n40205 = n32180 & n40204 ;
  assign n40206 = n15970 ^ n638 ^ 1'b0 ;
  assign n40207 = n375 & ~n28598 ;
  assign n40208 = n40207 ^ n36297 ^ 1'b0 ;
  assign n40209 = n38677 | n40208 ;
  assign n40210 = ~n4770 & n12319 ;
  assign n40211 = n1585 & ~n40210 ;
  assign n40212 = ~n22803 & n40211 ;
  assign n40213 = n3044 & n40212 ;
  assign n40214 = n23996 ^ n11128 ^ 1'b0 ;
  assign n40215 = ~n21285 & n40214 ;
  assign n40216 = n38799 & n40215 ;
  assign n40217 = n40216 ^ n432 ^ 1'b0 ;
  assign n40218 = n13497 | n16939 ;
  assign n40219 = n28629 ^ n26524 ^ 1'b0 ;
  assign n40220 = n40218 & ~n40219 ;
  assign n40221 = n27574 ^ n4876 ^ n4192 ;
  assign n40222 = n8363 ^ n5420 ^ 1'b0 ;
  assign n40223 = n2961 & ~n8473 ;
  assign n40224 = ~n6415 & n40223 ;
  assign n40225 = ( n6851 & ~n19155 ) | ( n6851 & n24317 ) | ( ~n19155 & n24317 ) ;
  assign n40226 = n15059 ^ n13309 ^ 1'b0 ;
  assign n40227 = n4649 | n40226 ;
  assign n40228 = n3855 & n14787 ;
  assign n40229 = ( ~n10611 & n40227 ) | ( ~n10611 & n40228 ) | ( n40227 & n40228 ) ;
  assign n40230 = n35755 ^ n7702 ^ 1'b0 ;
  assign n40231 = n6164 | n18776 ;
  assign n40232 = n23355 | n40231 ;
  assign n40233 = n3564 & ~n37168 ;
  assign n40234 = n40233 ^ n10502 ^ 1'b0 ;
  assign n40235 = n18145 ^ n15790 ^ 1'b0 ;
  assign n40236 = ~n18928 & n40235 ;
  assign n40237 = n4190 | n33247 ;
  assign n40238 = n40236 | n40237 ;
  assign n40239 = n2925 | n10445 ;
  assign n40240 = n35547 | n40239 ;
  assign n40241 = n40240 ^ n40178 ^ 1'b0 ;
  assign n40244 = ( ~n3329 & n9495 ) | ( ~n3329 & n20871 ) | ( n9495 & n20871 ) ;
  assign n40242 = n6121 & n22033 ;
  assign n40243 = n40242 ^ n19416 ^ n16805 ;
  assign n40245 = n40244 ^ n40243 ^ n12740 ;
  assign n40246 = ( ~n11883 & n18338 ) | ( ~n11883 & n32142 ) | ( n18338 & n32142 ) ;
  assign n40247 = x231 & n27800 ;
  assign n40248 = ( n1593 & n8072 ) | ( n1593 & ~n9801 ) | ( n8072 & ~n9801 ) ;
  assign n40249 = n835 & ~n40248 ;
  assign n40250 = n21037 & ~n29545 ;
  assign n40251 = n40249 & n40250 ;
  assign n40254 = ~n4462 & n24898 ;
  assign n40252 = n14538 | n27870 ;
  assign n40253 = n7831 & n40252 ;
  assign n40255 = n40254 ^ n40253 ^ 1'b0 ;
  assign n40256 = n20616 ^ n8654 ^ 1'b0 ;
  assign n40257 = n3972 | n40256 ;
  assign n40258 = n16559 | n40257 ;
  assign n40259 = n40255 & n40258 ;
  assign n40260 = n21496 ^ n8739 ^ 1'b0 ;
  assign n40261 = n9146 | n40260 ;
  assign n40262 = n7828 & ~n34814 ;
  assign n40263 = n22228 & n40262 ;
  assign n40264 = n17341 ^ n4323 ^ 1'b0 ;
  assign n40265 = n27958 & n35280 ;
  assign n40266 = n40265 ^ n21291 ^ 1'b0 ;
  assign n40267 = n10014 ^ n2202 ^ 1'b0 ;
  assign n40268 = n6751 ^ n1284 ^ 1'b0 ;
  assign n40269 = n8963 & ~n40268 ;
  assign n40270 = n40269 ^ n14749 ^ 1'b0 ;
  assign n40271 = n19138 & ~n40270 ;
  assign n40272 = n3912 | n12940 ;
  assign n40273 = n40272 ^ n21198 ^ 1'b0 ;
  assign n40274 = n11017 & n40273 ;
  assign n40275 = ~n8105 & n40274 ;
  assign n40276 = n5490 & n5668 ;
  assign n40277 = n40275 & n40276 ;
  assign n40280 = n1369 & n6131 ;
  assign n40281 = n16569 & ~n18181 ;
  assign n40282 = ~n40280 & n40281 ;
  assign n40278 = n4345 & ~n27763 ;
  assign n40279 = ~x154 & n40278 ;
  assign n40283 = n40282 ^ n40279 ^ 1'b0 ;
  assign n40284 = n14872 ^ n5379 ^ 1'b0 ;
  assign n40285 = n11762 & n40284 ;
  assign n40286 = n40285 ^ n15137 ^ 1'b0 ;
  assign n40287 = ~n31282 & n40286 ;
  assign n40288 = n20834 ^ n13084 ^ 1'b0 ;
  assign n40289 = ~n33931 & n40288 ;
  assign n40290 = n40289 ^ n24276 ^ n19356 ;
  assign n40291 = n40135 ^ x73 ^ 1'b0 ;
  assign n40292 = ~n20014 & n40291 ;
  assign n40293 = n18310 ^ n2963 ^ 1'b0 ;
  assign n40294 = n40292 & ~n40293 ;
  assign n40295 = n20249 | n24825 ;
  assign n40296 = n8125 & ~n40295 ;
  assign n40297 = n33326 ^ n11725 ^ 1'b0 ;
  assign n40298 = n6974 | n24399 ;
  assign n40299 = n29243 | n40298 ;
  assign n40301 = ~n3022 & n14586 ;
  assign n40302 = n40301 ^ x25 ^ 1'b0 ;
  assign n40300 = n25287 ^ x194 ^ 1'b0 ;
  assign n40303 = n40302 ^ n40300 ^ n11231 ;
  assign n40309 = n5651 & n21795 ;
  assign n40310 = ~n9684 & n40309 ;
  assign n40304 = ~n6140 & n25789 ;
  assign n40305 = n27116 & ~n40304 ;
  assign n40306 = n40305 ^ n21254 ^ 1'b0 ;
  assign n40307 = ~n15506 & n40306 ;
  assign n40308 = ~n14067 & n40307 ;
  assign n40311 = n40310 ^ n40308 ^ 1'b0 ;
  assign n40312 = n1495 ^ n467 ^ 1'b0 ;
  assign n40313 = n3722 | n32269 ;
  assign n40314 = n40313 ^ n6430 ^ n4867 ;
  assign n40315 = n40314 ^ n31491 ^ 1'b0 ;
  assign n40316 = n12998 | n16532 ;
  assign n40317 = n16095 & ~n38398 ;
  assign n40318 = ~n3309 & n40317 ;
  assign n40319 = n828 | n4200 ;
  assign n40320 = n23506 & ~n40319 ;
  assign n40321 = n15290 & ~n36153 ;
  assign n40322 = n28472 ^ n28320 ^ n1856 ;
  assign n40323 = n19162 ^ n9814 ^ 1'b0 ;
  assign n40324 = ~n17279 & n28127 ;
  assign n40325 = n40324 ^ n3845 ^ 1'b0 ;
  assign n40326 = n33528 & ~n39800 ;
  assign n40327 = n15609 ^ n3099 ^ 1'b0 ;
  assign n40328 = n12168 & n19046 ;
  assign n40329 = n6834 & n29055 ;
  assign n40330 = ~n8276 & n40329 ;
  assign n40331 = x190 & ~n1503 ;
  assign n40332 = n40331 ^ n4086 ^ 1'b0 ;
  assign n40333 = ~n33008 & n40082 ;
  assign n40334 = ~n5596 & n40333 ;
  assign n40335 = n4532 & ~n8529 ;
  assign n40336 = n40335 ^ n2082 ^ 1'b0 ;
  assign n40337 = n20930 ^ n9438 ^ 1'b0 ;
  assign n40338 = ~n12288 & n40337 ;
  assign n40339 = ~n5619 & n13524 ;
  assign n40340 = ~n40338 & n40339 ;
  assign n40341 = n2725 & n5508 ;
  assign n40342 = ( n2154 & n31236 ) | ( n2154 & n40341 ) | ( n31236 & n40341 ) ;
  assign n40343 = ~n1750 & n8809 ;
  assign n40344 = n12831 & n31136 ;
  assign n40345 = n40344 ^ n10628 ^ 1'b0 ;
  assign n40346 = ( n1627 & n3496 ) | ( n1627 & n18713 ) | ( n3496 & n18713 ) ;
  assign n40347 = n40346 ^ n29712 ^ 1'b0 ;
  assign n40348 = n40347 ^ n2291 ^ 1'b0 ;
  assign n40349 = n2715 | n16358 ;
  assign n40350 = ~n1081 & n16424 ;
  assign n40351 = n40350 ^ n21655 ^ 1'b0 ;
  assign n40352 = ~n9362 & n40351 ;
  assign n40358 = n7237 & n8430 ;
  assign n40354 = n8009 & n25107 ;
  assign n40355 = n40354 ^ n8603 ^ 1'b0 ;
  assign n40356 = ( n5423 & n8829 ) | ( n5423 & n40355 ) | ( n8829 & n40355 ) ;
  assign n40357 = n40356 ^ n11462 ^ 1'b0 ;
  assign n40353 = ~n29517 & n32620 ;
  assign n40359 = n40358 ^ n40357 ^ n40353 ;
  assign n40361 = n20807 ^ n12794 ^ n1361 ;
  assign n40360 = n2184 | n19813 ;
  assign n40362 = n40361 ^ n40360 ^ 1'b0 ;
  assign n40363 = n40362 ^ n29326 ^ n13254 ;
  assign n40364 = n21752 ^ n14174 ^ 1'b0 ;
  assign n40365 = n4585 | n36198 ;
  assign n40366 = n4824 & n4911 ;
  assign n40367 = n40366 ^ n2248 ^ 1'b0 ;
  assign n40368 = n40367 ^ n11891 ^ 1'b0 ;
  assign n40369 = n5293 & ~n40368 ;
  assign n40370 = n15707 | n28248 ;
  assign n40371 = ~n7150 & n12873 ;
  assign n40372 = n40371 ^ n7773 ^ 1'b0 ;
  assign n40374 = ( n1338 & n3151 ) | ( n1338 & n14582 ) | ( n3151 & n14582 ) ;
  assign n40373 = ~n3210 & n7149 ;
  assign n40375 = n40374 ^ n40373 ^ 1'b0 ;
  assign n40376 = n2774 & n9416 ;
  assign n40377 = n40376 ^ n8396 ^ 1'b0 ;
  assign n40378 = n29187 & ~n34237 ;
  assign n40379 = ~n40377 & n40378 ;
  assign n40380 = n7149 & n40379 ;
  assign n40381 = ( n1968 & n6405 ) | ( n1968 & n11492 ) | ( n6405 & n11492 ) ;
  assign n40382 = n2137 | n22064 ;
  assign n40383 = n2219 | n40382 ;
  assign n40384 = n40383 ^ n17541 ^ 1'b0 ;
  assign n40385 = n15492 & ~n40384 ;
  assign n40386 = n2013 & n40385 ;
  assign n40387 = n1952 & ~n22935 ;
  assign n40388 = n15653 & n17244 ;
  assign n40389 = n11626 & ~n40388 ;
  assign n40390 = n2959 & ~n3054 ;
  assign n40391 = ~n9175 & n40390 ;
  assign n40392 = n39465 ^ n13580 ^ 1'b0 ;
  assign n40393 = n31805 & n40392 ;
  assign n40394 = n40393 ^ n37904 ^ 1'b0 ;
  assign n40395 = ( x253 & n14895 ) | ( x253 & n18248 ) | ( n14895 & n18248 ) ;
  assign n40396 = n40395 ^ n16439 ^ 1'b0 ;
  assign n40397 = n2097 | n16421 ;
  assign n40398 = ( ~n1854 & n12733 ) | ( ~n1854 & n40397 ) | ( n12733 & n40397 ) ;
  assign n40399 = n40398 ^ n27946 ^ 1'b0 ;
  assign n40400 = ~n14781 & n40399 ;
  assign n40404 = n28597 ^ n4712 ^ n3861 ;
  assign n40401 = n19837 ^ n4686 ^ 1'b0 ;
  assign n40402 = n28527 & n40401 ;
  assign n40403 = n40402 ^ n29420 ^ 1'b0 ;
  assign n40405 = n40404 ^ n40403 ^ 1'b0 ;
  assign n40406 = n5308 & n40405 ;
  assign n40407 = ~n10364 & n25109 ;
  assign n40408 = n15260 & n40407 ;
  assign n40409 = n11344 ^ n5642 ^ 1'b0 ;
  assign n40410 = ~n18246 & n40409 ;
  assign n40411 = n2349 | n10272 ;
  assign n40412 = n11838 ^ n4927 ^ 1'b0 ;
  assign n40413 = n2297 | n40412 ;
  assign n40414 = ~n13647 & n16128 ;
  assign n40415 = n40414 ^ n28661 ^ 1'b0 ;
  assign n40416 = n9659 & n21177 ;
  assign n40417 = n16674 & n40416 ;
  assign n40418 = n40417 ^ n17672 ^ 1'b0 ;
  assign n40419 = n36029 ^ n1008 ^ 1'b0 ;
  assign n40420 = n2362 & n40419 ;
  assign n40421 = ( n12584 & ~n12804 ) | ( n12584 & n40420 ) | ( ~n12804 & n40420 ) ;
  assign n40422 = n3819 | n6977 ;
  assign n40423 = n2203 | n15989 ;
  assign n40424 = n40423 ^ n3699 ^ 1'b0 ;
  assign n40425 = n40424 ^ n24632 ^ 1'b0 ;
  assign n40426 = n7349 & ~n40425 ;
  assign n40427 = n3678 & ~n13267 ;
  assign n40428 = n39549 ^ n28574 ^ 1'b0 ;
  assign n40429 = n9985 & ~n40428 ;
  assign n40430 = ~n40427 & n40429 ;
  assign n40431 = n33739 ^ n13940 ^ 1'b0 ;
  assign n40432 = n6250 & ~n40431 ;
  assign n40433 = ~n4933 & n40432 ;
  assign n40434 = ~n8923 & n33667 ;
  assign n40435 = n40433 & n40434 ;
  assign n40439 = n5250 | n19534 ;
  assign n40436 = n9140 | n16346 ;
  assign n40437 = n1244 | n40436 ;
  assign n40438 = n40437 ^ n33027 ^ 1'b0 ;
  assign n40440 = n40439 ^ n40438 ^ n39938 ;
  assign n40441 = ( n20291 & ~n34195 ) | ( n20291 & n38915 ) | ( ~n34195 & n38915 ) ;
  assign n40442 = n32535 & n40441 ;
  assign n40443 = n13318 & ~n31520 ;
  assign n40444 = n3990 & n40443 ;
  assign n40446 = n11542 ^ n815 ^ 1'b0 ;
  assign n40445 = n26501 | n29873 ;
  assign n40447 = n40446 ^ n40445 ^ 1'b0 ;
  assign n40448 = ~n5091 & n32431 ;
  assign n40449 = n12649 ^ n10272 ^ 1'b0 ;
  assign n40450 = n6506 | n21755 ;
  assign n40451 = ~n40449 & n40450 ;
  assign n40452 = ~n23213 & n33191 ;
  assign n40453 = n27695 ^ n2993 ^ 1'b0 ;
  assign n40454 = n21050 & n40453 ;
  assign n40455 = n2576 & n16546 ;
  assign n40456 = n40455 ^ n21382 ^ n2209 ;
  assign n40457 = n5418 & n31818 ;
  assign n40458 = n40457 ^ n27872 ^ 1'b0 ;
  assign n40459 = n6470 & ~n40428 ;
  assign n40460 = n22447 & n40459 ;
  assign n40461 = n40460 ^ n4360 ^ 1'b0 ;
  assign n40462 = n15196 ^ n3739 ^ 1'b0 ;
  assign n40463 = n10928 & n40462 ;
  assign n40464 = n37928 ^ n16987 ^ 1'b0 ;
  assign n40465 = ~n26257 & n31860 ;
  assign n40466 = n14492 & n40465 ;
  assign n40467 = n1048 | n9289 ;
  assign n40468 = ~n13557 & n26393 ;
  assign n40469 = n17700 ^ n15249 ^ 1'b0 ;
  assign n40470 = n4807 ^ x100 ^ 1'b0 ;
  assign n40471 = n40470 ^ n14198 ^ 1'b0 ;
  assign n40476 = n22609 | n31994 ;
  assign n40477 = n40476 ^ n32778 ^ 1'b0 ;
  assign n40472 = n33754 ^ n756 ^ 1'b0 ;
  assign n40473 = n11856 & ~n27494 ;
  assign n40474 = ~n40472 & n40473 ;
  assign n40475 = n1746 & ~n40474 ;
  assign n40478 = n40477 ^ n40475 ^ 1'b0 ;
  assign n40479 = ~n2466 & n2739 ;
  assign n40480 = n14851 & n22015 ;
  assign n40481 = n20578 ^ n14846 ^ n14044 ;
  assign n40482 = n23763 & n40481 ;
  assign n40483 = n3942 & ~n10787 ;
  assign n40484 = n40483 ^ n922 ^ 1'b0 ;
  assign n40485 = n12937 & ~n16388 ;
  assign n40486 = ( n8804 & n14034 ) | ( n8804 & ~n36075 ) | ( n14034 & ~n36075 ) ;
  assign n40487 = n23641 ^ n12493 ^ 1'b0 ;
  assign n40488 = ( ~n30837 & n40486 ) | ( ~n30837 & n40487 ) | ( n40486 & n40487 ) ;
  assign n40489 = n1199 & ~n4200 ;
  assign n40490 = n40489 ^ n20188 ^ 1'b0 ;
  assign n40491 = n8429 & n40490 ;
  assign n40492 = n8782 & ~n21695 ;
  assign n40493 = ~n40491 & n40492 ;
  assign n40494 = n21739 | n40493 ;
  assign n40495 = n40494 ^ n4913 ^ 1'b0 ;
  assign n40496 = n10139 & ~n12217 ;
  assign n40497 = n21755 & n40496 ;
  assign n40498 = ~n40107 & n40497 ;
  assign n40499 = n37284 ^ n8414 ^ 1'b0 ;
  assign n40500 = n40498 & n40499 ;
  assign n40501 = ~n1475 & n8765 ;
  assign n40502 = n40501 ^ n13414 ^ 1'b0 ;
  assign n40503 = ~n40227 & n40502 ;
  assign n40504 = n10684 & n40503 ;
  assign n40505 = n40504 ^ n6294 ^ 1'b0 ;
  assign n40506 = ~n3086 & n17722 ;
  assign n40507 = ~n30409 & n40506 ;
  assign n40508 = ~n9237 & n40507 ;
  assign n40509 = ( n661 & n7513 ) | ( n661 & ~n26125 ) | ( n7513 & ~n26125 ) ;
  assign n40510 = n2493 & n18515 ;
  assign n40511 = ( n3614 & n8425 ) | ( n3614 & ~n40510 ) | ( n8425 & ~n40510 ) ;
  assign n40512 = n7028 | n9104 ;
  assign n40513 = n40512 ^ n3028 ^ 1'b0 ;
  assign n40514 = n40513 ^ n26389 ^ 1'b0 ;
  assign n40515 = n12781 & ~n40514 ;
  assign n40516 = n40515 ^ n38664 ^ 1'b0 ;
  assign n40518 = n5152 & n33331 ;
  assign n40519 = n17910 & n40518 ;
  assign n40517 = ~n1254 & n10880 ;
  assign n40520 = n40519 ^ n40517 ^ 1'b0 ;
  assign n40521 = n6154 | n36075 ;
  assign n40522 = n6730 & n40521 ;
  assign n40523 = n19624 & n22879 ;
  assign n40524 = n7510 & n29716 ;
  assign n40525 = n11734 & n37886 ;
  assign n40526 = n4595 | n6949 ;
  assign n40528 = n14269 ^ n3615 ^ 1'b0 ;
  assign n40527 = ~n496 & n18276 ;
  assign n40529 = n40528 ^ n40527 ^ 1'b0 ;
  assign n40530 = ( n20662 & n36153 ) | ( n20662 & n40529 ) | ( n36153 & n40529 ) ;
  assign n40531 = n14543 & ~n28416 ;
  assign n40532 = n40531 ^ n6479 ^ n1086 ;
  assign n40533 = n22902 | n34454 ;
  assign n40534 = n21018 & ~n26673 ;
  assign n40535 = n40534 ^ n31066 ^ 1'b0 ;
  assign n40536 = n33533 ^ n5722 ^ 1'b0 ;
  assign n40537 = n3994 | n32004 ;
  assign n40538 = n37974 & ~n40537 ;
  assign n40539 = n2643 & n11730 ;
  assign n40540 = ~n7541 & n40539 ;
  assign n40541 = n40540 ^ n28746 ^ 1'b0 ;
  assign n40542 = ~n2458 & n6204 ;
  assign n40543 = n18383 & n40542 ;
  assign n40544 = n40543 ^ n3504 ^ 1'b0 ;
  assign n40545 = n14448 & ~n40544 ;
  assign n40546 = n31716 ^ n30207 ^ 1'b0 ;
  assign n40547 = n32456 & ~n40546 ;
  assign n40548 = n40547 ^ n11895 ^ 1'b0 ;
  assign n40549 = n37101 ^ n11435 ^ 1'b0 ;
  assign n40550 = ( ~n4269 & n8026 ) | ( ~n4269 & n25880 ) | ( n8026 & n25880 ) ;
  assign n40551 = n8941 ^ n3203 ^ 1'b0 ;
  assign n40552 = n40550 | n40551 ;
  assign n40553 = ~n21409 & n40426 ;
  assign n40554 = n40553 ^ n12455 ^ 1'b0 ;
  assign n40555 = n3997 | n13523 ;
  assign n40556 = n32059 & ~n40555 ;
  assign n40557 = n40556 ^ n3312 ^ 1'b0 ;
  assign n40558 = n23703 ^ n7900 ^ 1'b0 ;
  assign n40559 = n34012 & n40558 ;
  assign n40560 = n9068 | n40559 ;
  assign n40561 = n40446 & n40560 ;
  assign n40562 = ( n3313 & n16932 ) | ( n3313 & ~n34518 ) | ( n16932 & ~n34518 ) ;
  assign n40563 = n30176 ^ n18796 ^ 1'b0 ;
  assign n40564 = n26378 ^ n2848 ^ 1'b0 ;
  assign n40565 = n14240 & ~n40564 ;
  assign n40566 = n22897 & n33516 ;
  assign n40567 = ~n40565 & n40566 ;
  assign n40568 = n11981 ^ n5508 ^ 1'b0 ;
  assign n40569 = ~n14346 & n40568 ;
  assign n40570 = n40569 ^ n3712 ^ 1'b0 ;
  assign n40571 = x155 & ~n40570 ;
  assign n40572 = n8024 | n11288 ;
  assign n40573 = ~n10696 & n25635 ;
  assign n40574 = n27101 & n40573 ;
  assign n40575 = ~n23065 & n40574 ;
  assign n40576 = n28176 ^ n9280 ^ 1'b0 ;
  assign n40577 = n31065 ^ n17596 ^ 1'b0 ;
  assign n40578 = n40576 | n40577 ;
  assign n40579 = ~n11531 & n23108 ;
  assign n40580 = n39070 & n40579 ;
  assign n40581 = ~n17045 & n40580 ;
  assign n40582 = ~n8397 & n28137 ;
  assign n40583 = n2097 & n40582 ;
  assign n40584 = n7336 | n40583 ;
  assign n40585 = n28356 & ~n40584 ;
  assign n40586 = ~n11551 & n13077 ;
  assign n40587 = n16313 | n20718 ;
  assign n40588 = n30397 ^ n25518 ^ 1'b0 ;
  assign n40589 = ~n40587 & n40588 ;
  assign n40590 = n20407 ^ n14358 ^ 1'b0 ;
  assign n40591 = ~n980 & n40590 ;
  assign n40592 = n2331 & ~n4675 ;
  assign n40593 = ~n9529 & n40258 ;
  assign n40594 = n40593 ^ n6805 ^ 1'b0 ;
  assign n40595 = ~n32470 & n40594 ;
  assign n40596 = ( n5093 & n12483 ) | ( n5093 & n28304 ) | ( n12483 & n28304 ) ;
  assign n40597 = ( n17228 & n23667 ) | ( n17228 & ~n40497 ) | ( n23667 & ~n40497 ) ;
  assign n40598 = n8163 & ~n12924 ;
  assign n40599 = n21030 ^ n15831 ^ 1'b0 ;
  assign n40600 = n40599 ^ n33669 ^ 1'b0 ;
  assign n40601 = n7319 & n22427 ;
  assign n40602 = n40601 ^ n25921 ^ 1'b0 ;
  assign n40603 = n4972 | n16612 ;
  assign n40604 = n3073 | n40603 ;
  assign n40605 = n2041 & n40604 ;
  assign n40606 = n2951 & n40605 ;
  assign n40607 = n2443 & ~n25517 ;
  assign n40608 = n21356 & n40607 ;
  assign n40609 = n40608 ^ n24132 ^ 1'b0 ;
  assign n40610 = n31109 ^ n4319 ^ 1'b0 ;
  assign n40611 = n1561 ^ n1048 ^ 1'b0 ;
  assign n40612 = n40611 ^ n28273 ^ n9814 ;
  assign n40613 = n1551 | n14715 ;
  assign n40614 = n24005 & ~n40613 ;
  assign n40615 = n21588 ^ n3012 ^ 1'b0 ;
  assign n40616 = n14994 & ~n40615 ;
  assign n40617 = ~n14372 & n37249 ;
  assign n40618 = n23404 & n40617 ;
  assign n40619 = n31090 & n33322 ;
  assign n40620 = n627 | n3389 ;
  assign n40621 = ~n6040 & n34245 ;
  assign n40622 = ~n10637 & n15569 ;
  assign n40623 = n40622 ^ n2408 ^ 1'b0 ;
  assign n40624 = n40623 ^ n20527 ^ n17008 ;
  assign n40625 = n15889 ^ n3874 ^ n483 ;
  assign n40626 = n37799 | n40625 ;
  assign n40627 = n8354 & ~n19550 ;
  assign n40628 = ~n30372 & n40627 ;
  assign n40629 = n1712 & ~n10783 ;
  assign n40630 = n14456 & n40629 ;
  assign n40633 = n38152 ^ n31437 ^ 1'b0 ;
  assign n40634 = n1841 & n40633 ;
  assign n40635 = ~n537 & n40634 ;
  assign n40631 = n6566 ^ n3617 ^ 1'b0 ;
  assign n40632 = n14175 & n40631 ;
  assign n40636 = n40635 ^ n40632 ^ 1'b0 ;
  assign n40637 = n15812 & ~n40098 ;
  assign n40638 = n28899 & n40637 ;
  assign n40639 = n40638 ^ n28433 ^ 1'b0 ;
  assign n40640 = n28143 & ~n40639 ;
  assign n40641 = n32274 ^ n22074 ^ 1'b0 ;
  assign n40642 = n7632 & n13315 ;
  assign n40643 = n40642 ^ n35597 ^ 1'b0 ;
  assign n40644 = n14867 ^ n2883 ^ 1'b0 ;
  assign n40645 = n11633 & n30787 ;
  assign n40646 = n13177 ^ n6687 ^ 1'b0 ;
  assign n40647 = n15292 & n16579 ;
  assign n40648 = ~n16244 & n40647 ;
  assign n40649 = n27444 ^ n1504 ^ 1'b0 ;
  assign n40650 = n11976 | n40649 ;
  assign n40651 = n40650 ^ n14052 ^ 1'b0 ;
  assign n40652 = ~n20705 & n40651 ;
  assign n40653 = n4906 ^ n1378 ^ 1'b0 ;
  assign n40654 = n40652 & n40653 ;
  assign n40655 = n2297 ^ n2055 ^ 1'b0 ;
  assign n40656 = n592 & ~n40655 ;
  assign n40657 = n34499 ^ n15359 ^ n1676 ;
  assign n40658 = n40657 ^ n24204 ^ 1'b0 ;
  assign n40659 = ~n21084 & n40658 ;
  assign n40660 = n9190 & n40659 ;
  assign n40661 = n23235 ^ n21623 ^ 1'b0 ;
  assign n40662 = n33688 & n40661 ;
  assign n40663 = n39603 ^ n11973 ^ n8249 ;
  assign n40664 = ~n2443 & n36826 ;
  assign n40665 = n8114 & ~n12260 ;
  assign n40666 = ~n11373 & n21440 ;
  assign n40667 = ~n492 & n40666 ;
  assign n40668 = ~n2679 & n18345 ;
  assign n40669 = n10408 & n40668 ;
  assign n40670 = n3643 | n11601 ;
  assign n40671 = n40670 ^ x45 ^ 1'b0 ;
  assign n40672 = n40671 ^ n7507 ^ 1'b0 ;
  assign n40673 = n40669 | n40672 ;
  assign n40674 = n10831 & n25211 ;
  assign n40675 = ~n10831 & n40674 ;
  assign n40676 = n12168 | n40675 ;
  assign n40677 = n40676 ^ n13054 ^ 1'b0 ;
  assign n40678 = n13725 & n34501 ;
  assign n40679 = n18252 ^ n2255 ^ 1'b0 ;
  assign n40680 = n15989 & n35737 ;
  assign n40681 = n8112 & n11504 ;
  assign n40682 = n40681 ^ n10698 ^ 1'b0 ;
  assign n40683 = n10900 ^ n8927 ^ 1'b0 ;
  assign n40684 = n10771 ^ n8950 ^ 1'b0 ;
  assign n40685 = ~n13617 & n40684 ;
  assign n40686 = n15418 & ~n27108 ;
  assign n40687 = ~n40685 & n40686 ;
  assign n40688 = n38508 ^ n6834 ^ 1'b0 ;
  assign n40689 = ~n3034 & n6639 ;
  assign n40690 = n19628 & ~n40689 ;
  assign n40691 = n1170 & ~n18371 ;
  assign n40692 = n3994 & ~n10737 ;
  assign n40693 = n40691 & n40692 ;
  assign n40694 = n13418 ^ n7663 ^ 1'b0 ;
  assign n40695 = n40693 | n40694 ;
  assign n40696 = ( n4964 & ~n23565 ) | ( n4964 & n40695 ) | ( ~n23565 & n40695 ) ;
  assign n40697 = n40696 ^ n31530 ^ 1'b0 ;
  assign n40698 = n649 | n40697 ;
  assign n40699 = n16348 ^ n4372 ^ 1'b0 ;
  assign n40700 = n21451 & n40699 ;
  assign n40701 = n19706 & ~n33857 ;
  assign n40702 = n20503 & n40701 ;
  assign n40703 = n25921 | n28096 ;
  assign n40704 = n2741 & ~n25151 ;
  assign n40705 = ( n1257 & n3397 ) | ( n1257 & n12238 ) | ( n3397 & n12238 ) ;
  assign n40706 = n11920 | n40705 ;
  assign n40707 = n22636 | n40706 ;
  assign n40708 = ( n4551 & n6373 ) | ( n4551 & ~n17278 ) | ( n6373 & ~n17278 ) ;
  assign n40709 = n40708 ^ n7624 ^ 1'b0 ;
  assign n40710 = ~n26168 & n40709 ;
  assign n40711 = n8336 & n12314 ;
  assign n40712 = n15579 ^ n4325 ^ 1'b0 ;
  assign n40713 = n40712 ^ n31431 ^ n3164 ;
  assign n40714 = n40711 & n40713 ;
  assign n40715 = ( n5560 & n31734 ) | ( n5560 & ~n36594 ) | ( n31734 & ~n36594 ) ;
  assign n40716 = n3939 & n4925 ;
  assign n40717 = ~n7600 & n28014 ;
  assign n40718 = n40717 ^ n11707 ^ 1'b0 ;
  assign n40719 = n900 & n35582 ;
  assign n40720 = n8185 & n40719 ;
  assign n40721 = n9619 & n24004 ;
  assign n40722 = n40721 ^ n1459 ^ 1'b0 ;
  assign n40723 = ( n11534 & n19881 ) | ( n11534 & ~n28893 ) | ( n19881 & ~n28893 ) ;
  assign n40724 = n15089 ^ n8499 ^ 1'b0 ;
  assign n40725 = n17874 & n24749 ;
  assign n40726 = ~n6987 & n9957 ;
  assign n40728 = n25725 ^ n15010 ^ 1'b0 ;
  assign n40729 = n31580 ^ n7312 ^ 1'b0 ;
  assign n40730 = ~n40728 & n40729 ;
  assign n40727 = n708 & n5237 ;
  assign n40731 = n40730 ^ n40727 ^ 1'b0 ;
  assign n40732 = n3805 | n17000 ;
  assign n40733 = n36024 ^ n33713 ^ 1'b0 ;
  assign n40734 = n32791 | n40733 ;
  assign n40735 = n14752 ^ n13919 ^ 1'b0 ;
  assign n40736 = n18661 | n40735 ;
  assign n40737 = n38430 ^ n6163 ^ 1'b0 ;
  assign n40738 = n40736 & n40737 ;
  assign n40739 = ( n15692 & n25472 ) | ( n15692 & n30228 ) | ( n25472 & n30228 ) ;
  assign n40740 = n29845 ^ n938 ^ 1'b0 ;
  assign n40741 = n40739 | n40740 ;
  assign n40742 = n19979 ^ n9935 ^ 1'b0 ;
  assign n40743 = n26056 & ~n40742 ;
  assign n40744 = n40743 ^ n1599 ^ 1'b0 ;
  assign n40745 = n3311 & ~n21739 ;
  assign n40746 = n23943 & n26968 ;
  assign n40747 = n643 & ~n19877 ;
  assign n40748 = n26393 & n32753 ;
  assign n40749 = n40748 ^ n12160 ^ 1'b0 ;
  assign n40750 = n27353 | n36955 ;
  assign n40752 = n31153 ^ n6184 ^ 1'b0 ;
  assign n40751 = n21320 & n40184 ;
  assign n40753 = n40752 ^ n40751 ^ 1'b0 ;
  assign n40754 = n38203 ^ n12123 ^ n5404 ;
  assign n40756 = n8495 & ~n15936 ;
  assign n40757 = ~n34727 & n40756 ;
  assign n40755 = n18453 | n22131 ;
  assign n40758 = n40757 ^ n40755 ^ 1'b0 ;
  assign n40759 = ~n16370 & n21220 ;
  assign n40760 = ~n2964 & n40759 ;
  assign n40761 = ~n5927 & n6531 ;
  assign n40762 = n40761 ^ n875 ^ 1'b0 ;
  assign n40763 = n12836 ^ n11659 ^ 1'b0 ;
  assign n40764 = ~n5151 & n40763 ;
  assign n40765 = n40764 ^ n11760 ^ 1'b0 ;
  assign n40766 = n18205 & ~n23238 ;
  assign n40767 = n40766 ^ n3884 ^ 1'b0 ;
  assign n40768 = n7810 | n13672 ;
  assign n40769 = n7620 | n40768 ;
  assign n40770 = n24601 ^ n15252 ^ n1782 ;
  assign n40771 = n40770 ^ n8440 ^ 1'b0 ;
  assign n40772 = n293 & n24508 ;
  assign n40773 = n2951 & n40772 ;
  assign n40774 = n29764 ^ n1101 ^ 1'b0 ;
  assign n40775 = n7711 & ~n39214 ;
  assign n40776 = ~n39230 & n40775 ;
  assign n40777 = n22077 & ~n40776 ;
  assign n40778 = ~n31010 & n40777 ;
  assign n40779 = n28330 ^ n23976 ^ 1'b0 ;
  assign n40780 = n7143 & ~n14617 ;
  assign n40781 = n291 & n40780 ;
  assign n40782 = n40781 ^ n15018 ^ 1'b0 ;
  assign n40783 = n18465 | n40782 ;
  assign n40784 = n40783 ^ n28129 ^ 1'b0 ;
  assign n40785 = n27862 ^ n10396 ^ 1'b0 ;
  assign n40786 = n25724 ^ n7231 ^ 1'b0 ;
  assign n40787 = ~n40785 & n40786 ;
  assign n40788 = n1680 | n4741 ;
  assign n40789 = n1680 & ~n40788 ;
  assign n40790 = n40789 ^ n15181 ^ n9931 ;
  assign n40791 = n29619 & ~n40790 ;
  assign n40792 = n40791 ^ n13972 ^ 1'b0 ;
  assign n40793 = n9590 & n40792 ;
  assign n40794 = ( n8026 & n39304 ) | ( n8026 & n40793 ) | ( n39304 & n40793 ) ;
  assign n40795 = n12247 | n32249 ;
  assign n40796 = n21315 ^ n12653 ^ 1'b0 ;
  assign n40797 = ~n1125 & n6413 ;
  assign n40798 = n40797 ^ n1463 ^ 1'b0 ;
  assign n40799 = n23671 | n31584 ;
  assign n40800 = n40799 ^ n27201 ^ 1'b0 ;
  assign n40801 = n21682 ^ n809 ^ 1'b0 ;
  assign n40802 = n11683 | n40801 ;
  assign n40803 = n7143 & n17843 ;
  assign n40804 = n39013 ^ x152 ^ 1'b0 ;
  assign n40805 = n7149 ^ n440 ^ 1'b0 ;
  assign n40806 = n40805 ^ n18875 ^ n17663 ;
  assign n40807 = n30050 ^ n20772 ^ 1'b0 ;
  assign n40808 = ~n4218 & n40807 ;
  assign n40809 = n40808 ^ n22759 ^ n6226 ;
  assign n40810 = n3588 & ~n16980 ;
  assign n40811 = n19365 & n40810 ;
  assign n40812 = n35810 ^ n26521 ^ 1'b0 ;
  assign n40813 = n17067 & ~n27712 ;
  assign n40814 = n16853 ^ n9353 ^ 1'b0 ;
  assign n40815 = ~n30328 & n40814 ;
  assign n40816 = n40815 ^ n16834 ^ 1'b0 ;
  assign n40817 = n40816 ^ n10829 ^ 1'b0 ;
  assign n40818 = n27045 | n40817 ;
  assign n40819 = n8842 & ~n15729 ;
  assign n40820 = n40819 ^ n38602 ^ 1'b0 ;
  assign n40821 = n14958 ^ n5087 ^ n359 ;
  assign n40822 = n33006 ^ n13327 ^ 1'b0 ;
  assign n40823 = ( n7200 & n40821 ) | ( n7200 & ~n40822 ) | ( n40821 & ~n40822 ) ;
  assign n40824 = n6066 | n24513 ;
  assign n40825 = n38872 ^ n12991 ^ 1'b0 ;
  assign n40826 = n27038 ^ n21406 ^ n12576 ;
  assign n40830 = n16150 | n17293 ;
  assign n40831 = n8332 & ~n19071 ;
  assign n40832 = ~n40830 & n40831 ;
  assign n40833 = n11943 | n40832 ;
  assign n40828 = n1449 | n17005 ;
  assign n40829 = n40828 ^ n16042 ^ 1'b0 ;
  assign n40827 = n39053 ^ n19769 ^ 1'b0 ;
  assign n40834 = n40833 ^ n40829 ^ n40827 ;
  assign n40835 = n11601 ^ n7632 ^ n3956 ;
  assign n40836 = n40835 ^ n858 ^ 1'b0 ;
  assign n40837 = n21973 & ~n40836 ;
  assign n40838 = ~n25326 & n40837 ;
  assign n40839 = n7810 ^ n5890 ^ 1'b0 ;
  assign n40840 = n7714 | n40839 ;
  assign n40841 = n16612 ^ n2741 ^ 1'b0 ;
  assign n40842 = n10028 & ~n10284 ;
  assign n40844 = n8529 ^ n4997 ^ 1'b0 ;
  assign n40845 = ~n10942 & n40844 ;
  assign n40843 = n22984 | n31697 ;
  assign n40846 = n40845 ^ n40843 ^ 1'b0 ;
  assign n40847 = n7196 ^ n1667 ^ 1'b0 ;
  assign n40848 = n15070 & ~n40847 ;
  assign n40849 = n13121 ^ n7476 ^ 1'b0 ;
  assign n40852 = n459 & ~n1613 ;
  assign n40853 = ~n7624 & n40852 ;
  assign n40850 = n8620 | n15953 ;
  assign n40851 = n40850 ^ n27382 ^ 1'b0 ;
  assign n40854 = n40853 ^ n40851 ^ n13432 ;
  assign n40855 = n12269 ^ n6233 ^ 1'b0 ;
  assign n40856 = n23247 & n40855 ;
  assign n40857 = ~n34094 & n40856 ;
  assign n40858 = n4508 & n7323 ;
  assign n40859 = ~n7654 & n21860 ;
  assign n40860 = n40859 ^ n28223 ^ 1'b0 ;
  assign n40861 = n11028 ^ n1671 ^ 1'b0 ;
  assign n40862 = ~n17397 & n40861 ;
  assign n40863 = n40860 & n40862 ;
  assign n40864 = n27953 | n39725 ;
  assign n40865 = n631 & n9622 ;
  assign n40868 = n9024 & n34335 ;
  assign n40866 = n1730 & n26238 ;
  assign n40867 = n40866 ^ n10148 ^ 1'b0 ;
  assign n40869 = n40868 ^ n40867 ^ 1'b0 ;
  assign n40870 = ( n3485 & n12632 ) | ( n3485 & ~n27427 ) | ( n12632 & ~n27427 ) ;
  assign n40871 = n1261 & n24554 ;
  assign n40872 = n5571 ^ n4456 ^ 1'b0 ;
  assign n40873 = ~n3885 & n11503 ;
  assign n40874 = ( n6931 & ~n9218 ) | ( n6931 & n33931 ) | ( ~n9218 & n33931 ) ;
  assign n40875 = n3168 & n24936 ;
  assign n40876 = n4747 & ~n40875 ;
  assign n40877 = n40874 & n40876 ;
  assign n40878 = ( ~n13424 & n22156 ) | ( ~n13424 & n34483 ) | ( n22156 & n34483 ) ;
  assign n40879 = n8322 & ~n12667 ;
  assign n40880 = n40879 ^ n8667 ^ 1'b0 ;
  assign n40881 = n8426 | n40880 ;
  assign n40882 = n6990 ^ x20 ^ 1'b0 ;
  assign n40883 = n34221 ^ n16926 ^ 1'b0 ;
  assign n40884 = n2559 | n12225 ;
  assign n40885 = ~n6510 & n11792 ;
  assign n40886 = n40885 ^ n8762 ^ 1'b0 ;
  assign n40887 = n40886 ^ n31700 ^ 1'b0 ;
  assign n40888 = n26644 ^ n4844 ^ 1'b0 ;
  assign n40889 = n24410 ^ n9256 ^ 1'b0 ;
  assign n40890 = x132 & n24241 ;
  assign n40891 = n6177 & n16609 ;
  assign n40892 = n40891 ^ n25344 ^ n7344 ;
  assign n40894 = n613 & n6023 ;
  assign n40895 = n16753 & n40894 ;
  assign n40896 = n13585 & ~n40895 ;
  assign n40897 = n40896 ^ n10401 ^ 1'b0 ;
  assign n40893 = n12526 & n14353 ;
  assign n40898 = n40897 ^ n40893 ^ 1'b0 ;
  assign n40899 = n3114 | n30837 ;
  assign n40900 = n26143 ^ n22658 ^ 1'b0 ;
  assign n40901 = n31308 ^ n15655 ^ 1'b0 ;
  assign n40902 = n13222 ^ n3529 ^ 1'b0 ;
  assign n40903 = n37968 ^ n19602 ^ 1'b0 ;
  assign n40904 = n40902 & n40903 ;
  assign n40905 = n30401 ^ n11973 ^ 1'b0 ;
  assign n40906 = n30653 | n40905 ;
  assign n40907 = n16508 ^ n14532 ^ 1'b0 ;
  assign n40909 = n11655 ^ x53 ^ 1'b0 ;
  assign n40908 = n10225 & n23322 ;
  assign n40910 = n40909 ^ n40908 ^ 1'b0 ;
  assign n40911 = n40910 ^ n7568 ^ 1'b0 ;
  assign n40912 = n40907 & n40911 ;
  assign n40913 = n710 ^ n426 ^ 1'b0 ;
  assign n40914 = n12123 | n40913 ;
  assign n40915 = n17529 & ~n19561 ;
  assign n40916 = ~n10627 & n40915 ;
  assign n40917 = n40916 ^ n26183 ^ n6075 ;
  assign n40918 = n39338 ^ n7974 ^ 1'b0 ;
  assign n40919 = n27173 ^ n4509 ^ 1'b0 ;
  assign n40920 = n15752 | n26230 ;
  assign n40921 = n40920 ^ n16615 ^ 1'b0 ;
  assign n40922 = n23111 ^ n3558 ^ 1'b0 ;
  assign n40923 = n14603 & n40922 ;
  assign n40924 = ( ~n27003 & n33096 ) | ( ~n27003 & n40923 ) | ( n33096 & n40923 ) ;
  assign n40925 = n31894 ^ n19527 ^ 1'b0 ;
  assign n40926 = n24399 | n40925 ;
  assign n40927 = n1748 & ~n40926 ;
  assign n40928 = ~n40924 & n40927 ;
  assign n40930 = n6160 & ~n17970 ;
  assign n40929 = n12339 | n24426 ;
  assign n40931 = n40930 ^ n40929 ^ 1'b0 ;
  assign n40932 = n5870 & n6152 ;
  assign n40933 = n40932 ^ n17614 ^ 1'b0 ;
  assign n40934 = n32833 | n40933 ;
  assign n40935 = n6987 ^ n5802 ^ n4555 ;
  assign n40936 = n17954 & n24007 ;
  assign n40937 = n40936 ^ n14099 ^ 1'b0 ;
  assign n40938 = ~n15279 & n40671 ;
  assign n40939 = n40938 ^ n653 ^ 1'b0 ;
  assign n40940 = n9314 & ~n9586 ;
  assign n40941 = n29428 | n40940 ;
  assign n40942 = ~n34625 & n37910 ;
  assign n40943 = n23662 ^ n18660 ^ n1439 ;
  assign n40944 = n40943 ^ n14598 ^ 1'b0 ;
  assign n40945 = n6916 ^ n3425 ^ n1138 ;
  assign n40946 = n14150 & ~n40923 ;
  assign n40947 = ~n21797 & n29808 ;
  assign n40948 = ~n8546 & n32948 ;
  assign n40949 = n40948 ^ n35887 ^ 1'b0 ;
  assign n40950 = n7283 ^ n6553 ^ 1'b0 ;
  assign n40951 = n40950 ^ n14705 ^ n2502 ;
  assign n40952 = n34004 ^ n21617 ^ n17889 ;
  assign n40953 = ( ~n2501 & n18082 ) | ( ~n2501 & n40952 ) | ( n18082 & n40952 ) ;
  assign n40954 = n5949 ^ n635 ^ 1'b0 ;
  assign n40955 = n26740 ^ n1013 ^ 1'b0 ;
  assign n40956 = n17181 & n40955 ;
  assign n40957 = n26868 & ~n40956 ;
  assign n40958 = ( n5780 & n7242 ) | ( n5780 & n10191 ) | ( n7242 & n10191 ) ;
  assign n40959 = n27405 & n36673 ;
  assign n40960 = n40958 & n40959 ;
  assign n40961 = n15153 ^ n8535 ^ 1'b0 ;
  assign n40962 = n6426 ^ n2116 ^ 1'b0 ;
  assign n40963 = n10983 ^ n1782 ^ n1614 ;
  assign n40964 = ~n11000 & n23455 ;
  assign n40965 = n40964 ^ n5855 ^ 1'b0 ;
  assign n40966 = n40965 ^ n15268 ^ n6844 ;
  assign n40967 = n40384 ^ n17427 ^ 1'b0 ;
  assign n40968 = n6765 & n40967 ;
  assign n40969 = n28381 & ~n40968 ;
  assign n40970 = n16888 | n25459 ;
  assign n40971 = n40970 ^ n19700 ^ 1'b0 ;
  assign n40972 = n10385 & ~n32529 ;
  assign n40973 = n18645 ^ n11453 ^ 1'b0 ;
  assign n40974 = x212 & ~n2464 ;
  assign n40975 = n856 | n40974 ;
  assign n40976 = n7624 ^ n1180 ^ 1'b0 ;
  assign n40977 = n1272 & n11534 ;
  assign n40978 = n16779 ^ n15805 ^ 1'b0 ;
  assign n40979 = n10578 & ~n40978 ;
  assign n40980 = n1667 | n16579 ;
  assign n40981 = n18229 & ~n40980 ;
  assign n40982 = n8424 & ~n17507 ;
  assign n40983 = n40982 ^ n39709 ^ 1'b0 ;
  assign n40984 = n17881 & ~n23972 ;
  assign n40985 = n314 | n5619 ;
  assign n40986 = n12275 | n40985 ;
  assign n40987 = n40984 & ~n40986 ;
  assign n40988 = n20877 ^ n9470 ^ 1'b0 ;
  assign n40989 = n1822 & n12638 ;
  assign n40990 = n1234 & n40989 ;
  assign n40991 = n1758 | n10959 ;
  assign n40992 = n40990 & ~n40991 ;
  assign n40993 = n16866 & ~n31850 ;
  assign n40994 = n7304 ^ n5602 ^ 1'b0 ;
  assign n40995 = n10996 & n16545 ;
  assign n40996 = ~n33529 & n40995 ;
  assign n40997 = ( ~n14805 & n40994 ) | ( ~n14805 & n40996 ) | ( n40994 & n40996 ) ;
  assign n40998 = ~n11901 & n14760 ;
  assign n40999 = n7054 & n11026 ;
  assign n41000 = n40999 ^ n699 ^ 1'b0 ;
  assign n41001 = n41000 ^ n14511 ^ 1'b0 ;
  assign n41002 = ~n675 & n41001 ;
  assign n41003 = ~x213 & n41002 ;
  assign n41004 = n5055 | n41003 ;
  assign n41005 = n15752 | n22128 ;
  assign n41006 = n8714 | n41005 ;
  assign n41007 = n41006 ^ n22451 ^ 1'b0 ;
  assign n41008 = n37128 & n41007 ;
  assign n41009 = ~n15614 & n31036 ;
  assign n41010 = n2477 | n10118 ;
  assign n41011 = n17717 ^ n4473 ^ 1'b0 ;
  assign n41012 = n28123 ^ n14408 ^ 1'b0 ;
  assign n41013 = n41011 & ~n41012 ;
  assign n41014 = n7603 & n39421 ;
  assign n41015 = n41014 ^ n19328 ^ 1'b0 ;
  assign n41016 = ~n5366 & n8336 ;
  assign n41017 = n41016 ^ n24413 ^ 1'b0 ;
  assign n41018 = n41017 ^ n39070 ^ n3866 ;
  assign n41019 = n41018 ^ n40907 ^ n10420 ;
  assign n41020 = n25729 & n31694 ;
  assign n41021 = ~n13449 & n36654 ;
  assign n41022 = n41021 ^ n457 ^ 1'b0 ;
  assign n41023 = n14436 ^ n7920 ^ 1'b0 ;
  assign n41024 = n7959 | n38099 ;
  assign n41025 = n32180 ^ n21057 ^ 1'b0 ;
  assign n41026 = n8273 ^ n1002 ^ 1'b0 ;
  assign n41027 = ~n710 & n41026 ;
  assign n41028 = n36023 & ~n41027 ;
  assign n41029 = n534 & n38306 ;
  assign n41030 = ( ~n9195 & n9912 ) | ( ~n9195 & n19210 ) | ( n9912 & n19210 ) ;
  assign n41031 = ~n11980 & n32057 ;
  assign n41032 = ~n41030 & n41031 ;
  assign n41033 = n6994 & n22310 ;
  assign n41034 = ( ~n2946 & n7532 ) | ( ~n2946 & n29558 ) | ( n7532 & n29558 ) ;
  assign n41035 = n5590 | n27440 ;
  assign n41036 = n4551 | n30103 ;
  assign n41037 = n17994 ^ n7511 ^ 1'b0 ;
  assign n41038 = ~n1932 & n41037 ;
  assign n41039 = n39338 & n41038 ;
  assign n41040 = n18926 ^ n2733 ^ 1'b0 ;
  assign n41041 = n20953 & ~n38436 ;
  assign n41042 = n19346 ^ n5697 ^ 1'b0 ;
  assign n41043 = ~n9930 & n38196 ;
  assign n41044 = n31996 ^ n10039 ^ n1671 ;
  assign n41045 = n6678 ^ n4035 ^ 1'b0 ;
  assign n41046 = n41045 ^ n19719 ^ n5067 ;
  assign n41047 = n5291 ^ x74 ^ 1'b0 ;
  assign n41048 = ~n16327 & n31410 ;
  assign n41049 = ~n6606 & n41048 ;
  assign n41050 = ~n41047 & n41049 ;
  assign n41051 = n36084 ^ n2343 ^ 1'b0 ;
  assign n41052 = ( n18307 & n21790 ) | ( n18307 & ~n23299 ) | ( n21790 & ~n23299 ) ;
  assign n41053 = n19441 ^ n2085 ^ 1'b0 ;
  assign n41054 = ~n41052 & n41053 ;
  assign n41055 = n14815 ^ n1851 ^ 1'b0 ;
  assign n41057 = n15206 ^ n6536 ^ 1'b0 ;
  assign n41058 = n9868 | n16740 ;
  assign n41059 = n41057 | n41058 ;
  assign n41056 = n35833 & ~n39524 ;
  assign n41060 = n41059 ^ n41056 ^ 1'b0 ;
  assign n41061 = n3898 | n28090 ;
  assign n41062 = n41061 ^ n13542 ^ 1'b0 ;
  assign n41063 = n11623 & n41062 ;
  assign n41064 = ~n3750 & n13860 ;
  assign n41065 = n2879 & n7084 ;
  assign n41066 = n12840 ^ n8491 ^ 1'b0 ;
  assign n41067 = n41066 ^ n32379 ^ 1'b0 ;
  assign n41068 = n1859 & n15148 ;
  assign n41069 = n28174 | n41068 ;
  assign n41070 = n21179 ^ n12336 ^ 1'b0 ;
  assign n41071 = n7543 & ~n41070 ;
  assign n41072 = n13409 & n41071 ;
  assign n41073 = n9213 & n41072 ;
  assign n41074 = n6228 & ~n41073 ;
  assign n41075 = ~n16861 & n37396 ;
  assign n41076 = n9538 & n41075 ;
  assign n41077 = n41076 ^ n6533 ^ 1'b0 ;
  assign n41078 = ~n8365 & n28242 ;
  assign n41079 = n41078 ^ n8052 ^ 1'b0 ;
  assign n41080 = n21643 & n38092 ;
  assign n41081 = n36743 ^ n2584 ^ 1'b0 ;
  assign n41082 = ( ~n1997 & n7271 ) | ( ~n1997 & n24973 ) | ( n7271 & n24973 ) ;
  assign n41083 = n4369 & n41082 ;
  assign n41084 = ~n10627 & n41083 ;
  assign n41085 = n31793 | n41084 ;
  assign n41086 = n14971 ^ n4569 ^ 1'b0 ;
  assign n41087 = n5678 | n21790 ;
  assign n41088 = n20220 ^ n7385 ^ 1'b0 ;
  assign n41089 = ~n13449 & n41088 ;
  assign n41090 = n18184 ^ n2249 ^ 1'b0 ;
  assign n41091 = n7150 | n41090 ;
  assign n41092 = n2056 | n41091 ;
  assign n41093 = ( ~n6496 & n19621 ) | ( ~n6496 & n22064 ) | ( n19621 & n22064 ) ;
  assign n41094 = ~n12232 & n39812 ;
  assign n41095 = ~n5339 & n41094 ;
  assign n41096 = n1095 | n11760 ;
  assign n41097 = n41096 ^ n23114 ^ 1'b0 ;
  assign n41098 = n5540 | n41097 ;
  assign n41099 = n22265 & ~n32381 ;
  assign n41100 = n14715 ^ n491 ^ 1'b0 ;
  assign n41101 = ~n9548 & n41100 ;
  assign n41102 = n10445 & ~n35218 ;
  assign n41103 = n22423 | n41102 ;
  assign n41104 = n40730 ^ n7312 ^ 1'b0 ;
  assign n41105 = ~n992 & n3458 ;
  assign n41106 = n992 & n41105 ;
  assign n41107 = n8309 & ~n41106 ;
  assign n41108 = n41106 & n41107 ;
  assign n41109 = n10352 & n41108 ;
  assign n41110 = n8424 & n41109 ;
  assign n41111 = n25985 | n41110 ;
  assign n41112 = n41111 ^ n24934 ^ 1'b0 ;
  assign n41113 = n41112 ^ n11717 ^ n8365 ;
  assign n41114 = n2456 | n36236 ;
  assign n41115 = n37863 ^ n8216 ^ n1712 ;
  assign n41116 = ~n24239 & n41115 ;
  assign n41117 = n8134 | n39056 ;
  assign n41118 = n36319 | n41117 ;
  assign n41119 = n40426 ^ n844 ^ 1'b0 ;
  assign n41120 = n10551 ^ n2263 ^ 1'b0 ;
  assign n41121 = n15574 & n41120 ;
  assign n41122 = n10862 & ~n41121 ;
  assign n41123 = n41122 ^ n14487 ^ 1'b0 ;
  assign n41124 = n26401 & ~n41123 ;
  assign n41125 = ( n2646 & n9260 ) | ( n2646 & n10008 ) | ( n9260 & n10008 ) ;
  assign n41126 = n26200 & ~n41125 ;
  assign n41127 = ( ~n3066 & n17914 ) | ( ~n3066 & n30029 ) | ( n17914 & n30029 ) ;
  assign n41128 = n41127 ^ n1624 ^ 1'b0 ;
  assign n41129 = ~n2272 & n41128 ;
  assign n41130 = n33189 ^ n9043 ^ 1'b0 ;
  assign n41131 = n5849 & ~n36618 ;
  assign n41133 = n25125 ^ n6844 ^ 1'b0 ;
  assign n41132 = n26033 & ~n33347 ;
  assign n41134 = n41133 ^ n41132 ^ 1'b0 ;
  assign n41135 = n25423 ^ n1786 ^ n1149 ;
  assign n41136 = n15239 & ~n41135 ;
  assign n41137 = n41136 ^ n37298 ^ 1'b0 ;
  assign n41138 = n905 & ~n15477 ;
  assign n41139 = ~n9970 & n41138 ;
  assign n41143 = n21262 ^ n10086 ^ 1'b0 ;
  assign n41144 = n7643 & ~n41143 ;
  assign n41140 = ~n4913 & n14196 ;
  assign n41141 = n2320 & n41140 ;
  assign n41142 = ~n34398 & n41141 ;
  assign n41145 = n41144 ^ n41142 ^ 1'b0 ;
  assign n41146 = ~n9993 & n37525 ;
  assign n41147 = n1782 & n41146 ;
  assign n41148 = n8886 & ~n12128 ;
  assign n41149 = n4617 & n41148 ;
  assign n41150 = n22198 & ~n41149 ;
  assign n41151 = n14153 ^ n2831 ^ 1'b0 ;
  assign n41152 = n15314 & n25010 ;
  assign n41153 = n41152 ^ n2781 ^ 1'b0 ;
  assign n41154 = ~n31723 & n41153 ;
  assign n41155 = n2638 & n41154 ;
  assign n41156 = n13630 ^ n13239 ^ 1'b0 ;
  assign n41157 = n32427 | n41156 ;
  assign n41158 = n36758 & ~n41157 ;
  assign n41159 = n4694 | n12947 ;
  assign n41160 = n6121 & ~n14543 ;
  assign n41161 = n41160 ^ n29311 ^ n25530 ;
  assign n41162 = n2286 & ~n4813 ;
  assign n41163 = n41162 ^ n27911 ^ 1'b0 ;
  assign n41164 = n27569 ^ n26161 ^ 1'b0 ;
  assign n41165 = ~n26257 & n34730 ;
  assign n41166 = n35339 & n41165 ;
  assign n41167 = n12728 & n18582 ;
  assign n41168 = n41167 ^ n23523 ^ 1'b0 ;
  assign n41169 = n18692 ^ n12216 ^ 1'b0 ;
  assign n41170 = n2091 & ~n41169 ;
  assign n41171 = ~n20043 & n41170 ;
  assign n41172 = n41171 ^ n38624 ^ 1'b0 ;
  assign n41173 = ~n19284 & n41172 ;
  assign n41174 = n13080 | n15834 ;
  assign n41175 = n17065 | n41174 ;
  assign n41176 = n11292 | n11734 ;
  assign n41177 = n35585 ^ n15840 ^ n2081 ;
  assign n41178 = n41176 & n41177 ;
  assign n41179 = ~n14199 & n19003 ;
  assign n41180 = n1316 & ~n41179 ;
  assign n41181 = n41180 ^ n4834 ^ 1'b0 ;
  assign n41182 = n41181 ^ n38170 ^ n29139 ;
  assign n41183 = n9574 ^ n6412 ^ 1'b0 ;
  assign n41184 = n25569 | n41183 ;
  assign n41185 = n39401 ^ n2774 ^ 1'b0 ;
  assign n41187 = n25328 ^ n22832 ^ n2107 ;
  assign n41186 = n3850 & n15825 ;
  assign n41188 = n41187 ^ n41186 ^ n35835 ;
  assign n41189 = n9573 ^ x197 ^ 1'b0 ;
  assign n41190 = n14879 & ~n36231 ;
  assign n41193 = n17763 & n20186 ;
  assign n41194 = n41193 ^ n9773 ^ 1'b0 ;
  assign n41191 = n7990 | n13844 ;
  assign n41192 = n15745 | n41191 ;
  assign n41195 = n41194 ^ n41192 ^ n29162 ;
  assign n41196 = n15337 ^ n2622 ^ 1'b0 ;
  assign n41197 = ~n41195 & n41196 ;
  assign n41198 = n39078 ^ n12494 ^ n10212 ;
  assign n41199 = n16537 & n32933 ;
  assign n41200 = n41199 ^ n26676 ^ 1'b0 ;
  assign n41201 = n41200 ^ n24343 ^ 1'b0 ;
  assign n41202 = n17443 ^ n9538 ^ 1'b0 ;
  assign n41203 = x195 | n34633 ;
  assign n41204 = n41203 ^ n6387 ^ 1'b0 ;
  assign n41205 = n2382 & ~n15549 ;
  assign n41206 = n9352 & n13975 ;
  assign n41207 = n41206 ^ x123 ^ 1'b0 ;
  assign n41208 = n17906 | n41207 ;
  assign n41209 = n1958 | n41208 ;
  assign n41210 = n41209 ^ n40384 ^ 1'b0 ;
  assign n41211 = n30949 ^ n847 ^ n624 ;
  assign n41212 = n21053 ^ n20389 ^ 1'b0 ;
  assign n41213 = n41212 ^ n38047 ^ 1'b0 ;
  assign n41214 = n8799 & ~n40439 ;
  assign n41215 = ~n5646 & n41214 ;
  assign n41216 = n40979 & n41215 ;
  assign n41217 = ~n41213 & n41216 ;
  assign n41218 = n12817 & n31526 ;
  assign n41219 = n24871 ^ n4660 ^ 1'b0 ;
  assign n41220 = n16366 & ~n41219 ;
  assign n41221 = n2157 & n38000 ;
  assign n41223 = ( ~n1521 & n4498 ) | ( ~n1521 & n24433 ) | ( n4498 & n24433 ) ;
  assign n41222 = ~n2211 & n3666 ;
  assign n41224 = n41223 ^ n41222 ^ 1'b0 ;
  assign n41226 = n16187 ^ n6033 ^ 1'b0 ;
  assign n41227 = ~n24063 & n41226 ;
  assign n41228 = ~n28732 & n41227 ;
  assign n41225 = n10894 & n27593 ;
  assign n41229 = n41228 ^ n41225 ^ 1'b0 ;
  assign n41230 = ( n32034 & n36330 ) | ( n32034 & n37537 ) | ( n36330 & n37537 ) ;
  assign n41231 = x152 & ~n587 ;
  assign n41232 = ~x152 & n41231 ;
  assign n41233 = n41232 ^ n2158 ^ 1'b0 ;
  assign n41234 = n2142 | n8094 ;
  assign n41235 = n41233 & ~n41234 ;
  assign n41236 = ~n12460 & n33663 ;
  assign n41237 = n41236 ^ n5001 ^ 1'b0 ;
  assign n41238 = n41235 & n41237 ;
  assign n41239 = ~n4251 & n14703 ;
  assign n41240 = ~x60 & n41239 ;
  assign n41241 = x167 | n41240 ;
  assign n41245 = n14830 ^ n14504 ^ 1'b0 ;
  assign n41246 = n5455 & ~n41245 ;
  assign n41244 = n3049 & ~n8558 ;
  assign n41242 = n3349 | n6116 ;
  assign n41243 = n26718 & ~n41242 ;
  assign n41247 = n41246 ^ n41244 ^ n41243 ;
  assign n41248 = n32846 ^ n2348 ^ 1'b0 ;
  assign n41249 = ~n41247 & n41248 ;
  assign n41250 = n7502 ^ n6621 ^ 1'b0 ;
  assign n41251 = n41249 & ~n41250 ;
  assign n41253 = n17427 ^ n1303 ^ 1'b0 ;
  assign n41254 = ~n6173 & n41253 ;
  assign n41252 = n8694 | n29445 ;
  assign n41255 = n41254 ^ n41252 ^ 1'b0 ;
  assign n41256 = ~n3704 & n34004 ;
  assign n41257 = n2746 & n13255 ;
  assign n41258 = n20998 & n41257 ;
  assign n41259 = n33473 & n41258 ;
  assign n41260 = n2887 & ~n7173 ;
  assign n41261 = n41260 ^ n4510 ^ 1'b0 ;
  assign n41262 = n4379 | n21802 ;
  assign n41263 = n22552 & n41262 ;
  assign n41264 = n34175 ^ n16693 ^ 1'b0 ;
  assign n41265 = n41263 & n41264 ;
  assign n41266 = ~n10157 & n10337 ;
  assign n41267 = ~n4608 & n41266 ;
  assign n41268 = n928 & ~n31116 ;
  assign n41269 = ~n12381 & n41268 ;
  assign n41270 = n41269 ^ n11891 ^ 1'b0 ;
  assign n41274 = n20153 & ~n34809 ;
  assign n41275 = n27546 & n41274 ;
  assign n41271 = n8456 ^ n1070 ^ 1'b0 ;
  assign n41272 = ~n6335 & n41271 ;
  assign n41273 = ~n4648 & n41272 ;
  assign n41276 = n41275 ^ n41273 ^ 1'b0 ;
  assign n41277 = n9919 | n28164 ;
  assign n41278 = ( ~n5391 & n7541 ) | ( ~n5391 & n41277 ) | ( n7541 & n41277 ) ;
  assign n41279 = n16271 ^ n2058 ^ 1'b0 ;
  assign n41280 = n14651 | n41279 ;
  assign n41281 = ( n25622 & ~n27871 ) | ( n25622 & n38399 ) | ( ~n27871 & n38399 ) ;
  assign n41282 = n31341 ^ n26819 ^ 1'b0 ;
  assign n41283 = n41281 | n41282 ;
  assign n41284 = n11414 ^ n1990 ^ 1'b0 ;
  assign n41285 = n7908 & ~n33993 ;
  assign n41286 = n41285 ^ n21745 ^ 1'b0 ;
  assign n41287 = n14206 | n19663 ;
  assign n41288 = ~n1805 & n9970 ;
  assign n41289 = n25269 ^ n20888 ^ 1'b0 ;
  assign n41290 = n1508 & ~n41289 ;
  assign n41291 = n41290 ^ n39599 ^ n28754 ;
  assign n41292 = ( n2077 & n6335 ) | ( n2077 & n11551 ) | ( n6335 & n11551 ) ;
  assign n41293 = n3326 | n41292 ;
  assign n41294 = n27712 & ~n41293 ;
  assign n41295 = n10397 & ~n11449 ;
  assign n41296 = ( n18586 & ~n32305 ) | ( n18586 & n41295 ) | ( ~n32305 & n41295 ) ;
  assign n41297 = n4770 ^ n4381 ^ 1'b0 ;
  assign n41298 = ~n4367 & n41297 ;
  assign n41299 = n34861 ^ n3895 ^ 1'b0 ;
  assign n41300 = ~n4792 & n41299 ;
  assign n41301 = n4226 & ~n17617 ;
  assign n41302 = n888 & ~n12287 ;
  assign n41303 = n1887 & n6981 ;
  assign n41304 = n31125 ^ n9513 ^ 1'b0 ;
  assign n41305 = n41303 | n41304 ;
  assign n41306 = n41305 ^ n6783 ^ n5932 ;
  assign n41309 = n13699 ^ n9958 ^ 1'b0 ;
  assign n41310 = n41309 ^ n20063 ^ x0 ;
  assign n41307 = n2511 & n3678 ;
  assign n41308 = n4670 & ~n41307 ;
  assign n41311 = n41310 ^ n41308 ^ 1'b0 ;
  assign n41312 = n8239 ^ n6490 ^ 1'b0 ;
  assign n41313 = n14875 & n15961 ;
  assign n41314 = n3823 & n4039 ;
  assign n41315 = n41314 ^ n1649 ^ 1'b0 ;
  assign n41316 = ~n15524 & n41315 ;
  assign n41317 = n41316 ^ n18262 ^ 1'b0 ;
  assign n41319 = n12007 | n12703 ;
  assign n41318 = ~n11277 & n20914 ;
  assign n41320 = n41319 ^ n41318 ^ 1'b0 ;
  assign n41321 = n9929 & n17321 ;
  assign n41322 = n41321 ^ n1802 ^ 1'b0 ;
  assign n41323 = n16695 & ~n41322 ;
  assign n41324 = n13292 & n41323 ;
  assign n41325 = n33653 | n37303 ;
  assign n41326 = ~n5733 & n9032 ;
  assign n41327 = n6324 & n14949 ;
  assign n41328 = n7961 & n41327 ;
  assign n41329 = n4452 & ~n4493 ;
  assign n41330 = n19091 & n41329 ;
  assign n41331 = n2165 & n41330 ;
  assign n41332 = ( n41326 & n41328 ) | ( n41326 & ~n41331 ) | ( n41328 & ~n41331 ) ;
  assign n41333 = n37368 ^ n26809 ^ 1'b0 ;
  assign n41334 = n5602 | n29760 ;
  assign n41335 = n36742 | n41334 ;
  assign n41336 = ~n5341 & n39048 ;
  assign n41337 = n3408 | n23042 ;
  assign n41338 = ~n1943 & n16739 ;
  assign n41339 = n36056 ^ n19543 ^ 1'b0 ;
  assign n41340 = ~n41338 & n41339 ;
  assign n41341 = n17836 | n37560 ;
  assign n41342 = n41341 ^ n3265 ^ 1'b0 ;
  assign n41343 = n8025 & ~n14971 ;
  assign n41344 = n41343 ^ n23659 ^ 1'b0 ;
  assign n41345 = ~n26562 & n41344 ;
  assign n41346 = n23011 & n41345 ;
  assign n41347 = n26366 ^ n13239 ^ 1'b0 ;
  assign n41348 = n2951 | n10999 ;
  assign n41349 = n25626 | n41348 ;
  assign n41350 = n41349 ^ n1733 ^ 1'b0 ;
  assign n41351 = n41347 | n41350 ;
  assign n41352 = ( n1250 & n9076 ) | ( n1250 & n14531 ) | ( n9076 & n14531 ) ;
  assign n41353 = n2055 | n34820 ;
  assign n41354 = n41353 ^ n37284 ^ n19723 ;
  assign n41355 = n25481 ^ n2934 ^ 1'b0 ;
  assign n41356 = n31044 | n41355 ;
  assign n41357 = n23830 & ~n41356 ;
  assign n41358 = n4619 | n26718 ;
  assign n41359 = n24465 & n41358 ;
  assign n41360 = ~n1387 & n33932 ;
  assign n41361 = n23726 & n41360 ;
  assign n41362 = ~x195 & n34908 ;
  assign n41363 = ~n26200 & n41362 ;
  assign n41364 = n11272 ^ n1100 ^ 1'b0 ;
  assign n41365 = n13917 | n41364 ;
  assign n41366 = n41365 ^ n32254 ^ 1'b0 ;
  assign n41367 = n29926 | n41366 ;
  assign n41368 = n7748 ^ n2415 ^ 1'b0 ;
  assign n41369 = n8888 & n41368 ;
  assign n41370 = n39787 & n41369 ;
  assign n41371 = n5621 & n15668 ;
  assign n41372 = n41371 ^ n29562 ^ n10015 ;
  assign n41373 = n2982 | n41372 ;
  assign n41374 = ~n16730 & n19727 ;
  assign n41375 = n14196 & n41374 ;
  assign n41376 = n27050 & ~n41375 ;
  assign n41377 = ~n543 & n41376 ;
  assign n41378 = n6879 | n40035 ;
  assign n41379 = n4039 | n41378 ;
  assign n41380 = ~n3579 & n8371 ;
  assign n41381 = n4180 | n5680 ;
  assign n41383 = n16857 & n24932 ;
  assign n41384 = n41383 ^ n12367 ^ 1'b0 ;
  assign n41385 = n41384 ^ n5313 ^ 1'b0 ;
  assign n41386 = n29866 & ~n41385 ;
  assign n41382 = n30778 ^ n20702 ^ 1'b0 ;
  assign n41387 = n41386 ^ n41382 ^ 1'b0 ;
  assign n41388 = n23063 & n28777 ;
  assign n41389 = n5311 & ~n41388 ;
  assign n41390 = n6492 & ~n10913 ;
  assign n41391 = n1259 | n5637 ;
  assign n41392 = n37980 | n41391 ;
  assign n41395 = n13620 ^ n10853 ^ n4409 ;
  assign n41393 = n12270 & n15507 ;
  assign n41394 = n41393 ^ n33624 ^ 1'b0 ;
  assign n41396 = n41395 ^ n41394 ^ 1'b0 ;
  assign n41397 = n9986 | n17526 ;
  assign n41398 = ~n19213 & n41397 ;
  assign n41399 = n34418 ^ n15500 ^ 1'b0 ;
  assign n41400 = n16899 ^ n5917 ^ 1'b0 ;
  assign n41401 = n3879 ^ n289 ^ 1'b0 ;
  assign n41402 = n41400 & n41401 ;
  assign n41403 = n41402 ^ n16429 ^ 1'b0 ;
  assign n41404 = n8658 | n16370 ;
  assign n41405 = n1746 & ~n38699 ;
  assign n41406 = n35711 ^ n23890 ^ 1'b0 ;
  assign n41407 = n2051 & ~n20524 ;
  assign n41408 = ~n6417 & n40252 ;
  assign n41409 = ~n41407 & n41408 ;
  assign n41410 = n41409 ^ n11053 ^ 1'b0 ;
  assign n41411 = n13774 & n41410 ;
  assign n41412 = n33182 ^ n6138 ^ 1'b0 ;
  assign n41413 = n26469 & ~n38272 ;
  assign n41414 = ~n4632 & n41413 ;
  assign n41415 = n41412 & n41414 ;
  assign n41416 = n2926 & n15392 ;
  assign n41417 = n33223 & n41416 ;
  assign n41418 = ~n17796 & n26963 ;
  assign n41419 = n41417 | n41418 ;
  assign n41420 = n25323 ^ n2287 ^ 1'b0 ;
  assign n41421 = n22118 & ~n27089 ;
  assign n41422 = n37369 ^ n25633 ^ 1'b0 ;
  assign n41423 = n28472 ^ n8830 ^ n856 ;
  assign n41424 = n41423 ^ n7257 ^ 1'b0 ;
  assign n41426 = n10493 & ~n40736 ;
  assign n41427 = n41426 ^ n25104 ^ 1'b0 ;
  assign n41425 = n6272 & n20714 ;
  assign n41428 = n41427 ^ n41425 ^ 1'b0 ;
  assign n41429 = n6358 & ~n6591 ;
  assign n41430 = n21984 & n41429 ;
  assign n41431 = n41430 ^ n39741 ^ 1'b0 ;
  assign n41432 = n25377 ^ n18425 ^ 1'b0 ;
  assign n41433 = ~n19534 & n41432 ;
  assign n41434 = n26739 ^ n13748 ^ 1'b0 ;
  assign n41435 = n41433 & ~n41434 ;
  assign n41436 = n9180 & n11749 ;
  assign n41437 = n41436 ^ n30081 ^ 1'b0 ;
  assign n41438 = n12288 | n41437 ;
  assign n41439 = n41438 ^ n34469 ^ 1'b0 ;
  assign n41440 = n9317 & n26243 ;
  assign n41441 = n2306 | n41440 ;
  assign n41442 = n21291 & ~n37402 ;
  assign n41443 = n38450 ^ n6350 ^ 1'b0 ;
  assign n41445 = n22321 ^ n11124 ^ 1'b0 ;
  assign n41444 = n18369 & ~n30228 ;
  assign n41446 = n41445 ^ n41444 ^ 1'b0 ;
  assign n41447 = n4263 | n31061 ;
  assign n41448 = n18856 & ~n41447 ;
  assign n41449 = n40833 & ~n41448 ;
  assign n41450 = n28627 ^ n6471 ^ 1'b0 ;
  assign n41451 = n36179 | n41450 ;
  assign n41452 = n27828 ^ n19082 ^ 1'b0 ;
  assign n41453 = ~n18254 & n41452 ;
  assign n41454 = n41453 ^ n39141 ^ 1'b0 ;
  assign n41455 = n23102 | n35103 ;
  assign n41456 = ~n1730 & n7069 ;
  assign n41457 = ~n15014 & n39486 ;
  assign n41458 = ~n41456 & n41457 ;
  assign n41459 = n6155 ^ n5302 ^ 1'b0 ;
  assign n41460 = n6206 & n41459 ;
  assign n41461 = n2755 & ~n41460 ;
  assign n41462 = n10854 & ~n13530 ;
  assign n41463 = n41462 ^ n18679 ^ 1'b0 ;
  assign n41464 = n20247 | n41463 ;
  assign n41465 = n28877 | n41464 ;
  assign n41466 = ~n25415 & n41465 ;
  assign n41467 = n26244 ^ n13675 ^ 1'b0 ;
  assign n41468 = n22826 ^ n19021 ^ n3040 ;
  assign n41469 = n41468 ^ n20675 ^ n500 ;
  assign n41471 = ~n4541 & n10387 ;
  assign n41472 = n27419 & ~n41471 ;
  assign n41473 = ~n8108 & n41472 ;
  assign n41470 = n8794 & ~n14640 ;
  assign n41474 = n41473 ^ n41470 ^ 1'b0 ;
  assign n41475 = ~n14956 & n32162 ;
  assign n41476 = n11479 | n20362 ;
  assign n41477 = n10399 & ~n41476 ;
  assign n41478 = n7752 ^ n6897 ^ 1'b0 ;
  assign n41479 = n12809 & n41478 ;
  assign n41480 = n41477 | n41479 ;
  assign n41481 = n13427 ^ n3329 ^ 1'b0 ;
  assign n41482 = n41480 | n41481 ;
  assign n41483 = ( n17779 & n31046 ) | ( n17779 & ~n41482 ) | ( n31046 & ~n41482 ) ;
  assign n41484 = n22083 ^ n19325 ^ 1'b0 ;
  assign n41485 = n41483 & n41484 ;
  assign n41486 = ~x116 & n597 ;
  assign n41487 = n6430 | n10845 ;
  assign n41488 = ~n11467 & n18016 ;
  assign n41489 = n41488 ^ n3845 ^ 1'b0 ;
  assign n41490 = n35404 & ~n41489 ;
  assign n41491 = n19552 & n41490 ;
  assign n41492 = n33182 ^ n20616 ^ 1'b0 ;
  assign n41493 = n858 & ~n41492 ;
  assign n41494 = n21881 ^ n18267 ^ 1'b0 ;
  assign n41495 = ( n9332 & n41493 ) | ( n9332 & ~n41494 ) | ( n41493 & ~n41494 ) ;
  assign n41496 = n1377 & ~n18070 ;
  assign n41497 = n33912 ^ n29036 ^ 1'b0 ;
  assign n41498 = n41305 ^ n916 ^ 1'b0 ;
  assign n41499 = n9345 | n41498 ;
  assign n41500 = n1025 & ~n20006 ;
  assign n41501 = n41499 & n41500 ;
  assign n41502 = n17499 ^ n3333 ^ 1'b0 ;
  assign n41503 = n780 | n41502 ;
  assign n41504 = n8351 & n8907 ;
  assign n41505 = n41503 & n41504 ;
  assign n41506 = n523 & ~n2044 ;
  assign n41507 = n25163 | n41506 ;
  assign n41508 = n36133 | n41507 ;
  assign n41509 = n11749 & ~n13800 ;
  assign n41510 = n41509 ^ n10289 ^ 1'b0 ;
  assign n41511 = n41510 ^ n16521 ^ 1'b0 ;
  assign n41512 = ( n28570 & n31471 ) | ( n28570 & n32150 ) | ( n31471 & n32150 ) ;
  assign n41513 = ~n7246 & n12096 ;
  assign n41514 = n41513 ^ n4682 ^ 1'b0 ;
  assign n41515 = n7332 | n8820 ;
  assign n41516 = n41514 & ~n41515 ;
  assign n41517 = n5276 & n16320 ;
  assign n41518 = n41517 ^ n4718 ^ 1'b0 ;
  assign n41519 = n13912 & n36848 ;
  assign n41520 = ~n41518 & n41519 ;
  assign n41521 = n24932 ^ n16428 ^ 1'b0 ;
  assign n41522 = n16846 | n41521 ;
  assign n41523 = n41522 ^ n21741 ^ 1'b0 ;
  assign n41524 = n10729 | n22460 ;
  assign n41525 = ( n2615 & n23689 ) | ( n2615 & n34116 ) | ( n23689 & n34116 ) ;
  assign n41526 = n10357 ^ n3615 ^ 1'b0 ;
  assign n41527 = n8585 & n41526 ;
  assign n41528 = n1384 & ~n5535 ;
  assign n41529 = ~n41527 & n41528 ;
  assign n41530 = n3300 | n7771 ;
  assign n41531 = n18976 & ~n30346 ;
  assign n41532 = n36798 ^ n3156 ^ 1'b0 ;
  assign n41533 = n287 & n28889 ;
  assign n41534 = n41533 ^ n20400 ^ n17109 ;
  assign n41535 = n2745 & ~n20614 ;
  assign n41536 = n1911 | n10429 ;
  assign n41537 = ~n41535 & n41536 ;
  assign n41538 = n41537 ^ n17521 ^ 1'b0 ;
  assign n41539 = n20726 & n41538 ;
  assign n41540 = n16113 & n41539 ;
  assign n41541 = ~n4285 & n41540 ;
  assign n41542 = x176 & ~n8016 ;
  assign n41543 = ~n9817 & n33601 ;
  assign n41545 = n9401 & n11272 ;
  assign n41546 = n41545 ^ n35075 ^ 1'b0 ;
  assign n41547 = n11665 | n41546 ;
  assign n41548 = n34025 ^ n17427 ^ 1'b0 ;
  assign n41549 = ~n41547 & n41548 ;
  assign n41544 = n18894 & ~n36295 ;
  assign n41550 = n41549 ^ n41544 ^ 1'b0 ;
  assign n41551 = n27265 ^ n2158 ^ 1'b0 ;
  assign n41552 = n35896 | n39105 ;
  assign n41553 = n41552 ^ n14952 ^ n1471 ;
  assign n41554 = ~n1341 & n38510 ;
  assign n41555 = n7205 & n29295 ;
  assign n41556 = n4298 & ~n7287 ;
  assign n41557 = n34373 ^ n4040 ^ n3747 ;
  assign n41558 = n41557 ^ n14092 ^ 1'b0 ;
  assign n41559 = n8710 & ~n10819 ;
  assign n41560 = n41559 ^ n1912 ^ 1'b0 ;
  assign n41561 = n9664 & n41560 ;
  assign n41562 = ~n20974 & n41561 ;
  assign n41563 = n41562 ^ n8408 ^ 1'b0 ;
  assign n41564 = n26515 ^ n23073 ^ 1'b0 ;
  assign n41565 = n28342 | n41564 ;
  assign n41566 = n4887 & ~n41565 ;
  assign n41567 = ~n41563 & n41566 ;
  assign n41568 = n36318 ^ n10405 ^ 1'b0 ;
  assign n41569 = n18024 & n19528 ;
  assign n41570 = n10657 & n41569 ;
  assign n41571 = ~n41315 & n41570 ;
  assign n41572 = n9113 & n41571 ;
  assign n41576 = n7746 & n11649 ;
  assign n41577 = n16068 & n41576 ;
  assign n41573 = x136 & ~n291 ;
  assign n41574 = n41573 ^ n22123 ^ 1'b0 ;
  assign n41575 = ~n813 & n41574 ;
  assign n41578 = n41577 ^ n41575 ^ 1'b0 ;
  assign n41579 = ( n4935 & ~n10068 ) | ( n4935 & n41578 ) | ( ~n10068 & n41578 ) ;
  assign n41580 = n29154 ^ n18551 ^ 1'b0 ;
  assign n41581 = n16273 ^ n11968 ^ 1'b0 ;
  assign n41582 = n9031 & n19813 ;
  assign n41583 = n15689 & n41582 ;
  assign n41584 = n1458 | n16975 ;
  assign n41585 = n9873 | n14846 ;
  assign n41586 = n41584 | n41585 ;
  assign n41587 = n16269 | n41156 ;
  assign n41588 = n27795 | n33233 ;
  assign n41589 = n19960 ^ n18482 ^ n3635 ;
  assign n41590 = n38205 ^ n22519 ^ 1'b0 ;
  assign n41591 = n3412 & n41590 ;
  assign n41592 = ( n5442 & n9758 ) | ( n5442 & ~n28203 ) | ( n9758 & ~n28203 ) ;
  assign n41593 = n21683 ^ n6984 ^ 1'b0 ;
  assign n41594 = n41593 ^ n30366 ^ 1'b0 ;
  assign n41595 = ~n41592 & n41594 ;
  assign n41596 = n4470 & ~n37792 ;
  assign n41597 = n36198 ^ n4031 ^ 1'b0 ;
  assign n41598 = n5668 & n13513 ;
  assign n41599 = n35161 ^ n27485 ^ 1'b0 ;
  assign n41600 = n8591 ^ n858 ^ 1'b0 ;
  assign n41601 = ( n1815 & n10570 ) | ( n1815 & ~n41600 ) | ( n10570 & ~n41600 ) ;
  assign n41602 = n24845 & ~n41601 ;
  assign n41603 = n41602 ^ n3050 ^ 1'b0 ;
  assign n41604 = ~n35775 & n41603 ;
  assign n41605 = n3985 & ~n4758 ;
  assign n41606 = n23135 & n23521 ;
  assign n41607 = n4080 & ~n26148 ;
  assign n41608 = n2227 & ~n41607 ;
  assign n41609 = n41608 ^ n8496 ^ 1'b0 ;
  assign n41610 = n16082 & n38661 ;
  assign n41611 = n19576 ^ n10805 ^ 1'b0 ;
  assign n41612 = n9667 | n41611 ;
  assign n41613 = n4970 & ~n15321 ;
  assign n41614 = ( n7107 & ~n33222 ) | ( n7107 & n40103 ) | ( ~n33222 & n40103 ) ;
  assign n41615 = ( ~n33648 & n41613 ) | ( ~n33648 & n41614 ) | ( n41613 & n41614 ) ;
  assign n41616 = n41615 ^ n39975 ^ n6502 ;
  assign n41617 = n2369 ^ n2245 ^ 1'b0 ;
  assign n41618 = ~n2710 & n41617 ;
  assign n41619 = n11815 & ~n41618 ;
  assign n41620 = ( n23489 & ~n31817 ) | ( n23489 & n41619 ) | ( ~n31817 & n41619 ) ;
  assign n41621 = n16304 ^ n15600 ^ 1'b0 ;
  assign n41622 = ~n8216 & n33253 ;
  assign n41623 = ~n41621 & n41622 ;
  assign n41624 = n19665 ^ x129 ^ 1'b0 ;
  assign n41625 = n274 & n894 ;
  assign n41626 = ~n41624 & n41625 ;
  assign n41627 = ~n8545 & n17241 ;
  assign n41628 = n6786 ^ n400 ^ 1'b0 ;
  assign n41629 = n41627 | n41628 ;
  assign n41630 = ~n8434 & n22332 ;
  assign n41631 = n41630 ^ n25610 ^ n5835 ;
  assign n41632 = n2615 | n17517 ;
  assign n41633 = x167 & ~n14852 ;
  assign n41634 = n41633 ^ n19830 ^ 1'b0 ;
  assign n41635 = n6271 ^ n5328 ^ 1'b0 ;
  assign n41636 = n41634 | n41635 ;
  assign n41637 = ~n2489 & n41560 ;
  assign n41638 = n41637 ^ n2246 ^ 1'b0 ;
  assign n41639 = n25386 ^ n21503 ^ 1'b0 ;
  assign n41640 = ~n22801 & n41639 ;
  assign n41641 = n6454 | n40576 ;
  assign n41642 = n11199 & n29329 ;
  assign n41643 = n1624 & n13897 ;
  assign n41644 = ~n41642 & n41643 ;
  assign n41645 = n41641 | n41644 ;
  assign n41646 = n10172 ^ n8548 ^ n922 ;
  assign n41647 = n535 & n41646 ;
  assign n41648 = n7918 ^ n1402 ^ 1'b0 ;
  assign n41649 = n8096 & ~n41648 ;
  assign n41650 = n41649 ^ n38801 ^ n30662 ;
  assign n41651 = n35475 ^ n27321 ^ n16446 ;
  assign n41670 = n7449 | n16187 ;
  assign n41671 = n41670 ^ n28559 ^ 1'b0 ;
  assign n41652 = x15 & ~n6632 ;
  assign n41653 = n6632 & n41652 ;
  assign n41654 = x97 & ~n509 ;
  assign n41655 = n509 & n41654 ;
  assign n41656 = x249 & ~n1345 ;
  assign n41657 = n1345 & n41656 ;
  assign n41658 = n41655 | n41657 ;
  assign n41659 = n41655 & ~n41658 ;
  assign n41660 = n8365 & ~n41659 ;
  assign n41661 = ~n8365 & n41660 ;
  assign n41662 = n10466 | n41661 ;
  assign n41663 = n10466 & ~n41662 ;
  assign n41664 = n41663 ^ n19390 ^ 1'b0 ;
  assign n41665 = ~n41653 & n41664 ;
  assign n41666 = ~n20805 & n41665 ;
  assign n41667 = n18079 & ~n41666 ;
  assign n41668 = ~n21479 & n41667 ;
  assign n41669 = n8248 | n41668 ;
  assign n41672 = n41671 ^ n41669 ^ 1'b0 ;
  assign n41673 = n10619 & ~n26370 ;
  assign n41674 = n41673 ^ n39477 ^ 1'b0 ;
  assign n41675 = n41674 ^ n1544 ^ 1'b0 ;
  assign n41676 = n10268 & n41675 ;
  assign n41677 = n16657 & ~n31462 ;
  assign n41678 = n16309 & ~n22396 ;
  assign n41679 = n3312 & ~n4430 ;
  assign n41680 = n41679 ^ n2657 ^ 1'b0 ;
  assign n41681 = n36142 & ~n41680 ;
  assign n41684 = n13761 ^ n12104 ^ n4169 ;
  assign n41685 = n1180 & ~n19482 ;
  assign n41686 = ~n41684 & n41685 ;
  assign n41682 = n6666 & n9371 ;
  assign n41683 = ~n5195 & n41682 ;
  assign n41687 = n41686 ^ n41683 ^ 1'b0 ;
  assign n41688 = n9487 | n40027 ;
  assign n41689 = n41688 ^ n10743 ^ 1'b0 ;
  assign n41690 = n5530 & n41689 ;
  assign n41691 = n41690 ^ n25386 ^ 1'b0 ;
  assign n41692 = n25183 ^ n883 ^ 1'b0 ;
  assign n41693 = ~n41691 & n41692 ;
  assign n41694 = n35951 ^ n3067 ^ 1'b0 ;
  assign n41695 = n8403 | n41694 ;
  assign n41698 = ( ~n2828 & n5125 ) | ( ~n2828 & n20030 ) | ( n5125 & n20030 ) ;
  assign n41696 = n18615 & ~n21361 ;
  assign n41697 = ~x86 & n41696 ;
  assign n41699 = n41698 ^ n41697 ^ 1'b0 ;
  assign n41700 = n2224 & ~n24132 ;
  assign n41701 = n41700 ^ n18226 ^ 1'b0 ;
  assign n41702 = n33931 ^ n5320 ^ 1'b0 ;
  assign n41703 = ~n4076 & n41702 ;
  assign n41704 = n28662 ^ n3615 ^ 1'b0 ;
  assign n41705 = n471 & n13340 ;
  assign n41706 = n12656 | n12737 ;
  assign n41707 = n41706 ^ n13466 ^ n13099 ;
  assign n41708 = n29578 ^ n28161 ^ n911 ;
  assign n41709 = ~n10731 & n41708 ;
  assign n41711 = n5478 & ~n27058 ;
  assign n41712 = n41711 ^ n37388 ^ n10515 ;
  assign n41710 = x168 & n14203 ;
  assign n41713 = n41712 ^ n41710 ^ 1'b0 ;
  assign n41714 = n9836 | n15312 ;
  assign n41715 = n34572 ^ n15131 ^ 1'b0 ;
  assign n41716 = n7742 & n22399 ;
  assign n41717 = ( n32550 & n36388 ) | ( n32550 & ~n41677 ) | ( n36388 & ~n41677 ) ;
  assign n41718 = n375 & n11870 ;
  assign n41720 = n16775 ^ n15297 ^ 1'b0 ;
  assign n41721 = n6525 ^ n4325 ^ 1'b0 ;
  assign n41722 = n41720 & n41721 ;
  assign n41719 = n2970 | n8609 ;
  assign n41723 = n41722 ^ n41719 ^ 1'b0 ;
  assign n41724 = n38904 ^ n14956 ^ 1'b0 ;
  assign n41725 = n3654 & n14984 ;
  assign n41726 = n29025 & n41725 ;
  assign n41727 = n1545 ^ n1398 ^ 1'b0 ;
  assign n41728 = n41727 ^ n30942 ^ 1'b0 ;
  assign n41729 = n28574 & ~n41728 ;
  assign n41730 = n9415 ^ n1862 ^ 1'b0 ;
  assign n41731 = n2887 & ~n41730 ;
  assign n41732 = n35844 ^ n5525 ^ 1'b0 ;
  assign n41733 = n41731 & ~n41732 ;
  assign n41734 = n22804 ^ n19218 ^ 1'b0 ;
  assign n41735 = n41539 ^ n9280 ^ 1'b0 ;
  assign n41736 = ~n11475 & n23411 ;
  assign n41737 = n16350 & ~n27063 ;
  assign n41738 = ~n16129 & n20439 ;
  assign n41739 = ~n41737 & n41738 ;
  assign n41740 = n35896 & n36440 ;
  assign n41741 = n38769 & n41740 ;
  assign n41742 = n3257 & n12357 ;
  assign n41743 = n41742 ^ n9100 ^ 1'b0 ;
  assign n41744 = n22817 & ~n30594 ;
  assign n41745 = n20023 & n41744 ;
  assign n41746 = ( n21131 & ~n37591 ) | ( n21131 & n41745 ) | ( ~n37591 & n41745 ) ;
  assign n41747 = ( n12862 & n13848 ) | ( n12862 & ~n18034 ) | ( n13848 & ~n18034 ) ;
  assign n41748 = n27640 & n41747 ;
  assign n41749 = ~n34845 & n41748 ;
  assign n41750 = n41749 ^ n29920 ^ n19475 ;
  assign n41751 = n18688 ^ n17641 ^ 1'b0 ;
  assign n41752 = n1765 & ~n41751 ;
  assign n41753 = n40642 ^ n5302 ^ 1'b0 ;
  assign n41754 = n5761 | n41753 ;
  assign n41755 = n9466 ^ n6906 ^ 1'b0 ;
  assign n41756 = n41755 ^ n38452 ^ n6844 ;
  assign n41757 = ~n35505 & n41756 ;
  assign n41758 = n11344 | n18054 ;
  assign n41759 = n11941 & n40874 ;
  assign n41760 = n41759 ^ n31736 ^ 1'b0 ;
  assign n41761 = n16695 & n18205 ;
  assign n41762 = ~n41760 & n41761 ;
  assign n41763 = ~n14807 & n24254 ;
  assign n41764 = n21198 ^ n6817 ^ 1'b0 ;
  assign n41765 = n7000 ^ n3395 ^ 1'b0 ;
  assign n41766 = n2602 & ~n2891 ;
  assign n41767 = n29852 & n41766 ;
  assign n41768 = n9100 & n27030 ;
  assign n41769 = n2755 | n41768 ;
  assign n41770 = n41769 ^ n11671 ^ 1'b0 ;
  assign n41771 = n16647 | n41770 ;
  assign n41772 = ~n2343 & n16509 ;
  assign n41773 = n41772 ^ n13954 ^ 1'b0 ;
  assign n41774 = ~n41771 & n41773 ;
  assign n41775 = n3670 | n13954 ;
  assign n41776 = n14844 ^ n5110 ^ n3518 ;
  assign n41777 = n10709 & n41776 ;
  assign n41778 = n23025 & n41777 ;
  assign n41779 = n15832 | n41778 ;
  assign n41780 = n35019 ^ n3689 ^ 1'b0 ;
  assign n41781 = n28418 & ~n41780 ;
  assign n41782 = n23579 | n31743 ;
  assign n41783 = n2356 & ~n41782 ;
  assign n41784 = n769 & ~n41783 ;
  assign n41785 = ~n41781 & n41784 ;
  assign n41786 = ~n7731 & n15600 ;
  assign n41787 = n1129 & n7711 ;
  assign n41788 = n41787 ^ n13291 ^ n5371 ;
  assign n41789 = n3716 | n31550 ;
  assign n41790 = n2400 & n7222 ;
  assign n41791 = n41789 & n41790 ;
  assign n41792 = n12793 ^ x140 ^ 1'b0 ;
  assign n41793 = ~n3639 & n16915 ;
  assign n41794 = n36274 ^ n30025 ^ 1'b0 ;
  assign n41795 = ~n2776 & n41794 ;
  assign n41796 = n41793 & n41795 ;
  assign n41798 = n12306 ^ n2338 ^ 1'b0 ;
  assign n41797 = ( ~n1177 & n23078 ) | ( ~n1177 & n29400 ) | ( n23078 & n29400 ) ;
  assign n41799 = n41798 ^ n41797 ^ n8454 ;
  assign n41800 = n41799 ^ n21578 ^ 1'b0 ;
  assign n41801 = ~n19068 & n33117 ;
  assign n41802 = n2155 & ~n5072 ;
  assign n41803 = n17928 & n41802 ;
  assign n41804 = ~n7974 & n40407 ;
  assign n41805 = n41803 & n41804 ;
  assign n41806 = ~n3137 & n29213 ;
  assign n41807 = ~n16857 & n41806 ;
  assign n41808 = ~n5021 & n5130 ;
  assign n41809 = n13362 ^ n406 ^ 1'b0 ;
  assign n41810 = n5203 | n41809 ;
  assign n41811 = n16522 ^ n1720 ^ 1'b0 ;
  assign n41812 = n41810 | n41811 ;
  assign n41813 = n1977 & n3245 ;
  assign n41814 = ~n31732 & n41813 ;
  assign n41815 = ~n24293 & n26238 ;
  assign n41816 = n22636 ^ n6272 ^ 1'b0 ;
  assign n41817 = n7449 ^ x49 ^ 1'b0 ;
  assign n41818 = n22039 & ~n41817 ;
  assign n41819 = n41818 ^ n38028 ^ 1'b0 ;
  assign n41820 = n14361 ^ n5754 ^ 1'b0 ;
  assign n41821 = n3822 & n7466 ;
  assign n41822 = ~n15750 & n41821 ;
  assign n41823 = ~n41820 & n41822 ;
  assign n41824 = ~n22270 & n33038 ;
  assign n41825 = n41824 ^ n3196 ^ 1'b0 ;
  assign n41826 = n16404 & n41825 ;
  assign n41827 = n16438 & n41826 ;
  assign n41828 = n10231 & n10706 ;
  assign n41829 = ~n6694 & n22476 ;
  assign n41830 = n31973 & n41829 ;
  assign n41831 = ~n22768 & n33815 ;
  assign n41832 = n41831 ^ n38007 ^ 1'b0 ;
  assign n41833 = ~n7999 & n23408 ;
  assign n41834 = ~n41832 & n41833 ;
  assign n41835 = ( n15493 & n17274 ) | ( n15493 & n29976 ) | ( n17274 & n29976 ) ;
  assign n41836 = ( n15607 & ~n19692 ) | ( n15607 & n21666 ) | ( ~n19692 & n21666 ) ;
  assign n41837 = ~n35202 & n37908 ;
  assign n41838 = n15051 ^ n11416 ^ 1'b0 ;
  assign n41839 = n7266 & ~n11096 ;
  assign n41840 = n22059 & n41839 ;
  assign n41841 = n6263 | n12064 ;
  assign n41842 = n41841 ^ n19798 ^ 1'b0 ;
  assign n41843 = n34101 & n41842 ;
  assign n41844 = ~n3014 & n41843 ;
  assign n41845 = n24290 ^ n263 ^ 1'b0 ;
  assign n41846 = n17179 | n41845 ;
  assign n41847 = n16712 ^ n9009 ^ n6117 ;
  assign n41848 = n5700 | n18777 ;
  assign n41849 = n41848 ^ n3291 ^ 1'b0 ;
  assign n41850 = ( n15507 & n17575 ) | ( n15507 & n41849 ) | ( n17575 & n41849 ) ;
  assign n41851 = n32571 ^ n1521 ^ 1'b0 ;
  assign n41852 = n41851 ^ n6177 ^ 1'b0 ;
  assign n41853 = n4306 & ~n14939 ;
  assign n41854 = n28168 & n41853 ;
  assign n41855 = n7976 | n41854 ;
  assign n41856 = n29000 | n41855 ;
  assign n41857 = n24159 & ~n34253 ;
  assign n41858 = n8974 & ~n9855 ;
  assign n41859 = ~n41857 & n41858 ;
  assign n41860 = n34526 ^ n21741 ^ 1'b0 ;
  assign n41861 = n14010 | n36129 ;
  assign n41862 = n5975 | n41861 ;
  assign n41863 = n16642 & ~n25877 ;
  assign n41864 = ~n41862 & n41863 ;
  assign n41865 = n16116 ^ n11268 ^ 1'b0 ;
  assign n41866 = n25205 & n41865 ;
  assign n41867 = n18601 & n32004 ;
  assign n41868 = n41866 & ~n41867 ;
  assign n41869 = n25296 ^ n9034 ^ 1'b0 ;
  assign n41870 = n41869 ^ n26554 ^ n26367 ;
  assign n41871 = n7365 & n17561 ;
  assign n41872 = n41871 ^ n17286 ^ 1'b0 ;
  assign n41873 = n7000 & n41872 ;
  assign n41874 = n3021 & ~n9173 ;
  assign n41875 = n879 & ~n24870 ;
  assign n41876 = n36862 ^ n18187 ^ n17222 ;
  assign n41877 = n29169 | n41876 ;
  assign n41878 = n15550 | n24819 ;
  assign n41879 = n19899 ^ n18526 ^ 1'b0 ;
  assign n41880 = n6521 & n30296 ;
  assign n41881 = ~n41879 & n41880 ;
  assign n41882 = n41881 ^ n27146 ^ n4252 ;
  assign n41883 = n41882 ^ n40306 ^ 1'b0 ;
  assign n41884 = n1680 ^ n1558 ^ 1'b0 ;
  assign n41885 = n41884 ^ n9389 ^ n7944 ;
  assign n41886 = n9013 & n12564 ;
  assign n41887 = n16058 ^ n10243 ^ 1'b0 ;
  assign n41888 = n13091 & n40327 ;
  assign n41889 = n2450 & n34672 ;
  assign n41890 = ~x171 & n17395 ;
  assign n41891 = n41890 ^ n13699 ^ n12778 ;
  assign n41892 = ~n14651 & n41891 ;
  assign n41893 = n41892 ^ n5318 ^ 1'b0 ;
  assign n41894 = n26954 ^ n22523 ^ 1'b0 ;
  assign n41895 = n6810 & n41894 ;
  assign n41896 = n14272 ^ n11692 ^ 1'b0 ;
  assign n41897 = ( n9478 & n11201 ) | ( n9478 & ~n23312 ) | ( n11201 & ~n23312 ) ;
  assign n41898 = n1439 & n8742 ;
  assign n41899 = n29050 & n41898 ;
  assign n41900 = n2509 | n15079 ;
  assign n41901 = n41900 ^ n28901 ^ 1'b0 ;
  assign n41902 = n2397 | n20365 ;
  assign n41903 = ~n19818 & n39091 ;
  assign n41904 = n7759 & n41903 ;
  assign n41905 = n3291 | n26322 ;
  assign n41906 = n11331 ^ n7089 ^ 1'b0 ;
  assign n41907 = ~n41905 & n41906 ;
  assign n41908 = ~n7643 & n41907 ;
  assign n41909 = ( n31721 & n37769 ) | ( n31721 & ~n41908 ) | ( n37769 & ~n41908 ) ;
  assign n41910 = n267 | n8724 ;
  assign n41911 = n16105 & ~n41910 ;
  assign n41912 = ( ~n1853 & n6626 ) | ( ~n1853 & n41911 ) | ( n6626 & n41911 ) ;
  assign n41913 = n26814 ^ n20933 ^ 1'b0 ;
  assign n41914 = n16366 ^ n4004 ^ 1'b0 ;
  assign n41915 = n17671 ^ n5257 ^ 1'b0 ;
  assign n41916 = n17285 & n41915 ;
  assign n41917 = n3007 & ~n26388 ;
  assign n41918 = n32121 ^ n24302 ^ n10747 ;
  assign n41919 = n41917 | n41918 ;
  assign n41920 = ~n2180 & n15192 ;
  assign n41921 = n33661 ^ n18222 ^ 1'b0 ;
  assign n41922 = n1231 ^ n289 ^ 1'b0 ;
  assign n41923 = n36543 ^ n21050 ^ 1'b0 ;
  assign n41924 = n11369 ^ n10968 ^ n10770 ;
  assign n41925 = n28794 & n41924 ;
  assign n41926 = n16423 & n41925 ;
  assign n41927 = n5529 ^ n2372 ^ n2182 ;
  assign n41931 = n24187 ^ n17456 ^ 1'b0 ;
  assign n41928 = n11490 ^ n7207 ^ 1'b0 ;
  assign n41929 = ~n9114 & n41928 ;
  assign n41930 = ~n5084 & n41929 ;
  assign n41932 = n41931 ^ n41930 ^ 1'b0 ;
  assign n41933 = n18319 ^ n1251 ^ 1'b0 ;
  assign n41934 = n32249 ^ n9628 ^ 1'b0 ;
  assign n41935 = n41934 ^ n30977 ^ 1'b0 ;
  assign n41936 = n16718 & n41935 ;
  assign n41937 = n11805 ^ n9754 ^ 1'b0 ;
  assign n41938 = n16023 & n41937 ;
  assign n41939 = ( n4638 & n8964 ) | ( n4638 & n23881 ) | ( n8964 & n23881 ) ;
  assign n41940 = ( n1148 & ~n6639 ) | ( n1148 & n7417 ) | ( ~n6639 & n7417 ) ;
  assign n41941 = x199 & n3258 ;
  assign n41942 = n2905 & ~n41941 ;
  assign n41943 = n38016 ^ n1749 ^ 1'b0 ;
  assign n41944 = ~n481 & n2668 ;
  assign n41945 = n41944 ^ n19109 ^ 1'b0 ;
  assign n41946 = n6005 & n41945 ;
  assign n41947 = n830 | n13228 ;
  assign n41948 = n41947 ^ n21985 ^ 1'b0 ;
  assign n41949 = n13058 & n41948 ;
  assign n41950 = ~n8944 & n15765 ;
  assign n41951 = n41950 ^ n11514 ^ 1'b0 ;
  assign n41952 = n41949 & ~n41951 ;
  assign n41953 = n1200 & ~n4818 ;
  assign n41954 = n30041 ^ n12939 ^ 1'b0 ;
  assign n41955 = ~n41953 & n41954 ;
  assign n41956 = n39368 & n41955 ;
  assign n41957 = n6834 & n41956 ;
  assign n41958 = n1856 & ~n4348 ;
  assign n41959 = n3400 & n41958 ;
  assign n41960 = n7522 ^ n5229 ^ 1'b0 ;
  assign n41961 = ~n22894 & n41960 ;
  assign n41962 = n41959 & n41961 ;
  assign n41963 = n4350 & n20519 ;
  assign n41964 = n41963 ^ n26209 ^ 1'b0 ;
  assign n41965 = n2286 & n10126 ;
  assign n41966 = n38546 ^ n19336 ^ n12603 ;
  assign n41967 = n3509 & n11182 ;
  assign n41969 = n6444 | n9746 ;
  assign n41968 = n14522 & ~n14737 ;
  assign n41970 = n41969 ^ n41968 ^ 1'b0 ;
  assign n41971 = ~n4555 & n9383 ;
  assign n41972 = n27546 ^ n26167 ^ 1'b0 ;
  assign n41974 = x64 & n2740 ;
  assign n41973 = n4642 | n14371 ;
  assign n41975 = n41974 ^ n41973 ^ 1'b0 ;
  assign n41976 = ( n1010 & n3985 ) | ( n1010 & n35218 ) | ( n3985 & n35218 ) ;
  assign n41977 = n15895 | n23871 ;
  assign n41978 = n41976 & ~n41977 ;
  assign n41979 = n29506 ^ n16891 ^ n1393 ;
  assign n41980 = n402 | n41979 ;
  assign n41981 = n31471 ^ n16963 ^ 1'b0 ;
  assign n41982 = n17824 ^ n2121 ^ 1'b0 ;
  assign n41983 = n25374 & ~n41982 ;
  assign n41984 = ~n21598 & n28297 ;
  assign n41985 = ~n41983 & n41984 ;
  assign n41986 = n10301 & ~n35606 ;
  assign n41987 = n591 & n19644 ;
  assign n41988 = n26640 ^ n7513 ^ 1'b0 ;
  assign n41989 = ~n18938 & n41988 ;
  assign n41990 = n2872 ^ n2039 ^ 1'b0 ;
  assign n41991 = n10305 & n41990 ;
  assign n41992 = n25023 | n26573 ;
  assign n41993 = ~n21537 & n41992 ;
  assign n41994 = ( n5023 & ~n7494 ) | ( n5023 & n25327 ) | ( ~n7494 & n25327 ) ;
  assign n41995 = n28662 | n41994 ;
  assign n41996 = n31836 ^ n21482 ^ 1'b0 ;
  assign n41997 = x185 & n18712 ;
  assign n41998 = ~n41996 & n41997 ;
  assign n41999 = n1451 & n23304 ;
  assign n42000 = n41999 ^ n13006 ^ 1'b0 ;
  assign n42001 = n13391 | n13437 ;
  assign n42002 = n42000 & ~n42001 ;
  assign n42003 = n8165 | n42002 ;
  assign n42004 = n42003 ^ n25029 ^ 1'b0 ;
  assign n42005 = n9495 & n11450 ;
  assign n42006 = ~n7199 & n42005 ;
  assign n42007 = n42006 ^ n2297 ^ 1'b0 ;
  assign n42008 = n29162 & ~n42007 ;
  assign n42009 = n34297 ^ n18892 ^ n5759 ;
  assign n42010 = n42009 ^ n4602 ^ 1'b0 ;
  assign n42011 = n579 & ~n12216 ;
  assign n42012 = n42011 ^ n26089 ^ 1'b0 ;
  assign n42013 = n19459 | n42012 ;
  assign n42014 = n42010 | n42013 ;
  assign n42015 = ( n18026 & ~n35174 ) | ( n18026 & n42014 ) | ( ~n35174 & n42014 ) ;
  assign n42016 = n12817 ^ n8728 ^ 1'b0 ;
  assign n42017 = n970 | n42016 ;
  assign n42018 = n2458 ^ n1261 ^ 1'b0 ;
  assign n42019 = n10094 | n42018 ;
  assign n42020 = n42019 ^ n2903 ^ 1'b0 ;
  assign n42021 = n5719 & n38883 ;
  assign n42022 = n38236 ^ n923 ^ 1'b0 ;
  assign n42023 = n35276 ^ n15571 ^ 1'b0 ;
  assign n42024 = n3654 ^ n894 ^ 1'b0 ;
  assign n42025 = n42024 ^ n8196 ^ 1'b0 ;
  assign n42026 = n19708 & n42025 ;
  assign n42027 = n20913 ^ n15914 ^ 1'b0 ;
  assign n42032 = n14059 & n28668 ;
  assign n42033 = n4748 & n42032 ;
  assign n42031 = n1244 | n2216 ;
  assign n42034 = n42033 ^ n42031 ^ 1'b0 ;
  assign n42028 = n814 | n34168 ;
  assign n42029 = n42028 ^ n26593 ^ 1'b0 ;
  assign n42030 = n4404 | n42029 ;
  assign n42035 = n42034 ^ n42030 ^ 1'b0 ;
  assign n42036 = ~n3560 & n26787 ;
  assign n42037 = n16241 | n28321 ;
  assign n42038 = n12138 ^ n4642 ^ 1'b0 ;
  assign n42039 = n2214 & n42038 ;
  assign n42040 = n42039 ^ n17843 ^ 1'b0 ;
  assign n42041 = n42037 & n42040 ;
  assign n42042 = x27 & n7222 ;
  assign n42043 = n23130 & n42042 ;
  assign n42044 = n14044 | n42043 ;
  assign n42045 = n3725 | n42044 ;
  assign n42046 = n20480 ^ n12165 ^ 1'b0 ;
  assign n42047 = ~n9074 & n42046 ;
  assign n42048 = n42047 ^ n36838 ^ n10408 ;
  assign n42049 = n9758 | n15518 ;
  assign n42050 = n16989 & n42049 ;
  assign n42051 = n591 & ~n13630 ;
  assign n42052 = ~x146 & n42051 ;
  assign n42053 = n42052 ^ n40278 ^ 1'b0 ;
  assign n42054 = n27419 & n40656 ;
  assign n42055 = n6742 & n42054 ;
  assign n42056 = n29979 ^ n2848 ^ 1'b0 ;
  assign n42057 = n20175 & ~n42056 ;
  assign n42058 = n18629 & n28421 ;
  assign n42059 = ~n42057 & n42058 ;
  assign n42060 = n8174 & n28333 ;
  assign n42061 = ~n9098 & n42060 ;
  assign n42062 = n42059 & n42061 ;
  assign n42063 = n29517 ^ n16615 ^ 1'b0 ;
  assign n42064 = n5919 | n42063 ;
  assign n42065 = ( ~n20156 & n32623 ) | ( ~n20156 & n37415 ) | ( n32623 & n37415 ) ;
  assign n42071 = n7670 & ~n16943 ;
  assign n42072 = ~n3296 & n42071 ;
  assign n42073 = n6789 & ~n42072 ;
  assign n42074 = n10250 & n42073 ;
  assign n42067 = ( n4115 & n5175 ) | ( n4115 & ~n6632 ) | ( n5175 & ~n6632 ) ;
  assign n42068 = ( n15300 & ~n27968 ) | ( n15300 & n42067 ) | ( ~n27968 & n42067 ) ;
  assign n42066 = ~n21623 & n29040 ;
  assign n42069 = n42068 ^ n42066 ^ 1'b0 ;
  assign n42070 = n42069 ^ n30723 ^ n2936 ;
  assign n42075 = n42074 ^ n42070 ^ 1'b0 ;
  assign n42076 = n293 | n6555 ;
  assign n42077 = n32933 | n42076 ;
  assign n42078 = n12554 & ~n20896 ;
  assign n42079 = n4983 & ~n26880 ;
  assign n42080 = n7849 | n15937 ;
  assign n42081 = n904 & n42080 ;
  assign n42082 = ~n10103 & n27715 ;
  assign n42083 = n42082 ^ n5754 ^ 1'b0 ;
  assign n42084 = n31150 | n42083 ;
  assign n42085 = n42084 ^ n24941 ^ 1'b0 ;
  assign n42086 = n40910 ^ n13327 ^ 1'b0 ;
  assign n42087 = n8114 & n8302 ;
  assign n42088 = n42087 ^ n13020 ^ 1'b0 ;
  assign n42089 = n42088 ^ n29972 ^ 1'b0 ;
  assign n42090 = n42089 ^ n26520 ^ x208 ;
  assign n42091 = ~n14961 & n22685 ;
  assign n42092 = ( ~n12891 & n20450 ) | ( ~n12891 & n42091 ) | ( n20450 & n42091 ) ;
  assign n42093 = ~n7298 & n42092 ;
  assign n42094 = n1333 & ~n1803 ;
  assign n42095 = n22905 ^ n13995 ^ 1'b0 ;
  assign n42096 = n1665 & n8004 ;
  assign n42097 = n3785 | n42096 ;
  assign n42098 = n42097 ^ n11014 ^ 1'b0 ;
  assign n42099 = ~n12524 & n31911 ;
  assign n42100 = ~n42098 & n42099 ;
  assign n42101 = n24702 ^ n1501 ^ 1'b0 ;
  assign n42102 = ( n25497 & n35358 ) | ( n25497 & ~n42101 ) | ( n35358 & ~n42101 ) ;
  assign n42103 = n3054 & n38167 ;
  assign n42104 = n860 & ~n42103 ;
  assign n42105 = ~n15637 & n38647 ;
  assign n42106 = n33446 ^ n18444 ^ 1'b0 ;
  assign n42107 = n26400 ^ n2184 ^ 1'b0 ;
  assign n42108 = n21749 | n42107 ;
  assign n42109 = n1590 & n8914 ;
  assign n42110 = n31593 ^ n1801 ^ 1'b0 ;
  assign n42111 = n34957 | n42110 ;
  assign n42112 = n34728 ^ n312 ^ 1'b0 ;
  assign n42113 = ~n2506 & n34941 ;
  assign n42114 = n42113 ^ n35450 ^ 1'b0 ;
  assign n42115 = n13003 & n42114 ;
  assign n42116 = n42115 ^ n9964 ^ 1'b0 ;
  assign n42117 = n5704 & ~n21994 ;
  assign n42118 = n40444 ^ n35979 ^ 1'b0 ;
  assign n42119 = n12222 & n32305 ;
  assign n42120 = ~n29904 & n42119 ;
  assign n42121 = n1105 | n13636 ;
  assign n42122 = ( ~n20293 & n33788 ) | ( ~n20293 & n38811 ) | ( n33788 & n38811 ) ;
  assign n42123 = n1795 & ~n42122 ;
  assign n42124 = ~n13448 & n42123 ;
  assign n42125 = n2643 & ~n13960 ;
  assign n42126 = ( n8495 & ~n12874 ) | ( n8495 & n42125 ) | ( ~n12874 & n42125 ) ;
  assign n42127 = n26243 ^ n5992 ^ 1'b0 ;
  assign n42128 = n21949 & n42127 ;
  assign n42129 = n5775 & n38599 ;
  assign n42130 = n11905 ^ n794 ^ 1'b0 ;
  assign n42131 = n42130 ^ n23005 ^ n10961 ;
  assign n42132 = n7877 ^ n4898 ^ 1'b0 ;
  assign n42133 = n4632 | n42132 ;
  assign n42134 = n6998 & n31205 ;
  assign n42135 = n42134 ^ n1903 ^ 1'b0 ;
  assign n42136 = n18673 | n42135 ;
  assign n42137 = n9205 | n31303 ;
  assign n42138 = n9059 & n29902 ;
  assign n42139 = n17919 | n24969 ;
  assign n42140 = n20737 | n42139 ;
  assign n42141 = n42140 ^ n16791 ^ 1'b0 ;
  assign n42142 = n13972 | n31836 ;
  assign n42143 = n42142 ^ n5509 ^ 1'b0 ;
  assign n42144 = n42143 ^ n12059 ^ 1'b0 ;
  assign n42145 = n42144 ^ n24032 ^ 1'b0 ;
  assign n42146 = n12476 ^ n1557 ^ 1'b0 ;
  assign n42147 = n9014 ^ n2043 ^ 1'b0 ;
  assign n42148 = n13679 & n42147 ;
  assign n42149 = n14812 & n38179 ;
  assign n42150 = n15773 ^ n8835 ^ x254 ;
  assign n42151 = n20998 ^ n20220 ^ n2170 ;
  assign n42152 = n15119 & n40988 ;
  assign n42153 = n42152 ^ x163 ^ 1'b0 ;
  assign n42155 = n15385 ^ n3195 ^ 1'b0 ;
  assign n42156 = n8867 & ~n42155 ;
  assign n42154 = n16006 & ~n40178 ;
  assign n42157 = n42156 ^ n42154 ^ 1'b0 ;
  assign n42158 = n3768 | n11467 ;
  assign n42159 = n40950 | n42158 ;
  assign n42160 = n11747 | n16068 ;
  assign n42161 = n42160 ^ n12320 ^ 1'b0 ;
  assign n42162 = n19983 ^ n5522 ^ 1'b0 ;
  assign n42163 = n42161 | n42162 ;
  assign n42164 = n5259 & ~n37606 ;
  assign n42165 = n42164 ^ n38845 ^ 1'b0 ;
  assign n42166 = n11134 ^ n4008 ^ 1'b0 ;
  assign n42167 = n42165 | n42166 ;
  assign n42168 = n42167 ^ n25776 ^ 1'b0 ;
  assign n42169 = n2618 & ~n26458 ;
  assign n42170 = n29922 ^ n2463 ^ 1'b0 ;
  assign n42171 = n36601 & ~n42170 ;
  assign n42172 = n11691 | n16934 ;
  assign n42173 = ~n4258 & n7580 ;
  assign n42174 = n20362 ^ n8551 ^ n3873 ;
  assign n42175 = n14816 ^ n1269 ^ 1'b0 ;
  assign n42176 = n2167 & ~n42175 ;
  assign n42177 = n42176 ^ n20585 ^ n3866 ;
  assign n42178 = ~n37249 & n42177 ;
  assign n42179 = n3674 & ~n41228 ;
  assign n42180 = x218 & ~n13941 ;
  assign n42181 = n38417 ^ n12287 ^ n6836 ;
  assign n42182 = n8312 ^ n8145 ^ 1'b0 ;
  assign n42183 = n9885 | n42182 ;
  assign n42184 = n6415 | n28897 ;
  assign n42185 = n1624 & ~n15798 ;
  assign n42186 = n42185 ^ n7036 ^ 1'b0 ;
  assign n42187 = ( n12903 & n19258 ) | ( n12903 & n42186 ) | ( n19258 & n42186 ) ;
  assign n42188 = n19915 | n25739 ;
  assign n42189 = ~n14014 & n38372 ;
  assign n42190 = ~n8251 & n14311 ;
  assign n42191 = ~n37995 & n42190 ;
  assign n42192 = n23331 ^ n10731 ^ 1'b0 ;
  assign n42193 = n19186 & n42192 ;
  assign n42194 = n15337 ^ n4843 ^ 1'b0 ;
  assign n42195 = n4914 & ~n42194 ;
  assign n42196 = n8116 ^ n1095 ^ 1'b0 ;
  assign n42197 = n11803 & n29886 ;
  assign n42198 = n2537 & ~n34231 ;
  assign n42199 = n42198 ^ n8691 ^ 1'b0 ;
  assign n42200 = n24139 & n25246 ;
  assign n42201 = n42199 | n42200 ;
  assign n42202 = ~n3873 & n25457 ;
  assign n42203 = n4688 | n21304 ;
  assign n42204 = n19310 & ~n42203 ;
  assign n42205 = n19822 & n29866 ;
  assign n42206 = n3560 | n42205 ;
  assign n42207 = n42204 & ~n42206 ;
  assign n42208 = n1208 | n33524 ;
  assign n42209 = n16791 & ~n42208 ;
  assign n42210 = n42209 ^ n19207 ^ 1'b0 ;
  assign n42211 = ~n12804 & n34076 ;
  assign n42212 = n20505 ^ n5232 ^ n4976 ;
  assign n42213 = n28643 & ~n34285 ;
  assign n42214 = x52 | n18828 ;
  assign n42215 = n1328 & n13222 ;
  assign n42216 = n42214 & n42215 ;
  assign n42217 = n32045 | n37300 ;
  assign n42218 = n30465 | n42217 ;
  assign n42219 = ~n7867 & n42218 ;
  assign n42220 = n42219 ^ n7627 ^ 1'b0 ;
  assign n42221 = n3823 & ~n13142 ;
  assign n42222 = ~n32822 & n42221 ;
  assign n42223 = n31595 ^ n19383 ^ 1'b0 ;
  assign n42224 = n42222 | n42223 ;
  assign n42225 = n6968 ^ n3446 ^ 1'b0 ;
  assign n42226 = ~n12961 & n42225 ;
  assign n42227 = n34317 ^ n12736 ^ 1'b0 ;
  assign n42228 = n9958 & n42227 ;
  assign n42229 = n9635 & ~n10744 ;
  assign n42230 = n7515 | n15733 ;
  assign n42231 = n17323 & ~n42230 ;
  assign n42232 = n42229 & n42231 ;
  assign n42233 = n1525 | n19011 ;
  assign n42234 = n42233 ^ n23017 ^ n2324 ;
  assign n42235 = ~n9603 & n31977 ;
  assign n42236 = n42235 ^ n41121 ^ 1'b0 ;
  assign n42237 = n30333 ^ n1778 ^ 1'b0 ;
  assign n42238 = ~n6632 & n42237 ;
  assign n42239 = ~n7803 & n14014 ;
  assign n42240 = n11804 ^ n558 ^ 1'b0 ;
  assign n42241 = n35957 & ~n42240 ;
  assign n42242 = n12150 & n42241 ;
  assign n42243 = n14423 ^ n2436 ^ 1'b0 ;
  assign n42244 = n8219 | n21244 ;
  assign n42245 = n42244 ^ n30778 ^ 1'b0 ;
  assign n42246 = n18478 ^ n4069 ^ 1'b0 ;
  assign n42247 = n29489 & n42246 ;
  assign n42248 = n42245 & n42247 ;
  assign n42249 = n42248 ^ n24399 ^ 1'b0 ;
  assign n42250 = ~n2249 & n23898 ;
  assign n42251 = n4626 & n42250 ;
  assign n42252 = n39759 ^ n5341 ^ 1'b0 ;
  assign n42253 = n5802 & n41489 ;
  assign n42254 = n42253 ^ n411 ^ 1'b0 ;
  assign n42255 = x154 & ~n42254 ;
  assign y0 = x3 ;
  assign y1 = x6 ;
  assign y2 = x8 ;
  assign y3 = x9 ;
  assign y4 = x11 ;
  assign y5 = x13 ;
  assign y6 = x16 ;
  assign y7 = x19 ;
  assign y8 = x21 ;
  assign y9 = x27 ;
  assign y10 = x28 ;
  assign y11 = x30 ;
  assign y12 = x32 ;
  assign y13 = x33 ;
  assign y14 = x37 ;
  assign y15 = x39 ;
  assign y16 = x41 ;
  assign y17 = x45 ;
  assign y18 = x46 ;
  assign y19 = x52 ;
  assign y20 = x55 ;
  assign y21 = x58 ;
  assign y22 = x61 ;
  assign y23 = x65 ;
  assign y24 = x67 ;
  assign y25 = x74 ;
  assign y26 = x76 ;
  assign y27 = x83 ;
  assign y28 = x86 ;
  assign y29 = x88 ;
  assign y30 = x89 ;
  assign y31 = x90 ;
  assign y32 = x109 ;
  assign y33 = x120 ;
  assign y34 = x122 ;
  assign y35 = x123 ;
  assign y36 = x127 ;
  assign y37 = x128 ;
  assign y38 = x129 ;
  assign y39 = x131 ;
  assign y40 = x132 ;
  assign y41 = x135 ;
  assign y42 = x136 ;
  assign y43 = x137 ;
  assign y44 = x149 ;
  assign y45 = x160 ;
  assign y46 = x162 ;
  assign y47 = x166 ;
  assign y48 = x171 ;
  assign y49 = x172 ;
  assign y50 = x174 ;
  assign y51 = x179 ;
  assign y52 = x186 ;
  assign y53 = x188 ;
  assign y54 = x190 ;
  assign y55 = x197 ;
  assign y56 = x201 ;
  assign y57 = x202 ;
  assign y58 = x206 ;
  assign y59 = x207 ;
  assign y60 = x210 ;
  assign y61 = x211 ;
  assign y62 = x215 ;
  assign y63 = x218 ;
  assign y64 = x221 ;
  assign y65 = x222 ;
  assign y66 = x227 ;
  assign y67 = x228 ;
  assign y68 = x230 ;
  assign y69 = x231 ;
  assign y70 = x248 ;
  assign y71 = x250 ;
  assign y72 = x251 ;
  assign y73 = x253 ;
  assign y74 = ~n256 ;
  assign y75 = ~n258 ;
  assign y76 = n260 ;
  assign y77 = n262 ;
  assign y78 = n263 ;
  assign y79 = ~1'b0 ;
  assign y80 = n266 ;
  assign y81 = ~n267 ;
  assign y82 = ~1'b0 ;
  assign y83 = n268 ;
  assign y84 = ~n270 ;
  assign y85 = n271 ;
  assign y86 = n272 ;
  assign y87 = ~n274 ;
  assign y88 = ~n277 ;
  assign y89 = n279 ;
  assign y90 = ~1'b0 ;
  assign y91 = ~n281 ;
  assign y92 = n283 ;
  assign y93 = n289 ;
  assign y94 = ~n291 ;
  assign y95 = n294 ;
  assign y96 = ~n296 ;
  assign y97 = ~n298 ;
  assign y98 = n302 ;
  assign y99 = ~1'b0 ;
  assign y100 = ~n306 ;
  assign y101 = ~1'b0 ;
  assign y102 = n310 ;
  assign y103 = ~n312 ;
  assign y104 = ~n314 ;
  assign y105 = ~n315 ;
  assign y106 = 1'b0 ;
  assign y107 = ~n317 ;
  assign y108 = ~n320 ;
  assign y109 = ~n329 ;
  assign y110 = ~n332 ;
  assign y111 = ~1'b0 ;
  assign y112 = ~n334 ;
  assign y113 = n336 ;
  assign y114 = ~n338 ;
  assign y115 = ~1'b0 ;
  assign y116 = ~n340 ;
  assign y117 = ~n344 ;
  assign y118 = ~n348 ;
  assign y119 = ~1'b0 ;
  assign y120 = ~1'b0 ;
  assign y121 = ~n349 ;
  assign y122 = n351 ;
  assign y123 = n355 ;
  assign y124 = n359 ;
  assign y125 = ~n361 ;
  assign y126 = ~n364 ;
  assign y127 = ~1'b0 ;
  assign y128 = n366 ;
  assign y129 = ~1'b0 ;
  assign y130 = ~1'b0 ;
  assign y131 = n367 ;
  assign y132 = ~n369 ;
  assign y133 = ~1'b0 ;
  assign y134 = ~n370 ;
  assign y135 = ~n376 ;
  assign y136 = n378 ;
  assign y137 = n387 ;
  assign y138 = ~n389 ;
  assign y139 = n395 ;
  assign y140 = ~n397 ;
  assign y141 = ~n399 ;
  assign y142 = n406 ;
  assign y143 = n409 ;
  assign y144 = ~n411 ;
  assign y145 = n415 ;
  assign y146 = n417 ;
  assign y147 = ~n419 ;
  assign y148 = n420 ;
  assign y149 = ~n423 ;
  assign y150 = ~1'b0 ;
  assign y151 = n424 ;
  assign y152 = ~1'b0 ;
  assign y153 = ~n426 ;
  assign y154 = n431 ;
  assign y155 = ~1'b0 ;
  assign y156 = n433 ;
  assign y157 = ~n437 ;
  assign y158 = n445 ;
  assign y159 = ~n446 ;
  assign y160 = ~1'b0 ;
  assign y161 = n449 ;
  assign y162 = n453 ;
  assign y163 = n459 ;
  assign y164 = ~1'b0 ;
  assign y165 = ~n461 ;
  assign y166 = ~n469 ;
  assign y167 = ~n475 ;
  assign y168 = ~n483 ;
  assign y169 = ~n490 ;
  assign y170 = ~1'b0 ;
  assign y171 = ~1'b0 ;
  assign y172 = ~1'b0 ;
  assign y173 = ~n491 ;
  assign y174 = ~n494 ;
  assign y175 = ~n505 ;
  assign y176 = n510 ;
  assign y177 = ~1'b0 ;
  assign y178 = ~n511 ;
  assign y179 = ~n514 ;
  assign y180 = ~n520 ;
  assign y181 = ~n522 ;
  assign y182 = ~1'b0 ;
  assign y183 = n523 ;
  assign y184 = n530 ;
  assign y185 = n534 ;
  assign y186 = ~x6 ;
  assign y187 = ~n535 ;
  assign y188 = n537 ;
  assign y189 = ~1'b0 ;
  assign y190 = ~1'b0 ;
  assign y191 = ~1'b0 ;
  assign y192 = n545 ;
  assign y193 = ~1'b0 ;
  assign y194 = n547 ;
  assign y195 = ~n548 ;
  assign y196 = ~n552 ;
  assign y197 = ~1'b0 ;
  assign y198 = ~n555 ;
  assign y199 = n558 ;
  assign y200 = ~n564 ;
  assign y201 = n572 ;
  assign y202 = ~1'b0 ;
  assign y203 = ~n574 ;
  assign y204 = ~n577 ;
  assign y205 = n580 ;
  assign y206 = ~1'b0 ;
  assign y207 = ~1'b0 ;
  assign y208 = ~n587 ;
  assign y209 = ~1'b0 ;
  assign y210 = ~n589 ;
  assign y211 = n592 ;
  assign y212 = ~n596 ;
  assign y213 = n597 ;
  assign y214 = ~1'b0 ;
  assign y215 = ~n606 ;
  assign y216 = ~n618 ;
  assign y217 = ~n622 ;
  assign y218 = ~n624 ;
  assign y219 = n625 ;
  assign y220 = ~n627 ;
  assign y221 = n634 ;
  assign y222 = ~n637 ;
  assign y223 = ~n638 ;
  assign y224 = ~1'b0 ;
  assign y225 = ~n643 ;
  assign y226 = ~n645 ;
  assign y227 = ~n651 ;
  assign y228 = ~n655 ;
  assign y229 = n659 ;
  assign y230 = n663 ;
  assign y231 = ~1'b0 ;
  assign y232 = n666 ;
  assign y233 = ~1'b0 ;
  assign y234 = ~n668 ;
  assign y235 = ~n673 ;
  assign y236 = ~1'b0 ;
  assign y237 = ~n679 ;
  assign y238 = ~1'b0 ;
  assign y239 = n703 ;
  assign y240 = ~n705 ;
  assign y241 = ~1'b0 ;
  assign y242 = ~1'b0 ;
  assign y243 = n707 ;
  assign y244 = ~n709 ;
  assign y245 = ~n710 ;
  assign y246 = ~1'b0 ;
  assign y247 = n713 ;
  assign y248 = ~n714 ;
  assign y249 = n518 ;
  assign y250 = n718 ;
  assign y251 = ~1'b0 ;
  assign y252 = ~n720 ;
  assign y253 = ~n723 ;
  assign y254 = ~n725 ;
  assign y255 = ~1'b0 ;
  assign y256 = n729 ;
  assign y257 = n732 ;
  assign y258 = n735 ;
  assign y259 = n737 ;
  assign y260 = ~1'b0 ;
  assign y261 = ~1'b0 ;
  assign y262 = n739 ;
  assign y263 = ~1'b0 ;
  assign y264 = n742 ;
  assign y265 = ~1'b0 ;
  assign y266 = ~1'b0 ;
  assign y267 = n747 ;
  assign y268 = ~n751 ;
  assign y269 = ~n754 ;
  assign y270 = ~n755 ;
  assign y271 = n757 ;
  assign y272 = n763 ;
  assign y273 = ~1'b0 ;
  assign y274 = ~n765 ;
  assign y275 = n769 ;
  assign y276 = n772 ;
  assign y277 = ~1'b0 ;
  assign y278 = ~n787 ;
  assign y279 = ~n792 ;
  assign y280 = ~n797 ;
  assign y281 = n808 ;
  assign y282 = ~n466 ;
  assign y283 = ~n810 ;
  assign y284 = ~n812 ;
  assign y285 = ~n813 ;
  assign y286 = n815 ;
  assign y287 = n821 ;
  assign y288 = ~1'b0 ;
  assign y289 = n826 ;
  assign y290 = ~n828 ;
  assign y291 = ~n830 ;
  assign y292 = n836 ;
  assign y293 = n839 ;
  assign y294 = ~1'b0 ;
  assign y295 = ~n851 ;
  assign y296 = ~n858 ;
  assign y297 = n862 ;
  assign y298 = ~n863 ;
  assign y299 = ~1'b0 ;
  assign y300 = ~n871 ;
  assign y301 = n705 ;
  assign y302 = ~n874 ;
  assign y303 = ~1'b0 ;
  assign y304 = ~n876 ;
  assign y305 = n877 ;
  assign y306 = ~n879 ;
  assign y307 = ~n882 ;
  assign y308 = ~n886 ;
  assign y309 = n789 ;
  assign y310 = ~n888 ;
  assign y311 = n890 ;
  assign y312 = n891 ;
  assign y313 = n894 ;
  assign y314 = ~n897 ;
  assign y315 = n906 ;
  assign y316 = n909 ;
  assign y317 = ~1'b0 ;
  assign y318 = ~1'b0 ;
  assign y319 = n914 ;
  assign y320 = n915 ;
  assign y321 = n921 ;
  assign y322 = n925 ;
  assign y323 = n930 ;
  assign y324 = ~n932 ;
  assign y325 = n937 ;
  assign y326 = ~n941 ;
  assign y327 = ~1'b0 ;
  assign y328 = n946 ;
  assign y329 = n949 ;
  assign y330 = n951 ;
  assign y331 = ~1'b0 ;
  assign y332 = ~1'b0 ;
  assign y333 = ~n953 ;
  assign y334 = ~n547 ;
  assign y335 = n954 ;
  assign y336 = ~1'b0 ;
  assign y337 = ~1'b0 ;
  assign y338 = ~1'b0 ;
  assign y339 = n958 ;
  assign y340 = ~n959 ;
  assign y341 = ~n964 ;
  assign y342 = n968 ;
  assign y343 = ~n969 ;
  assign y344 = n970 ;
  assign y345 = n971 ;
  assign y346 = ~n977 ;
  assign y347 = ~1'b0 ;
  assign y348 = ~n978 ;
  assign y349 = n982 ;
  assign y350 = ~n986 ;
  assign y351 = n987 ;
  assign y352 = ~n988 ;
  assign y353 = ~1'b0 ;
  assign y354 = n991 ;
  assign y355 = ~n992 ;
  assign y356 = ~1'b0 ;
  assign y357 = ~1'b0 ;
  assign y358 = ~n994 ;
  assign y359 = ~1'b0 ;
  assign y360 = ~1'b0 ;
  assign y361 = ~1'b0 ;
  assign y362 = ~n995 ;
  assign y363 = ~n997 ;
  assign y364 = ~1'b0 ;
  assign y365 = ~n589 ;
  assign y366 = ~n998 ;
  assign y367 = ~n1004 ;
  assign y368 = ~n1014 ;
  assign y369 = ~1'b0 ;
  assign y370 = ~n1021 ;
  assign y371 = n1023 ;
  assign y372 = n1025 ;
  assign y373 = ~1'b0 ;
  assign y374 = ~1'b0 ;
  assign y375 = ~1'b0 ;
  assign y376 = ~n1036 ;
  assign y377 = n1037 ;
  assign y378 = ~1'b0 ;
  assign y379 = n1045 ;
  assign y380 = ~n1051 ;
  assign y381 = ~1'b0 ;
  assign y382 = ~n1059 ;
  assign y383 = ~n1062 ;
  assign y384 = n1070 ;
  assign y385 = ~1'b0 ;
  assign y386 = ~n1071 ;
  assign y387 = ~n1075 ;
  assign y388 = ~n1078 ;
  assign y389 = n1088 ;
  assign y390 = n1091 ;
  assign y391 = n1092 ;
  assign y392 = n1093 ;
  assign y393 = ~1'b0 ;
  assign y394 = ~n1096 ;
  assign y395 = ~1'b0 ;
  assign y396 = ~n1098 ;
  assign y397 = ~1'b0 ;
  assign y398 = ~n1099 ;
  assign y399 = ~n1105 ;
  assign y400 = ~n1114 ;
  assign y401 = ~n1116 ;
  assign y402 = n1123 ;
  assign y403 = ~1'b0 ;
  assign y404 = n1124 ;
  assign y405 = ~1'b0 ;
  assign y406 = ~n1125 ;
  assign y407 = ~n1130 ;
  assign y408 = ~1'b0 ;
  assign y409 = n1133 ;
  assign y410 = n1134 ;
  assign y411 = n1135 ;
  assign y412 = ~n1140 ;
  assign y413 = x162 ;
  assign y414 = ~n1149 ;
  assign y415 = ~n1153 ;
  assign y416 = ~n1159 ;
  assign y417 = ~n1163 ;
  assign y418 = n1168 ;
  assign y419 = n1174 ;
  assign y420 = ~n1175 ;
  assign y421 = ~1'b0 ;
  assign y422 = ~n1176 ;
  assign y423 = ~n1177 ;
  assign y424 = n1182 ;
  assign y425 = n1186 ;
  assign y426 = ~1'b0 ;
  assign y427 = n1190 ;
  assign y428 = ~n1192 ;
  assign y429 = ~n1197 ;
  assign y430 = ~1'b0 ;
  assign y431 = ~1'b0 ;
  assign y432 = n631 ;
  assign y433 = ~1'b0 ;
  assign y434 = ~n1199 ;
  assign y435 = ~n1204 ;
  assign y436 = ~n1206 ;
  assign y437 = n1213 ;
  assign y438 = n1217 ;
  assign y439 = n1223 ;
  assign y440 = ~n1227 ;
  assign y441 = n1230 ;
  assign y442 = n1231 ;
  assign y443 = ~1'b0 ;
  assign y444 = ~1'b0 ;
  assign y445 = n1238 ;
  assign y446 = n1245 ;
  assign y447 = ~x247 ;
  assign y448 = n445 ;
  assign y449 = n1249 ;
  assign y450 = ~1'b0 ;
  assign y451 = n1252 ;
  assign y452 = ~1'b0 ;
  assign y453 = ~n1255 ;
  assign y454 = ~n1261 ;
  assign y455 = n1262 ;
  assign y456 = ~1'b0 ;
  assign y457 = ~1'b0 ;
  assign y458 = ~n1267 ;
  assign y459 = ~n1271 ;
  assign y460 = ~n1276 ;
  assign y461 = ~n938 ;
  assign y462 = n1278 ;
  assign y463 = ~n1279 ;
  assign y464 = ~1'b0 ;
  assign y465 = ~n1284 ;
  assign y466 = ~1'b0 ;
  assign y467 = ~1'b0 ;
  assign y468 = ~1'b0 ;
  assign y469 = ~1'b0 ;
  assign y470 = ~1'b0 ;
  assign y471 = ~n1288 ;
  assign y472 = n1290 ;
  assign y473 = n1294 ;
  assign y474 = ~1'b0 ;
  assign y475 = n1298 ;
  assign y476 = n1300 ;
  assign y477 = ~1'b0 ;
  assign y478 = ~n1301 ;
  assign y479 = ~n1303 ;
  assign y480 = ~1'b0 ;
  assign y481 = n1311 ;
  assign y482 = n1316 ;
  assign y483 = ~n1317 ;
  assign y484 = n1318 ;
  assign y485 = n1319 ;
  assign y486 = n1322 ;
  assign y487 = ~n1332 ;
  assign y488 = n1333 ;
  assign y489 = n1338 ;
  assign y490 = ~n1340 ;
  assign y491 = ~n908 ;
  assign y492 = n1344 ;
  assign y493 = n1346 ;
  assign y494 = ~n1349 ;
  assign y495 = ~1'b0 ;
  assign y496 = ~n1352 ;
  assign y497 = ~n1354 ;
  assign y498 = n1358 ;
  assign y499 = ~n1328 ;
  assign y500 = ~1'b0 ;
  assign y501 = ~n1361 ;
  assign y502 = ~n1362 ;
  assign y503 = ~n1276 ;
  assign y504 = ~n1364 ;
  assign y505 = ~1'b0 ;
  assign y506 = n1366 ;
  assign y507 = ~n1368 ;
  assign y508 = ~n1369 ;
  assign y509 = ~1'b0 ;
  assign y510 = ~1'b0 ;
  assign y511 = ~n1378 ;
  assign y512 = ~1'b0 ;
  assign y513 = n1379 ;
  assign y514 = n1383 ;
  assign y515 = n1384 ;
  assign y516 = ~n1385 ;
  assign y517 = ~1'b0 ;
  assign y518 = n1387 ;
  assign y519 = n1388 ;
  assign y520 = n1389 ;
  assign y521 = n1392 ;
  assign y522 = n1395 ;
  assign y523 = ~1'b0 ;
  assign y524 = ~1'b0 ;
  assign y525 = ~n1400 ;
  assign y526 = ~n1402 ;
  assign y527 = ~n1404 ;
  assign y528 = ~n1254 ;
  assign y529 = ~n1405 ;
  assign y530 = n1406 ;
  assign y531 = n1413 ;
  assign y532 = ~n1422 ;
  assign y533 = ~n1428 ;
  assign y534 = ~n1432 ;
  assign y535 = n1435 ;
  assign y536 = ~n1439 ;
  assign y537 = ~n1440 ;
  assign y538 = n1456 ;
  assign y539 = n1457 ;
  assign y540 = ~n1458 ;
  assign y541 = 1'b0 ;
  assign y542 = ~n1463 ;
  assign y543 = n1039 ;
  assign y544 = ~n1465 ;
  assign y545 = n1466 ;
  assign y546 = n1249 ;
  assign y547 = ~n1467 ;
  assign y548 = n1470 ;
  assign y549 = ~n1473 ;
  assign y550 = ~1'b0 ;
  assign y551 = ~n1474 ;
  assign y552 = ~n627 ;
  assign y553 = ~n1475 ;
  assign y554 = n1478 ;
  assign y555 = n1328 ;
  assign y556 = ~n1480 ;
  assign y557 = ~1'b0 ;
  assign y558 = n1481 ;
  assign y559 = ~1'b0 ;
  assign y560 = 1'b0 ;
  assign y561 = ~n1489 ;
  assign y562 = ~1'b0 ;
  assign y563 = ~n1492 ;
  assign y564 = ~n1504 ;
  assign y565 = ~n1505 ;
  assign y566 = n1506 ;
  assign y567 = n1510 ;
  assign y568 = n1513 ;
  assign y569 = n1517 ;
  assign y570 = n1219 ;
  assign y571 = ~1'b0 ;
  assign y572 = ~n1519 ;
  assign y573 = n1528 ;
  assign y574 = ~1'b0 ;
  assign y575 = n1536 ;
  assign y576 = ~1'b0 ;
  assign y577 = n1543 ;
  assign y578 = ~n1544 ;
  assign y579 = ~n1547 ;
  assign y580 = ~1'b0 ;
  assign y581 = n1548 ;
  assign y582 = n1550 ;
  assign y583 = ~n1295 ;
  assign y584 = ~n1553 ;
  assign y585 = ~n1562 ;
  assign y586 = n1563 ;
  assign y587 = ~1'b0 ;
  assign y588 = n1568 ;
  assign y589 = ~n1569 ;
  assign y590 = ~n276 ;
  assign y591 = n1573 ;
  assign y592 = ~n1575 ;
  assign y593 = ~n1586 ;
  assign y594 = n1369 ;
  assign y595 = n1588 ;
  assign y596 = n1591 ;
  assign y597 = ~n1592 ;
  assign y598 = n1596 ;
  assign y599 = n1600 ;
  assign y600 = n1608 ;
  assign y601 = ~1'b0 ;
  assign y602 = n1611 ;
  assign y603 = n1612 ;
  assign y604 = ~1'b0 ;
  assign y605 = ~1'b0 ;
  assign y606 = n1613 ;
  assign y607 = n1615 ;
  assign y608 = ~1'b0 ;
  assign y609 = ~1'b0 ;
  assign y610 = ~n1617 ;
  assign y611 = ~1'b0 ;
  assign y612 = n1622 ;
  assign y613 = ~1'b0 ;
  assign y614 = n1624 ;
  assign y615 = ~n1628 ;
  assign y616 = ~1'b0 ;
  assign y617 = ~n1630 ;
  assign y618 = n1634 ;
  assign y619 = n1635 ;
  assign y620 = ~1'b0 ;
  assign y621 = n1638 ;
  assign y622 = ~n1639 ;
  assign y623 = ~n1641 ;
  assign y624 = n1645 ;
  assign y625 = ~1'b0 ;
  assign y626 = ~n1654 ;
  assign y627 = ~1'b0 ;
  assign y628 = ~n1656 ;
  assign y629 = n1662 ;
  assign y630 = ~n1665 ;
  assign y631 = ~1'b0 ;
  assign y632 = n1669 ;
  assign y633 = ~1'b0 ;
  assign y634 = n1672 ;
  assign y635 = n1680 ;
  assign y636 = ~1'b0 ;
  assign y637 = n1682 ;
  assign y638 = ~1'b0 ;
  assign y639 = ~1'b0 ;
  assign y640 = n1623 ;
  assign y641 = ~1'b0 ;
  assign y642 = n604 ;
  assign y643 = ~1'b0 ;
  assign y644 = n1688 ;
  assign y645 = ~n1690 ;
  assign y646 = ~n1694 ;
  assign y647 = n1696 ;
  assign y648 = ~n1699 ;
  assign y649 = ~n1701 ;
  assign y650 = ~1'b0 ;
  assign y651 = ~n1048 ;
  assign y652 = ~n1709 ;
  assign y653 = ~n1718 ;
  assign y654 = n1721 ;
  assign y655 = n1726 ;
  assign y656 = ~n1727 ;
  assign y657 = ~n1729 ;
  assign y658 = n1730 ;
  assign y659 = ~n1731 ;
  assign y660 = ~n1733 ;
  assign y661 = ~1'b0 ;
  assign y662 = ~n1736 ;
  assign y663 = ~1'b0 ;
  assign y664 = ~n1741 ;
  assign y665 = n1742 ;
  assign y666 = ~n1744 ;
  assign y667 = n1746 ;
  assign y668 = n1748 ;
  assign y669 = ~1'b0 ;
  assign y670 = n1749 ;
  assign y671 = n1753 ;
  assign y672 = n1756 ;
  assign y673 = n1757 ;
  assign y674 = ~1'b0 ;
  assign y675 = n1759 ;
  assign y676 = ~1'b0 ;
  assign y677 = ~n1760 ;
  assign y678 = ~n1772 ;
  assign y679 = ~n1777 ;
  assign y680 = ~1'b0 ;
  assign y681 = ~n1780 ;
  assign y682 = ~1'b0 ;
  assign y683 = n1784 ;
  assign y684 = ~1'b0 ;
  assign y685 = ~n1789 ;
  assign y686 = ~n1791 ;
  assign y687 = n1793 ;
  assign y688 = ~1'b0 ;
  assign y689 = ~1'b0 ;
  assign y690 = n1796 ;
  assign y691 = n1798 ;
  assign y692 = ~n1801 ;
  assign y693 = n1807 ;
  assign y694 = x192 ;
  assign y695 = ~n1809 ;
  assign y696 = n1810 ;
  assign y697 = ~1'b0 ;
  assign y698 = ~1'b0 ;
  assign y699 = ~1'b0 ;
  assign y700 = ~1'b0 ;
  assign y701 = ~1'b0 ;
  assign y702 = ~n973 ;
  assign y703 = ~1'b0 ;
  assign y704 = n1814 ;
  assign y705 = ~n1820 ;
  assign y706 = n1822 ;
  assign y707 = ~n1826 ;
  assign y708 = n1832 ;
  assign y709 = n1843 ;
  assign y710 = ~1'b0 ;
  assign y711 = ~n1844 ;
  assign y712 = n1845 ;
  assign y713 = ~n1846 ;
  assign y714 = ~n1848 ;
  assign y715 = n1861 ;
  assign y716 = n1862 ;
  assign y717 = n1866 ;
  assign y718 = n1870 ;
  assign y719 = ~1'b0 ;
  assign y720 = ~1'b0 ;
  assign y721 = ~1'b0 ;
  assign y722 = ~n1873 ;
  assign y723 = ~1'b0 ;
  assign y724 = ~n1875 ;
  assign y725 = ~n1877 ;
  assign y726 = n1878 ;
  assign y727 = n1879 ;
  assign y728 = ~1'b0 ;
  assign y729 = ~1'b0 ;
  assign y730 = n1885 ;
  assign y731 = n1889 ;
  assign y732 = ~n1891 ;
  assign y733 = n1893 ;
  assign y734 = ~n1894 ;
  assign y735 = n1896 ;
  assign y736 = ~x175 ;
  assign y737 = ~n1898 ;
  assign y738 = ~1'b0 ;
  assign y739 = n1900 ;
  assign y740 = ~1'b0 ;
  assign y741 = ~1'b0 ;
  assign y742 = n1901 ;
  assign y743 = ~n1911 ;
  assign y744 = ~n1917 ;
  assign y745 = ~1'b0 ;
  assign y746 = ~1'b0 ;
  assign y747 = ~1'b0 ;
  assign y748 = ~1'b0 ;
  assign y749 = n1926 ;
  assign y750 = ~x172 ;
  assign y751 = ~n1929 ;
  assign y752 = ~n1933 ;
  assign y753 = ~n1936 ;
  assign y754 = n1944 ;
  assign y755 = n1947 ;
  assign y756 = ~1'b0 ;
  assign y757 = ~n1948 ;
  assign y758 = ~n1950 ;
  assign y759 = ~n1954 ;
  assign y760 = n1965 ;
  assign y761 = n1966 ;
  assign y762 = ~n905 ;
  assign y763 = ~1'b0 ;
  assign y764 = n1971 ;
  assign y765 = n1980 ;
  assign y766 = ~1'b0 ;
  assign y767 = n1983 ;
  assign y768 = n1856 ;
  assign y769 = ~1'b0 ;
  assign y770 = ~n1985 ;
  assign y771 = ~n1986 ;
  assign y772 = ~n1990 ;
  assign y773 = n1995 ;
  assign y774 = ~n1998 ;
  assign y775 = ~n2001 ;
  assign y776 = ~n2003 ;
  assign y777 = n2006 ;
  assign y778 = n2007 ;
  assign y779 = n2014 ;
  assign y780 = n2015 ;
  assign y781 = ~n2018 ;
  assign y782 = ~n2024 ;
  assign y783 = n2030 ;
  assign y784 = ~1'b0 ;
  assign y785 = ~1'b0 ;
  assign y786 = n2041 ;
  assign y787 = n2043 ;
  assign y788 = ~n2045 ;
  assign y789 = n2048 ;
  assign y790 = n2050 ;
  assign y791 = ~n2053 ;
  assign y792 = ~n627 ;
  assign y793 = ~n2054 ;
  assign y794 = ~1'b0 ;
  assign y795 = ~n2058 ;
  assign y796 = ~n2062 ;
  assign y797 = n2064 ;
  assign y798 = ~1'b0 ;
  assign y799 = ~1'b0 ;
  assign y800 = ~n2065 ;
  assign y801 = n2069 ;
  assign y802 = ~n2070 ;
  assign y803 = ~n2072 ;
  assign y804 = ~1'b0 ;
  assign y805 = ~n1376 ;
  assign y806 = ~x204 ;
  assign y807 = ~n2078 ;
  assign y808 = ~1'b0 ;
  assign y809 = n2082 ;
  assign y810 = n2083 ;
  assign y811 = ~1'b0 ;
  assign y812 = ~1'b0 ;
  assign y813 = n2091 ;
  assign y814 = ~n2093 ;
  assign y815 = ~1'b0 ;
  assign y816 = ~n2098 ;
  assign y817 = ~n2101 ;
  assign y818 = ~1'b0 ;
  assign y819 = n2102 ;
  assign y820 = ~n2103 ;
  assign y821 = ~n2105 ;
  assign y822 = ~1'b0 ;
  assign y823 = n2107 ;
  assign y824 = n2110 ;
  assign y825 = ~n2112 ;
  assign y826 = ~n2113 ;
  assign y827 = ~1'b0 ;
  assign y828 = n2114 ;
  assign y829 = n2116 ;
  assign y830 = n2123 ;
  assign y831 = ~n2137 ;
  assign y832 = ~1'b0 ;
  assign y833 = n2141 ;
  assign y834 = ~1'b0 ;
  assign y835 = ~1'b0 ;
  assign y836 = ~1'b0 ;
  assign y837 = ~1'b0 ;
  assign y838 = ~1'b0 ;
  assign y839 = ~n2142 ;
  assign y840 = ~1'b0 ;
  assign y841 = ~n2143 ;
  assign y842 = ~1'b0 ;
  assign y843 = n2146 ;
  assign y844 = ~n2149 ;
  assign y845 = n2155 ;
  assign y846 = n2159 ;
  assign y847 = ~1'b0 ;
  assign y848 = n2164 ;
  assign y849 = n2167 ;
  assign y850 = 1'b0 ;
  assign y851 = ~n2171 ;
  assign y852 = n2172 ;
  assign y853 = ~n2178 ;
  assign y854 = ~n2184 ;
  assign y855 = n2191 ;
  assign y856 = ~1'b0 ;
  assign y857 = ~1'b0 ;
  assign y858 = 1'b0 ;
  assign y859 = ~n2193 ;
  assign y860 = n2198 ;
  assign y861 = ~n1185 ;
  assign y862 = ~n1416 ;
  assign y863 = ~n2199 ;
  assign y864 = ~1'b0 ;
  assign y865 = n2200 ;
  assign y866 = ~n2203 ;
  assign y867 = n2214 ;
  assign y868 = ~n2215 ;
  assign y869 = ~n2216 ;
  assign y870 = ~n2221 ;
  assign y871 = n2224 ;
  assign y872 = ~1'b0 ;
  assign y873 = ~x107 ;
  assign y874 = ~n2225 ;
  assign y875 = ~n2226 ;
  assign y876 = n2227 ;
  assign y877 = n2228 ;
  assign y878 = n2231 ;
  assign y879 = ~n2237 ;
  assign y880 = ~n2242 ;
  assign y881 = ~n2243 ;
  assign y882 = ~n2244 ;
  assign y883 = n2245 ;
  assign y884 = ~n2249 ;
  assign y885 = n2256 ;
  assign y886 = n2257 ;
  assign y887 = n2258 ;
  assign y888 = ~1'b0 ;
  assign y889 = n2259 ;
  assign y890 = 1'b0 ;
  assign y891 = ~1'b0 ;
  assign y892 = ~1'b0 ;
  assign y893 = ~n2263 ;
  assign y894 = ~1'b0 ;
  assign y895 = ~1'b0 ;
  assign y896 = ~1'b0 ;
  assign y897 = ~1'b0 ;
  assign y898 = ~n2264 ;
  assign y899 = ~n2265 ;
  assign y900 = ~1'b0 ;
  assign y901 = n2268 ;
  assign y902 = ~1'b0 ;
  assign y903 = ~n2275 ;
  assign y904 = n2276 ;
  assign y905 = ~n2277 ;
  assign y906 = ~n2279 ;
  assign y907 = ~n2281 ;
  assign y908 = n2283 ;
  assign y909 = ~n2286 ;
  assign y910 = ~n2289 ;
  assign y911 = n2299 ;
  assign y912 = ~n2301 ;
  assign y913 = ~n2302 ;
  assign y914 = n2309 ;
  assign y915 = ~n2310 ;
  assign y916 = ~n2316 ;
  assign y917 = ~n2192 ;
  assign y918 = ~x107 ;
  assign y919 = n2317 ;
  assign y920 = ~1'b0 ;
  assign y921 = ~n1244 ;
  assign y922 = ~1'b0 ;
  assign y923 = n2320 ;
  assign y924 = ~n2322 ;
  assign y925 = ~x241 ;
  assign y926 = ~n2323 ;
  assign y927 = ~n2325 ;
  assign y928 = n2328 ;
  assign y929 = ~n2330 ;
  assign y930 = n2335 ;
  assign y931 = ~1'b0 ;
  assign y932 = ~n2343 ;
  assign y933 = ~1'b0 ;
  assign y934 = ~n2345 ;
  assign y935 = ~1'b0 ;
  assign y936 = ~1'b0 ;
  assign y937 = n2347 ;
  assign y938 = ~n2348 ;
  assign y939 = ~n2351 ;
  assign y940 = ~1'b0 ;
  assign y941 = ~n2355 ;
  assign y942 = n274 ;
  assign y943 = ~1'b0 ;
  assign y944 = ~n2357 ;
  assign y945 = n2358 ;
  assign y946 = n2362 ;
  assign y947 = ~n2367 ;
  assign y948 = ~1'b0 ;
  assign y949 = ~1'b0 ;
  assign y950 = ~n2368 ;
  assign y951 = ~1'b0 ;
  assign y952 = n2369 ;
  assign y953 = ~x169 ;
  assign y954 = ~n2370 ;
  assign y955 = ~n2371 ;
  assign y956 = n2372 ;
  assign y957 = ~n2374 ;
  assign y958 = n2375 ;
  assign y959 = ~1'b0 ;
  assign y960 = ~1'b0 ;
  assign y961 = ~n2376 ;
  assign y962 = n2378 ;
  assign y963 = n2380 ;
  assign y964 = ~n2387 ;
  assign y965 = ~n2389 ;
  assign y966 = ~n2395 ;
  assign y967 = n1958 ;
  assign y968 = ~n2399 ;
  assign y969 = ~1'b0 ;
  assign y970 = ~1'b0 ;
  assign y971 = 1'b0 ;
  assign y972 = ~1'b0 ;
  assign y973 = ~1'b0 ;
  assign y974 = ~n2400 ;
  assign y975 = ~1'b0 ;
  assign y976 = ~1'b0 ;
  assign y977 = ~1'b0 ;
  assign y978 = n428 ;
  assign y979 = ~1'b0 ;
  assign y980 = n2401 ;
  assign y981 = n2404 ;
  assign y982 = ~n2406 ;
  assign y983 = n2407 ;
  assign y984 = n2408 ;
  assign y985 = ~1'b0 ;
  assign y986 = ~n2411 ;
  assign y987 = n2332 ;
  assign y988 = ~1'b0 ;
  assign y989 = ~n2418 ;
  assign y990 = n2420 ;
  assign y991 = ~n2422 ;
  assign y992 = ~n2426 ;
  assign y993 = ~1'b0 ;
  assign y994 = ~1'b0 ;
  assign y995 = ~1'b0 ;
  assign y996 = n2433 ;
  assign y997 = n2438 ;
  assign y998 = n2439 ;
  assign y999 = ~1'b0 ;
  assign y1000 = n1813 ;
  assign y1001 = ~n2441 ;
  assign y1002 = n2446 ;
  assign y1003 = ~1'b0 ;
  assign y1004 = ~n2452 ;
  assign y1005 = ~1'b0 ;
  assign y1006 = n2453 ;
  assign y1007 = ~n2456 ;
  assign y1008 = ~n2458 ;
  assign y1009 = ~n2460 ;
  assign y1010 = ~n1538 ;
  assign y1011 = n2463 ;
  assign y1012 = n2465 ;
  assign y1013 = n2468 ;
  assign y1014 = ~n2477 ;
  assign y1015 = 1'b0 ;
  assign y1016 = n2479 ;
  assign y1017 = ~1'b0 ;
  assign y1018 = ~1'b0 ;
  assign y1019 = ~1'b0 ;
  assign y1020 = n2481 ;
  assign y1021 = ~1'b0 ;
  assign y1022 = n2482 ;
  assign y1023 = ~n1981 ;
  assign y1024 = ~1'b0 ;
  assign y1025 = n2485 ;
  assign y1026 = ~n2489 ;
  assign y1027 = ~n2492 ;
  assign y1028 = n2494 ;
  assign y1029 = ~n2499 ;
  assign y1030 = ~n550 ;
  assign y1031 = ~1'b0 ;
  assign y1032 = n2500 ;
  assign y1033 = ~n2502 ;
  assign y1034 = ~x86 ;
  assign y1035 = ~n2506 ;
  assign y1036 = n2508 ;
  assign y1037 = n2511 ;
  assign y1038 = ~1'b0 ;
  assign y1039 = n2520 ;
  assign y1040 = ~n2521 ;
  assign y1041 = ~1'b0 ;
  assign y1042 = ~1'b0 ;
  assign y1043 = ~1'b0 ;
  assign y1044 = n2525 ;
  assign y1045 = n2526 ;
  assign y1046 = ~n2531 ;
  assign y1047 = ~1'b0 ;
  assign y1048 = n2532 ;
  assign y1049 = n2537 ;
  assign y1050 = n2541 ;
  assign y1051 = n2544 ;
  assign y1052 = n2545 ;
  assign y1053 = n569 ;
  assign y1054 = n2557 ;
  assign y1055 = n2564 ;
  assign y1056 = ~1'b0 ;
  assign y1057 = n2568 ;
  assign y1058 = ~1'b0 ;
  assign y1059 = ~1'b0 ;
  assign y1060 = n2570 ;
  assign y1061 = ~n2015 ;
  assign y1062 = n547 ;
  assign y1063 = ~1'b0 ;
  assign y1064 = ~1'b0 ;
  assign y1065 = n2572 ;
  assign y1066 = ~n2579 ;
  assign y1067 = ~1'b0 ;
  assign y1068 = n2580 ;
  assign y1069 = ~n2587 ;
  assign y1070 = 1'b0 ;
  assign y1071 = n2590 ;
  assign y1072 = ~n2600 ;
  assign y1073 = ~1'b0 ;
  assign y1074 = ~1'b0 ;
  assign y1075 = 1'b0 ;
  assign y1076 = ~1'b0 ;
  assign y1077 = 1'b0 ;
  assign y1078 = ~x100 ;
  assign y1079 = n2606 ;
  assign y1080 = ~n2608 ;
  assign y1081 = n2609 ;
  assign y1082 = ~n2617 ;
  assign y1083 = ~n2620 ;
  assign y1084 = n2624 ;
  assign y1085 = n2631 ;
  assign y1086 = ~n2633 ;
  assign y1087 = n2634 ;
  assign y1088 = ~1'b0 ;
  assign y1089 = n2636 ;
  assign y1090 = ~n2651 ;
  assign y1091 = ~n651 ;
  assign y1092 = n2654 ;
  assign y1093 = ~1'b0 ;
  assign y1094 = ~1'b0 ;
  assign y1095 = ~1'b0 ;
  assign y1096 = ~n2659 ;
  assign y1097 = ~n2661 ;
  assign y1098 = ~n2665 ;
  assign y1099 = n2668 ;
  assign y1100 = n2675 ;
  assign y1101 = ~n2681 ;
  assign y1102 = ~1'b0 ;
  assign y1103 = 1'b0 ;
  assign y1104 = n2685 ;
  assign y1105 = ~1'b0 ;
  assign y1106 = ~1'b0 ;
  assign y1107 = n2686 ;
  assign y1108 = n2687 ;
  assign y1109 = n2697 ;
  assign y1110 = n2699 ;
  assign y1111 = ~1'b0 ;
  assign y1112 = ~n2703 ;
  assign y1113 = n694 ;
  assign y1114 = n2705 ;
  assign y1115 = ~1'b0 ;
  assign y1116 = ~1'b0 ;
  assign y1117 = 1'b0 ;
  assign y1118 = 1'b0 ;
  assign y1119 = n2708 ;
  assign y1120 = ~n2711 ;
  assign y1121 = ~n2715 ;
  assign y1122 = ~1'b0 ;
  assign y1123 = ~n2716 ;
  assign y1124 = ~1'b0 ;
  assign y1125 = ~n2378 ;
  assign y1126 = ~n2719 ;
  assign y1127 = n2721 ;
  assign y1128 = n2739 ;
  assign y1129 = ~1'b0 ;
  assign y1130 = ~1'b0 ;
  assign y1131 = n2740 ;
  assign y1132 = n2746 ;
  assign y1133 = n2750 ;
  assign y1134 = n2755 ;
  assign y1135 = ~n2756 ;
  assign y1136 = ~1'b0 ;
  assign y1137 = n2761 ;
  assign y1138 = ~n2763 ;
  assign y1139 = ~1'b0 ;
  assign y1140 = n2764 ;
  assign y1141 = ~n2765 ;
  assign y1142 = n2767 ;
  assign y1143 = n2774 ;
  assign y1144 = ~n2776 ;
  assign y1145 = ~n2778 ;
  assign y1146 = n2779 ;
  assign y1147 = ~n2781 ;
  assign y1148 = ~1'b0 ;
  assign y1149 = ~n2783 ;
  assign y1150 = 1'b0 ;
  assign y1151 = ~1'b0 ;
  assign y1152 = ~n2788 ;
  assign y1153 = ~1'b0 ;
  assign y1154 = ~n710 ;
  assign y1155 = ~1'b0 ;
  assign y1156 = ~1'b0 ;
  assign y1157 = ~n2789 ;
  assign y1158 = ~n2792 ;
  assign y1159 = n2795 ;
  assign y1160 = ~n2796 ;
  assign y1161 = n2797 ;
  assign y1162 = n2798 ;
  assign y1163 = ~1'b0 ;
  assign y1164 = ~1'b0 ;
  assign y1165 = ~n2799 ;
  assign y1166 = ~n2815 ;
  assign y1167 = n2622 ;
  assign y1168 = n2817 ;
  assign y1169 = n2821 ;
  assign y1170 = n2827 ;
  assign y1171 = ~n2839 ;
  assign y1172 = ~1'b0 ;
  assign y1173 = ~1'b0 ;
  assign y1174 = ~1'b0 ;
  assign y1175 = ~n2843 ;
  assign y1176 = ~n2850 ;
  assign y1177 = n2855 ;
  assign y1178 = n2856 ;
  assign y1179 = ~1'b0 ;
  assign y1180 = n2858 ;
  assign y1181 = ~1'b0 ;
  assign y1182 = ~n2859 ;
  assign y1183 = ~n2867 ;
  assign y1184 = ~n2873 ;
  assign y1185 = n2875 ;
  assign y1186 = ~n2877 ;
  assign y1187 = ~n2885 ;
  assign y1188 = n2887 ;
  assign y1189 = ~n2889 ;
  assign y1190 = ~n2891 ;
  assign y1191 = ~n2895 ;
  assign y1192 = ~1'b0 ;
  assign y1193 = ~1'b0 ;
  assign y1194 = 1'b0 ;
  assign y1195 = n2896 ;
  assign y1196 = 1'b0 ;
  assign y1197 = ~n2897 ;
  assign y1198 = n2898 ;
  assign y1199 = n2905 ;
  assign y1200 = ~n2909 ;
  assign y1201 = ~n2916 ;
  assign y1202 = ~n2919 ;
  assign y1203 = ~1'b0 ;
  assign y1204 = ~n2920 ;
  assign y1205 = n2924 ;
  assign y1206 = n2926 ;
  assign y1207 = ~n2933 ;
  assign y1208 = ~n2934 ;
  assign y1209 = ~1'b0 ;
  assign y1210 = ~n2937 ;
  assign y1211 = ~n2939 ;
  assign y1212 = ~n2940 ;
  assign y1213 = n2942 ;
  assign y1214 = ~n2945 ;
  assign y1215 = 1'b0 ;
  assign y1216 = ~n2946 ;
  assign y1217 = ~n2948 ;
  assign y1218 = ~n2957 ;
  assign y1219 = ~n2958 ;
  assign y1220 = n2959 ;
  assign y1221 = ~1'b0 ;
  assign y1222 = ~n2960 ;
  assign y1223 = ~1'b0 ;
  assign y1224 = n2148 ;
  assign y1225 = n2978 ;
  assign y1226 = ~n2980 ;
  assign y1227 = n2986 ;
  assign y1228 = ~n2988 ;
  assign y1229 = ~1'b0 ;
  assign y1230 = n2992 ;
  assign y1231 = ~n2995 ;
  assign y1232 = ~n3000 ;
  assign y1233 = ~1'b0 ;
  assign y1234 = ~n3005 ;
  assign y1235 = ~n3009 ;
  assign y1236 = ~n3011 ;
  assign y1237 = n3012 ;
  assign y1238 = n3021 ;
  assign y1239 = ~1'b0 ;
  assign y1240 = ~1'b0 ;
  assign y1241 = ~1'b0 ;
  assign y1242 = ~n3023 ;
  assign y1243 = n3025 ;
  assign y1244 = ~1'b0 ;
  assign y1245 = ~1'b0 ;
  assign y1246 = ~1'b0 ;
  assign y1247 = ~n3028 ;
  assign y1248 = n3036 ;
  assign y1249 = ~n3037 ;
  assign y1250 = n3040 ;
  assign y1251 = ~1'b0 ;
  assign y1252 = ~1'b0 ;
  assign y1253 = n3041 ;
  assign y1254 = ~n3050 ;
  assign y1255 = ~n3052 ;
  assign y1256 = ~n3057 ;
  assign y1257 = n3062 ;
  assign y1258 = ~n3066 ;
  assign y1259 = n3067 ;
  assign y1260 = n858 ;
  assign y1261 = n3070 ;
  assign y1262 = ~n3074 ;
  assign y1263 = ~1'b0 ;
  assign y1264 = ~1'b0 ;
  assign y1265 = ~1'b0 ;
  assign y1266 = ~1'b0 ;
  assign y1267 = ~n3078 ;
  assign y1268 = ~n3080 ;
  assign y1269 = n3088 ;
  assign y1270 = ~n3090 ;
  assign y1271 = ~1'b0 ;
  assign y1272 = ~n3091 ;
  assign y1273 = ~1'b0 ;
  assign y1274 = n3100 ;
  assign y1275 = ~n3102 ;
  assign y1276 = ~n3104 ;
  assign y1277 = n3106 ;
  assign y1278 = ~1'b0 ;
  assign y1279 = n3115 ;
  assign y1280 = n3116 ;
  assign y1281 = ~1'b0 ;
  assign y1282 = ~1'b0 ;
  assign y1283 = ~n3117 ;
  assign y1284 = ~1'b0 ;
  assign y1285 = ~n3118 ;
  assign y1286 = ~n3119 ;
  assign y1287 = ~1'b0 ;
  assign y1288 = n3127 ;
  assign y1289 = n3131 ;
  assign y1290 = ~n3138 ;
  assign y1291 = ~n3140 ;
  assign y1292 = ~1'b0 ;
  assign y1293 = n3142 ;
  assign y1294 = n3144 ;
  assign y1295 = n3154 ;
  assign y1296 = ~1'b0 ;
  assign y1297 = ~1'b0 ;
  assign y1298 = ~n3155 ;
  assign y1299 = n3158 ;
  assign y1300 = ~n3159 ;
  assign y1301 = n3163 ;
  assign y1302 = ~1'b0 ;
  assign y1303 = ~n3169 ;
  assign y1304 = n3172 ;
  assign y1305 = n2942 ;
  assign y1306 = ~n3176 ;
  assign y1307 = ~x243 ;
  assign y1308 = ~n3184 ;
  assign y1309 = n3191 ;
  assign y1310 = n3195 ;
  assign y1311 = n3197 ;
  assign y1312 = ~n3198 ;
  assign y1313 = n3199 ;
  assign y1314 = n3202 ;
  assign y1315 = ~1'b0 ;
  assign y1316 = ~n3205 ;
  assign y1317 = n1219 ;
  assign y1318 = n3206 ;
  assign y1319 = ~1'b0 ;
  assign y1320 = ~n3209 ;
  assign y1321 = n3210 ;
  assign y1322 = n3211 ;
  assign y1323 = n3217 ;
  assign y1324 = n3218 ;
  assign y1325 = n3222 ;
  assign y1326 = ~n3231 ;
  assign y1327 = n3232 ;
  assign y1328 = ~1'b0 ;
  assign y1329 = n3233 ;
  assign y1330 = ~n3234 ;
  assign y1331 = n3235 ;
  assign y1332 = n3238 ;
  assign y1333 = ~1'b0 ;
  assign y1334 = ~1'b0 ;
  assign y1335 = ~1'b0 ;
  assign y1336 = n3240 ;
  assign y1337 = ~1'b0 ;
  assign y1338 = ~1'b0 ;
  assign y1339 = ~n3243 ;
  assign y1340 = n3245 ;
  assign y1341 = n3246 ;
  assign y1342 = ~n3251 ;
  assign y1343 = ~n3256 ;
  assign y1344 = n3263 ;
  assign y1345 = n3264 ;
  assign y1346 = ~1'b0 ;
  assign y1347 = ~1'b0 ;
  assign y1348 = ~1'b0 ;
  assign y1349 = ~n3266 ;
  assign y1350 = n3267 ;
  assign y1351 = n3269 ;
  assign y1352 = ~1'b0 ;
  assign y1353 = n3274 ;
  assign y1354 = ~1'b0 ;
  assign y1355 = ~1'b0 ;
  assign y1356 = ~1'b0 ;
  assign y1357 = n3275 ;
  assign y1358 = ~n3279 ;
  assign y1359 = n3281 ;
  assign y1360 = ~n3284 ;
  assign y1361 = ~1'b0 ;
  assign y1362 = ~n3291 ;
  assign y1363 = n1404 ;
  assign y1364 = ~1'b0 ;
  assign y1365 = ~1'b0 ;
  assign y1366 = ~1'b0 ;
  assign y1367 = ~n3297 ;
  assign y1368 = ~n3304 ;
  assign y1369 = n3308 ;
  assign y1370 = ~1'b0 ;
  assign y1371 = ~n3311 ;
  assign y1372 = n3312 ;
  assign y1373 = ~1'b0 ;
  assign y1374 = n3313 ;
  assign y1375 = n2706 ;
  assign y1376 = ~n3315 ;
  assign y1377 = ~n3319 ;
  assign y1378 = n3321 ;
  assign y1379 = ~n3325 ;
  assign y1380 = ~n3327 ;
  assign y1381 = ~1'b0 ;
  assign y1382 = ~n2158 ;
  assign y1383 = ~n3332 ;
  assign y1384 = ~1'b0 ;
  assign y1385 = x225 ;
  assign y1386 = ~n3333 ;
  assign y1387 = n3335 ;
  assign y1388 = ~n1775 ;
  assign y1389 = ~1'b0 ;
  assign y1390 = n3339 ;
  assign y1391 = ~n3340 ;
  assign y1392 = ~n3344 ;
  assign y1393 = n3352 ;
  assign y1394 = n3370 ;
  assign y1395 = n3371 ;
  assign y1396 = n3372 ;
  assign y1397 = ~1'b0 ;
  assign y1398 = ~1'b0 ;
  assign y1399 = ~n3375 ;
  assign y1400 = n3378 ;
  assign y1401 = n3380 ;
  assign y1402 = n3383 ;
  assign y1403 = ~n3386 ;
  assign y1404 = n3389 ;
  assign y1405 = ~1'b0 ;
  assign y1406 = ~n3393 ;
  assign y1407 = n3396 ;
  assign y1408 = n3399 ;
  assign y1409 = ~1'b0 ;
  assign y1410 = ~n3400 ;
  assign y1411 = ~n3410 ;
  assign y1412 = ~1'b0 ;
  assign y1413 = ~1'b0 ;
  assign y1414 = ~1'b0 ;
  assign y1415 = n3412 ;
  assign y1416 = n3417 ;
  assign y1417 = ~1'b0 ;
  assign y1418 = ~n3424 ;
  assign y1419 = ~n3427 ;
  assign y1420 = ~1'b0 ;
  assign y1421 = n3429 ;
  assign y1422 = ~1'b0 ;
  assign y1423 = ~n3432 ;
  assign y1424 = n3435 ;
  assign y1425 = ~n3439 ;
  assign y1426 = n3440 ;
  assign y1427 = n3442 ;
  assign y1428 = n3446 ;
  assign y1429 = ~n3457 ;
  assign y1430 = n3460 ;
  assign y1431 = ~1'b0 ;
  assign y1432 = ~n3461 ;
  assign y1433 = n3468 ;
  assign y1434 = ~1'b0 ;
  assign y1435 = ~n3478 ;
  assign y1436 = n2936 ;
  assign y1437 = ~n3481 ;
  assign y1438 = ~n3486 ;
  assign y1439 = n3488 ;
  assign y1440 = ~n3490 ;
  assign y1441 = n3498 ;
  assign y1442 = ~1'b0 ;
  assign y1443 = ~1'b0 ;
  assign y1444 = ~1'b0 ;
  assign y1445 = ~n3502 ;
  assign y1446 = n3504 ;
  assign y1447 = n3508 ;
  assign y1448 = ~1'b0 ;
  assign y1449 = ~n3513 ;
  assign y1450 = ~n3514 ;
  assign y1451 = n3518 ;
  assign y1452 = ~n3527 ;
  assign y1453 = n3532 ;
  assign y1454 = ~n3534 ;
  assign y1455 = ~n3535 ;
  assign y1456 = n3537 ;
  assign y1457 = n3541 ;
  assign y1458 = ~1'b0 ;
  assign y1459 = n3542 ;
  assign y1460 = ~1'b0 ;
  assign y1461 = n3547 ;
  assign y1462 = ~n3554 ;
  assign y1463 = ~1'b0 ;
  assign y1464 = 1'b0 ;
  assign y1465 = ~1'b0 ;
  assign y1466 = ~n3362 ;
  assign y1467 = ~n3558 ;
  assign y1468 = ~n3560 ;
  assign y1469 = ~n3561 ;
  assign y1470 = ~n3563 ;
  assign y1471 = n3564 ;
  assign y1472 = n3565 ;
  assign y1473 = ~n3571 ;
  assign y1474 = n3573 ;
  assign y1475 = ~1'b0 ;
  assign y1476 = n3574 ;
  assign y1477 = n3576 ;
  assign y1478 = ~1'b0 ;
  assign y1479 = ~1'b0 ;
  assign y1480 = n3584 ;
  assign y1481 = ~1'b0 ;
  assign y1482 = ~n3590 ;
  assign y1483 = ~n3592 ;
  assign y1484 = ~n3594 ;
  assign y1485 = ~1'b0 ;
  assign y1486 = n3596 ;
  assign y1487 = ~1'b0 ;
  assign y1488 = n3606 ;
  assign y1489 = n3608 ;
  assign y1490 = n3611 ;
  assign y1491 = n3616 ;
  assign y1492 = ~n3617 ;
  assign y1493 = ~1'b0 ;
  assign y1494 = n3619 ;
  assign y1495 = ~n3622 ;
  assign y1496 = ~1'b0 ;
  assign y1497 = n3624 ;
  assign y1498 = ~n3626 ;
  assign y1499 = ~1'b0 ;
  assign y1500 = ~1'b0 ;
  assign y1501 = ~n3627 ;
  assign y1502 = ~1'b0 ;
  assign y1503 = ~n3628 ;
  assign y1504 = ~1'b0 ;
  assign y1505 = n3631 ;
  assign y1506 = ~1'b0 ;
  assign y1507 = ~n3639 ;
  assign y1508 = n3641 ;
  assign y1509 = ~1'b0 ;
  assign y1510 = ~1'b0 ;
  assign y1511 = ~n3012 ;
  assign y1512 = ~n3643 ;
  assign y1513 = n3649 ;
  assign y1514 = ~1'b0 ;
  assign y1515 = n3651 ;
  assign y1516 = ~n3654 ;
  assign y1517 = ~n3656 ;
  assign y1518 = ~1'b0 ;
  assign y1519 = n3665 ;
  assign y1520 = n3666 ;
  assign y1521 = n3668 ;
  assign y1522 = n749 ;
  assign y1523 = ~n3676 ;
  assign y1524 = n3684 ;
  assign y1525 = n3694 ;
  assign y1526 = ~1'b0 ;
  assign y1527 = n3695 ;
  assign y1528 = ~1'b0 ;
  assign y1529 = ~n3698 ;
  assign y1530 = ~1'b0 ;
  assign y1531 = ~n3705 ;
  assign y1532 = n3707 ;
  assign y1533 = ~n3709 ;
  assign y1534 = n3710 ;
  assign y1535 = ~n3712 ;
  assign y1536 = ~n3717 ;
  assign y1537 = ~n2287 ;
  assign y1538 = ~1'b0 ;
  assign y1539 = ~n3721 ;
  assign y1540 = ~1'b0 ;
  assign y1541 = ~1'b0 ;
  assign y1542 = ~1'b0 ;
  assign y1543 = ~1'b0 ;
  assign y1544 = ~n3722 ;
  assign y1545 = n3726 ;
  assign y1546 = ~1'b0 ;
  assign y1547 = ~1'b0 ;
  assign y1548 = n3729 ;
  assign y1549 = ~n617 ;
  assign y1550 = ~n3736 ;
  assign y1551 = ~n3739 ;
  assign y1552 = ~n3740 ;
  assign y1553 = n3742 ;
  assign y1554 = n3745 ;
  assign y1555 = ~1'b0 ;
  assign y1556 = n1519 ;
  assign y1557 = ~1'b0 ;
  assign y1558 = ~n3749 ;
  assign y1559 = ~1'b0 ;
  assign y1560 = n3750 ;
  assign y1561 = ~n3754 ;
  assign y1562 = ~n3757 ;
  assign y1563 = ~1'b0 ;
  assign y1564 = ~1'b0 ;
  assign y1565 = n3760 ;
  assign y1566 = ~1'b0 ;
  assign y1567 = ~n3763 ;
  assign y1568 = 1'b0 ;
  assign y1569 = 1'b0 ;
  assign y1570 = ~n3771 ;
  assign y1571 = n3777 ;
  assign y1572 = n3783 ;
  assign y1573 = n3786 ;
  assign y1574 = ~n3788 ;
  assign y1575 = ~n3793 ;
  assign y1576 = ~1'b0 ;
  assign y1577 = ~n2070 ;
  assign y1578 = ~1'b0 ;
  assign y1579 = ~1'b0 ;
  assign y1580 = ~n3795 ;
  assign y1581 = n3796 ;
  assign y1582 = n3797 ;
  assign y1583 = n3799 ;
  assign y1584 = ~1'b0 ;
  assign y1585 = ~n3802 ;
  assign y1586 = n3805 ;
  assign y1587 = n3810 ;
  assign y1588 = ~1'b0 ;
  assign y1589 = ~n3812 ;
  assign y1590 = ~1'b0 ;
  assign y1591 = ~1'b0 ;
  assign y1592 = ~1'b0 ;
  assign y1593 = ~n3821 ;
  assign y1594 = ~1'b0 ;
  assign y1595 = ~1'b0 ;
  assign y1596 = n3825 ;
  assign y1597 = n3829 ;
  assign y1598 = ~n3835 ;
  assign y1599 = ~1'b0 ;
  assign y1600 = ~n3839 ;
  assign y1601 = n3840 ;
  assign y1602 = ~n3843 ;
  assign y1603 = n3844 ;
  assign y1604 = n3845 ;
  assign y1605 = n3850 ;
  assign y1606 = ~1'b0 ;
  assign y1607 = n3853 ;
  assign y1608 = n3861 ;
  assign y1609 = n883 ;
  assign y1610 = n2472 ;
  assign y1611 = n3867 ;
  assign y1612 = ~n3868 ;
  assign y1613 = ~n3874 ;
  assign y1614 = n3875 ;
  assign y1615 = n3876 ;
  assign y1616 = ~n3877 ;
  assign y1617 = ~1'b0 ;
  assign y1618 = ~n3878 ;
  assign y1619 = ~n3881 ;
  assign y1620 = ~n3882 ;
  assign y1621 = ~n3885 ;
  assign y1622 = 1'b0 ;
  assign y1623 = ~1'b0 ;
  assign y1624 = ~n1591 ;
  assign y1625 = n3887 ;
  assign y1626 = n3889 ;
  assign y1627 = ~n3893 ;
  assign y1628 = n3895 ;
  assign y1629 = n3899 ;
  assign y1630 = ~n3904 ;
  assign y1631 = ~n3908 ;
  assign y1632 = ~1'b0 ;
  assign y1633 = ~n3912 ;
  assign y1634 = n1968 ;
  assign y1635 = ~n3913 ;
  assign y1636 = ~1'b0 ;
  assign y1637 = n3915 ;
  assign y1638 = n3930 ;
  assign y1639 = ~n3934 ;
  assign y1640 = ~n3935 ;
  assign y1641 = n3936 ;
  assign y1642 = n3939 ;
  assign y1643 = n3945 ;
  assign y1644 = ~1'b0 ;
  assign y1645 = ~n3946 ;
  assign y1646 = n3950 ;
  assign y1647 = n3952 ;
  assign y1648 = ~1'b0 ;
  assign y1649 = n3957 ;
  assign y1650 = n3958 ;
  assign y1651 = n3963 ;
  assign y1652 = n3966 ;
  assign y1653 = ~n3967 ;
  assign y1654 = 1'b0 ;
  assign y1655 = ~1'b0 ;
  assign y1656 = ~1'b0 ;
  assign y1657 = ~1'b0 ;
  assign y1658 = ~n3969 ;
  assign y1659 = ~1'b0 ;
  assign y1660 = ~1'b0 ;
  assign y1661 = ~n3972 ;
  assign y1662 = n3975 ;
  assign y1663 = ~n3977 ;
  assign y1664 = ~1'b0 ;
  assign y1665 = n3978 ;
  assign y1666 = ~1'b0 ;
  assign y1667 = n3981 ;
  assign y1668 = n3982 ;
  assign y1669 = ~n3984 ;
  assign y1670 = ~n3985 ;
  assign y1671 = ~n3996 ;
  assign y1672 = n3999 ;
  assign y1673 = ~1'b0 ;
  assign y1674 = n4001 ;
  assign y1675 = n4005 ;
  assign y1676 = n4009 ;
  assign y1677 = n4014 ;
  assign y1678 = ~1'b0 ;
  assign y1679 = ~n4018 ;
  assign y1680 = ~1'b0 ;
  assign y1681 = ~n4020 ;
  assign y1682 = ~1'b0 ;
  assign y1683 = ~n4023 ;
  assign y1684 = ~n4032 ;
  assign y1685 = n4037 ;
  assign y1686 = n4040 ;
  assign y1687 = ~n4042 ;
  assign y1688 = ~n4045 ;
  assign y1689 = ~n4046 ;
  assign y1690 = n4047 ;
  assign y1691 = ~1'b0 ;
  assign y1692 = n4062 ;
  assign y1693 = ~1'b0 ;
  assign y1694 = ~1'b0 ;
  assign y1695 = ~n4066 ;
  assign y1696 = ~n4067 ;
  assign y1697 = n4080 ;
  assign y1698 = ~1'b0 ;
  assign y1699 = ~1'b0 ;
  assign y1700 = ~n3319 ;
  assign y1701 = ~n4083 ;
  assign y1702 = ~1'b0 ;
  assign y1703 = ~n4091 ;
  assign y1704 = n4092 ;
  assign y1705 = ~1'b0 ;
  assign y1706 = ~1'b0 ;
  assign y1707 = n4093 ;
  assign y1708 = n4095 ;
  assign y1709 = n4096 ;
  assign y1710 = ~1'b0 ;
  assign y1711 = n4102 ;
  assign y1712 = n4105 ;
  assign y1713 = ~n4117 ;
  assign y1714 = ~n4119 ;
  assign y1715 = ~n4122 ;
  assign y1716 = n4123 ;
  assign y1717 = ~1'b0 ;
  assign y1718 = ~1'b0 ;
  assign y1719 = n4125 ;
  assign y1720 = ~1'b0 ;
  assign y1721 = ~1'b0 ;
  assign y1722 = n4128 ;
  assign y1723 = n4135 ;
  assign y1724 = ~n4136 ;
  assign y1725 = ~n4138 ;
  assign y1726 = ~n4139 ;
  assign y1727 = ~n3425 ;
  assign y1728 = 1'b0 ;
  assign y1729 = n4142 ;
  assign y1730 = n4144 ;
  assign y1731 = ~1'b0 ;
  assign y1732 = ~1'b0 ;
  assign y1733 = ~n4145 ;
  assign y1734 = ~1'b0 ;
  assign y1735 = ~n3554 ;
  assign y1736 = n4146 ;
  assign y1737 = ~1'b0 ;
  assign y1738 = n4148 ;
  assign y1739 = n4149 ;
  assign y1740 = n4152 ;
  assign y1741 = ~1'b0 ;
  assign y1742 = ~1'b0 ;
  assign y1743 = ~n4165 ;
  assign y1744 = ~n4166 ;
  assign y1745 = n4172 ;
  assign y1746 = ~n4175 ;
  assign y1747 = n4178 ;
  assign y1748 = n4180 ;
  assign y1749 = ~1'b0 ;
  assign y1750 = ~n4184 ;
  assign y1751 = ~n4185 ;
  assign y1752 = n4186 ;
  assign y1753 = ~n4187 ;
  assign y1754 = ~n4189 ;
  assign y1755 = ~1'b0 ;
  assign y1756 = ~n4192 ;
  assign y1757 = ~n4193 ;
  assign y1758 = n4196 ;
  assign y1759 = ~n4202 ;
  assign y1760 = ~1'b0 ;
  assign y1761 = ~n4203 ;
  assign y1762 = ~n4206 ;
  assign y1763 = ~n4207 ;
  assign y1764 = n4208 ;
  assign y1765 = ~1'b0 ;
  assign y1766 = ~n4209 ;
  assign y1767 = ~1'b0 ;
  assign y1768 = n4212 ;
  assign y1769 = n4214 ;
  assign y1770 = n4222 ;
  assign y1771 = ~1'b0 ;
  assign y1772 = ~n4227 ;
  assign y1773 = n4229 ;
  assign y1774 = ~x118 ;
  assign y1775 = n4236 ;
  assign y1776 = ~1'b0 ;
  assign y1777 = ~n4238 ;
  assign y1778 = n4244 ;
  assign y1779 = ~n4248 ;
  assign y1780 = n4249 ;
  assign y1781 = ~1'b0 ;
  assign y1782 = ~n4252 ;
  assign y1783 = ~n4257 ;
  assign y1784 = ~1'b0 ;
  assign y1785 = ~1'b0 ;
  assign y1786 = ~1'b0 ;
  assign y1787 = n4259 ;
  assign y1788 = ~1'b0 ;
  assign y1789 = n4268 ;
  assign y1790 = n1600 ;
  assign y1791 = n4270 ;
  assign y1792 = ~1'b0 ;
  assign y1793 = n4276 ;
  assign y1794 = n4280 ;
  assign y1795 = ~1'b0 ;
  assign y1796 = ~n4284 ;
  assign y1797 = n4286 ;
  assign y1798 = n4287 ;
  assign y1799 = ~1'b0 ;
  assign y1800 = ~n2919 ;
  assign y1801 = ~1'b0 ;
  assign y1802 = ~1'b0 ;
  assign y1803 = ~1'b0 ;
  assign y1804 = ~n4288 ;
  assign y1805 = ~n4292 ;
  assign y1806 = ~n4294 ;
  assign y1807 = ~n4295 ;
  assign y1808 = n4296 ;
  assign y1809 = ~1'b0 ;
  assign y1810 = n4298 ;
  assign y1811 = n4300 ;
  assign y1812 = ~n4302 ;
  assign y1813 = n4303 ;
  assign y1814 = ~n4305 ;
  assign y1815 = ~n3325 ;
  assign y1816 = ~1'b0 ;
  assign y1817 = n4306 ;
  assign y1818 = n4309 ;
  assign y1819 = ~n387 ;
  assign y1820 = ~n634 ;
  assign y1821 = ~n4316 ;
  assign y1822 = ~1'b0 ;
  assign y1823 = ~1'b0 ;
  assign y1824 = n4317 ;
  assign y1825 = n4321 ;
  assign y1826 = n4323 ;
  assign y1827 = n4326 ;
  assign y1828 = ~n4333 ;
  assign y1829 = ~n4335 ;
  assign y1830 = n4338 ;
  assign y1831 = ~1'b0 ;
  assign y1832 = ~1'b0 ;
  assign y1833 = ~1'b0 ;
  assign y1834 = 1'b0 ;
  assign y1835 = n4341 ;
  assign y1836 = ~n4342 ;
  assign y1837 = ~1'b0 ;
  assign y1838 = ~1'b0 ;
  assign y1839 = ~n4343 ;
  assign y1840 = ~1'b0 ;
  assign y1841 = n3258 ;
  assign y1842 = ~1'b0 ;
  assign y1843 = ~n4346 ;
  assign y1844 = ~n4352 ;
  assign y1845 = ~n4355 ;
  assign y1846 = ~1'b0 ;
  assign y1847 = ~1'b0 ;
  assign y1848 = ~n4356 ;
  assign y1849 = ~1'b0 ;
  assign y1850 = ~1'b0 ;
  assign y1851 = n4364 ;
  assign y1852 = n4368 ;
  assign y1853 = n4369 ;
  assign y1854 = ~n4370 ;
  assign y1855 = ~n4372 ;
  assign y1856 = ~n4379 ;
  assign y1857 = n4380 ;
  assign y1858 = ~n4381 ;
  assign y1859 = ~n686 ;
  assign y1860 = n537 ;
  assign y1861 = ~n4383 ;
  assign y1862 = n4384 ;
  assign y1863 = n4386 ;
  assign y1864 = ~n4387 ;
  assign y1865 = ~n4391 ;
  assign y1866 = ~n4393 ;
  assign y1867 = ~1'b0 ;
  assign y1868 = ~n4395 ;
  assign y1869 = ~n4404 ;
  assign y1870 = ~n4407 ;
  assign y1871 = n4411 ;
  assign y1872 = n4416 ;
  assign y1873 = n3508 ;
  assign y1874 = ~1'b0 ;
  assign y1875 = n4417 ;
  assign y1876 = n4420 ;
  assign y1877 = n2317 ;
  assign y1878 = n4424 ;
  assign y1879 = ~1'b0 ;
  assign y1880 = n4425 ;
  assign y1881 = n4428 ;
  assign y1882 = ~n4433 ;
  assign y1883 = ~n4437 ;
  assign y1884 = ~n4438 ;
  assign y1885 = ~n4439 ;
  assign y1886 = ~n4442 ;
  assign y1887 = n4452 ;
  assign y1888 = 1'b0 ;
  assign y1889 = n4454 ;
  assign y1890 = n4456 ;
  assign y1891 = ~1'b0 ;
  assign y1892 = n4459 ;
  assign y1893 = n4460 ;
  assign y1894 = n4463 ;
  assign y1895 = n4470 ;
  assign y1896 = ~1'b0 ;
  assign y1897 = n4474 ;
  assign y1898 = n4476 ;
  assign y1899 = ~1'b0 ;
  assign y1900 = ~1'b0 ;
  assign y1901 = n4478 ;
  assign y1902 = ~n4481 ;
  assign y1903 = n4482 ;
  assign y1904 = ~n4487 ;
  assign y1905 = ~n4488 ;
  assign y1906 = ~n4497 ;
  assign y1907 = ~n4498 ;
  assign y1908 = ~1'b0 ;
  assign y1909 = ~n4500 ;
  assign y1910 = ~n4501 ;
  assign y1911 = ~1'b0 ;
  assign y1912 = n4506 ;
  assign y1913 = ~1'b0 ;
  assign y1914 = n4509 ;
  assign y1915 = ~1'b0 ;
  assign y1916 = ~1'b0 ;
  assign y1917 = ~n3961 ;
  assign y1918 = ~n4510 ;
  assign y1919 = ~1'b0 ;
  assign y1920 = n4514 ;
  assign y1921 = ~n4516 ;
  assign y1922 = ~1'b0 ;
  assign y1923 = n4519 ;
  assign y1924 = ~1'b0 ;
  assign y1925 = ~n4522 ;
  assign y1926 = ~n4524 ;
  assign y1927 = ~1'b0 ;
  assign y1928 = ~n4534 ;
  assign y1929 = 1'b0 ;
  assign y1930 = n4539 ;
  assign y1931 = ~n4541 ;
  assign y1932 = n4547 ;
  assign y1933 = n4557 ;
  assign y1934 = ~n4559 ;
  assign y1935 = ~n4562 ;
  assign y1936 = n2529 ;
  assign y1937 = ~1'b0 ;
  assign y1938 = n2622 ;
  assign y1939 = n4566 ;
  assign y1940 = n4567 ;
  assign y1941 = ~n4569 ;
  assign y1942 = ~n4571 ;
  assign y1943 = n4572 ;
  assign y1944 = ~1'b0 ;
  assign y1945 = ~n4574 ;
  assign y1946 = n4575 ;
  assign y1947 = ~n890 ;
  assign y1948 = ~1'b0 ;
  assign y1949 = n4576 ;
  assign y1950 = ~n4578 ;
  assign y1951 = n4585 ;
  assign y1952 = n4596 ;
  assign y1953 = ~n4598 ;
  assign y1954 = ~1'b0 ;
  assign y1955 = n4599 ;
  assign y1956 = ~n4605 ;
  assign y1957 = ~1'b0 ;
  assign y1958 = ~1'b0 ;
  assign y1959 = n4615 ;
  assign y1960 = ~n4617 ;
  assign y1961 = ~n4624 ;
  assign y1962 = ~1'b0 ;
  assign y1963 = ~1'b0 ;
  assign y1964 = n4631 ;
  assign y1965 = n4633 ;
  assign y1966 = n4638 ;
  assign y1967 = ~n4639 ;
  assign y1968 = ~1'b0 ;
  assign y1969 = ~1'b0 ;
  assign y1970 = n4640 ;
  assign y1971 = ~1'b0 ;
  assign y1972 = ~n4645 ;
  assign y1973 = ~1'b0 ;
  assign y1974 = ~n4648 ;
  assign y1975 = ~n4654 ;
  assign y1976 = ~n4660 ;
  assign y1977 = ~n2203 ;
  assign y1978 = ~n4663 ;
  assign y1979 = ~1'b0 ;
  assign y1980 = ~n4668 ;
  assign y1981 = n4669 ;
  assign y1982 = n4670 ;
  assign y1983 = n4676 ;
  assign y1984 = ~1'b0 ;
  assign y1985 = n4677 ;
  assign y1986 = ~1'b0 ;
  assign y1987 = n4682 ;
  assign y1988 = n4685 ;
  assign y1989 = ~1'b0 ;
  assign y1990 = n4686 ;
  assign y1991 = ~n4691 ;
  assign y1992 = n4693 ;
  assign y1993 = n4696 ;
  assign y1994 = ~n4704 ;
  assign y1995 = ~1'b0 ;
  assign y1996 = n4706 ;
  assign y1997 = n4710 ;
  assign y1998 = n4712 ;
  assign y1999 = ~1'b0 ;
  assign y2000 = ~n4718 ;
  assign y2001 = n917 ;
  assign y2002 = ~1'b0 ;
  assign y2003 = ~n4720 ;
  assign y2004 = ~n4723 ;
  assign y2005 = n4724 ;
  assign y2006 = 1'b0 ;
  assign y2007 = ~1'b0 ;
  assign y2008 = ~1'b0 ;
  assign y2009 = ~1'b0 ;
  assign y2010 = ~n4725 ;
  assign y2011 = ~n4726 ;
  assign y2012 = n4728 ;
  assign y2013 = ~n4732 ;
  assign y2014 = n4742 ;
  assign y2015 = ~1'b0 ;
  assign y2016 = ~1'b0 ;
  assign y2017 = ~n2735 ;
  assign y2018 = ~n4744 ;
  assign y2019 = ~1'b0 ;
  assign y2020 = ~1'b0 ;
  assign y2021 = n4747 ;
  assign y2022 = ~n4757 ;
  assign y2023 = ~n4766 ;
  assign y2024 = ~1'b0 ;
  assign y2025 = ~n3600 ;
  assign y2026 = n4770 ;
  assign y2027 = ~1'b0 ;
  assign y2028 = n4773 ;
  assign y2029 = ~n4780 ;
  assign y2030 = n4783 ;
  assign y2031 = n4790 ;
  assign y2032 = n3588 ;
  assign y2033 = ~1'b0 ;
  assign y2034 = ~1'b0 ;
  assign y2035 = ~n4791 ;
  assign y2036 = ~n4793 ;
  assign y2037 = n4795 ;
  assign y2038 = ~n4797 ;
  assign y2039 = n4802 ;
  assign y2040 = ~n4806 ;
  assign y2041 = ~1'b0 ;
  assign y2042 = n4809 ;
  assign y2043 = n4815 ;
  assign y2044 = ~n3777 ;
  assign y2045 = ~1'b0 ;
  assign y2046 = ~1'b0 ;
  assign y2047 = ~1'b0 ;
  assign y2048 = ~1'b0 ;
  assign y2049 = ~n4818 ;
  assign y2050 = ~1'b0 ;
  assign y2051 = ~1'b0 ;
  assign y2052 = n4819 ;
  assign y2053 = n4828 ;
  assign y2054 = n4830 ;
  assign y2055 = ~1'b0 ;
  assign y2056 = ~n4836 ;
  assign y2057 = n4838 ;
  assign y2058 = n4840 ;
  assign y2059 = ~n4842 ;
  assign y2060 = n4843 ;
  assign y2061 = ~1'b0 ;
  assign y2062 = ~n4848 ;
  assign y2063 = n4849 ;
  assign y2064 = n4852 ;
  assign y2065 = n4853 ;
  assign y2066 = ~1'b0 ;
  assign y2067 = n4857 ;
  assign y2068 = n4859 ;
  assign y2069 = 1'b0 ;
  assign y2070 = ~n4860 ;
  assign y2071 = ~1'b0 ;
  assign y2072 = ~n4867 ;
  assign y2073 = ~1'b0 ;
  assign y2074 = ~n4872 ;
  assign y2075 = ~1'b0 ;
  assign y2076 = ~n4875 ;
  assign y2077 = ~n4876 ;
  assign y2078 = ~n4878 ;
  assign y2079 = ~1'b0 ;
  assign y2080 = 1'b0 ;
  assign y2081 = ~n4880 ;
  assign y2082 = n4881 ;
  assign y2083 = n4885 ;
  assign y2084 = n4887 ;
  assign y2085 = n4890 ;
  assign y2086 = ~n4892 ;
  assign y2087 = n4895 ;
  assign y2088 = n4900 ;
  assign y2089 = ~n4909 ;
  assign y2090 = n4910 ;
  assign y2091 = n4916 ;
  assign y2092 = n4921 ;
  assign y2093 = ~1'b0 ;
  assign y2094 = n4922 ;
  assign y2095 = ~n4927 ;
  assign y2096 = n4931 ;
  assign y2097 = ~n4934 ;
  assign y2098 = n4936 ;
  assign y2099 = n4941 ;
  assign y2100 = ~1'b0 ;
  assign y2101 = n4944 ;
  assign y2102 = ~1'b0 ;
  assign y2103 = ~1'b0 ;
  assign y2104 = ~n4949 ;
  assign y2105 = ~1'b0 ;
  assign y2106 = ~1'b0 ;
  assign y2107 = n4953 ;
  assign y2108 = n4954 ;
  assign y2109 = ~n4956 ;
  assign y2110 = ~1'b0 ;
  assign y2111 = ~1'b0 ;
  assign y2112 = ~n4958 ;
  assign y2113 = ~1'b0 ;
  assign y2114 = 1'b0 ;
  assign y2115 = 1'b0 ;
  assign y2116 = n4959 ;
  assign y2117 = ~n4965 ;
  assign y2118 = n4966 ;
  assign y2119 = ~n4094 ;
  assign y2120 = ~n1545 ;
  assign y2121 = ~1'b0 ;
  assign y2122 = n4974 ;
  assign y2123 = n4981 ;
  assign y2124 = n4986 ;
  assign y2125 = ~n4988 ;
  assign y2126 = ~n4989 ;
  assign y2127 = n1585 ;
  assign y2128 = ~n4992 ;
  assign y2129 = ~n4998 ;
  assign y2130 = n5001 ;
  assign y2131 = n5008 ;
  assign y2132 = ~n5014 ;
  assign y2133 = n5017 ;
  assign y2134 = ~n5018 ;
  assign y2135 = ~n5020 ;
  assign y2136 = n5021 ;
  assign y2137 = ~1'b0 ;
  assign y2138 = ~n5022 ;
  assign y2139 = ~1'b0 ;
  assign y2140 = ~n5023 ;
  assign y2141 = ~n5031 ;
  assign y2142 = ~1'b0 ;
  assign y2143 = ~n5033 ;
  assign y2144 = ~1'b0 ;
  assign y2145 = ~n5034 ;
  assign y2146 = n1879 ;
  assign y2147 = n5036 ;
  assign y2148 = ~n5041 ;
  assign y2149 = n5047 ;
  assign y2150 = ~1'b0 ;
  assign y2151 = n5049 ;
  assign y2152 = ~1'b0 ;
  assign y2153 = ~1'b0 ;
  assign y2154 = n5052 ;
  assign y2155 = ~n5059 ;
  assign y2156 = n5062 ;
  assign y2157 = ~n5063 ;
  assign y2158 = n5065 ;
  assign y2159 = ~n5066 ;
  assign y2160 = ~n5074 ;
  assign y2161 = ~1'b0 ;
  assign y2162 = ~n5075 ;
  assign y2163 = ~1'b0 ;
  assign y2164 = ~n5076 ;
  assign y2165 = n5078 ;
  assign y2166 = ~n5079 ;
  assign y2167 = ~n5080 ;
  assign y2168 = ~n5082 ;
  assign y2169 = ~n5084 ;
  assign y2170 = ~1'b0 ;
  assign y2171 = n5086 ;
  assign y2172 = ~n5089 ;
  assign y2173 = n5091 ;
  assign y2174 = ~n5099 ;
  assign y2175 = n5103 ;
  assign y2176 = n5104 ;
  assign y2177 = ~1'b0 ;
  assign y2178 = n5105 ;
  assign y2179 = n5108 ;
  assign y2180 = ~1'b0 ;
  assign y2181 = ~n5110 ;
  assign y2182 = n5111 ;
  assign y2183 = n5113 ;
  assign y2184 = ~1'b0 ;
  assign y2185 = n5114 ;
  assign y2186 = ~n5116 ;
  assign y2187 = n5118 ;
  assign y2188 = n5123 ;
  assign y2189 = ~n5125 ;
  assign y2190 = n5134 ;
  assign y2191 = ~1'b0 ;
  assign y2192 = n5135 ;
  assign y2193 = 1'b0 ;
  assign y2194 = ~1'b0 ;
  assign y2195 = ~n5139 ;
  assign y2196 = n5140 ;
  assign y2197 = ~n5148 ;
  assign y2198 = ~1'b0 ;
  assign y2199 = ~n5151 ;
  assign y2200 = n5152 ;
  assign y2201 = ~1'b0 ;
  assign y2202 = n5153 ;
  assign y2203 = ~1'b0 ;
  assign y2204 = ~n5156 ;
  assign y2205 = ~n5167 ;
  assign y2206 = ~n5168 ;
  assign y2207 = n5170 ;
  assign y2208 = ~n5175 ;
  assign y2209 = ~1'b0 ;
  assign y2210 = n5180 ;
  assign y2211 = n5181 ;
  assign y2212 = n5182 ;
  assign y2213 = ~1'b0 ;
  assign y2214 = n5186 ;
  assign y2215 = n5187 ;
  assign y2216 = ~n5192 ;
  assign y2217 = ~1'b0 ;
  assign y2218 = ~n5193 ;
  assign y2219 = ~1'b0 ;
  assign y2220 = ~n5195 ;
  assign y2221 = ~n5199 ;
  assign y2222 = ~n5203 ;
  assign y2223 = ~1'b0 ;
  assign y2224 = ~n5207 ;
  assign y2225 = n5212 ;
  assign y2226 = ~n5214 ;
  assign y2227 = n5216 ;
  assign y2228 = ~n5223 ;
  assign y2229 = ~n4520 ;
  assign y2230 = ~1'b0 ;
  assign y2231 = ~1'b0 ;
  assign y2232 = ~n5225 ;
  assign y2233 = ~n2383 ;
  assign y2234 = ~1'b0 ;
  assign y2235 = ~n5227 ;
  assign y2236 = ~1'b0 ;
  assign y2237 = ~n5231 ;
  assign y2238 = n3929 ;
  assign y2239 = ~n5234 ;
  assign y2240 = ~1'b0 ;
  assign y2241 = ~n5236 ;
  assign y2242 = ~n5240 ;
  assign y2243 = ~n5241 ;
  assign y2244 = ~n5242 ;
  assign y2245 = ~n5245 ;
  assign y2246 = ~n5252 ;
  assign y2247 = n5253 ;
  assign y2248 = 1'b0 ;
  assign y2249 = n5256 ;
  assign y2250 = n5259 ;
  assign y2251 = n5262 ;
  assign y2252 = ~n5269 ;
  assign y2253 = n5270 ;
  assign y2254 = n5272 ;
  assign y2255 = ~1'b0 ;
  assign y2256 = ~1'b0 ;
  assign y2257 = ~1'b0 ;
  assign y2258 = ~1'b0 ;
  assign y2259 = ~1'b0 ;
  assign y2260 = n5273 ;
  assign y2261 = ~1'b0 ;
  assign y2262 = 1'b0 ;
  assign y2263 = ~1'b0 ;
  assign y2264 = n5276 ;
  assign y2265 = ~1'b0 ;
  assign y2266 = n5286 ;
  assign y2267 = ~n5288 ;
  assign y2268 = n5292 ;
  assign y2269 = ~1'b0 ;
  assign y2270 = ~n5295 ;
  assign y2271 = ~n5298 ;
  assign y2272 = ~1'b0 ;
  assign y2273 = ~1'b0 ;
  assign y2274 = n5301 ;
  assign y2275 = ~n5302 ;
  assign y2276 = ~n5303 ;
  assign y2277 = n1522 ;
  assign y2278 = ~n5305 ;
  assign y2279 = n5313 ;
  assign y2280 = ~n5317 ;
  assign y2281 = ~n5320 ;
  assign y2282 = n5322 ;
  assign y2283 = ~1'b0 ;
  assign y2284 = n5325 ;
  assign y2285 = n3440 ;
  assign y2286 = ~1'b0 ;
  assign y2287 = ~n5326 ;
  assign y2288 = ~n5328 ;
  assign y2289 = ~n5330 ;
  assign y2290 = ~1'b0 ;
  assign y2291 = ~n5334 ;
  assign y2292 = n5335 ;
  assign y2293 = n5336 ;
  assign y2294 = n5340 ;
  assign y2295 = n5341 ;
  assign y2296 = ~n5347 ;
  assign y2297 = ~1'b0 ;
  assign y2298 = n5349 ;
  assign y2299 = n5355 ;
  assign y2300 = n5356 ;
  assign y2301 = n5357 ;
  assign y2302 = ~1'b0 ;
  assign y2303 = n5360 ;
  assign y2304 = n5364 ;
  assign y2305 = ~1'b0 ;
  assign y2306 = ~1'b0 ;
  assign y2307 = ~n5366 ;
  assign y2308 = ~n5369 ;
  assign y2309 = ~n5371 ;
  assign y2310 = ~1'b0 ;
  assign y2311 = ~1'b0 ;
  assign y2312 = n5375 ;
  assign y2313 = ~n5380 ;
  assign y2314 = ~1'b0 ;
  assign y2315 = ~1'b0 ;
  assign y2316 = n5386 ;
  assign y2317 = ~1'b0 ;
  assign y2318 = ~n5388 ;
  assign y2319 = ~n5392 ;
  assign y2320 = n5393 ;
  assign y2321 = n5400 ;
  assign y2322 = ~1'b0 ;
  assign y2323 = n4428 ;
  assign y2324 = ~1'b0 ;
  assign y2325 = ~n5401 ;
  assign y2326 = ~1'b0 ;
  assign y2327 = ~n5403 ;
  assign y2328 = n5406 ;
  assign y2329 = n5409 ;
  assign y2330 = ~n5412 ;
  assign y2331 = ~n5414 ;
  assign y2332 = ~n5416 ;
  assign y2333 = n5421 ;
  assign y2334 = ~n5422 ;
  assign y2335 = ~n5423 ;
  assign y2336 = ~1'b0 ;
  assign y2337 = ~n5427 ;
  assign y2338 = n5428 ;
  assign y2339 = ~n302 ;
  assign y2340 = n5431 ;
  assign y2341 = n4065 ;
  assign y2342 = n5432 ;
  assign y2343 = ~1'b0 ;
  assign y2344 = ~1'b0 ;
  assign y2345 = n1997 ;
  assign y2346 = n5437 ;
  assign y2347 = ~n5438 ;
  assign y2348 = ~n2065 ;
  assign y2349 = ~1'b0 ;
  assign y2350 = ~1'b0 ;
  assign y2351 = ~n5163 ;
  assign y2352 = n5440 ;
  assign y2353 = ~n5442 ;
  assign y2354 = ~1'b0 ;
  assign y2355 = ~n5446 ;
  assign y2356 = ~n5458 ;
  assign y2357 = ~n5471 ;
  assign y2358 = ~1'b0 ;
  assign y2359 = ~1'b0 ;
  assign y2360 = ~n4770 ;
  assign y2361 = n2819 ;
  assign y2362 = n5473 ;
  assign y2363 = n5474 ;
  assign y2364 = ~1'b0 ;
  assign y2365 = n5476 ;
  assign y2366 = 1'b0 ;
  assign y2367 = ~1'b0 ;
  assign y2368 = ~n2944 ;
  assign y2369 = n5479 ;
  assign y2370 = ~n5481 ;
  assign y2371 = n5482 ;
  assign y2372 = ~1'b0 ;
  assign y2373 = ~1'b0 ;
  assign y2374 = ~n5485 ;
  assign y2375 = ~1'b0 ;
  assign y2376 = ~n5494 ;
  assign y2377 = n5497 ;
  assign y2378 = ~1'b0 ;
  assign y2379 = n5507 ;
  assign y2380 = n5509 ;
  assign y2381 = ~n5510 ;
  assign y2382 = ~1'b0 ;
  assign y2383 = ~n5512 ;
  assign y2384 = n5515 ;
  assign y2385 = ~1'b0 ;
  assign y2386 = n5517 ;
  assign y2387 = n5522 ;
  assign y2388 = 1'b0 ;
  assign y2389 = n5529 ;
  assign y2390 = ~1'b0 ;
  assign y2391 = n5530 ;
  assign y2392 = ~1'b0 ;
  assign y2393 = n5535 ;
  assign y2394 = n5536 ;
  assign y2395 = ~1'b0 ;
  assign y2396 = ~1'b0 ;
  assign y2397 = n943 ;
  assign y2398 = ~n2322 ;
  assign y2399 = ~n5539 ;
  assign y2400 = n5540 ;
  assign y2401 = ~1'b0 ;
  assign y2402 = ~1'b0 ;
  assign y2403 = ~n2625 ;
  assign y2404 = ~n5542 ;
  assign y2405 = n5549 ;
  assign y2406 = n5553 ;
  assign y2407 = ~1'b0 ;
  assign y2408 = 1'b0 ;
  assign y2409 = ~n5554 ;
  assign y2410 = n5556 ;
  assign y2411 = ~n5559 ;
  assign y2412 = n5568 ;
  assign y2413 = ~1'b0 ;
  assign y2414 = ~1'b0 ;
  assign y2415 = ~n5573 ;
  assign y2416 = ~1'b0 ;
  assign y2417 = ~1'b0 ;
  assign y2418 = ~n5574 ;
  assign y2419 = n5576 ;
  assign y2420 = n5578 ;
  assign y2421 = ~n5583 ;
  assign y2422 = ~n5585 ;
  assign y2423 = ~n5594 ;
  assign y2424 = n5595 ;
  assign y2425 = ~1'b0 ;
  assign y2426 = 1'b0 ;
  assign y2427 = ~n2622 ;
  assign y2428 = n5598 ;
  assign y2429 = ~1'b0 ;
  assign y2430 = ~n5605 ;
  assign y2431 = ~1'b0 ;
  assign y2432 = ~1'b0 ;
  assign y2433 = ~1'b0 ;
  assign y2434 = ~1'b0 ;
  assign y2435 = ~n5606 ;
  assign y2436 = ~1'b0 ;
  assign y2437 = n5607 ;
  assign y2438 = ~1'b0 ;
  assign y2439 = n5613 ;
  assign y2440 = ~n5614 ;
  assign y2441 = 1'b0 ;
  assign y2442 = ~n5617 ;
  assign y2443 = n5622 ;
  assign y2444 = n5625 ;
  assign y2445 = n5628 ;
  assign y2446 = ~1'b0 ;
  assign y2447 = ~1'b0 ;
  assign y2448 = n5632 ;
  assign y2449 = ~1'b0 ;
  assign y2450 = 1'b0 ;
  assign y2451 = n5634 ;
  assign y2452 = ~n5637 ;
  assign y2453 = ~1'b0 ;
  assign y2454 = ~1'b0 ;
  assign y2455 = ~n5642 ;
  assign y2456 = ~1'b0 ;
  assign y2457 = ~x20 ;
  assign y2458 = ~1'b0 ;
  assign y2459 = ~n5649 ;
  assign y2460 = ~n5650 ;
  assign y2461 = ~1'b0 ;
  assign y2462 = ~1'b0 ;
  assign y2463 = ~n5654 ;
  assign y2464 = n5659 ;
  assign y2465 = ~1'b0 ;
  assign y2466 = ~1'b0 ;
  assign y2467 = n5664 ;
  assign y2468 = ~n5665 ;
  assign y2469 = n5668 ;
  assign y2470 = ~n5675 ;
  assign y2471 = ~1'b0 ;
  assign y2472 = ~n5683 ;
  assign y2473 = ~1'b0 ;
  assign y2474 = ~1'b0 ;
  assign y2475 = ~n5685 ;
  assign y2476 = n5686 ;
  assign y2477 = n5697 ;
  assign y2478 = n5698 ;
  assign y2479 = ~n5700 ;
  assign y2480 = n5703 ;
  assign y2481 = ~n5708 ;
  assign y2482 = n5713 ;
  assign y2483 = n5717 ;
  assign y2484 = ~n5719 ;
  assign y2485 = ~n890 ;
  assign y2486 = ~1'b0 ;
  assign y2487 = ~n5727 ;
  assign y2488 = ~n5728 ;
  assign y2489 = n5729 ;
  assign y2490 = ~1'b0 ;
  assign y2491 = ~n2715 ;
  assign y2492 = ~n5733 ;
  assign y2493 = ~n5735 ;
  assign y2494 = ~1'b0 ;
  assign y2495 = ~1'b0 ;
  assign y2496 = ~1'b0 ;
  assign y2497 = ~n5745 ;
  assign y2498 = n5746 ;
  assign y2499 = n5748 ;
  assign y2500 = n5749 ;
  assign y2501 = 1'b0 ;
  assign y2502 = ~n5763 ;
  assign y2503 = ~1'b0 ;
  assign y2504 = ~1'b0 ;
  assign y2505 = ~n5765 ;
  assign y2506 = 1'b0 ;
  assign y2507 = ~1'b0 ;
  assign y2508 = ~n2901 ;
  assign y2509 = ~n5768 ;
  assign y2510 = ~1'b0 ;
  assign y2511 = ~n5769 ;
  assign y2512 = ~n5771 ;
  assign y2513 = n5772 ;
  assign y2514 = ~1'b0 ;
  assign y2515 = n5773 ;
  assign y2516 = ~n5774 ;
  assign y2517 = ~n5780 ;
  assign y2518 = n5783 ;
  assign y2519 = n5788 ;
  assign y2520 = ~1'b0 ;
  assign y2521 = n5794 ;
  assign y2522 = n5795 ;
  assign y2523 = ~1'b0 ;
  assign y2524 = ~n5797 ;
  assign y2525 = n5802 ;
  assign y2526 = ~1'b0 ;
  assign y2527 = n5803 ;
  assign y2528 = ~1'b0 ;
  assign y2529 = n4442 ;
  assign y2530 = ~n5806 ;
  assign y2531 = ~1'b0 ;
  assign y2532 = ~n5813 ;
  assign y2533 = ~n5816 ;
  assign y2534 = ~n5823 ;
  assign y2535 = ~1'b0 ;
  assign y2536 = n5825 ;
  assign y2537 = ~1'b0 ;
  assign y2538 = n5827 ;
  assign y2539 = ~n5829 ;
  assign y2540 = ~1'b0 ;
  assign y2541 = ~1'b0 ;
  assign y2542 = ~n4027 ;
  assign y2543 = n5208 ;
  assign y2544 = ~n5835 ;
  assign y2545 = ~1'b0 ;
  assign y2546 = n5836 ;
  assign y2547 = ~1'b0 ;
  assign y2548 = n5837 ;
  assign y2549 = n5838 ;
  assign y2550 = ~1'b0 ;
  assign y2551 = ~n5839 ;
  assign y2552 = n5849 ;
  assign y2553 = ~n5851 ;
  assign y2554 = ~n5862 ;
  assign y2555 = n5864 ;
  assign y2556 = ~1'b0 ;
  assign y2557 = ~n5865 ;
  assign y2558 = n708 ;
  assign y2559 = n5866 ;
  assign y2560 = ~1'b0 ;
  assign y2561 = n5869 ;
  assign y2562 = n5870 ;
  assign y2563 = ~1'b0 ;
  assign y2564 = ~n5879 ;
  assign y2565 = n5883 ;
  assign y2566 = ~1'b0 ;
  assign y2567 = ~1'b0 ;
  assign y2568 = ~1'b0 ;
  assign y2569 = n5890 ;
  assign y2570 = ~n5891 ;
  assign y2571 = ~n5894 ;
  assign y2572 = ~n5895 ;
  assign y2573 = ~n5896 ;
  assign y2574 = ~n5900 ;
  assign y2575 = ~n5905 ;
  assign y2576 = ~x48 ;
  assign y2577 = n5908 ;
  assign y2578 = ~n5911 ;
  assign y2579 = n3710 ;
  assign y2580 = ~n5913 ;
  assign y2581 = ~1'b0 ;
  assign y2582 = n5917 ;
  assign y2583 = n5924 ;
  assign y2584 = ~1'b0 ;
  assign y2585 = ~1'b0 ;
  assign y2586 = ~1'b0 ;
  assign y2587 = ~n3646 ;
  assign y2588 = ~n3326 ;
  assign y2589 = ~n5927 ;
  assign y2590 = n5928 ;
  assign y2591 = ~1'b0 ;
  assign y2592 = ~1'b0 ;
  assign y2593 = ~n1048 ;
  assign y2594 = ~1'b0 ;
  assign y2595 = n5930 ;
  assign y2596 = n845 ;
  assign y2597 = n5934 ;
  assign y2598 = ~1'b0 ;
  assign y2599 = ~n5936 ;
  assign y2600 = n5939 ;
  assign y2601 = n5941 ;
  assign y2602 = n5943 ;
  assign y2603 = ~1'b0 ;
  assign y2604 = n5944 ;
  assign y2605 = ~n5951 ;
  assign y2606 = ~n5957 ;
  assign y2607 = ~n5959 ;
  assign y2608 = n5961 ;
  assign y2609 = ~n5962 ;
  assign y2610 = n5966 ;
  assign y2611 = ~n5967 ;
  assign y2612 = ~n5971 ;
  assign y2613 = n5975 ;
  assign y2614 = ~n5034 ;
  assign y2615 = n5976 ;
  assign y2616 = ~1'b0 ;
  assign y2617 = n5978 ;
  assign y2618 = ~1'b0 ;
  assign y2619 = ~n5980 ;
  assign y2620 = ~1'b0 ;
  assign y2621 = ~n5984 ;
  assign y2622 = ~1'b0 ;
  assign y2623 = n5986 ;
  assign y2624 = ~n5992 ;
  assign y2625 = n5995 ;
  assign y2626 = n5996 ;
  assign y2627 = ~1'b0 ;
  assign y2628 = ~1'b0 ;
  assign y2629 = ~n1369 ;
  assign y2630 = n5999 ;
  assign y2631 = n6005 ;
  assign y2632 = ~n6006 ;
  assign y2633 = n6009 ;
  assign y2634 = ~n6010 ;
  assign y2635 = ~1'b0 ;
  assign y2636 = ~n6014 ;
  assign y2637 = n6015 ;
  assign y2638 = n4503 ;
  assign y2639 = ~1'b0 ;
  assign y2640 = 1'b0 ;
  assign y2641 = ~n6018 ;
  assign y2642 = ~1'b0 ;
  assign y2643 = ~1'b0 ;
  assign y2644 = ~x112 ;
  assign y2645 = ~1'b0 ;
  assign y2646 = n6019 ;
  assign y2647 = ~1'b0 ;
  assign y2648 = ~1'b0 ;
  assign y2649 = n6024 ;
  assign y2650 = ~n6025 ;
  assign y2651 = ~1'b0 ;
  assign y2652 = ~n6027 ;
  assign y2653 = ~1'b0 ;
  assign y2654 = n6035 ;
  assign y2655 = n453 ;
  assign y2656 = n6036 ;
  assign y2657 = ~n6040 ;
  assign y2658 = ~n6042 ;
  assign y2659 = ~1'b0 ;
  assign y2660 = ~n6043 ;
  assign y2661 = ~1'b0 ;
  assign y2662 = ~1'b0 ;
  assign y2663 = ~1'b0 ;
  assign y2664 = ~1'b0 ;
  assign y2665 = 1'b0 ;
  assign y2666 = ~n6046 ;
  assign y2667 = ~1'b0 ;
  assign y2668 = ~1'b0 ;
  assign y2669 = n6055 ;
  assign y2670 = n6058 ;
  assign y2671 = n6061 ;
  assign y2672 = n6066 ;
  assign y2673 = ~1'b0 ;
  assign y2674 = ~n6072 ;
  assign y2675 = ~n5540 ;
  assign y2676 = ~n6073 ;
  assign y2677 = ~n6075 ;
  assign y2678 = ~n6081 ;
  assign y2679 = ~n6085 ;
  assign y2680 = ~n6086 ;
  assign y2681 = ~n6091 ;
  assign y2682 = ~n6097 ;
  assign y2683 = n6098 ;
  assign y2684 = ~n3411 ;
  assign y2685 = ~1'b0 ;
  assign y2686 = ~1'b0 ;
  assign y2687 = n6102 ;
  assign y2688 = n6114 ;
  assign y2689 = ~1'b0 ;
  assign y2690 = n957 ;
  assign y2691 = ~n6115 ;
  assign y2692 = ~1'b0 ;
  assign y2693 = n6117 ;
  assign y2694 = ~n4905 ;
  assign y2695 = ~1'b0 ;
  assign y2696 = n6120 ;
  assign y2697 = n6121 ;
  assign y2698 = ~n6125 ;
  assign y2699 = ~n6128 ;
  assign y2700 = ~1'b0 ;
  assign y2701 = ~1'b0 ;
  assign y2702 = n6134 ;
  assign y2703 = ~n6137 ;
  assign y2704 = n6139 ;
  assign y2705 = ~1'b0 ;
  assign y2706 = ~n6144 ;
  assign y2707 = n6146 ;
  assign y2708 = n6148 ;
  assign y2709 = n6152 ;
  assign y2710 = ~1'b0 ;
  assign y2711 = ~n6154 ;
  assign y2712 = ~1'b0 ;
  assign y2713 = n6158 ;
  assign y2714 = ~1'b0 ;
  assign y2715 = ~1'b0 ;
  assign y2716 = ~n6160 ;
  assign y2717 = n6163 ;
  assign y2718 = ~n6164 ;
  assign y2719 = n6166 ;
  assign y2720 = ~n6173 ;
  assign y2721 = ~n6175 ;
  assign y2722 = ~1'b0 ;
  assign y2723 = ~n6177 ;
  assign y2724 = n6180 ;
  assign y2725 = n6184 ;
  assign y2726 = ~n6197 ;
  assign y2727 = n6112 ;
  assign y2728 = ~1'b0 ;
  assign y2729 = ~n6198 ;
  assign y2730 = ~n6199 ;
  assign y2731 = n6200 ;
  assign y2732 = n6203 ;
  assign y2733 = n6204 ;
  assign y2734 = ~x180 ;
  assign y2735 = ~n6207 ;
  assign y2736 = ~1'b0 ;
  assign y2737 = n1111 ;
  assign y2738 = n6208 ;
  assign y2739 = ~n6210 ;
  assign y2740 = ~n6212 ;
  assign y2741 = ~n6218 ;
  assign y2742 = ~1'b0 ;
  assign y2743 = ~n6219 ;
  assign y2744 = n6222 ;
  assign y2745 = ~n6225 ;
  assign y2746 = ~1'b0 ;
  assign y2747 = n6238 ;
  assign y2748 = ~n6241 ;
  assign y2749 = ~n865 ;
  assign y2750 = n6243 ;
  assign y2751 = ~1'b0 ;
  assign y2752 = ~n6251 ;
  assign y2753 = ~1'b0 ;
  assign y2754 = ~1'b0 ;
  assign y2755 = n6254 ;
  assign y2756 = ~1'b0 ;
  assign y2757 = ~n6255 ;
  assign y2758 = ~n6263 ;
  assign y2759 = ~n6265 ;
  assign y2760 = n6267 ;
  assign y2761 = ~n6268 ;
  assign y2762 = ~n6278 ;
  assign y2763 = ~n6280 ;
  assign y2764 = ~1'b0 ;
  assign y2765 = ~1'b0 ;
  assign y2766 = ~n6281 ;
  assign y2767 = ~n6289 ;
  assign y2768 = n6293 ;
  assign y2769 = ~1'b0 ;
  assign y2770 = ~n6297 ;
  assign y2771 = ~1'b0 ;
  assign y2772 = n4260 ;
  assign y2773 = n6299 ;
  assign y2774 = n6300 ;
  assign y2775 = ~1'b0 ;
  assign y2776 = n1129 ;
  assign y2777 = ~1'b0 ;
  assign y2778 = ~n6305 ;
  assign y2779 = n6307 ;
  assign y2780 = ~n6309 ;
  assign y2781 = ~n6315 ;
  assign y2782 = ~1'b0 ;
  assign y2783 = n2286 ;
  assign y2784 = ~1'b0 ;
  assign y2785 = ~n625 ;
  assign y2786 = ~1'b0 ;
  assign y2787 = n6318 ;
  assign y2788 = ~1'b0 ;
  assign y2789 = ~1'b0 ;
  assign y2790 = n4516 ;
  assign y2791 = n6319 ;
  assign y2792 = ~1'b0 ;
  assign y2793 = ~1'b0 ;
  assign y2794 = ~1'b0 ;
  assign y2795 = ~n6321 ;
  assign y2796 = n6325 ;
  assign y2797 = ~1'b0 ;
  assign y2798 = ~n6326 ;
  assign y2799 = ~1'b0 ;
  assign y2800 = ~1'b0 ;
  assign y2801 = n6177 ;
  assign y2802 = ~n6327 ;
  assign y2803 = n6331 ;
  assign y2804 = ~n6335 ;
  assign y2805 = n6337 ;
  assign y2806 = ~n6338 ;
  assign y2807 = n6340 ;
  assign y2808 = n6341 ;
  assign y2809 = ~1'b0 ;
  assign y2810 = ~n6345 ;
  assign y2811 = ~1'b0 ;
  assign y2812 = ~n6347 ;
  assign y2813 = n6350 ;
  assign y2814 = ~1'b0 ;
  assign y2815 = ~n6353 ;
  assign y2816 = ~1'b0 ;
  assign y2817 = ~1'b0 ;
  assign y2818 = ~n6354 ;
  assign y2819 = n6355 ;
  assign y2820 = n6361 ;
  assign y2821 = ~n6363 ;
  assign y2822 = ~n6369 ;
  assign y2823 = ~1'b0 ;
  assign y2824 = ~1'b0 ;
  assign y2825 = ~1'b0 ;
  assign y2826 = ~n6378 ;
  assign y2827 = ~n6386 ;
  assign y2828 = ~n6389 ;
  assign y2829 = ~n6393 ;
  assign y2830 = ~n6399 ;
  assign y2831 = 1'b0 ;
  assign y2832 = ~1'b0 ;
  assign y2833 = n6405 ;
  assign y2834 = ~n6406 ;
  assign y2835 = ~n6409 ;
  assign y2836 = n6411 ;
  assign y2837 = n6412 ;
  assign y2838 = ~1'b0 ;
  assign y2839 = ~n6416 ;
  assign y2840 = ~n6417 ;
  assign y2841 = ~n6419 ;
  assign y2842 = n464 ;
  assign y2843 = ~n6423 ;
  assign y2844 = 1'b0 ;
  assign y2845 = ~1'b0 ;
  assign y2846 = ~1'b0 ;
  assign y2847 = n6428 ;
  assign y2848 = ~n6429 ;
  assign y2849 = n6433 ;
  assign y2850 = ~n6434 ;
  assign y2851 = ~n6436 ;
  assign y2852 = ~n6440 ;
  assign y2853 = ~n6441 ;
  assign y2854 = n3202 ;
  assign y2855 = ~n6446 ;
  assign y2856 = ~n6450 ;
  assign y2857 = n4610 ;
  assign y2858 = ~1'b0 ;
  assign y2859 = ~n6462 ;
  assign y2860 = 1'b0 ;
  assign y2861 = ~n2525 ;
  assign y2862 = ~n6464 ;
  assign y2863 = n2249 ;
  assign y2864 = ~n6409 ;
  assign y2865 = n6467 ;
  assign y2866 = ~n6471 ;
  assign y2867 = n274 ;
  assign y2868 = n6473 ;
  assign y2869 = n6475 ;
  assign y2870 = ~n6479 ;
  assign y2871 = ~n6481 ;
  assign y2872 = n6489 ;
  assign y2873 = ~1'b0 ;
  assign y2874 = n6495 ;
  assign y2875 = n6496 ;
  assign y2876 = n6499 ;
  assign y2877 = ~1'b0 ;
  assign y2878 = ~n6500 ;
  assign y2879 = n6504 ;
  assign y2880 = ~1'b0 ;
  assign y2881 = ~n6510 ;
  assign y2882 = ~n6512 ;
  assign y2883 = ~1'b0 ;
  assign y2884 = ~n6514 ;
  assign y2885 = ~1'b0 ;
  assign y2886 = ~1'b0 ;
  assign y2887 = ~1'b0 ;
  assign y2888 = n6522 ;
  assign y2889 = ~1'b0 ;
  assign y2890 = n6525 ;
  assign y2891 = n6526 ;
  assign y2892 = ~n6527 ;
  assign y2893 = ~n6537 ;
  assign y2894 = ~1'b0 ;
  assign y2895 = ~n6539 ;
  assign y2896 = n6542 ;
  assign y2897 = ~1'b0 ;
  assign y2898 = n6547 ;
  assign y2899 = n6553 ;
  assign y2900 = ~n6555 ;
  assign y2901 = ~n6559 ;
  assign y2902 = ~1'b0 ;
  assign y2903 = ~n6560 ;
  assign y2904 = ~n6566 ;
  assign y2905 = ~n6571 ;
  assign y2906 = ~1'b0 ;
  assign y2907 = ~1'b0 ;
  assign y2908 = ~1'b0 ;
  assign y2909 = ~n6574 ;
  assign y2910 = n6576 ;
  assign y2911 = n6580 ;
  assign y2912 = ~1'b0 ;
  assign y2913 = ~1'b0 ;
  assign y2914 = ~n6581 ;
  assign y2915 = n6583 ;
  assign y2916 = ~n6591 ;
  assign y2917 = n6592 ;
  assign y2918 = ~1'b0 ;
  assign y2919 = ~n6593 ;
  assign y2920 = ~1'b0 ;
  assign y2921 = n6597 ;
  assign y2922 = ~1'b0 ;
  assign y2923 = ~1'b0 ;
  assign y2924 = ~1'b0 ;
  assign y2925 = n3707 ;
  assign y2926 = ~n6603 ;
  assign y2927 = ~1'b0 ;
  assign y2928 = ~n6604 ;
  assign y2929 = ~1'b0 ;
  assign y2930 = n6605 ;
  assign y2931 = ~n6606 ;
  assign y2932 = ~n6607 ;
  assign y2933 = ~1'b0 ;
  assign y2934 = ~n6615 ;
  assign y2935 = ~n1261 ;
  assign y2936 = ~1'b0 ;
  assign y2937 = ~n6618 ;
  assign y2938 = n6619 ;
  assign y2939 = n6621 ;
  assign y2940 = n6626 ;
  assign y2941 = n6636 ;
  assign y2942 = ~1'b0 ;
  assign y2943 = ~1'b0 ;
  assign y2944 = ~1'b0 ;
  assign y2945 = n6640 ;
  assign y2946 = ~1'b0 ;
  assign y2947 = n6648 ;
  assign y2948 = ~n6652 ;
  assign y2949 = ~n6653 ;
  assign y2950 = ~n6654 ;
  assign y2951 = n6657 ;
  assign y2952 = ~1'b0 ;
  assign y2953 = ~1'b0 ;
  assign y2954 = ~n6660 ;
  assign y2955 = ~n6662 ;
  assign y2956 = ~n6666 ;
  assign y2957 = ~n6668 ;
  assign y2958 = n6670 ;
  assign y2959 = ~1'b0 ;
  assign y2960 = n6672 ;
  assign y2961 = ~1'b0 ;
  assign y2962 = n6674 ;
  assign y2963 = ~n6676 ;
  assign y2964 = ~1'b0 ;
  assign y2965 = n6677 ;
  assign y2966 = ~1'b0 ;
  assign y2967 = n6679 ;
  assign y2968 = ~n6688 ;
  assign y2969 = n6690 ;
  assign y2970 = ~n6694 ;
  assign y2971 = n6699 ;
  assign y2972 = n6701 ;
  assign y2973 = ~n6705 ;
  assign y2974 = n2831 ;
  assign y2975 = n6709 ;
  assign y2976 = n6714 ;
  assign y2977 = ~n6718 ;
  assign y2978 = ~1'b0 ;
  assign y2979 = ~n6719 ;
  assign y2980 = ~n6722 ;
  assign y2981 = ~n6723 ;
  assign y2982 = n6730 ;
  assign y2983 = ~x192 ;
  assign y2984 = ~n6731 ;
  assign y2985 = n6735 ;
  assign y2986 = ~1'b0 ;
  assign y2987 = ~1'b0 ;
  assign y2988 = ~n6741 ;
  assign y2989 = ~1'b0 ;
  assign y2990 = 1'b0 ;
  assign y2991 = ~n6750 ;
  assign y2992 = n6751 ;
  assign y2993 = ~1'b0 ;
  assign y2994 = ~n6753 ;
  assign y2995 = ~1'b0 ;
  assign y2996 = ~1'b0 ;
  assign y2997 = n6755 ;
  assign y2998 = ~1'b0 ;
  assign y2999 = n6759 ;
  assign y3000 = ~n6763 ;
  assign y3001 = 1'b0 ;
  assign y3002 = n6769 ;
  assign y3003 = ~1'b0 ;
  assign y3004 = 1'b0 ;
  assign y3005 = n6772 ;
  assign y3006 = ~1'b0 ;
  assign y3007 = n6776 ;
  assign y3008 = ~n6778 ;
  assign y3009 = n6781 ;
  assign y3010 = ~1'b0 ;
  assign y3011 = n6783 ;
  assign y3012 = ~1'b0 ;
  assign y3013 = 1'b0 ;
  assign y3014 = ~n6788 ;
  assign y3015 = n1815 ;
  assign y3016 = ~1'b0 ;
  assign y3017 = n6789 ;
  assign y3018 = ~n6793 ;
  assign y3019 = n6797 ;
  assign y3020 = ~1'b0 ;
  assign y3021 = ~n6800 ;
  assign y3022 = ~1'b0 ;
  assign y3023 = ~1'b0 ;
  assign y3024 = ~n6807 ;
  assign y3025 = ~n6809 ;
  assign y3026 = n4031 ;
  assign y3027 = ~1'b0 ;
  assign y3028 = n6812 ;
  assign y3029 = 1'b0 ;
  assign y3030 = n911 ;
  assign y3031 = ~n6818 ;
  assign y3032 = 1'b0 ;
  assign y3033 = ~n6820 ;
  assign y3034 = ~n6821 ;
  assign y3035 = ~1'b0 ;
  assign y3036 = ~1'b0 ;
  assign y3037 = ~n6831 ;
  assign y3038 = ~n6833 ;
  assign y3039 = ~1'b0 ;
  assign y3040 = ~n6840 ;
  assign y3041 = ~n2708 ;
  assign y3042 = ~1'b0 ;
  assign y3043 = ~n6844 ;
  assign y3044 = n6850 ;
  assign y3045 = ~n1890 ;
  assign y3046 = ~n6853 ;
  assign y3047 = ~1'b0 ;
  assign y3048 = ~n6854 ;
  assign y3049 = ~n6859 ;
  assign y3050 = n2903 ;
  assign y3051 = ~1'b0 ;
  assign y3052 = ~1'b0 ;
  assign y3053 = ~n6861 ;
  assign y3054 = ~1'b0 ;
  assign y3055 = ~1'b0 ;
  assign y3056 = ~1'b0 ;
  assign y3057 = ~1'b0 ;
  assign y3058 = ~n6862 ;
  assign y3059 = n6865 ;
  assign y3060 = ~n6868 ;
  assign y3061 = n6874 ;
  assign y3062 = n6875 ;
  assign y3063 = ~1'b0 ;
  assign y3064 = ~n6879 ;
  assign y3065 = n6881 ;
  assign y3066 = 1'b0 ;
  assign y3067 = ~1'b0 ;
  assign y3068 = 1'b0 ;
  assign y3069 = ~1'b0 ;
  assign y3070 = n6889 ;
  assign y3071 = ~1'b0 ;
  assign y3072 = 1'b0 ;
  assign y3073 = n6891 ;
  assign y3074 = ~n6893 ;
  assign y3075 = n6896 ;
  assign y3076 = ~n6900 ;
  assign y3077 = ~n6902 ;
  assign y3078 = n6903 ;
  assign y3079 = n6907 ;
  assign y3080 = n5690 ;
  assign y3081 = ~1'b0 ;
  assign y3082 = n1338 ;
  assign y3083 = ~n6908 ;
  assign y3084 = n6914 ;
  assign y3085 = ~n6916 ;
  assign y3086 = ~1'b0 ;
  assign y3087 = ~n6919 ;
  assign y3088 = n6925 ;
  assign y3089 = n6930 ;
  assign y3090 = ~n6933 ;
  assign y3091 = ~1'b0 ;
  assign y3092 = ~n6935 ;
  assign y3093 = 1'b0 ;
  assign y3094 = ~1'b0 ;
  assign y3095 = n6941 ;
  assign y3096 = ~n6951 ;
  assign y3097 = n6956 ;
  assign y3098 = n6960 ;
  assign y3099 = ~1'b0 ;
  assign y3100 = ~n6964 ;
  assign y3101 = ~n6965 ;
  assign y3102 = n6971 ;
  assign y3103 = n6972 ;
  assign y3104 = ~n6974 ;
  assign y3105 = ~1'b0 ;
  assign y3106 = ~n6976 ;
  assign y3107 = n3265 ;
  assign y3108 = n6978 ;
  assign y3109 = n6982 ;
  assign y3110 = n6983 ;
  assign y3111 = n6986 ;
  assign y3112 = n6989 ;
  assign y3113 = n6990 ;
  assign y3114 = n6992 ;
  assign y3115 = n6998 ;
  assign y3116 = ~n432 ;
  assign y3117 = ~n6999 ;
  assign y3118 = ~1'b0 ;
  assign y3119 = ~n7000 ;
  assign y3120 = ~n7002 ;
  assign y3121 = ~1'b0 ;
  assign y3122 = n7005 ;
  assign y3123 = ~1'b0 ;
  assign y3124 = n7006 ;
  assign y3125 = ~1'b0 ;
  assign y3126 = n7018 ;
  assign y3127 = n7019 ;
  assign y3128 = ~n7020 ;
  assign y3129 = n7025 ;
  assign y3130 = n7027 ;
  assign y3131 = ~1'b0 ;
  assign y3132 = ~n7029 ;
  assign y3133 = ~1'b0 ;
  assign y3134 = ~n7032 ;
  assign y3135 = n7038 ;
  assign y3136 = n7041 ;
  assign y3137 = n7045 ;
  assign y3138 = ~n7046 ;
  assign y3139 = 1'b0 ;
  assign y3140 = ~n7048 ;
  assign y3141 = ~1'b0 ;
  assign y3142 = ~n3805 ;
  assign y3143 = n7050 ;
  assign y3144 = n7051 ;
  assign y3145 = ~1'b0 ;
  assign y3146 = ~n7057 ;
  assign y3147 = ~n7063 ;
  assign y3148 = n1055 ;
  assign y3149 = ~n585 ;
  assign y3150 = n7066 ;
  assign y3151 = n7067 ;
  assign y3152 = ~n7073 ;
  assign y3153 = ~n7075 ;
  assign y3154 = ~n7078 ;
  assign y3155 = ~1'b0 ;
  assign y3156 = ~n7084 ;
  assign y3157 = n7086 ;
  assign y3158 = ~n7087 ;
  assign y3159 = n7089 ;
  assign y3160 = ~n7090 ;
  assign y3161 = ~n7093 ;
  assign y3162 = ~n7094 ;
  assign y3163 = ~1'b0 ;
  assign y3164 = ~1'b0 ;
  assign y3165 = ~1'b0 ;
  assign y3166 = ~1'b0 ;
  assign y3167 = n7096 ;
  assign y3168 = n7101 ;
  assign y3169 = n7104 ;
  assign y3170 = n7105 ;
  assign y3171 = ~n7107 ;
  assign y3172 = ~1'b0 ;
  assign y3173 = ~x143 ;
  assign y3174 = ~n7110 ;
  assign y3175 = n7113 ;
  assign y3176 = n7117 ;
  assign y3177 = ~n7122 ;
  assign y3178 = ~1'b0 ;
  assign y3179 = ~n7134 ;
  assign y3180 = ~1'b0 ;
  assign y3181 = ~1'b0 ;
  assign y3182 = n7137 ;
  assign y3183 = n7140 ;
  assign y3184 = n7143 ;
  assign y3185 = ~1'b0 ;
  assign y3186 = n7148 ;
  assign y3187 = ~n7150 ;
  assign y3188 = ~1'b0 ;
  assign y3189 = n7152 ;
  assign y3190 = n7154 ;
  assign y3191 = ~n7156 ;
  assign y3192 = ~n7157 ;
  assign y3193 = n7158 ;
  assign y3194 = n7160 ;
  assign y3195 = ~n7161 ;
  assign y3196 = ~n7165 ;
  assign y3197 = ~1'b0 ;
  assign y3198 = ~1'b0 ;
  assign y3199 = 1'b0 ;
  assign y3200 = ~n7168 ;
  assign y3201 = ~n7173 ;
  assign y3202 = 1'b0 ;
  assign y3203 = ~n7175 ;
  assign y3204 = ~n7177 ;
  assign y3205 = ~n7179 ;
  assign y3206 = ~1'b0 ;
  assign y3207 = n7180 ;
  assign y3208 = ~1'b0 ;
  assign y3209 = n6943 ;
  assign y3210 = ~n7183 ;
  assign y3211 = n7190 ;
  assign y3212 = n7191 ;
  assign y3213 = n7193 ;
  assign y3214 = n7195 ;
  assign y3215 = n7196 ;
  assign y3216 = ~n2900 ;
  assign y3217 = ~1'b0 ;
  assign y3218 = ~n7199 ;
  assign y3219 = n7202 ;
  assign y3220 = ~1'b0 ;
  assign y3221 = ~1'b0 ;
  assign y3222 = ~1'b0 ;
  assign y3223 = ~n7203 ;
  assign y3224 = ~n7204 ;
  assign y3225 = n7205 ;
  assign y3226 = n7212 ;
  assign y3227 = n7218 ;
  assign y3228 = ~1'b0 ;
  assign y3229 = n7220 ;
  assign y3230 = ~1'b0 ;
  assign y3231 = n7224 ;
  assign y3232 = ~1'b0 ;
  assign y3233 = ~1'b0 ;
  assign y3234 = n7226 ;
  assign y3235 = n7229 ;
  assign y3236 = ~n7231 ;
  assign y3237 = ~n7232 ;
  assign y3238 = ~1'b0 ;
  assign y3239 = ~n7234 ;
  assign y3240 = ~n7239 ;
  assign y3241 = ~n7243 ;
  assign y3242 = ~1'b0 ;
  assign y3243 = ~n7246 ;
  assign y3244 = ~n6359 ;
  assign y3245 = ~1'b0 ;
  assign y3246 = ~1'b0 ;
  assign y3247 = n7250 ;
  assign y3248 = ~n7265 ;
  assign y3249 = ~1'b0 ;
  assign y3250 = ~1'b0 ;
  assign y3251 = n7270 ;
  assign y3252 = ~1'b0 ;
  assign y3253 = ~1'b0 ;
  assign y3254 = ~1'b0 ;
  assign y3255 = ~1'b0 ;
  assign y3256 = ~n7271 ;
  assign y3257 = ~1'b0 ;
  assign y3258 = ~n7272 ;
  assign y3259 = n7275 ;
  assign y3260 = ~n7283 ;
  assign y3261 = ~1'b0 ;
  assign y3262 = n7285 ;
  assign y3263 = n7286 ;
  assign y3264 = ~n7290 ;
  assign y3265 = ~1'b0 ;
  assign y3266 = ~n7292 ;
  assign y3267 = ~n7294 ;
  assign y3268 = ~1'b0 ;
  assign y3269 = ~n4997 ;
  assign y3270 = n7296 ;
  assign y3271 = ~1'b0 ;
  assign y3272 = ~1'b0 ;
  assign y3273 = n7301 ;
  assign y3274 = n7304 ;
  assign y3275 = ~n7306 ;
  assign y3276 = n7307 ;
  assign y3277 = n7308 ;
  assign y3278 = ~n7314 ;
  assign y3279 = n7315 ;
  assign y3280 = x82 ;
  assign y3281 = ~1'b0 ;
  assign y3282 = n7318 ;
  assign y3283 = n7329 ;
  assign y3284 = n7331 ;
  assign y3285 = ~n7336 ;
  assign y3286 = ~n7345 ;
  assign y3287 = ~n7349 ;
  assign y3288 = n7355 ;
  assign y3289 = n7363 ;
  assign y3290 = ~1'b0 ;
  assign y3291 = ~1'b0 ;
  assign y3292 = ~1'b0 ;
  assign y3293 = n7364 ;
  assign y3294 = n7365 ;
  assign y3295 = ~n7366 ;
  assign y3296 = ~1'b0 ;
  assign y3297 = n7371 ;
  assign y3298 = n7373 ;
  assign y3299 = ~1'b0 ;
  assign y3300 = n7375 ;
  assign y3301 = ~n7383 ;
  assign y3302 = ~n7384 ;
  assign y3303 = ~n7385 ;
  assign y3304 = ~1'b0 ;
  assign y3305 = ~n7386 ;
  assign y3306 = ~n7389 ;
  assign y3307 = ~1'b0 ;
  assign y3308 = n7392 ;
  assign y3309 = ~1'b0 ;
  assign y3310 = n7395 ;
  assign y3311 = ~n7396 ;
  assign y3312 = ~1'b0 ;
  assign y3313 = ~1'b0 ;
  assign y3314 = ~1'b0 ;
  assign y3315 = n7397 ;
  assign y3316 = n7398 ;
  assign y3317 = ~n7399 ;
  assign y3318 = n7401 ;
  assign y3319 = n7402 ;
  assign y3320 = ~1'b0 ;
  assign y3321 = ~n7405 ;
  assign y3322 = n7412 ;
  assign y3323 = ~1'b0 ;
  assign y3324 = n7416 ;
  assign y3325 = ~1'b0 ;
  assign y3326 = ~1'b0 ;
  assign y3327 = n7418 ;
  assign y3328 = ~1'b0 ;
  assign y3329 = ~n7419 ;
  assign y3330 = n7420 ;
  assign y3331 = n7423 ;
  assign y3332 = ~n7424 ;
  assign y3333 = ~1'b0 ;
  assign y3334 = n7426 ;
  assign y3335 = n7427 ;
  assign y3336 = ~1'b0 ;
  assign y3337 = ~n7430 ;
  assign y3338 = n7431 ;
  assign y3339 = ~n7437 ;
  assign y3340 = ~n7442 ;
  assign y3341 = n7443 ;
  assign y3342 = ~n1557 ;
  assign y3343 = n7450 ;
  assign y3344 = ~n7452 ;
  assign y3345 = n7455 ;
  assign y3346 = ~n7463 ;
  assign y3347 = ~1'b0 ;
  assign y3348 = n7469 ;
  assign y3349 = n7472 ;
  assign y3350 = ~1'b0 ;
  assign y3351 = ~n7474 ;
  assign y3352 = n7480 ;
  assign y3353 = n7487 ;
  assign y3354 = n5410 ;
  assign y3355 = ~n7490 ;
  assign y3356 = ~1'b0 ;
  assign y3357 = ~1'b0 ;
  assign y3358 = n7492 ;
  assign y3359 = n7493 ;
  assign y3360 = ~n4993 ;
  assign y3361 = ~n7494 ;
  assign y3362 = ~n7499 ;
  assign y3363 = ~1'b0 ;
  assign y3364 = ~1'b0 ;
  assign y3365 = n7501 ;
  assign y3366 = n7504 ;
  assign y3367 = ~1'b0 ;
  assign y3368 = n7511 ;
  assign y3369 = ~1'b0 ;
  assign y3370 = n7513 ;
  assign y3371 = ~1'b0 ;
  assign y3372 = n7515 ;
  assign y3373 = ~1'b0 ;
  assign y3374 = n7516 ;
  assign y3375 = ~1'b0 ;
  assign y3376 = ~n7522 ;
  assign y3377 = ~n344 ;
  assign y3378 = ~1'b0 ;
  assign y3379 = ~n7523 ;
  assign y3380 = ~1'b0 ;
  assign y3381 = n7524 ;
  assign y3382 = ~n7528 ;
  assign y3383 = ~1'b0 ;
  assign y3384 = n7530 ;
  assign y3385 = ~1'b0 ;
  assign y3386 = ~n7538 ;
  assign y3387 = ~1'b0 ;
  assign y3388 = ~n2988 ;
  assign y3389 = ~n7539 ;
  assign y3390 = ~n3344 ;
  assign y3391 = ~n7541 ;
  assign y3392 = ~n7542 ;
  assign y3393 = ~1'b0 ;
  assign y3394 = ~1'b0 ;
  assign y3395 = ~n7550 ;
  assign y3396 = n2995 ;
  assign y3397 = ~1'b0 ;
  assign y3398 = ~1'b0 ;
  assign y3399 = n7553 ;
  assign y3400 = n7554 ;
  assign y3401 = ~n7557 ;
  assign y3402 = ~n7558 ;
  assign y3403 = ~n2291 ;
  assign y3404 = ~1'b0 ;
  assign y3405 = ~n7561 ;
  assign y3406 = n7563 ;
  assign y3407 = n7564 ;
  assign y3408 = n7565 ;
  assign y3409 = n7568 ;
  assign y3410 = n7569 ;
  assign y3411 = ~1'b0 ;
  assign y3412 = n7570 ;
  assign y3413 = ~n7575 ;
  assign y3414 = ~1'b0 ;
  assign y3415 = ~1'b0 ;
  assign y3416 = n7576 ;
  assign y3417 = n7579 ;
  assign y3418 = n7581 ;
  assign y3419 = ~n7584 ;
  assign y3420 = ~n4803 ;
  assign y3421 = ~1'b0 ;
  assign y3422 = n7587 ;
  assign y3423 = n7593 ;
  assign y3424 = ~1'b0 ;
  assign y3425 = n7596 ;
  assign y3426 = n7605 ;
  assign y3427 = ~1'b0 ;
  assign y3428 = ~1'b0 ;
  assign y3429 = n7608 ;
  assign y3430 = n4757 ;
  assign y3431 = n7611 ;
  assign y3432 = n7038 ;
  assign y3433 = ~n7613 ;
  assign y3434 = n7615 ;
  assign y3435 = ~n7623 ;
  assign y3436 = ~1'b0 ;
  assign y3437 = n7629 ;
  assign y3438 = ~n7634 ;
  assign y3439 = ~n7638 ;
  assign y3440 = n7641 ;
  assign y3441 = ~n7646 ;
  assign y3442 = ~n7651 ;
  assign y3443 = ~n7653 ;
  assign y3444 = ~n7654 ;
  assign y3445 = n7659 ;
  assign y3446 = ~1'b0 ;
  assign y3447 = n7663 ;
  assign y3448 = n7665 ;
  assign y3449 = ~1'b0 ;
  assign y3450 = ~n5754 ;
  assign y3451 = ~n7666 ;
  assign y3452 = ~1'b0 ;
  assign y3453 = n7668 ;
  assign y3454 = ~1'b0 ;
  assign y3455 = ~1'b0 ;
  assign y3456 = ~n7674 ;
  assign y3457 = ~n7676 ;
  assign y3458 = ~1'b0 ;
  assign y3459 = n7681 ;
  assign y3460 = ~1'b0 ;
  assign y3461 = ~1'b0 ;
  assign y3462 = ~n7687 ;
  assign y3463 = ~n7691 ;
  assign y3464 = n7693 ;
  assign y3465 = ~n7699 ;
  assign y3466 = ~1'b0 ;
  assign y3467 = 1'b0 ;
  assign y3468 = ~n7701 ;
  assign y3469 = ~1'b0 ;
  assign y3470 = ~1'b0 ;
  assign y3471 = n7702 ;
  assign y3472 = ~1'b0 ;
  assign y3473 = n7703 ;
  assign y3474 = ~1'b0 ;
  assign y3475 = ~1'b0 ;
  assign y3476 = n7704 ;
  assign y3477 = n5696 ;
  assign y3478 = ~n7707 ;
  assign y3479 = n7711 ;
  assign y3480 = ~n7712 ;
  assign y3481 = ~n7716 ;
  assign y3482 = ~n7722 ;
  assign y3483 = ~n7555 ;
  assign y3484 = n7726 ;
  assign y3485 = n7729 ;
  assign y3486 = n7734 ;
  assign y3487 = n7736 ;
  assign y3488 = ~n7738 ;
  assign y3489 = n7739 ;
  assign y3490 = ~1'b0 ;
  assign y3491 = ~n7741 ;
  assign y3492 = ~1'b0 ;
  assign y3493 = ~1'b0 ;
  assign y3494 = ~n7745 ;
  assign y3495 = n7746 ;
  assign y3496 = ~n7752 ;
  assign y3497 = ~n7754 ;
  assign y3498 = ~1'b0 ;
  assign y3499 = n7766 ;
  assign y3500 = ~n7768 ;
  assign y3501 = ~1'b0 ;
  assign y3502 = ~1'b0 ;
  assign y3503 = ~n7769 ;
  assign y3504 = ~n7770 ;
  assign y3505 = ~1'b0 ;
  assign y3506 = ~n7772 ;
  assign y3507 = n7776 ;
  assign y3508 = ~1'b0 ;
  assign y3509 = ~1'b0 ;
  assign y3510 = ~n7778 ;
  assign y3511 = n7788 ;
  assign y3512 = ~n7789 ;
  assign y3513 = ~n7796 ;
  assign y3514 = ~1'b0 ;
  assign y3515 = x51 ;
  assign y3516 = ~1'b0 ;
  assign y3517 = n7799 ;
  assign y3518 = ~n7803 ;
  assign y3519 = ~1'b0 ;
  assign y3520 = n7805 ;
  assign y3521 = ~n7809 ;
  assign y3522 = ~n7811 ;
  assign y3523 = ~1'b0 ;
  assign y3524 = n7812 ;
  assign y3525 = ~n7814 ;
  assign y3526 = n7818 ;
  assign y3527 = ~n7821 ;
  assign y3528 = n7826 ;
  assign y3529 = ~n3213 ;
  assign y3530 = ~1'b0 ;
  assign y3531 = n7831 ;
  assign y3532 = ~n7832 ;
  assign y3533 = ~1'b0 ;
  assign y3534 = ~1'b0 ;
  assign y3535 = n2301 ;
  assign y3536 = n7834 ;
  assign y3537 = ~1'b0 ;
  assign y3538 = n7836 ;
  assign y3539 = ~n3704 ;
  assign y3540 = ~n407 ;
  assign y3541 = n7838 ;
  assign y3542 = n7840 ;
  assign y3543 = n7844 ;
  assign y3544 = n7856 ;
  assign y3545 = n7859 ;
  assign y3546 = ~n7861 ;
  assign y3547 = n7866 ;
  assign y3548 = ~n5136 ;
  assign y3549 = ~n7867 ;
  assign y3550 = ~n7869 ;
  assign y3551 = ~n7873 ;
  assign y3552 = n7879 ;
  assign y3553 = ~n7880 ;
  assign y3554 = ~1'b0 ;
  assign y3555 = ~1'b0 ;
  assign y3556 = n7882 ;
  assign y3557 = ~1'b0 ;
  assign y3558 = ~1'b0 ;
  assign y3559 = ~1'b0 ;
  assign y3560 = ~n7886 ;
  assign y3561 = n7887 ;
  assign y3562 = ~n7891 ;
  assign y3563 = n7897 ;
  assign y3564 = ~n7898 ;
  assign y3565 = n7899 ;
  assign y3566 = ~1'b0 ;
  assign y3567 = ~1'b0 ;
  assign y3568 = n7908 ;
  assign y3569 = ~n7911 ;
  assign y3570 = n7916 ;
  assign y3571 = n7917 ;
  assign y3572 = ~n7918 ;
  assign y3573 = ~1'b0 ;
  assign y3574 = ~1'b0 ;
  assign y3575 = ~n7922 ;
  assign y3576 = ~1'b0 ;
  assign y3577 = x182 ;
  assign y3578 = 1'b0 ;
  assign y3579 = ~n2701 ;
  assign y3580 = n7925 ;
  assign y3581 = ~n4001 ;
  assign y3582 = ~1'b0 ;
  assign y3583 = n7927 ;
  assign y3584 = n7930 ;
  assign y3585 = ~1'b0 ;
  assign y3586 = n7933 ;
  assign y3587 = ~1'b0 ;
  assign y3588 = ~n7934 ;
  assign y3589 = ~n7938 ;
  assign y3590 = ~1'b0 ;
  assign y3591 = n7940 ;
  assign y3592 = ~1'b0 ;
  assign y3593 = ~1'b0 ;
  assign y3594 = n7941 ;
  assign y3595 = ~n5580 ;
  assign y3596 = ~n7942 ;
  assign y3597 = ~1'b0 ;
  assign y3598 = ~n7947 ;
  assign y3599 = ~n7948 ;
  assign y3600 = ~n6655 ;
  assign y3601 = n7954 ;
  assign y3602 = n7958 ;
  assign y3603 = n7959 ;
  assign y3604 = ~n7962 ;
  assign y3605 = ~n7964 ;
  assign y3606 = n3416 ;
  assign y3607 = n7969 ;
  assign y3608 = n7971 ;
  assign y3609 = 1'b0 ;
  assign y3610 = ~n7973 ;
  assign y3611 = ~1'b0 ;
  assign y3612 = ~n7974 ;
  assign y3613 = ~1'b0 ;
  assign y3614 = n7975 ;
  assign y3615 = ~n7976 ;
  assign y3616 = ~n7979 ;
  assign y3617 = 1'b0 ;
  assign y3618 = n7987 ;
  assign y3619 = n7989 ;
  assign y3620 = ~1'b0 ;
  assign y3621 = ~1'b0 ;
  assign y3622 = ~n7990 ;
  assign y3623 = n7992 ;
  assign y3624 = n7996 ;
  assign y3625 = ~n7998 ;
  assign y3626 = n8000 ;
  assign y3627 = n8002 ;
  assign y3628 = ~1'b0 ;
  assign y3629 = n8004 ;
  assign y3630 = ~n8005 ;
  assign y3631 = ~1'b0 ;
  assign y3632 = n8008 ;
  assign y3633 = ~1'b0 ;
  assign y3634 = n8009 ;
  assign y3635 = n8020 ;
  assign y3636 = ~n8022 ;
  assign y3637 = n8025 ;
  assign y3638 = n8029 ;
  assign y3639 = n8030 ;
  assign y3640 = ~n8031 ;
  assign y3641 = n8036 ;
  assign y3642 = n8039 ;
  assign y3643 = n8044 ;
  assign y3644 = ~1'b0 ;
  assign y3645 = ~1'b0 ;
  assign y3646 = ~n8046 ;
  assign y3647 = n8048 ;
  assign y3648 = ~n8049 ;
  assign y3649 = n8053 ;
  assign y3650 = n8054 ;
  assign y3651 = n8056 ;
  assign y3652 = ~1'b0 ;
  assign y3653 = n8059 ;
  assign y3654 = ~n8063 ;
  assign y3655 = ~1'b0 ;
  assign y3656 = ~n8068 ;
  assign y3657 = ~1'b0 ;
  assign y3658 = ~n8075 ;
  assign y3659 = n8077 ;
  assign y3660 = n8081 ;
  assign y3661 = ~n8083 ;
  assign y3662 = ~n8084 ;
  assign y3663 = n8096 ;
  assign y3664 = ~n8097 ;
  assign y3665 = ~n2400 ;
  assign y3666 = n8098 ;
  assign y3667 = ~n8101 ;
  assign y3668 = ~n8109 ;
  assign y3669 = ~n8110 ;
  assign y3670 = ~1'b0 ;
  assign y3671 = ~1'b0 ;
  assign y3672 = n8114 ;
  assign y3673 = n8115 ;
  assign y3674 = ~n8129 ;
  assign y3675 = ~n8130 ;
  assign y3676 = ~n8131 ;
  assign y3677 = ~n8133 ;
  assign y3678 = ~1'b0 ;
  assign y3679 = ~n8134 ;
  assign y3680 = n8135 ;
  assign y3681 = ~1'b0 ;
  assign y3682 = n8137 ;
  assign y3683 = ~n8138 ;
  assign y3684 = ~n8147 ;
  assign y3685 = ~n8149 ;
  assign y3686 = n8151 ;
  assign y3687 = n8153 ;
  assign y3688 = n8155 ;
  assign y3689 = n8157 ;
  assign y3690 = ~1'b0 ;
  assign y3691 = ~n8162 ;
  assign y3692 = ~n8164 ;
  assign y3693 = ~n8165 ;
  assign y3694 = ~n8167 ;
  assign y3695 = ~n8180 ;
  assign y3696 = ~n8185 ;
  assign y3697 = ~n8189 ;
  assign y3698 = ~n8191 ;
  assign y3699 = n8194 ;
  assign y3700 = ~n8196 ;
  assign y3701 = ~n8197 ;
  assign y3702 = n8198 ;
  assign y3703 = ~1'b0 ;
  assign y3704 = n8202 ;
  assign y3705 = ~n8205 ;
  assign y3706 = ~1'b0 ;
  assign y3707 = ~n8207 ;
  assign y3708 = n8210 ;
  assign y3709 = ~n8211 ;
  assign y3710 = ~1'b0 ;
  assign y3711 = ~1'b0 ;
  assign y3712 = ~n8217 ;
  assign y3713 = ~n8219 ;
  assign y3714 = ~1'b0 ;
  assign y3715 = n8228 ;
  assign y3716 = ~1'b0 ;
  assign y3717 = n8230 ;
  assign y3718 = ~n8233 ;
  assign y3719 = n8235 ;
  assign y3720 = ~n8237 ;
  assign y3721 = ~n8239 ;
  assign y3722 = ~1'b0 ;
  assign y3723 = n8242 ;
  assign y3724 = ~1'b0 ;
  assign y3725 = ~n1718 ;
  assign y3726 = n3496 ;
  assign y3727 = ~n8244 ;
  assign y3728 = ~1'b0 ;
  assign y3729 = ~n8248 ;
  assign y3730 = ~n8250 ;
  assign y3731 = 1'b0 ;
  assign y3732 = 1'b0 ;
  assign y3733 = ~1'b0 ;
  assign y3734 = ~1'b0 ;
  assign y3735 = ~1'b0 ;
  assign y3736 = ~n8251 ;
  assign y3737 = ~n8253 ;
  assign y3738 = ~1'b0 ;
  assign y3739 = ~1'b0 ;
  assign y3740 = ~1'b0 ;
  assign y3741 = ~1'b0 ;
  assign y3742 = n8260 ;
  assign y3743 = ~n8262 ;
  assign y3744 = ~1'b0 ;
  assign y3745 = n8264 ;
  assign y3746 = n8265 ;
  assign y3747 = ~n8267 ;
  assign y3748 = ~n8273 ;
  assign y3749 = n4315 ;
  assign y3750 = ~1'b0 ;
  assign y3751 = ~n8276 ;
  assign y3752 = ~1'b0 ;
  assign y3753 = n8277 ;
  assign y3754 = n8278 ;
  assign y3755 = n8279 ;
  assign y3756 = ~1'b0 ;
  assign y3757 = n8281 ;
  assign y3758 = ~1'b0 ;
  assign y3759 = n8286 ;
  assign y3760 = n8287 ;
  assign y3761 = ~n8289 ;
  assign y3762 = n1387 ;
  assign y3763 = n8291 ;
  assign y3764 = ~1'b0 ;
  assign y3765 = ~n8298 ;
  assign y3766 = n8302 ;
  assign y3767 = ~n8303 ;
  assign y3768 = n8308 ;
  assign y3769 = ~n8311 ;
  assign y3770 = ~1'b0 ;
  assign y3771 = ~n8312 ;
  assign y3772 = ~n8317 ;
  assign y3773 = ~n2282 ;
  assign y3774 = ~n8323 ;
  assign y3775 = ~n8325 ;
  assign y3776 = ~1'b0 ;
  assign y3777 = ~n8327 ;
  assign y3778 = ~1'b0 ;
  assign y3779 = ~1'b0 ;
  assign y3780 = 1'b0 ;
  assign y3781 = n8328 ;
  assign y3782 = n8330 ;
  assign y3783 = n8333 ;
  assign y3784 = ~1'b0 ;
  assign y3785 = ~1'b0 ;
  assign y3786 = n8340 ;
  assign y3787 = ~n3266 ;
  assign y3788 = ~n3744 ;
  assign y3789 = ~n8342 ;
  assign y3790 = ~1'b0 ;
  assign y3791 = ~1'b0 ;
  assign y3792 = n8346 ;
  assign y3793 = n8351 ;
  assign y3794 = ~1'b0 ;
  assign y3795 = n8354 ;
  assign y3796 = ~1'b0 ;
  assign y3797 = n8359 ;
  assign y3798 = 1'b0 ;
  assign y3799 = ~1'b0 ;
  assign y3800 = ~1'b0 ;
  assign y3801 = n8368 ;
  assign y3802 = ~n8369 ;
  assign y3803 = ~1'b0 ;
  assign y3804 = n8373 ;
  assign y3805 = ~n3590 ;
  assign y3806 = ~n8381 ;
  assign y3807 = ~1'b0 ;
  assign y3808 = ~n8384 ;
  assign y3809 = ~n8393 ;
  assign y3810 = ~1'b0 ;
  assign y3811 = ~n8397 ;
  assign y3812 = ~n8399 ;
  assign y3813 = ~n8403 ;
  assign y3814 = ~n8408 ;
  assign y3815 = ~n8411 ;
  assign y3816 = ~1'b0 ;
  assign y3817 = ~1'b0 ;
  assign y3818 = n5091 ;
  assign y3819 = ~n8413 ;
  assign y3820 = ~n8414 ;
  assign y3821 = ~n8415 ;
  assign y3822 = ~1'b0 ;
  assign y3823 = ~n8419 ;
  assign y3824 = n8421 ;
  assign y3825 = ~1'b0 ;
  assign y3826 = ~n8422 ;
  assign y3827 = ~n8423 ;
  assign y3828 = ~1'b0 ;
  assign y3829 = ~1'b0 ;
  assign y3830 = 1'b0 ;
  assign y3831 = ~n8426 ;
  assign y3832 = n8428 ;
  assign y3833 = ~n8430 ;
  assign y3834 = ~1'b0 ;
  assign y3835 = n8431 ;
  assign y3836 = ~n8434 ;
  assign y3837 = ~n8435 ;
  assign y3838 = n8438 ;
  assign y3839 = ~n8444 ;
  assign y3840 = ~1'b0 ;
  assign y3841 = ~n8450 ;
  assign y3842 = ~n8452 ;
  assign y3843 = n6633 ;
  assign y3844 = ~1'b0 ;
  assign y3845 = ~1'b0 ;
  assign y3846 = n8456 ;
  assign y3847 = ~1'b0 ;
  assign y3848 = ~n8459 ;
  assign y3849 = ~n8460 ;
  assign y3850 = n8462 ;
  assign y3851 = ~1'b0 ;
  assign y3852 = ~n8468 ;
  assign y3853 = n8475 ;
  assign y3854 = ~n8479 ;
  assign y3855 = n8481 ;
  assign y3856 = n8482 ;
  assign y3857 = n8483 ;
  assign y3858 = 1'b0 ;
  assign y3859 = ~n8485 ;
  assign y3860 = n8488 ;
  assign y3861 = ~n8489 ;
  assign y3862 = n8490 ;
  assign y3863 = ~n8491 ;
  assign y3864 = n8493 ;
  assign y3865 = ~1'b0 ;
  assign y3866 = ~n8498 ;
  assign y3867 = ~1'b0 ;
  assign y3868 = ~n8502 ;
  assign y3869 = ~1'b0 ;
  assign y3870 = ~1'b0 ;
  assign y3871 = ~1'b0 ;
  assign y3872 = ~n8503 ;
  assign y3873 = ~n8504 ;
  assign y3874 = ~n8506 ;
  assign y3875 = ~n3386 ;
  assign y3876 = ~n1138 ;
  assign y3877 = ~n8510 ;
  assign y3878 = ~1'b0 ;
  assign y3879 = 1'b0 ;
  assign y3880 = n8514 ;
  assign y3881 = ~n8515 ;
  assign y3882 = ~n8517 ;
  assign y3883 = ~1'b0 ;
  assign y3884 = ~1'b0 ;
  assign y3885 = ~n8519 ;
  assign y3886 = ~n8520 ;
  assign y3887 = n8524 ;
  assign y3888 = ~n8527 ;
  assign y3889 = ~n8530 ;
  assign y3890 = n8532 ;
  assign y3891 = ~1'b0 ;
  assign y3892 = ~1'b0 ;
  assign y3893 = n8535 ;
  assign y3894 = ~1'b0 ;
  assign y3895 = n8540 ;
  assign y3896 = n8543 ;
  assign y3897 = n8545 ;
  assign y3898 = ~n8546 ;
  assign y3899 = ~1'b0 ;
  assign y3900 = 1'b0 ;
  assign y3901 = ~1'b0 ;
  assign y3902 = ~n4638 ;
  assign y3903 = n8547 ;
  assign y3904 = ~n8550 ;
  assign y3905 = n8553 ;
  assign y3906 = ~1'b0 ;
  assign y3907 = ~n8556 ;
  assign y3908 = n8557 ;
  assign y3909 = ~1'b0 ;
  assign y3910 = n8558 ;
  assign y3911 = ~1'b0 ;
  assign y3912 = ~1'b0 ;
  assign y3913 = ~1'b0 ;
  assign y3914 = n8559 ;
  assign y3915 = ~n8561 ;
  assign y3916 = ~n4430 ;
  assign y3917 = n8565 ;
  assign y3918 = n8570 ;
  assign y3919 = n8573 ;
  assign y3920 = n8574 ;
  assign y3921 = n8582 ;
  assign y3922 = ~n8584 ;
  assign y3923 = n8585 ;
  assign y3924 = ~n8597 ;
  assign y3925 = ~n8602 ;
  assign y3926 = ~1'b0 ;
  assign y3927 = n8604 ;
  assign y3928 = ~1'b0 ;
  assign y3929 = ~n8605 ;
  assign y3930 = ~n6619 ;
  assign y3931 = ~1'b0 ;
  assign y3932 = n8606 ;
  assign y3933 = ~n8609 ;
  assign y3934 = ~n8610 ;
  assign y3935 = n8613 ;
  assign y3936 = ~n8614 ;
  assign y3937 = ~n8616 ;
  assign y3938 = ~n8618 ;
  assign y3939 = n8622 ;
  assign y3940 = ~1'b0 ;
  assign y3941 = ~n8624 ;
  assign y3942 = ~1'b0 ;
  assign y3943 = ~n8625 ;
  assign y3944 = n8626 ;
  assign y3945 = n8629 ;
  assign y3946 = n8639 ;
  assign y3947 = ~1'b0 ;
  assign y3948 = ~n8641 ;
  assign y3949 = ~1'b0 ;
  assign y3950 = ~n8646 ;
  assign y3951 = ~n8647 ;
  assign y3952 = ~1'b0 ;
  assign y3953 = ~n8651 ;
  assign y3954 = ~1'b0 ;
  assign y3955 = ~n8653 ;
  assign y3956 = ~n8657 ;
  assign y3957 = ~n8658 ;
  assign y3958 = n8659 ;
  assign y3959 = ~1'b0 ;
  assign y3960 = n8663 ;
  assign y3961 = ~1'b0 ;
  assign y3962 = n8664 ;
  assign y3963 = n2569 ;
  assign y3964 = ~n8670 ;
  assign y3965 = ~1'b0 ;
  assign y3966 = ~n8673 ;
  assign y3967 = ~1'b0 ;
  assign y3968 = n8677 ;
  assign y3969 = n8678 ;
  assign y3970 = n8679 ;
  assign y3971 = n8681 ;
  assign y3972 = ~1'b0 ;
  assign y3973 = ~1'b0 ;
  assign y3974 = ~1'b0 ;
  assign y3975 = n8683 ;
  assign y3976 = ~1'b0 ;
  assign y3977 = ~1'b0 ;
  assign y3978 = ~1'b0 ;
  assign y3979 = n8687 ;
  assign y3980 = n378 ;
  assign y3981 = n8691 ;
  assign y3982 = ~n1557 ;
  assign y3983 = ~n6429 ;
  assign y3984 = ~n8693 ;
  assign y3985 = ~n8694 ;
  assign y3986 = ~n8695 ;
  assign y3987 = ~n8698 ;
  assign y3988 = ~n8700 ;
  assign y3989 = n8702 ;
  assign y3990 = ~1'b0 ;
  assign y3991 = n8710 ;
  assign y3992 = n8720 ;
  assign y3993 = ~n8722 ;
  assign y3994 = n8723 ;
  assign y3995 = ~n8724 ;
  assign y3996 = n8726 ;
  assign y3997 = n8729 ;
  assign y3998 = ~1'b0 ;
  assign y3999 = ~n8731 ;
  assign y4000 = n8735 ;
  assign y4001 = ~1'b0 ;
  assign y4002 = ~n8739 ;
  assign y4003 = ~1'b0 ;
  assign y4004 = n8740 ;
  assign y4005 = ~1'b0 ;
  assign y4006 = n8742 ;
  assign y4007 = n8745 ;
  assign y4008 = ~n8749 ;
  assign y4009 = ~1'b0 ;
  assign y4010 = n8754 ;
  assign y4011 = ~1'b0 ;
  assign y4012 = ~1'b0 ;
  assign y4013 = n8755 ;
  assign y4014 = ~1'b0 ;
  assign y4015 = n8756 ;
  assign y4016 = ~1'b0 ;
  assign y4017 = ~1'b0 ;
  assign y4018 = ~n2799 ;
  assign y4019 = n8764 ;
  assign y4020 = n8766 ;
  assign y4021 = ~n8770 ;
  assign y4022 = ~n8772 ;
  assign y4023 = n8774 ;
  assign y4024 = n8777 ;
  assign y4025 = ~n8778 ;
  assign y4026 = ~1'b0 ;
  assign y4027 = n8780 ;
  assign y4028 = ~1'b0 ;
  assign y4029 = ~1'b0 ;
  assign y4030 = n8788 ;
  assign y4031 = ~n8789 ;
  assign y4032 = n8794 ;
  assign y4033 = ~1'b0 ;
  assign y4034 = n8796 ;
  assign y4035 = ~1'b0 ;
  assign y4036 = ~n3686 ;
  assign y4037 = ~1'b0 ;
  assign y4038 = ~1'b0 ;
  assign y4039 = ~n8798 ;
  assign y4040 = ~1'b0 ;
  assign y4041 = ~1'b0 ;
  assign y4042 = ~1'b0 ;
  assign y4043 = n8799 ;
  assign y4044 = ~1'b0 ;
  assign y4045 = ~n8802 ;
  assign y4046 = ~1'b0 ;
  assign y4047 = ~n8806 ;
  assign y4048 = ~1'b0 ;
  assign y4049 = n8807 ;
  assign y4050 = n8811 ;
  assign y4051 = 1'b0 ;
  assign y4052 = ~1'b0 ;
  assign y4053 = n8814 ;
  assign y4054 = ~1'b0 ;
  assign y4055 = n8816 ;
  assign y4056 = ~1'b0 ;
  assign y4057 = ~1'b0 ;
  assign y4058 = ~n8820 ;
  assign y4059 = n8825 ;
  assign y4060 = ~1'b0 ;
  assign y4061 = ~n8829 ;
  assign y4062 = ~1'b0 ;
  assign y4063 = ~n8830 ;
  assign y4064 = ~1'b0 ;
  assign y4065 = ~1'b0 ;
  assign y4066 = x96 ;
  assign y4067 = ~n8834 ;
  assign y4068 = n8837 ;
  assign y4069 = ~1'b0 ;
  assign y4070 = n8839 ;
  assign y4071 = ~1'b0 ;
  assign y4072 = ~n8841 ;
  assign y4073 = n5317 ;
  assign y4074 = n8849 ;
  assign y4075 = ~1'b0 ;
  assign y4076 = n8851 ;
  assign y4077 = n8857 ;
  assign y4078 = n8860 ;
  assign y4079 = n8862 ;
  assign y4080 = ~n8864 ;
  assign y4081 = ~n300 ;
  assign y4082 = n8865 ;
  assign y4083 = ~1'b0 ;
  assign y4084 = ~1'b0 ;
  assign y4085 = n8866 ;
  assign y4086 = ~1'b0 ;
  assign y4087 = n8868 ;
  assign y4088 = n8878 ;
  assign y4089 = ~n8883 ;
  assign y4090 = ~1'b0 ;
  assign y4091 = n8885 ;
  assign y4092 = ~1'b0 ;
  assign y4093 = ~1'b0 ;
  assign y4094 = n8889 ;
  assign y4095 = ~1'b0 ;
  assign y4096 = n8891 ;
  assign y4097 = n5461 ;
  assign y4098 = ~n8892 ;
  assign y4099 = n8895 ;
  assign y4100 = 1'b0 ;
  assign y4101 = ~n8899 ;
  assign y4102 = n8904 ;
  assign y4103 = ~1'b0 ;
  assign y4104 = ~1'b0 ;
  assign y4105 = ~1'b0 ;
  assign y4106 = ~1'b0 ;
  assign y4107 = ~1'b0 ;
  assign y4108 = n708 ;
  assign y4109 = 1'b0 ;
  assign y4110 = ~n8905 ;
  assign y4111 = ~1'b0 ;
  assign y4112 = ~n8907 ;
  assign y4113 = ~n8909 ;
  assign y4114 = ~n8914 ;
  assign y4115 = ~1'b0 ;
  assign y4116 = n8916 ;
  assign y4117 = ~1'b0 ;
  assign y4118 = n8919 ;
  assign y4119 = ~n4325 ;
  assign y4120 = ~n8923 ;
  assign y4121 = n8926 ;
  assign y4122 = ~n8928 ;
  assign y4123 = n8940 ;
  assign y4124 = ~n8941 ;
  assign y4125 = ~n8943 ;
  assign y4126 = n8945 ;
  assign y4127 = ~n8948 ;
  assign y4128 = n8950 ;
  assign y4129 = ~n8951 ;
  assign y4130 = ~n8954 ;
  assign y4131 = ~1'b0 ;
  assign y4132 = ~1'b0 ;
  assign y4133 = n8959 ;
  assign y4134 = ~n8963 ;
  assign y4135 = ~n8966 ;
  assign y4136 = n8969 ;
  assign y4137 = n8971 ;
  assign y4138 = 1'b0 ;
  assign y4139 = ~n8973 ;
  assign y4140 = n8981 ;
  assign y4141 = n8984 ;
  assign y4142 = n8990 ;
  assign y4143 = n8998 ;
  assign y4144 = n9007 ;
  assign y4145 = n9009 ;
  assign y4146 = ~n9017 ;
  assign y4147 = n9019 ;
  assign y4148 = n9021 ;
  assign y4149 = n9024 ;
  assign y4150 = ~1'b0 ;
  assign y4151 = ~1'b0 ;
  assign y4152 = ~1'b0 ;
  assign y4153 = n9027 ;
  assign y4154 = ~1'b0 ;
  assign y4155 = ~n9031 ;
  assign y4156 = n9038 ;
  assign y4157 = ~n9045 ;
  assign y4158 = ~n9046 ;
  assign y4159 = ~n9053 ;
  assign y4160 = ~1'b0 ;
  assign y4161 = n9057 ;
  assign y4162 = ~1'b0 ;
  assign y4163 = n9059 ;
  assign y4164 = ~1'b0 ;
  assign y4165 = n9060 ;
  assign y4166 = n3474 ;
  assign y4167 = ~1'b0 ;
  assign y4168 = ~1'b0 ;
  assign y4169 = ~1'b0 ;
  assign y4170 = ~n9062 ;
  assign y4171 = ~1'b0 ;
  assign y4172 = ~n9064 ;
  assign y4173 = ~n9065 ;
  assign y4174 = n9075 ;
  assign y4175 = n9088 ;
  assign y4176 = ~n9096 ;
  assign y4177 = ~1'b0 ;
  assign y4178 = ~n9098 ;
  assign y4179 = ~1'b0 ;
  assign y4180 = ~n635 ;
  assign y4181 = ~n9104 ;
  assign y4182 = ~n9107 ;
  assign y4183 = ~n9109 ;
  assign y4184 = ~n9115 ;
  assign y4185 = 1'b0 ;
  assign y4186 = ~1'b0 ;
  assign y4187 = ~1'b0 ;
  assign y4188 = n9119 ;
  assign y4189 = ~n9130 ;
  assign y4190 = ~n9138 ;
  assign y4191 = n9142 ;
  assign y4192 = ~n9149 ;
  assign y4193 = ~n9151 ;
  assign y4194 = ~n9159 ;
  assign y4195 = ~1'b0 ;
  assign y4196 = ~1'b0 ;
  assign y4197 = ~n9162 ;
  assign y4198 = n9171 ;
  assign y4199 = n9179 ;
  assign y4200 = ~n9180 ;
  assign y4201 = ~n9181 ;
  assign y4202 = ~n9183 ;
  assign y4203 = ~1'b0 ;
  assign y4204 = ~n1828 ;
  assign y4205 = ~n9186 ;
  assign y4206 = ~n9190 ;
  assign y4207 = ~1'b0 ;
  assign y4208 = 1'b0 ;
  assign y4209 = n9192 ;
  assign y4210 = ~1'b0 ;
  assign y4211 = n3265 ;
  assign y4212 = n9193 ;
  assign y4213 = n9198 ;
  assign y4214 = n9202 ;
  assign y4215 = n9206 ;
  assign y4216 = ~n9210 ;
  assign y4217 = ~n9211 ;
  assign y4218 = n9215 ;
  assign y4219 = n9219 ;
  assign y4220 = ~1'b0 ;
  assign y4221 = n9223 ;
  assign y4222 = n9225 ;
  assign y4223 = ~1'b0 ;
  assign y4224 = n9226 ;
  assign y4225 = n6433 ;
  assign y4226 = ~n9228 ;
  assign y4227 = ~1'b0 ;
  assign y4228 = n9230 ;
  assign y4229 = ~1'b0 ;
  assign y4230 = n9232 ;
  assign y4231 = n9236 ;
  assign y4232 = ~n9237 ;
  assign y4233 = ~n9239 ;
  assign y4234 = ~1'b0 ;
  assign y4235 = n9241 ;
  assign y4236 = n9246 ;
  assign y4237 = ~1'b0 ;
  assign y4238 = ~n9248 ;
  assign y4239 = n9250 ;
  assign y4240 = ~n9252 ;
  assign y4241 = ~n9255 ;
  assign y4242 = ~1'b0 ;
  assign y4243 = n9256 ;
  assign y4244 = ~n9258 ;
  assign y4245 = n9259 ;
  assign y4246 = ~1'b0 ;
  assign y4247 = ~n9263 ;
  assign y4248 = ~n9276 ;
  assign y4249 = n9283 ;
  assign y4250 = 1'b0 ;
  assign y4251 = ~1'b0 ;
  assign y4252 = ~n9287 ;
  assign y4253 = ~1'b0 ;
  assign y4254 = ~1'b0 ;
  assign y4255 = 1'b0 ;
  assign y4256 = ~n8678 ;
  assign y4257 = n9288 ;
  assign y4258 = n9289 ;
  assign y4259 = ~1'b0 ;
  assign y4260 = ~n9293 ;
  assign y4261 = ~1'b0 ;
  assign y4262 = n9294 ;
  assign y4263 = ~n9295 ;
  assign y4264 = n9299 ;
  assign y4265 = 1'b0 ;
  assign y4266 = n9302 ;
  assign y4267 = n9304 ;
  assign y4268 = n9307 ;
  assign y4269 = n9314 ;
  assign y4270 = ~1'b0 ;
  assign y4271 = ~n9319 ;
  assign y4272 = ~n9321 ;
  assign y4273 = ~n9325 ;
  assign y4274 = ~1'b0 ;
  assign y4275 = n9327 ;
  assign y4276 = n9335 ;
  assign y4277 = ~n9343 ;
  assign y4278 = ~1'b0 ;
  assign y4279 = ~n9345 ;
  assign y4280 = n9353 ;
  assign y4281 = ~1'b0 ;
  assign y4282 = ~1'b0 ;
  assign y4283 = ~n7383 ;
  assign y4284 = ~1'b0 ;
  assign y4285 = ~1'b0 ;
  assign y4286 = n772 ;
  assign y4287 = ~n9354 ;
  assign y4288 = ~1'b0 ;
  assign y4289 = ~n9355 ;
  assign y4290 = ~1'b0 ;
  assign y4291 = ~n9360 ;
  assign y4292 = n9367 ;
  assign y4293 = ~n9370 ;
  assign y4294 = ~n9378 ;
  assign y4295 = n9382 ;
  assign y4296 = ~n9386 ;
  assign y4297 = n6616 ;
  assign y4298 = ~1'b0 ;
  assign y4299 = n9388 ;
  assign y4300 = ~1'b0 ;
  assign y4301 = n9391 ;
  assign y4302 = ~1'b0 ;
  assign y4303 = 1'b0 ;
  assign y4304 = ~n9398 ;
  assign y4305 = n9400 ;
  assign y4306 = ~n4546 ;
  assign y4307 = n9401 ;
  assign y4308 = ~1'b0 ;
  assign y4309 = ~n9406 ;
  assign y4310 = n9408 ;
  assign y4311 = ~n9413 ;
  assign y4312 = n9416 ;
  assign y4313 = ~1'b0 ;
  assign y4314 = ~1'b0 ;
  assign y4315 = n9418 ;
  assign y4316 = n9419 ;
  assign y4317 = ~1'b0 ;
  assign y4318 = ~1'b0 ;
  assign y4319 = ~n9072 ;
  assign y4320 = n9420 ;
  assign y4321 = n9422 ;
  assign y4322 = ~n9423 ;
  assign y4323 = ~n9432 ;
  assign y4324 = ~n8578 ;
  assign y4325 = ~1'b0 ;
  assign y4326 = n9433 ;
  assign y4327 = ~1'b0 ;
  assign y4328 = ~n9434 ;
  assign y4329 = n9444 ;
  assign y4330 = n9446 ;
  assign y4331 = ~n9447 ;
  assign y4332 = ~n9448 ;
  assign y4333 = ~n9452 ;
  assign y4334 = ~n9454 ;
  assign y4335 = n9459 ;
  assign y4336 = ~n9463 ;
  assign y4337 = n9465 ;
  assign y4338 = n9466 ;
  assign y4339 = ~n9468 ;
  assign y4340 = n9473 ;
  assign y4341 = 1'b0 ;
  assign y4342 = n9477 ;
  assign y4343 = ~n9481 ;
  assign y4344 = n9483 ;
  assign y4345 = ~n9486 ;
  assign y4346 = n9489 ;
  assign y4347 = ~1'b0 ;
  assign y4348 = n9493 ;
  assign y4349 = ~1'b0 ;
  assign y4350 = ~n9495 ;
  assign y4351 = ~n9496 ;
  assign y4352 = ~n9502 ;
  assign y4353 = ~n9505 ;
  assign y4354 = n9510 ;
  assign y4355 = ~1'b0 ;
  assign y4356 = n9512 ;
  assign y4357 = ~1'b0 ;
  assign y4358 = n9513 ;
  assign y4359 = ~n9514 ;
  assign y4360 = n9518 ;
  assign y4361 = ~n9521 ;
  assign y4362 = n9522 ;
  assign y4363 = n9523 ;
  assign y4364 = ~1'b0 ;
  assign y4365 = n9525 ;
  assign y4366 = ~n8622 ;
  assign y4367 = n9527 ;
  assign y4368 = ~n9531 ;
  assign y4369 = n9532 ;
  assign y4370 = ~n9534 ;
  assign y4371 = n9538 ;
  assign y4372 = ~n9539 ;
  assign y4373 = n9540 ;
  assign y4374 = ~1'b0 ;
  assign y4375 = n6731 ;
  assign y4376 = ~1'b0 ;
  assign y4377 = ~n9544 ;
  assign y4378 = ~n9546 ;
  assign y4379 = ~1'b0 ;
  assign y4380 = ~n9554 ;
  assign y4381 = ~n9556 ;
  assign y4382 = ~n9566 ;
  assign y4383 = n9571 ;
  assign y4384 = n9572 ;
  assign y4385 = ~1'b0 ;
  assign y4386 = n9576 ;
  assign y4387 = n9577 ;
  assign y4388 = ~1'b0 ;
  assign y4389 = n9580 ;
  assign y4390 = n9584 ;
  assign y4391 = n9587 ;
  assign y4392 = n9590 ;
  assign y4393 = ~1'b0 ;
  assign y4394 = ~1'b0 ;
  assign y4395 = ~1'b0 ;
  assign y4396 = ~1'b0 ;
  assign y4397 = n3019 ;
  assign y4398 = 1'b0 ;
  assign y4399 = ~n9595 ;
  assign y4400 = ~n9599 ;
  assign y4401 = n9600 ;
  assign y4402 = ~n9607 ;
  assign y4403 = n7677 ;
  assign y4404 = ~n9608 ;
  assign y4405 = ~1'b0 ;
  assign y4406 = n9618 ;
  assign y4407 = ~n9620 ;
  assign y4408 = n9623 ;
  assign y4409 = ~1'b0 ;
  assign y4410 = ~n9624 ;
  assign y4411 = n9625 ;
  assign y4412 = ~1'b0 ;
  assign y4413 = n9628 ;
  assign y4414 = ~n9634 ;
  assign y4415 = ~1'b0 ;
  assign y4416 = n9636 ;
  assign y4417 = n8114 ;
  assign y4418 = n9640 ;
  assign y4419 = n9641 ;
  assign y4420 = ~1'b0 ;
  assign y4421 = ~1'b0 ;
  assign y4422 = ~1'b0 ;
  assign y4423 = n9643 ;
  assign y4424 = ~1'b0 ;
  assign y4425 = n9646 ;
  assign y4426 = ~n9651 ;
  assign y4427 = ~n9654 ;
  assign y4428 = ~n9657 ;
  assign y4429 = ~n8219 ;
  assign y4430 = ~1'b0 ;
  assign y4431 = n9661 ;
  assign y4432 = ~n9662 ;
  assign y4433 = n9664 ;
  assign y4434 = n9665 ;
  assign y4435 = n9670 ;
  assign y4436 = ~n9674 ;
  assign y4437 = ~n9688 ;
  assign y4438 = n9691 ;
  assign y4439 = ~1'b0 ;
  assign y4440 = n9692 ;
  assign y4441 = ~n9693 ;
  assign y4442 = ~n9694 ;
  assign y4443 = ~n9698 ;
  assign y4444 = n9699 ;
  assign y4445 = ~n9700 ;
  assign y4446 = ~n9702 ;
  assign y4447 = ~1'b0 ;
  assign y4448 = n5685 ;
  assign y4449 = n9703 ;
  assign y4450 = n9704 ;
  assign y4451 = n9705 ;
  assign y4452 = ~1'b0 ;
  assign y4453 = n9709 ;
  assign y4454 = ~1'b0 ;
  assign y4455 = n9711 ;
  assign y4456 = ~1'b0 ;
  assign y4457 = n9717 ;
  assign y4458 = ~1'b0 ;
  assign y4459 = ~1'b0 ;
  assign y4460 = n9724 ;
  assign y4461 = ~1'b0 ;
  assign y4462 = n9728 ;
  assign y4463 = n9729 ;
  assign y4464 = ~1'b0 ;
  assign y4465 = n9730 ;
  assign y4466 = ~1'b0 ;
  assign y4467 = n9736 ;
  assign y4468 = n9738 ;
  assign y4469 = ~n9739 ;
  assign y4470 = n9744 ;
  assign y4471 = n9745 ;
  assign y4472 = ~n9749 ;
  assign y4473 = ~1'b0 ;
  assign y4474 = n9759 ;
  assign y4475 = ~1'b0 ;
  assign y4476 = ~1'b0 ;
  assign y4477 = ~n9761 ;
  assign y4478 = n9764 ;
  assign y4479 = ~1'b0 ;
  assign y4480 = ~n9769 ;
  assign y4481 = n3114 ;
  assign y4482 = ~n9770 ;
  assign y4483 = ~1'b0 ;
  assign y4484 = ~1'b0 ;
  assign y4485 = ~n9774 ;
  assign y4486 = ~n9778 ;
  assign y4487 = ~n9780 ;
  assign y4488 = ~1'b0 ;
  assign y4489 = n9781 ;
  assign y4490 = n9782 ;
  assign y4491 = n9791 ;
  assign y4492 = ~1'b0 ;
  assign y4493 = n9793 ;
  assign y4494 = 1'b0 ;
  assign y4495 = n9794 ;
  assign y4496 = ~n9799 ;
  assign y4497 = n9801 ;
  assign y4498 = ~n9802 ;
  assign y4499 = ~n9808 ;
  assign y4500 = n9815 ;
  assign y4501 = ~1'b0 ;
  assign y4502 = n9819 ;
  assign y4503 = ~n9821 ;
  assign y4504 = ~1'b0 ;
  assign y4505 = ~n9826 ;
  assign y4506 = ~1'b0 ;
  assign y4507 = ~1'b0 ;
  assign y4508 = ~1'b0 ;
  assign y4509 = n9827 ;
  assign y4510 = ~n9828 ;
  assign y4511 = ~1'b0 ;
  assign y4512 = ~n9829 ;
  assign y4513 = ~n9830 ;
  assign y4514 = ~1'b0 ;
  assign y4515 = n9832 ;
  assign y4516 = ~1'b0 ;
  assign y4517 = ~n9835 ;
  assign y4518 = ~n9837 ;
  assign y4519 = n9840 ;
  assign y4520 = ~n1833 ;
  assign y4521 = ~1'b0 ;
  assign y4522 = n9841 ;
  assign y4523 = ~n9847 ;
  assign y4524 = n9848 ;
  assign y4525 = ~n9850 ;
  assign y4526 = ~1'b0 ;
  assign y4527 = ~1'b0 ;
  assign y4528 = n9852 ;
  assign y4529 = 1'b0 ;
  assign y4530 = ~n9855 ;
  assign y4531 = n6780 ;
  assign y4532 = ~1'b0 ;
  assign y4533 = ~1'b0 ;
  assign y4534 = ~1'b0 ;
  assign y4535 = ~1'b0 ;
  assign y4536 = ~n9859 ;
  assign y4537 = ~n9862 ;
  assign y4538 = ~1'b0 ;
  assign y4539 = ~1'b0 ;
  assign y4540 = n9864 ;
  assign y4541 = n9865 ;
  assign y4542 = ~n9867 ;
  assign y4543 = ~1'b0 ;
  assign y4544 = n9872 ;
  assign y4545 = ~1'b0 ;
  assign y4546 = ~n9873 ;
  assign y4547 = n6121 ;
  assign y4548 = ~1'b0 ;
  assign y4549 = n9874 ;
  assign y4550 = n9879 ;
  assign y4551 = ~n9885 ;
  assign y4552 = n9887 ;
  assign y4553 = ~n9889 ;
  assign y4554 = ~n9890 ;
  assign y4555 = ~1'b0 ;
  assign y4556 = ~n9892 ;
  assign y4557 = n9894 ;
  assign y4558 = n9406 ;
  assign y4559 = ~n9900 ;
  assign y4560 = ~n9904 ;
  assign y4561 = ~n8740 ;
  assign y4562 = ~n9906 ;
  assign y4563 = ~1'b0 ;
  assign y4564 = n9909 ;
  assign y4565 = ~n9911 ;
  assign y4566 = ~1'b0 ;
  assign y4567 = n9912 ;
  assign y4568 = ~n9917 ;
  assign y4569 = n9920 ;
  assign y4570 = ~n6510 ;
  assign y4571 = ~n8219 ;
  assign y4572 = n9921 ;
  assign y4573 = ~n9922 ;
  assign y4574 = ~1'b0 ;
  assign y4575 = ~n9924 ;
  assign y4576 = ~n9926 ;
  assign y4577 = ~n9927 ;
  assign y4578 = n9929 ;
  assign y4579 = n9935 ;
  assign y4580 = n9936 ;
  assign y4581 = n9942 ;
  assign y4582 = n9944 ;
  assign y4583 = ~1'b0 ;
  assign y4584 = n9948 ;
  assign y4585 = n9949 ;
  assign y4586 = n9950 ;
  assign y4587 = ~1'b0 ;
  assign y4588 = ~n9953 ;
  assign y4589 = ~n9957 ;
  assign y4590 = ~n9963 ;
  assign y4591 = ~n9965 ;
  assign y4592 = ~1'b0 ;
  assign y4593 = ~1'b0 ;
  assign y4594 = ~n9971 ;
  assign y4595 = ~1'b0 ;
  assign y4596 = n9984 ;
  assign y4597 = ~1'b0 ;
  assign y4598 = n9985 ;
  assign y4599 = ~n9986 ;
  assign y4600 = ~n4003 ;
  assign y4601 = ~n9989 ;
  assign y4602 = n9990 ;
  assign y4603 = ~1'b0 ;
  assign y4604 = ~n9995 ;
  assign y4605 = ~n9998 ;
  assign y4606 = ~1'b0 ;
  assign y4607 = ~1'b0 ;
  assign y4608 = n9999 ;
  assign y4609 = n10001 ;
  assign y4610 = n10003 ;
  assign y4611 = ~n10004 ;
  assign y4612 = ~1'b0 ;
  assign y4613 = ~n8627 ;
  assign y4614 = ~1'b0 ;
  assign y4615 = ~1'b0 ;
  assign y4616 = ~n7351 ;
  assign y4617 = n10009 ;
  assign y4618 = ~n10015 ;
  assign y4619 = ~n10019 ;
  assign y4620 = ~n10026 ;
  assign y4621 = ~1'b0 ;
  assign y4622 = n10028 ;
  assign y4623 = ~n10033 ;
  assign y4624 = ~1'b0 ;
  assign y4625 = ~1'b0 ;
  assign y4626 = ~1'b0 ;
  assign y4627 = n10034 ;
  assign y4628 = n10040 ;
  assign y4629 = ~1'b0 ;
  assign y4630 = 1'b0 ;
  assign y4631 = ~1'b0 ;
  assign y4632 = ~1'b0 ;
  assign y4633 = ~n5368 ;
  assign y4634 = n10044 ;
  assign y4635 = n5309 ;
  assign y4636 = n10047 ;
  assign y4637 = ~n10049 ;
  assign y4638 = n10063 ;
  assign y4639 = n10064 ;
  assign y4640 = ~1'b0 ;
  assign y4641 = ~n10065 ;
  assign y4642 = n10066 ;
  assign y4643 = ~1'b0 ;
  assign y4644 = n10070 ;
  assign y4645 = ~n10075 ;
  assign y4646 = ~n10081 ;
  assign y4647 = ~n10084 ;
  assign y4648 = ~1'b0 ;
  assign y4649 = ~n10086 ;
  assign y4650 = n10088 ;
  assign y4651 = ~n10094 ;
  assign y4652 = ~1'b0 ;
  assign y4653 = ~n10095 ;
  assign y4654 = n10096 ;
  assign y4655 = ~n10099 ;
  assign y4656 = ~n10100 ;
  assign y4657 = ~n10101 ;
  assign y4658 = ~1'b0 ;
  assign y4659 = ~1'b0 ;
  assign y4660 = ~1'b0 ;
  assign y4661 = n10102 ;
  assign y4662 = ~1'b0 ;
  assign y4663 = ~1'b0 ;
  assign y4664 = ~n10105 ;
  assign y4665 = ~n10106 ;
  assign y4666 = ~1'b0 ;
  assign y4667 = n10111 ;
  assign y4668 = n10113 ;
  assign y4669 = n10114 ;
  assign y4670 = ~n10122 ;
  assign y4671 = ~n10124 ;
  assign y4672 = ~1'b0 ;
  assign y4673 = n10127 ;
  assign y4674 = ~1'b0 ;
  assign y4675 = ~1'b0 ;
  assign y4676 = 1'b0 ;
  assign y4677 = ~1'b0 ;
  assign y4678 = ~n10129 ;
  assign y4679 = n10133 ;
  assign y4680 = ~n10135 ;
  assign y4681 = ~n10137 ;
  assign y4682 = ~n10143 ;
  assign y4683 = n10147 ;
  assign y4684 = n10167 ;
  assign y4685 = ~n10169 ;
  assign y4686 = ~1'b0 ;
  assign y4687 = n6506 ;
  assign y4688 = ~n2735 ;
  assign y4689 = ~1'b0 ;
  assign y4690 = ~1'b0 ;
  assign y4691 = n10175 ;
  assign y4692 = ~n10177 ;
  assign y4693 = n10178 ;
  assign y4694 = ~n10179 ;
  assign y4695 = ~n10180 ;
  assign y4696 = ~n9679 ;
  assign y4697 = n1820 ;
  assign y4698 = ~n6097 ;
  assign y4699 = n10190 ;
  assign y4700 = ~n10194 ;
  assign y4701 = ~n10205 ;
  assign y4702 = n10207 ;
  assign y4703 = ~n10209 ;
  assign y4704 = n10218 ;
  assign y4705 = ~n10221 ;
  assign y4706 = ~n10223 ;
  assign y4707 = n10232 ;
  assign y4708 = ~n10237 ;
  assign y4709 = ~n6817 ;
  assign y4710 = ~n9456 ;
  assign y4711 = n10240 ;
  assign y4712 = ~1'b0 ;
  assign y4713 = ~1'b0 ;
  assign y4714 = ~1'b0 ;
  assign y4715 = ~1'b0 ;
  assign y4716 = ~n10243 ;
  assign y4717 = ~n10096 ;
  assign y4718 = n5221 ;
  assign y4719 = ~1'b0 ;
  assign y4720 = ~n10248 ;
  assign y4721 = n10253 ;
  assign y4722 = n10254 ;
  assign y4723 = ~n10256 ;
  assign y4724 = 1'b0 ;
  assign y4725 = n10258 ;
  assign y4726 = n10259 ;
  assign y4727 = ~n10262 ;
  assign y4728 = ~1'b0 ;
  assign y4729 = ~n10267 ;
  assign y4730 = ~n10272 ;
  assign y4731 = n10275 ;
  assign y4732 = ~1'b0 ;
  assign y4733 = ~1'b0 ;
  assign y4734 = n10277 ;
  assign y4735 = n10279 ;
  assign y4736 = ~1'b0 ;
  assign y4737 = ~1'b0 ;
  assign y4738 = ~n10292 ;
  assign y4739 = n10294 ;
  assign y4740 = n10295 ;
  assign y4741 = n10296 ;
  assign y4742 = n10297 ;
  assign y4743 = ~1'b0 ;
  assign y4744 = ~1'b0 ;
  assign y4745 = ~n10298 ;
  assign y4746 = n10299 ;
  assign y4747 = n10305 ;
  assign y4748 = ~n10307 ;
  assign y4749 = n10308 ;
  assign y4750 = n10309 ;
  assign y4751 = n10312 ;
  assign y4752 = n10313 ;
  assign y4753 = ~1'b0 ;
  assign y4754 = ~n10315 ;
  assign y4755 = ~1'b0 ;
  assign y4756 = ~1'b0 ;
  assign y4757 = ~n10317 ;
  assign y4758 = ~n10318 ;
  assign y4759 = ~1'b0 ;
  assign y4760 = ~n10320 ;
  assign y4761 = ~n10324 ;
  assign y4762 = n10329 ;
  assign y4763 = ~1'b0 ;
  assign y4764 = ~n10331 ;
  assign y4765 = ~n10335 ;
  assign y4766 = ~1'b0 ;
  assign y4767 = n10336 ;
  assign y4768 = n10337 ;
  assign y4769 = 1'b0 ;
  assign y4770 = n10340 ;
  assign y4771 = n10342 ;
  assign y4772 = ~1'b0 ;
  assign y4773 = ~n5619 ;
  assign y4774 = ~n10343 ;
  assign y4775 = n10345 ;
  assign y4776 = n10351 ;
  assign y4777 = n10352 ;
  assign y4778 = n10353 ;
  assign y4779 = n10360 ;
  assign y4780 = ~1'b0 ;
  assign y4781 = n10363 ;
  assign y4782 = n10365 ;
  assign y4783 = n10367 ;
  assign y4784 = ~1'b0 ;
  assign y4785 = ~1'b0 ;
  assign y4786 = n10369 ;
  assign y4787 = ~n10371 ;
  assign y4788 = 1'b0 ;
  assign y4789 = n10373 ;
  assign y4790 = n10376 ;
  assign y4791 = n10378 ;
  assign y4792 = n10381 ;
  assign y4793 = ~n10383 ;
  assign y4794 = ~n10387 ;
  assign y4795 = n7181 ;
  assign y4796 = n10390 ;
  assign y4797 = n10397 ;
  assign y4798 = ~n10401 ;
  assign y4799 = x64 ;
  assign y4800 = ~n10410 ;
  assign y4801 = ~1'b0 ;
  assign y4802 = ~n810 ;
  assign y4803 = ~1'b0 ;
  assign y4804 = ~1'b0 ;
  assign y4805 = ~1'b0 ;
  assign y4806 = n8322 ;
  assign y4807 = n10412 ;
  assign y4808 = ~n10414 ;
  assign y4809 = ~n765 ;
  assign y4810 = ~1'b0 ;
  assign y4811 = ~1'b0 ;
  assign y4812 = ~n10418 ;
  assign y4813 = ~n10419 ;
  assign y4814 = ~1'b0 ;
  assign y4815 = ~n10425 ;
  assign y4816 = n10426 ;
  assign y4817 = ~n10429 ;
  assign y4818 = n10431 ;
  assign y4819 = ~n10433 ;
  assign y4820 = n10437 ;
  assign y4821 = n10441 ;
  assign y4822 = n10449 ;
  assign y4823 = ~n10451 ;
  assign y4824 = n10469 ;
  assign y4825 = ~1'b0 ;
  assign y4826 = n8963 ;
  assign y4827 = ~1'b0 ;
  assign y4828 = n10471 ;
  assign y4829 = n10472 ;
  assign y4830 = ~1'b0 ;
  assign y4831 = ~1'b0 ;
  assign y4832 = ~n10476 ;
  assign y4833 = ~n10483 ;
  assign y4834 = ~n10484 ;
  assign y4835 = ~1'b0 ;
  assign y4836 = ~1'b0 ;
  assign y4837 = ~n10485 ;
  assign y4838 = ~n10489 ;
  assign y4839 = n10490 ;
  assign y4840 = ~n10491 ;
  assign y4841 = ~n10492 ;
  assign y4842 = ~1'b0 ;
  assign y4843 = 1'b0 ;
  assign y4844 = ~1'b0 ;
  assign y4845 = n10493 ;
  assign y4846 = ~n10497 ;
  assign y4847 = ~1'b0 ;
  assign y4848 = ~1'b0 ;
  assign y4849 = ~n10498 ;
  assign y4850 = n10501 ;
  assign y4851 = ~n10507 ;
  assign y4852 = ~n997 ;
  assign y4853 = n10508 ;
  assign y4854 = n10509 ;
  assign y4855 = n10510 ;
  assign y4856 = n10512 ;
  assign y4857 = ~n10516 ;
  assign y4858 = n9067 ;
  assign y4859 = ~n10517 ;
  assign y4860 = ~n10518 ;
  assign y4861 = n10526 ;
  assign y4862 = ~n10535 ;
  assign y4863 = n10536 ;
  assign y4864 = ~n10537 ;
  assign y4865 = n10538 ;
  assign y4866 = ~1'b0 ;
  assign y4867 = n10542 ;
  assign y4868 = n10546 ;
  assign y4869 = ~n10549 ;
  assign y4870 = n10552 ;
  assign y4871 = ~n10554 ;
  assign y4872 = ~1'b0 ;
  assign y4873 = n7398 ;
  assign y4874 = ~n10556 ;
  assign y4875 = ~n10559 ;
  assign y4876 = ~n10561 ;
  assign y4877 = ~n10564 ;
  assign y4878 = n10567 ;
  assign y4879 = n10569 ;
  assign y4880 = ~1'b0 ;
  assign y4881 = n10571 ;
  assign y4882 = ~n10572 ;
  assign y4883 = n10574 ;
  assign y4884 = ~n10575 ;
  assign y4885 = ~n10586 ;
  assign y4886 = n10591 ;
  assign y4887 = ~n10598 ;
  assign y4888 = n10599 ;
  assign y4889 = ~n10601 ;
  assign y4890 = n6477 ;
  assign y4891 = ~n10603 ;
  assign y4892 = n10614 ;
  assign y4893 = n10618 ;
  assign y4894 = ~n10626 ;
  assign y4895 = ~1'b0 ;
  assign y4896 = n3806 ;
  assign y4897 = ~1'b0 ;
  assign y4898 = n10636 ;
  assign y4899 = ~n10637 ;
  assign y4900 = ~1'b0 ;
  assign y4901 = ~n10643 ;
  assign y4902 = n10644 ;
  assign y4903 = n10646 ;
  assign y4904 = n10651 ;
  assign y4905 = n10654 ;
  assign y4906 = n10655 ;
  assign y4907 = n10657 ;
  assign y4908 = ~n10659 ;
  assign y4909 = ~n10662 ;
  assign y4910 = ~1'b0 ;
  assign y4911 = ~n10663 ;
  assign y4912 = ~n10666 ;
  assign y4913 = ~n10668 ;
  assign y4914 = ~1'b0 ;
  assign y4915 = ~1'b0 ;
  assign y4916 = ~1'b0 ;
  assign y4917 = n10670 ;
  assign y4918 = ~n10672 ;
  assign y4919 = ~n10674 ;
  assign y4920 = n10676 ;
  assign y4921 = ~1'b0 ;
  assign y4922 = 1'b0 ;
  assign y4923 = ~n6830 ;
  assign y4924 = ~n10678 ;
  assign y4925 = n10679 ;
  assign y4926 = n10680 ;
  assign y4927 = ~n10682 ;
  assign y4928 = n10684 ;
  assign y4929 = ~1'b0 ;
  assign y4930 = 1'b0 ;
  assign y4931 = ~1'b0 ;
  assign y4932 = n10687 ;
  assign y4933 = n10691 ;
  assign y4934 = ~n10692 ;
  assign y4935 = ~1'b0 ;
  assign y4936 = ~1'b0 ;
  assign y4937 = n10695 ;
  assign y4938 = ~n3904 ;
  assign y4939 = n10699 ;
  assign y4940 = n10702 ;
  assign y4941 = ~n10705 ;
  assign y4942 = ~n10706 ;
  assign y4943 = ~n10710 ;
  assign y4944 = ~n10713 ;
  assign y4945 = ~1'b0 ;
  assign y4946 = ~1'b0 ;
  assign y4947 = ~n10714 ;
  assign y4948 = n10715 ;
  assign y4949 = ~n10719 ;
  assign y4950 = ~1'b0 ;
  assign y4951 = ~1'b0 ;
  assign y4952 = ~n10722 ;
  assign y4953 = ~n10724 ;
  assign y4954 = ~1'b0 ;
  assign y4955 = ~1'b0 ;
  assign y4956 = n10728 ;
  assign y4957 = n10732 ;
  assign y4958 = ~n10733 ;
  assign y4959 = ~1'b0 ;
  assign y4960 = ~n10737 ;
  assign y4961 = ~1'b0 ;
  assign y4962 = ~n10740 ;
  assign y4963 = n10741 ;
  assign y4964 = n10744 ;
  assign y4965 = ~1'b0 ;
  assign y4966 = ~n10746 ;
  assign y4967 = ~1'b0 ;
  assign y4968 = n10750 ;
  assign y4969 = n7002 ;
  assign y4970 = ~n10754 ;
  assign y4971 = ~n10755 ;
  assign y4972 = ~n10756 ;
  assign y4973 = ~n10758 ;
  assign y4974 = n10759 ;
  assign y4975 = ~n10762 ;
  assign y4976 = 1'b0 ;
  assign y4977 = ~1'b0 ;
  assign y4978 = ~1'b0 ;
  assign y4979 = 1'b0 ;
  assign y4980 = ~n10763 ;
  assign y4981 = ~n10766 ;
  assign y4982 = ~n10771 ;
  assign y4983 = n10777 ;
  assign y4984 = n10784 ;
  assign y4985 = ~1'b0 ;
  assign y4986 = ~1'b0 ;
  assign y4987 = ~n10785 ;
  assign y4988 = ~n10789 ;
  assign y4989 = n10790 ;
  assign y4990 = ~1'b0 ;
  assign y4991 = n1766 ;
  assign y4992 = ~n10792 ;
  assign y4993 = n10795 ;
  assign y4994 = ~1'b0 ;
  assign y4995 = ~n10797 ;
  assign y4996 = ~1'b0 ;
  assign y4997 = ~1'b0 ;
  assign y4998 = ~1'b0 ;
  assign y4999 = ~n10798 ;
  assign y5000 = ~1'b0 ;
  assign y5001 = ~n10803 ;
  assign y5002 = n10804 ;
  assign y5003 = n10808 ;
  assign y5004 = ~1'b0 ;
  assign y5005 = ~n10810 ;
  assign y5006 = ~n10813 ;
  assign y5007 = ~n10814 ;
  assign y5008 = ~n10820 ;
  assign y5009 = ~1'b0 ;
  assign y5010 = n10821 ;
  assign y5011 = ~n10822 ;
  assign y5012 = n10823 ;
  assign y5013 = n10826 ;
  assign y5014 = ~n10829 ;
  assign y5015 = ~1'b0 ;
  assign y5016 = n10832 ;
  assign y5017 = ~1'b0 ;
  assign y5018 = n6687 ;
  assign y5019 = ~1'b0 ;
  assign y5020 = ~n10834 ;
  assign y5021 = n3594 ;
  assign y5022 = ~1'b0 ;
  assign y5023 = ~n10840 ;
  assign y5024 = ~n10841 ;
  assign y5025 = n2830 ;
  assign y5026 = ~1'b0 ;
  assign y5027 = n10845 ;
  assign y5028 = ~n10847 ;
  assign y5029 = n10851 ;
  assign y5030 = ~n10852 ;
  assign y5031 = ~1'b0 ;
  assign y5032 = 1'b0 ;
  assign y5033 = n10854 ;
  assign y5034 = n10855 ;
  assign y5035 = n10862 ;
  assign y5036 = ~1'b0 ;
  assign y5037 = ~1'b0 ;
  assign y5038 = ~n10871 ;
  assign y5039 = ~n10877 ;
  assign y5040 = ~1'b0 ;
  assign y5041 = ~1'b0 ;
  assign y5042 = ~1'b0 ;
  assign y5043 = ~n10878 ;
  assign y5044 = ~n10886 ;
  assign y5045 = ~n10893 ;
  assign y5046 = n10894 ;
  assign y5047 = ~n10897 ;
  assign y5048 = ~1'b0 ;
  assign y5049 = ~1'b0 ;
  assign y5050 = ~n10900 ;
  assign y5051 = ~n10903 ;
  assign y5052 = ~1'b0 ;
  assign y5053 = ~n10907 ;
  assign y5054 = n10908 ;
  assign y5055 = ~1'b0 ;
  assign y5056 = ~n10913 ;
  assign y5057 = ~1'b0 ;
  assign y5058 = n10918 ;
  assign y5059 = n10922 ;
  assign y5060 = n10923 ;
  assign y5061 = ~1'b0 ;
  assign y5062 = ~n10926 ;
  assign y5063 = n2062 ;
  assign y5064 = ~n10930 ;
  assign y5065 = n10934 ;
  assign y5066 = ~1'b0 ;
  assign y5067 = ~1'b0 ;
  assign y5068 = n10935 ;
  assign y5069 = ~n10940 ;
  assign y5070 = ~1'b0 ;
  assign y5071 = n10947 ;
  assign y5072 = ~1'b0 ;
  assign y5073 = n10950 ;
  assign y5074 = ~n10955 ;
  assign y5075 = ~n10959 ;
  assign y5076 = ~1'b0 ;
  assign y5077 = n10960 ;
  assign y5078 = ~1'b0 ;
  assign y5079 = n10963 ;
  assign y5080 = ~1'b0 ;
  assign y5081 = n10966 ;
  assign y5082 = ~n10969 ;
  assign y5083 = n10971 ;
  assign y5084 = n10982 ;
  assign y5085 = ~n5047 ;
  assign y5086 = ~n10984 ;
  assign y5087 = n10986 ;
  assign y5088 = n10990 ;
  assign y5089 = ~1'b0 ;
  assign y5090 = n10994 ;
  assign y5091 = n10996 ;
  assign y5092 = ~n10999 ;
  assign y5093 = ~1'b0 ;
  assign y5094 = ~n11008 ;
  assign y5095 = n11010 ;
  assign y5096 = n11019 ;
  assign y5097 = ~n11020 ;
  assign y5098 = ~1'b0 ;
  assign y5099 = n11028 ;
  assign y5100 = ~n11029 ;
  assign y5101 = ~n11030 ;
  assign y5102 = ~n11034 ;
  assign y5103 = ~n11035 ;
  assign y5104 = ~n11044 ;
  assign y5105 = n11046 ;
  assign y5106 = ~1'b0 ;
  assign y5107 = ~n11047 ;
  assign y5108 = n11052 ;
  assign y5109 = ~1'b0 ;
  assign y5110 = ~n11053 ;
  assign y5111 = ~n11059 ;
  assign y5112 = ~1'b0 ;
  assign y5113 = ~n11071 ;
  assign y5114 = ~n11072 ;
  assign y5115 = n6049 ;
  assign y5116 = n11074 ;
  assign y5117 = ~1'b0 ;
  assign y5118 = ~1'b0 ;
  assign y5119 = n11077 ;
  assign y5120 = ~n11078 ;
  assign y5121 = ~n11080 ;
  assign y5122 = ~n11081 ;
  assign y5123 = n11083 ;
  assign y5124 = ~n11084 ;
  assign y5125 = ~1'b0 ;
  assign y5126 = n11017 ;
  assign y5127 = ~n11093 ;
  assign y5128 = ~n11094 ;
  assign y5129 = ~n11096 ;
  assign y5130 = ~1'b0 ;
  assign y5131 = n11103 ;
  assign y5132 = ~1'b0 ;
  assign y5133 = ~n11109 ;
  assign y5134 = ~n11110 ;
  assign y5135 = ~n7107 ;
  assign y5136 = n11112 ;
  assign y5137 = ~n11114 ;
  assign y5138 = ~1'b0 ;
  assign y5139 = n11118 ;
  assign y5140 = ~n11119 ;
  assign y5141 = ~n11122 ;
  assign y5142 = ~1'b0 ;
  assign y5143 = 1'b0 ;
  assign y5144 = ~n11125 ;
  assign y5145 = n11128 ;
  assign y5146 = ~n11130 ;
  assign y5147 = n11134 ;
  assign y5148 = ~n11135 ;
  assign y5149 = ~1'b0 ;
  assign y5150 = 1'b0 ;
  assign y5151 = ~n11138 ;
  assign y5152 = ~n11141 ;
  assign y5153 = ~n11142 ;
  assign y5154 = ~n11144 ;
  assign y5155 = ~1'b0 ;
  assign y5156 = n4721 ;
  assign y5157 = ~n11147 ;
  assign y5158 = ~1'b0 ;
  assign y5159 = ~n11148 ;
  assign y5160 = ~n11153 ;
  assign y5161 = n11158 ;
  assign y5162 = n4010 ;
  assign y5163 = n11164 ;
  assign y5164 = n11167 ;
  assign y5165 = ~1'b0 ;
  assign y5166 = ~n8233 ;
  assign y5167 = n11168 ;
  assign y5168 = ~n11172 ;
  assign y5169 = 1'b0 ;
  assign y5170 = n11174 ;
  assign y5171 = ~1'b0 ;
  assign y5172 = ~n11179 ;
  assign y5173 = ~1'b0 ;
  assign y5174 = ~n11182 ;
  assign y5175 = n11184 ;
  assign y5176 = ~n992 ;
  assign y5177 = ~n11186 ;
  assign y5178 = ~n11195 ;
  assign y5179 = n11203 ;
  assign y5180 = n11204 ;
  assign y5181 = ~n11208 ;
  assign y5182 = ~1'b0 ;
  assign y5183 = ~1'b0 ;
  assign y5184 = n11224 ;
  assign y5185 = ~n796 ;
  assign y5186 = n5143 ;
  assign y5187 = ~n11234 ;
  assign y5188 = n11235 ;
  assign y5189 = ~n11237 ;
  assign y5190 = ~n11239 ;
  assign y5191 = ~n11241 ;
  assign y5192 = n11244 ;
  assign y5193 = ~1'b0 ;
  assign y5194 = ~n11245 ;
  assign y5195 = ~n11247 ;
  assign y5196 = ~n11249 ;
  assign y5197 = ~1'b0 ;
  assign y5198 = ~1'b0 ;
  assign y5199 = ~n8843 ;
  assign y5200 = ~1'b0 ;
  assign y5201 = ~n5437 ;
  assign y5202 = ~n11253 ;
  assign y5203 = ~1'b0 ;
  assign y5204 = ~n11255 ;
  assign y5205 = n11256 ;
  assign y5206 = n11257 ;
  assign y5207 = ~1'b0 ;
  assign y5208 = n11260 ;
  assign y5209 = ~1'b0 ;
  assign y5210 = n11262 ;
  assign y5211 = ~1'b0 ;
  assign y5212 = n2319 ;
  assign y5213 = ~n11264 ;
  assign y5214 = ~1'b0 ;
  assign y5215 = ~1'b0 ;
  assign y5216 = ~n11269 ;
  assign y5217 = n11275 ;
  assign y5218 = n11276 ;
  assign y5219 = ~n11277 ;
  assign y5220 = n11279 ;
  assign y5221 = ~1'b0 ;
  assign y5222 = ~n11280 ;
  assign y5223 = ~n3210 ;
  assign y5224 = ~1'b0 ;
  assign y5225 = 1'b0 ;
  assign y5226 = ~n11284 ;
  assign y5227 = n11287 ;
  assign y5228 = ~n11288 ;
  assign y5229 = ~1'b0 ;
  assign y5230 = ~n5659 ;
  assign y5231 = n11291 ;
  assign y5232 = ~1'b0 ;
  assign y5233 = ~n6793 ;
  assign y5234 = n11299 ;
  assign y5235 = n11311 ;
  assign y5236 = ~n11314 ;
  assign y5237 = ~n5075 ;
  assign y5238 = ~n4169 ;
  assign y5239 = ~n11319 ;
  assign y5240 = ~1'b0 ;
  assign y5241 = ~1'b0 ;
  assign y5242 = ~n3479 ;
  assign y5243 = n11320 ;
  assign y5244 = n11324 ;
  assign y5245 = n11326 ;
  assign y5246 = ~1'b0 ;
  assign y5247 = n11327 ;
  assign y5248 = ~n9649 ;
  assign y5249 = ~n11328 ;
  assign y5250 = ~1'b0 ;
  assign y5251 = n11330 ;
  assign y5252 = ~1'b0 ;
  assign y5253 = ~1'b0 ;
  assign y5254 = ~n11333 ;
  assign y5255 = n11334 ;
  assign y5256 = n6471 ;
  assign y5257 = ~n11336 ;
  assign y5258 = ~1'b0 ;
  assign y5259 = ~n3986 ;
  assign y5260 = n11339 ;
  assign y5261 = ~n11340 ;
  assign y5262 = n11341 ;
  assign y5263 = ~n8178 ;
  assign y5264 = n11346 ;
  assign y5265 = n11347 ;
  assign y5266 = ~n11353 ;
  assign y5267 = ~1'b0 ;
  assign y5268 = ~1'b0 ;
  assign y5269 = ~1'b0 ;
  assign y5270 = ~1'b0 ;
  assign y5271 = ~n11355 ;
  assign y5272 = ~1'b0 ;
  assign y5273 = ~n11357 ;
  assign y5274 = ~1'b0 ;
  assign y5275 = ~1'b0 ;
  assign y5276 = n11358 ;
  assign y5277 = ~n11359 ;
  assign y5278 = n11361 ;
  assign y5279 = ~n11365 ;
  assign y5280 = n11369 ;
  assign y5281 = ~1'b0 ;
  assign y5282 = ~1'b0 ;
  assign y5283 = n11372 ;
  assign y5284 = ~n11373 ;
  assign y5285 = ~1'b0 ;
  assign y5286 = ~n11374 ;
  assign y5287 = ~n11377 ;
  assign y5288 = ~n11379 ;
  assign y5289 = ~n11382 ;
  assign y5290 = ~1'b0 ;
  assign y5291 = ~1'b0 ;
  assign y5292 = n11383 ;
  assign y5293 = ~1'b0 ;
  assign y5294 = ~n11384 ;
  assign y5295 = n11386 ;
  assign y5296 = ~1'b0 ;
  assign y5297 = ~n11388 ;
  assign y5298 = ~1'b0 ;
  assign y5299 = ~1'b0 ;
  assign y5300 = ~n11390 ;
  assign y5301 = ~n11392 ;
  assign y5302 = ~n11396 ;
  assign y5303 = ~1'b0 ;
  assign y5304 = ~n11399 ;
  assign y5305 = ~n8107 ;
  assign y5306 = ~n11401 ;
  assign y5307 = ~n11402 ;
  assign y5308 = n11405 ;
  assign y5309 = n11411 ;
  assign y5310 = ~n11415 ;
  assign y5311 = n11416 ;
  assign y5312 = 1'b0 ;
  assign y5313 = n11428 ;
  assign y5314 = ~1'b0 ;
  assign y5315 = ~1'b0 ;
  assign y5316 = n11431 ;
  assign y5317 = n11437 ;
  assign y5318 = ~n11443 ;
  assign y5319 = ~1'b0 ;
  assign y5320 = ~n11444 ;
  assign y5321 = ~n11447 ;
  assign y5322 = ~1'b0 ;
  assign y5323 = ~n11452 ;
  assign y5324 = n888 ;
  assign y5325 = 1'b0 ;
  assign y5326 = n11455 ;
  assign y5327 = ~1'b0 ;
  assign y5328 = n11457 ;
  assign y5329 = n11458 ;
  assign y5330 = n11459 ;
  assign y5331 = ~n11460 ;
  assign y5332 = ~1'b0 ;
  assign y5333 = ~1'b0 ;
  assign y5334 = n11461 ;
  assign y5335 = ~n11464 ;
  assign y5336 = ~1'b0 ;
  assign y5337 = ~1'b0 ;
  assign y5338 = ~n11467 ;
  assign y5339 = n11468 ;
  assign y5340 = ~n10554 ;
  assign y5341 = n11476 ;
  assign y5342 = n11482 ;
  assign y5343 = n11483 ;
  assign y5344 = ~1'b0 ;
  assign y5345 = ~n11487 ;
  assign y5346 = ~n11493 ;
  assign y5347 = ~1'b0 ;
  assign y5348 = n11498 ;
  assign y5349 = ~n11502 ;
  assign y5350 = n11504 ;
  assign y5351 = n11515 ;
  assign y5352 = ~n11531 ;
  assign y5353 = n11534 ;
  assign y5354 = ~1'b0 ;
  assign y5355 = ~n11541 ;
  assign y5356 = ~n11547 ;
  assign y5357 = n11548 ;
  assign y5358 = ~n11549 ;
  assign y5359 = ~n11552 ;
  assign y5360 = n11561 ;
  assign y5361 = ~n9218 ;
  assign y5362 = n11568 ;
  assign y5363 = ~n11576 ;
  assign y5364 = ~1'b0 ;
  assign y5365 = ~1'b0 ;
  assign y5366 = n11585 ;
  assign y5367 = ~n11592 ;
  assign y5368 = ~n11593 ;
  assign y5369 = ~n11594 ;
  assign y5370 = ~n11596 ;
  assign y5371 = ~n11602 ;
  assign y5372 = ~n11603 ;
  assign y5373 = n11606 ;
  assign y5374 = ~1'b0 ;
  assign y5375 = ~1'b0 ;
  assign y5376 = ~n11607 ;
  assign y5377 = ~1'b0 ;
  assign y5378 = ~n11608 ;
  assign y5379 = n11609 ;
  assign y5380 = n11613 ;
  assign y5381 = ~1'b0 ;
  assign y5382 = n11614 ;
  assign y5383 = ~1'b0 ;
  assign y5384 = ~n11619 ;
  assign y5385 = n11621 ;
  assign y5386 = ~n11622 ;
  assign y5387 = n11623 ;
  assign y5388 = n11625 ;
  assign y5389 = ~n11630 ;
  assign y5390 = n8073 ;
  assign y5391 = n11632 ;
  assign y5392 = n11633 ;
  assign y5393 = ~1'b0 ;
  assign y5394 = ~n11636 ;
  assign y5395 = n11640 ;
  assign y5396 = ~1'b0 ;
  assign y5397 = n11645 ;
  assign y5398 = ~n11650 ;
  assign y5399 = n11653 ;
  assign y5400 = n11655 ;
  assign y5401 = ~1'b0 ;
  assign y5402 = ~1'b0 ;
  assign y5403 = ~n11660 ;
  assign y5404 = n11663 ;
  assign y5405 = ~1'b0 ;
  assign y5406 = ~n11665 ;
  assign y5407 = n11666 ;
  assign y5408 = ~n11671 ;
  assign y5409 = ~n11674 ;
  assign y5410 = n11678 ;
  assign y5411 = ~1'b0 ;
  assign y5412 = n11685 ;
  assign y5413 = n11687 ;
  assign y5414 = ~1'b0 ;
  assign y5415 = n10247 ;
  assign y5416 = ~1'b0 ;
  assign y5417 = ~n11689 ;
  assign y5418 = n7663 ;
  assign y5419 = ~n11691 ;
  assign y5420 = ~n11699 ;
  assign y5421 = n11700 ;
  assign y5422 = ~n7877 ;
  assign y5423 = ~1'b0 ;
  assign y5424 = ~1'b0 ;
  assign y5425 = ~1'b0 ;
  assign y5426 = ~1'b0 ;
  assign y5427 = ~1'b0 ;
  assign y5428 = ~1'b0 ;
  assign y5429 = ~1'b0 ;
  assign y5430 = n11701 ;
  assign y5431 = ~1'b0 ;
  assign y5432 = ~n11709 ;
  assign y5433 = ~n11712 ;
  assign y5434 = n7623 ;
  assign y5435 = ~1'b0 ;
  assign y5436 = n11719 ;
  assign y5437 = n11721 ;
  assign y5438 = ~n11722 ;
  assign y5439 = ~n11723 ;
  assign y5440 = ~n11725 ;
  assign y5441 = ~n11730 ;
  assign y5442 = ~1'b0 ;
  assign y5443 = ~n11735 ;
  assign y5444 = ~1'b0 ;
  assign y5445 = n11741 ;
  assign y5446 = n11743 ;
  assign y5447 = ~n11745 ;
  assign y5448 = n11749 ;
  assign y5449 = ~1'b0 ;
  assign y5450 = n11754 ;
  assign y5451 = n11755 ;
  assign y5452 = n11757 ;
  assign y5453 = n11758 ;
  assign y5454 = ~n11763 ;
  assign y5455 = ~n1499 ;
  assign y5456 = ~n11766 ;
  assign y5457 = n11767 ;
  assign y5458 = n11769 ;
  assign y5459 = n11772 ;
  assign y5460 = ~n11773 ;
  assign y5461 = ~1'b0 ;
  assign y5462 = ~1'b0 ;
  assign y5463 = ~n10805 ;
  assign y5464 = ~1'b0 ;
  assign y5465 = n11775 ;
  assign y5466 = n11778 ;
  assign y5467 = ~n11780 ;
  assign y5468 = 1'b0 ;
  assign y5469 = 1'b0 ;
  assign y5470 = ~n11782 ;
  assign y5471 = ~n11788 ;
  assign y5472 = ~n11793 ;
  assign y5473 = ~1'b0 ;
  assign y5474 = ~n11796 ;
  assign y5475 = ~1'b0 ;
  assign y5476 = ~n11798 ;
  assign y5477 = n11804 ;
  assign y5478 = ~1'b0 ;
  assign y5479 = ~n11805 ;
  assign y5480 = n11807 ;
  assign y5481 = ~1'b0 ;
  assign y5482 = ~1'b0 ;
  assign y5483 = n11808 ;
  assign y5484 = ~1'b0 ;
  assign y5485 = n11811 ;
  assign y5486 = ~1'b0 ;
  assign y5487 = ~n11814 ;
  assign y5488 = n11815 ;
  assign y5489 = ~1'b0 ;
  assign y5490 = n11817 ;
  assign y5491 = n11821 ;
  assign y5492 = ~1'b0 ;
  assign y5493 = ~1'b0 ;
  assign y5494 = ~n11822 ;
  assign y5495 = ~n11836 ;
  assign y5496 = ~1'b0 ;
  assign y5497 = n11840 ;
  assign y5498 = ~n11842 ;
  assign y5499 = ~n9973 ;
  assign y5500 = ~1'b0 ;
  assign y5501 = n11843 ;
  assign y5502 = ~1'b0 ;
  assign y5503 = ~1'b0 ;
  assign y5504 = ~1'b0 ;
  assign y5505 = n11848 ;
  assign y5506 = ~n11849 ;
  assign y5507 = ~n11853 ;
  assign y5508 = n11856 ;
  assign y5509 = ~1'b0 ;
  assign y5510 = ~n11857 ;
  assign y5511 = ~n11858 ;
  assign y5512 = n11861 ;
  assign y5513 = ~1'b0 ;
  assign y5514 = ~n11864 ;
  assign y5515 = ~n11867 ;
  assign y5516 = n11870 ;
  assign y5517 = ~n11872 ;
  assign y5518 = ~n11873 ;
  assign y5519 = ~n11875 ;
  assign y5520 = ~1'b0 ;
  assign y5521 = ~n11885 ;
  assign y5522 = x171 ;
  assign y5523 = n11887 ;
  assign y5524 = ~1'b0 ;
  assign y5525 = ~n11891 ;
  assign y5526 = ~n11898 ;
  assign y5527 = n10733 ;
  assign y5528 = ~1'b0 ;
  assign y5529 = n11899 ;
  assign y5530 = 1'b0 ;
  assign y5531 = ~n11902 ;
  assign y5532 = n11909 ;
  assign y5533 = ~1'b0 ;
  assign y5534 = n11910 ;
  assign y5535 = ~n11911 ;
  assign y5536 = ~n11917 ;
  assign y5537 = n10169 ;
  assign y5538 = n11923 ;
  assign y5539 = n11924 ;
  assign y5540 = ~n11926 ;
  assign y5541 = ~1'b0 ;
  assign y5542 = 1'b0 ;
  assign y5543 = ~n11927 ;
  assign y5544 = ~1'b0 ;
  assign y5545 = n11929 ;
  assign y5546 = ~1'b0 ;
  assign y5547 = n11930 ;
  assign y5548 = ~1'b0 ;
  assign y5549 = ~1'b0 ;
  assign y5550 = ~n11933 ;
  assign y5551 = n11934 ;
  assign y5552 = ~n11935 ;
  assign y5553 = n11936 ;
  assign y5554 = n11939 ;
  assign y5555 = n11947 ;
  assign y5556 = ~1'b0 ;
  assign y5557 = ~n11952 ;
  assign y5558 = ~1'b0 ;
  assign y5559 = ~n11955 ;
  assign y5560 = ~n11957 ;
  assign y5561 = ~n11965 ;
  assign y5562 = ~n11968 ;
  assign y5563 = ~1'b0 ;
  assign y5564 = ~1'b0 ;
  assign y5565 = ~n11972 ;
  assign y5566 = n11974 ;
  assign y5567 = ~n11975 ;
  assign y5568 = ~1'b0 ;
  assign y5569 = ~n11979 ;
  assign y5570 = ~n11982 ;
  assign y5571 = n8087 ;
  assign y5572 = ~1'b0 ;
  assign y5573 = ~n11985 ;
  assign y5574 = n372 ;
  assign y5575 = ~1'b0 ;
  assign y5576 = n11994 ;
  assign y5577 = n11995 ;
  assign y5578 = ~1'b0 ;
  assign y5579 = ~n12000 ;
  assign y5580 = ~1'b0 ;
  assign y5581 = ~1'b0 ;
  assign y5582 = ~1'b0 ;
  assign y5583 = ~n12002 ;
  assign y5584 = n12006 ;
  assign y5585 = n12008 ;
  assign y5586 = n12015 ;
  assign y5587 = n12017 ;
  assign y5588 = ~n12019 ;
  assign y5589 = n12020 ;
  assign y5590 = n12022 ;
  assign y5591 = ~1'b0 ;
  assign y5592 = ~n6075 ;
  assign y5593 = n12024 ;
  assign y5594 = ~n12028 ;
  assign y5595 = n12029 ;
  assign y5596 = ~1'b0 ;
  assign y5597 = n12034 ;
  assign y5598 = n12038 ;
  assign y5599 = n12040 ;
  assign y5600 = n12041 ;
  assign y5601 = n12052 ;
  assign y5602 = n12053 ;
  assign y5603 = n12057 ;
  assign y5604 = ~n12058 ;
  assign y5605 = n12059 ;
  assign y5606 = ~1'b0 ;
  assign y5607 = n12063 ;
  assign y5608 = n12068 ;
  assign y5609 = ~1'b0 ;
  assign y5610 = ~n12075 ;
  assign y5611 = ~1'b0 ;
  assign y5612 = n12077 ;
  assign y5613 = ~n12079 ;
  assign y5614 = ~n12080 ;
  assign y5615 = n12083 ;
  assign y5616 = ~1'b0 ;
  assign y5617 = ~n12087 ;
  assign y5618 = ~n12090 ;
  assign y5619 = n4364 ;
  assign y5620 = n12099 ;
  assign y5621 = n12100 ;
  assign y5622 = ~n7022 ;
  assign y5623 = ~1'b0 ;
  assign y5624 = ~n12102 ;
  assign y5625 = ~n12105 ;
  assign y5626 = n12106 ;
  assign y5627 = ~n12107 ;
  assign y5628 = n2831 ;
  assign y5629 = n12109 ;
  assign y5630 = ~1'b0 ;
  assign y5631 = n12112 ;
  assign y5632 = n12113 ;
  assign y5633 = ~n12119 ;
  assign y5634 = ~1'b0 ;
  assign y5635 = n12120 ;
  assign y5636 = ~n12126 ;
  assign y5637 = n12129 ;
  assign y5638 = ~n12131 ;
  assign y5639 = ~n12133 ;
  assign y5640 = ~1'b0 ;
  assign y5641 = ~1'b0 ;
  assign y5642 = ~n12138 ;
  assign y5643 = ~n12139 ;
  assign y5644 = n12140 ;
  assign y5645 = n12145 ;
  assign y5646 = ~n12148 ;
  assign y5647 = ~n12153 ;
  assign y5648 = ~n12155 ;
  assign y5649 = ~n12157 ;
  assign y5650 = ~1'b0 ;
  assign y5651 = n3588 ;
  assign y5652 = ~1'b0 ;
  assign y5653 = ~n12159 ;
  assign y5654 = ~n12161 ;
  assign y5655 = ~1'b0 ;
  assign y5656 = ~n8216 ;
  assign y5657 = ~n12167 ;
  assign y5658 = ~1'b0 ;
  assign y5659 = ~n12180 ;
  assign y5660 = n12182 ;
  assign y5661 = ~1'b0 ;
  assign y5662 = ~1'b0 ;
  assign y5663 = ~1'b0 ;
  assign y5664 = n6046 ;
  assign y5665 = ~n12183 ;
  assign y5666 = n12186 ;
  assign y5667 = n12190 ;
  assign y5668 = ~n12192 ;
  assign y5669 = ~1'b0 ;
  assign y5670 = ~1'b0 ;
  assign y5671 = ~n12193 ;
  assign y5672 = ~n12197 ;
  assign y5673 = ~1'b0 ;
  assign y5674 = ~n12200 ;
  assign y5675 = n12201 ;
  assign y5676 = n12204 ;
  assign y5677 = ~1'b0 ;
  assign y5678 = ~n12205 ;
  assign y5679 = n1059 ;
  assign y5680 = n12210 ;
  assign y5681 = ~n12212 ;
  assign y5682 = ~n12214 ;
  assign y5683 = ~1'b0 ;
  assign y5684 = ~n12217 ;
  assign y5685 = ~n12220 ;
  assign y5686 = n12225 ;
  assign y5687 = ~1'b0 ;
  assign y5688 = ~n12228 ;
  assign y5689 = ~n12232 ;
  assign y5690 = ~1'b0 ;
  assign y5691 = ~n12234 ;
  assign y5692 = n12236 ;
  assign y5693 = ~n12240 ;
  assign y5694 = ~n12241 ;
  assign y5695 = n6616 ;
  assign y5696 = ~1'b0 ;
  assign y5697 = ~n12245 ;
  assign y5698 = ~n5961 ;
  assign y5699 = n12246 ;
  assign y5700 = n12253 ;
  assign y5701 = ~1'b0 ;
  assign y5702 = n12254 ;
  assign y5703 = ~1'b0 ;
  assign y5704 = ~n12256 ;
  assign y5705 = ~n12259 ;
  assign y5706 = ~n12262 ;
  assign y5707 = ~1'b0 ;
  assign y5708 = n12266 ;
  assign y5709 = ~n12267 ;
  assign y5710 = ~n12271 ;
  assign y5711 = ~x230 ;
  assign y5712 = n12274 ;
  assign y5713 = ~n12278 ;
  assign y5714 = ~n12280 ;
  assign y5715 = ~1'b0 ;
  assign y5716 = ~n12283 ;
  assign y5717 = ~n12287 ;
  assign y5718 = ~n12288 ;
  assign y5719 = n3565 ;
  assign y5720 = ~1'b0 ;
  assign y5721 = ~1'b0 ;
  assign y5722 = ~n12290 ;
  assign y5723 = ~1'b0 ;
  assign y5724 = ~1'b0 ;
  assign y5725 = ~n12292 ;
  assign y5726 = ~n12295 ;
  assign y5727 = n12297 ;
  assign y5728 = ~n2870 ;
  assign y5729 = ~1'b0 ;
  assign y5730 = n10731 ;
  assign y5731 = ~n12298 ;
  assign y5732 = ~n12301 ;
  assign y5733 = n2743 ;
  assign y5734 = n12306 ;
  assign y5735 = n12308 ;
  assign y5736 = ~n12309 ;
  assign y5737 = ~n12310 ;
  assign y5738 = n12312 ;
  assign y5739 = n12316 ;
  assign y5740 = n12319 ;
  assign y5741 = ~1'b0 ;
  assign y5742 = n12323 ;
  assign y5743 = ~1'b0 ;
  assign y5744 = ~1'b0 ;
  assign y5745 = ~1'b0 ;
  assign y5746 = n6733 ;
  assign y5747 = ~1'b0 ;
  assign y5748 = ~n12329 ;
  assign y5749 = n12332 ;
  assign y5750 = ~1'b0 ;
  assign y5751 = 1'b0 ;
  assign y5752 = n12333 ;
  assign y5753 = ~1'b0 ;
  assign y5754 = n12335 ;
  assign y5755 = ~n12337 ;
  assign y5756 = n12338 ;
  assign y5757 = n12342 ;
  assign y5758 = n12346 ;
  assign y5759 = ~n12352 ;
  assign y5760 = n12354 ;
  assign y5761 = ~1'b0 ;
  assign y5762 = n12357 ;
  assign y5763 = ~1'b0 ;
  assign y5764 = n12361 ;
  assign y5765 = n12363 ;
  assign y5766 = ~1'b0 ;
  assign y5767 = 1'b0 ;
  assign y5768 = ~n12364 ;
  assign y5769 = n12367 ;
  assign y5770 = n12369 ;
  assign y5771 = ~1'b0 ;
  assign y5772 = ~1'b0 ;
  assign y5773 = n12371 ;
  assign y5774 = ~n12372 ;
  assign y5775 = ~n12375 ;
  assign y5776 = ~n12379 ;
  assign y5777 = ~n12384 ;
  assign y5778 = ~x180 ;
  assign y5779 = n12386 ;
  assign y5780 = ~n12388 ;
  assign y5781 = ~n12393 ;
  assign y5782 = ~n12394 ;
  assign y5783 = ~1'b0 ;
  assign y5784 = n12395 ;
  assign y5785 = ~n12397 ;
  assign y5786 = ~1'b0 ;
  assign y5787 = ~1'b0 ;
  assign y5788 = n12398 ;
  assign y5789 = ~1'b0 ;
  assign y5790 = ~1'b0 ;
  assign y5791 = ~n12400 ;
  assign y5792 = ~1'b0 ;
  assign y5793 = ~1'b0 ;
  assign y5794 = n12410 ;
  assign y5795 = n12413 ;
  assign y5796 = n12417 ;
  assign y5797 = n12421 ;
  assign y5798 = n1521 ;
  assign y5799 = 1'b0 ;
  assign y5800 = ~n12422 ;
  assign y5801 = ~n12428 ;
  assign y5802 = n12429 ;
  assign y5803 = n12435 ;
  assign y5804 = ~1'b0 ;
  assign y5805 = ~1'b0 ;
  assign y5806 = n12439 ;
  assign y5807 = ~1'b0 ;
  assign y5808 = n12441 ;
  assign y5809 = ~1'b0 ;
  assign y5810 = ~n12444 ;
  assign y5811 = n12445 ;
  assign y5812 = ~n12447 ;
  assign y5813 = ~n12448 ;
  assign y5814 = n12449 ;
  assign y5815 = ~n12450 ;
  assign y5816 = ~1'b0 ;
  assign y5817 = ~1'b0 ;
  assign y5818 = 1'b0 ;
  assign y5819 = n12451 ;
  assign y5820 = ~1'b0 ;
  assign y5821 = ~1'b0 ;
  assign y5822 = ~1'b0 ;
  assign y5823 = n12461 ;
  assign y5824 = ~n12462 ;
  assign y5825 = n12464 ;
  assign y5826 = ~n12465 ;
  assign y5827 = ~1'b0 ;
  assign y5828 = ~1'b0 ;
  assign y5829 = ~1'b0 ;
  assign y5830 = ~n4072 ;
  assign y5831 = n12471 ;
  assign y5832 = n12473 ;
  assign y5833 = ~n12476 ;
  assign y5834 = ~1'b0 ;
  assign y5835 = ~n12479 ;
  assign y5836 = ~1'b0 ;
  assign y5837 = ~n12488 ;
  assign y5838 = n12490 ;
  assign y5839 = n375 ;
  assign y5840 = ~1'b0 ;
  assign y5841 = ~1'b0 ;
  assign y5842 = ~n12495 ;
  assign y5843 = n7586 ;
  assign y5844 = ~n12503 ;
  assign y5845 = n12509 ;
  assign y5846 = ~1'b0 ;
  assign y5847 = n12511 ;
  assign y5848 = n12514 ;
  assign y5849 = ~n12520 ;
  assign y5850 = ~n12522 ;
  assign y5851 = n12526 ;
  assign y5852 = ~n12528 ;
  assign y5853 = n12530 ;
  assign y5854 = ~n12531 ;
  assign y5855 = n5416 ;
  assign y5856 = ~1'b0 ;
  assign y5857 = ~1'b0 ;
  assign y5858 = ~1'b0 ;
  assign y5859 = ~n12533 ;
  assign y5860 = ~1'b0 ;
  assign y5861 = ~n12534 ;
  assign y5862 = ~1'b0 ;
  assign y5863 = n12535 ;
  assign y5864 = ~1'b0 ;
  assign y5865 = n12537 ;
  assign y5866 = ~n12544 ;
  assign y5867 = ~1'b0 ;
  assign y5868 = n12549 ;
  assign y5869 = n7379 ;
  assign y5870 = n12550 ;
  assign y5871 = ~1'b0 ;
  assign y5872 = n12552 ;
  assign y5873 = n12553 ;
  assign y5874 = ~1'b0 ;
  assign y5875 = ~1'b0 ;
  assign y5876 = n7462 ;
  assign y5877 = ~1'b0 ;
  assign y5878 = ~n12554 ;
  assign y5879 = ~n12559 ;
  assign y5880 = ~1'b0 ;
  assign y5881 = ~1'b0 ;
  assign y5882 = n12565 ;
  assign y5883 = ~n12567 ;
  assign y5884 = ~n12574 ;
  assign y5885 = ~n12578 ;
  assign y5886 = ~1'b0 ;
  assign y5887 = ~1'b0 ;
  assign y5888 = 1'b0 ;
  assign y5889 = n12580 ;
  assign y5890 = ~1'b0 ;
  assign y5891 = n12583 ;
  assign y5892 = 1'b0 ;
  assign y5893 = ~n8079 ;
  assign y5894 = n12585 ;
  assign y5895 = ~n12586 ;
  assign y5896 = ~n12591 ;
  assign y5897 = ~1'b0 ;
  assign y5898 = ~1'b0 ;
  assign y5899 = ~n12592 ;
  assign y5900 = n12596 ;
  assign y5901 = n12597 ;
  assign y5902 = ~1'b0 ;
  assign y5903 = n12599 ;
  assign y5904 = ~n12601 ;
  assign y5905 = ~n12607 ;
  assign y5906 = n12608 ;
  assign y5907 = ~1'b0 ;
  assign y5908 = ~1'b0 ;
  assign y5909 = ~1'b0 ;
  assign y5910 = ~1'b0 ;
  assign y5911 = ~n12609 ;
  assign y5912 = 1'b0 ;
  assign y5913 = ~n12610 ;
  assign y5914 = n12611 ;
  assign y5915 = ~1'b0 ;
  assign y5916 = n12614 ;
  assign y5917 = n12617 ;
  assign y5918 = ~n12619 ;
  assign y5919 = ~n12622 ;
  assign y5920 = n12623 ;
  assign y5921 = ~n12628 ;
  assign y5922 = 1'b0 ;
  assign y5923 = ~1'b0 ;
  assign y5924 = ~1'b0 ;
  assign y5925 = n12631 ;
  assign y5926 = ~n12633 ;
  assign y5927 = ~1'b0 ;
  assign y5928 = ~n12634 ;
  assign y5929 = ~1'b0 ;
  assign y5930 = ~1'b0 ;
  assign y5931 = n3704 ;
  assign y5932 = 1'b0 ;
  assign y5933 = ~1'b0 ;
  assign y5934 = n4387 ;
  assign y5935 = n12636 ;
  assign y5936 = ~n12639 ;
  assign y5937 = ~n12641 ;
  assign y5938 = ~n12651 ;
  assign y5939 = n12655 ;
  assign y5940 = ~n12656 ;
  assign y5941 = ~n12659 ;
  assign y5942 = n12660 ;
  assign y5943 = ~1'b0 ;
  assign y5944 = n12661 ;
  assign y5945 = ~1'b0 ;
  assign y5946 = n12663 ;
  assign y5947 = ~1'b0 ;
  assign y5948 = ~n12667 ;
  assign y5949 = ~n12669 ;
  assign y5950 = ~1'b0 ;
  assign y5951 = ~n12673 ;
  assign y5952 = n12674 ;
  assign y5953 = n12683 ;
  assign y5954 = ~1'b0 ;
  assign y5955 = n501 ;
  assign y5956 = n12684 ;
  assign y5957 = n12686 ;
  assign y5958 = ~1'b0 ;
  assign y5959 = ~1'b0 ;
  assign y5960 = ~1'b0 ;
  assign y5961 = ~n12687 ;
  assign y5962 = ~1'b0 ;
  assign y5963 = ~n12690 ;
  assign y5964 = n12692 ;
  assign y5965 = n12697 ;
  assign y5966 = ~n12699 ;
  assign y5967 = n12704 ;
  assign y5968 = ~1'b0 ;
  assign y5969 = n12092 ;
  assign y5970 = ~n12705 ;
  assign y5971 = ~1'b0 ;
  assign y5972 = ~n12706 ;
  assign y5973 = ~n12708 ;
  assign y5974 = ~n12709 ;
  assign y5975 = n12711 ;
  assign y5976 = ~1'b0 ;
  assign y5977 = n12712 ;
  assign y5978 = ~1'b0 ;
  assign y5979 = ~n12716 ;
  assign y5980 = ~n12718 ;
  assign y5981 = ~n12720 ;
  assign y5982 = n12722 ;
  assign y5983 = ~1'b0 ;
  assign y5984 = ~n12725 ;
  assign y5985 = n12730 ;
  assign y5986 = ~1'b0 ;
  assign y5987 = n10094 ;
  assign y5988 = ~n12732 ;
  assign y5989 = ~1'b0 ;
  assign y5990 = n12733 ;
  assign y5991 = ~n12736 ;
  assign y5992 = ~n12741 ;
  assign y5993 = ~n12742 ;
  assign y5994 = n12744 ;
  assign y5995 = 1'b0 ;
  assign y5996 = ~1'b0 ;
  assign y5997 = n4237 ;
  assign y5998 = ~n12745 ;
  assign y5999 = ~1'b0 ;
  assign y6000 = ~n12751 ;
  assign y6001 = ~n12752 ;
  assign y6002 = n12758 ;
  assign y6003 = ~1'b0 ;
  assign y6004 = ~1'b0 ;
  assign y6005 = n12762 ;
  assign y6006 = n12764 ;
  assign y6007 = n12769 ;
  assign y6008 = n12773 ;
  assign y6009 = ~n12775 ;
  assign y6010 = ~1'b0 ;
  assign y6011 = ~n7124 ;
  assign y6012 = n12778 ;
  assign y6013 = n12781 ;
  assign y6014 = ~1'b0 ;
  assign y6015 = n12782 ;
  assign y6016 = n12783 ;
  assign y6017 = n12786 ;
  assign y6018 = ~1'b0 ;
  assign y6019 = ~1'b0 ;
  assign y6020 = n9416 ;
  assign y6021 = ~1'b0 ;
  assign y6022 = n3447 ;
  assign y6023 = ~1'b0 ;
  assign y6024 = ~n12791 ;
  assign y6025 = ~1'b0 ;
  assign y6026 = ~n1793 ;
  assign y6027 = ~n12793 ;
  assign y6028 = ~n12797 ;
  assign y6029 = n12800 ;
  assign y6030 = n12804 ;
  assign y6031 = n2951 ;
  assign y6032 = n12806 ;
  assign y6033 = ~1'b0 ;
  assign y6034 = ~1'b0 ;
  assign y6035 = n3754 ;
  assign y6036 = n12807 ;
  assign y6037 = ~n4621 ;
  assign y6038 = n12810 ;
  assign y6039 = ~n12813 ;
  assign y6040 = n12818 ;
  assign y6041 = n12820 ;
  assign y6042 = ~n12822 ;
  assign y6043 = ~1'b0 ;
  assign y6044 = n12831 ;
  assign y6045 = n12832 ;
  assign y6046 = ~1'b0 ;
  assign y6047 = n12833 ;
  assign y6048 = ~n12836 ;
  assign y6049 = ~1'b0 ;
  assign y6050 = ~1'b0 ;
  assign y6051 = ~n12842 ;
  assign y6052 = ~n12846 ;
  assign y6053 = ~n12850 ;
  assign y6054 = n12853 ;
  assign y6055 = n12854 ;
  assign y6056 = ~n3100 ;
  assign y6057 = n12855 ;
  assign y6058 = ~n10096 ;
  assign y6059 = ~1'b0 ;
  assign y6060 = ~n12859 ;
  assign y6061 = n12862 ;
  assign y6062 = n12863 ;
  assign y6063 = ~n12867 ;
  assign y6064 = ~n12872 ;
  assign y6065 = n12875 ;
  assign y6066 = n12878 ;
  assign y6067 = n12879 ;
  assign y6068 = n12882 ;
  assign y6069 = ~n12884 ;
  assign y6070 = ~1'b0 ;
  assign y6071 = n12885 ;
  assign y6072 = n12890 ;
  assign y6073 = n12892 ;
  assign y6074 = n12897 ;
  assign y6075 = ~1'b0 ;
  assign y6076 = 1'b0 ;
  assign y6077 = ~n12898 ;
  assign y6078 = n12904 ;
  assign y6079 = n12911 ;
  assign y6080 = ~1'b0 ;
  assign y6081 = ~1'b0 ;
  assign y6082 = ~n12913 ;
  assign y6083 = n12919 ;
  assign y6084 = ~1'b0 ;
  assign y6085 = ~1'b0 ;
  assign y6086 = ~n12922 ;
  assign y6087 = n12923 ;
  assign y6088 = ~n12924 ;
  assign y6089 = ~1'b0 ;
  assign y6090 = ~n12928 ;
  assign y6091 = ~1'b0 ;
  assign y6092 = n12929 ;
  assign y6093 = ~n12933 ;
  assign y6094 = n8679 ;
  assign y6095 = ~1'b0 ;
  assign y6096 = ~1'b0 ;
  assign y6097 = ~1'b0 ;
  assign y6098 = n12938 ;
  assign y6099 = ~1'b0 ;
  assign y6100 = ~1'b0 ;
  assign y6101 = ~1'b0 ;
  assign y6102 = n12942 ;
  assign y6103 = ~n12945 ;
  assign y6104 = n12947 ;
  assign y6105 = ~n12952 ;
  assign y6106 = n12966 ;
  assign y6107 = ~n12967 ;
  assign y6108 = ~1'b0 ;
  assign y6109 = ~1'b0 ;
  assign y6110 = n12970 ;
  assign y6111 = n12974 ;
  assign y6112 = ~n12975 ;
  assign y6113 = n12980 ;
  assign y6114 = n12981 ;
  assign y6115 = ~n12983 ;
  assign y6116 = n12984 ;
  assign y6117 = n12991 ;
  assign y6118 = ~1'b0 ;
  assign y6119 = n12995 ;
  assign y6120 = n12996 ;
  assign y6121 = ~n12998 ;
  assign y6122 = ~1'b0 ;
  assign y6123 = ~1'b0 ;
  assign y6124 = ~n13005 ;
  assign y6125 = ~n4770 ;
  assign y6126 = n13008 ;
  assign y6127 = ~n13017 ;
  assign y6128 = ~1'b0 ;
  assign y6129 = n13018 ;
  assign y6130 = ~n12352 ;
  assign y6131 = ~1'b0 ;
  assign y6132 = ~n13019 ;
  assign y6133 = n13022 ;
  assign y6134 = ~n9803 ;
  assign y6135 = n13027 ;
  assign y6136 = n13034 ;
  assign y6137 = ~n13035 ;
  assign y6138 = ~1'b0 ;
  assign y6139 = n13038 ;
  assign y6140 = ~1'b0 ;
  assign y6141 = ~1'b0 ;
  assign y6142 = ~n13039 ;
  assign y6143 = n13041 ;
  assign y6144 = ~n13042 ;
  assign y6145 = 1'b0 ;
  assign y6146 = ~n4585 ;
  assign y6147 = n13044 ;
  assign y6148 = n6572 ;
  assign y6149 = n13048 ;
  assign y6150 = ~n13053 ;
  assign y6151 = ~n13055 ;
  assign y6152 = n13057 ;
  assign y6153 = ~n13060 ;
  assign y6154 = n13063 ;
  assign y6155 = ~n13064 ;
  assign y6156 = ~n13065 ;
  assign y6157 = ~n13070 ;
  assign y6158 = n13075 ;
  assign y6159 = ~n13080 ;
  assign y6160 = n13082 ;
  assign y6161 = ~n13083 ;
  assign y6162 = ~n13085 ;
  assign y6163 = ~1'b0 ;
  assign y6164 = ~1'b0 ;
  assign y6165 = ~n13088 ;
  assign y6166 = ~n13089 ;
  assign y6167 = ~1'b0 ;
  assign y6168 = ~n13090 ;
  assign y6169 = ~1'b0 ;
  assign y6170 = n13096 ;
  assign y6171 = ~1'b0 ;
  assign y6172 = n13097 ;
  assign y6173 = n13100 ;
  assign y6174 = ~n13104 ;
  assign y6175 = n13106 ;
  assign y6176 = n13107 ;
  assign y6177 = ~n13108 ;
  assign y6178 = ~n13111 ;
  assign y6179 = n13114 ;
  assign y6180 = ~1'b0 ;
  assign y6181 = ~n13116 ;
  assign y6182 = n12074 ;
  assign y6183 = 1'b0 ;
  assign y6184 = ~n13118 ;
  assign y6185 = ~1'b0 ;
  assign y6186 = ~1'b0 ;
  assign y6187 = ~1'b0 ;
  assign y6188 = ~1'b0 ;
  assign y6189 = n13119 ;
  assign y6190 = ~n13122 ;
  assign y6191 = ~n13131 ;
  assign y6192 = ~n13133 ;
  assign y6193 = n13136 ;
  assign y6194 = ~n13141 ;
  assign y6195 = ~n13152 ;
  assign y6196 = n13162 ;
  assign y6197 = n13163 ;
  assign y6198 = n13165 ;
  assign y6199 = ~1'b0 ;
  assign y6200 = ~n13167 ;
  assign y6201 = ~n13168 ;
  assign y6202 = ~1'b0 ;
  assign y6203 = n13170 ;
  assign y6204 = n13171 ;
  assign y6205 = ~n8375 ;
  assign y6206 = 1'b0 ;
  assign y6207 = ~n13172 ;
  assign y6208 = n13177 ;
  assign y6209 = ~1'b0 ;
  assign y6210 = n13179 ;
  assign y6211 = ~1'b0 ;
  assign y6212 = ~n13181 ;
  assign y6213 = n13182 ;
  assign y6214 = ~n13187 ;
  assign y6215 = ~n13192 ;
  assign y6216 = n13196 ;
  assign y6217 = ~1'b0 ;
  assign y6218 = n13198 ;
  assign y6219 = ~1'b0 ;
  assign y6220 = ~n13200 ;
  assign y6221 = ~n13207 ;
  assign y6222 = n13211 ;
  assign y6223 = ~n13214 ;
  assign y6224 = n13219 ;
  assign y6225 = ~1'b0 ;
  assign y6226 = ~1'b0 ;
  assign y6227 = n13222 ;
  assign y6228 = n13224 ;
  assign y6229 = ~1'b0 ;
  assign y6230 = n13227 ;
  assign y6231 = n13229 ;
  assign y6232 = ~n13230 ;
  assign y6233 = ~x46 ;
  assign y6234 = n13232 ;
  assign y6235 = n13233 ;
  assign y6236 = n13236 ;
  assign y6237 = ~1'b0 ;
  assign y6238 = n13239 ;
  assign y6239 = ~1'b0 ;
  assign y6240 = 1'b0 ;
  assign y6241 = ~n13244 ;
  assign y6242 = ~n13251 ;
  assign y6243 = n13255 ;
  assign y6244 = ~1'b0 ;
  assign y6245 = n13258 ;
  assign y6246 = ~n13261 ;
  assign y6247 = n13264 ;
  assign y6248 = ~n13266 ;
  assign y6249 = n10520 ;
  assign y6250 = ~n13268 ;
  assign y6251 = n5540 ;
  assign y6252 = ~1'b0 ;
  assign y6253 = n13273 ;
  assign y6254 = n13277 ;
  assign y6255 = ~1'b0 ;
  assign y6256 = n13279 ;
  assign y6257 = ~n12524 ;
  assign y6258 = n13281 ;
  assign y6259 = ~1'b0 ;
  assign y6260 = ~n13283 ;
  assign y6261 = n9511 ;
  assign y6262 = ~n13286 ;
  assign y6263 = ~1'b0 ;
  assign y6264 = ~1'b0 ;
  assign y6265 = ~1'b0 ;
  assign y6266 = n13288 ;
  assign y6267 = n13289 ;
  assign y6268 = n13292 ;
  assign y6269 = n13293 ;
  assign y6270 = ~1'b0 ;
  assign y6271 = ~n7179 ;
  assign y6272 = n13294 ;
  assign y6273 = n13296 ;
  assign y6274 = ~n13299 ;
  assign y6275 = ~n13304 ;
  assign y6276 = ~1'b0 ;
  assign y6277 = ~1'b0 ;
  assign y6278 = ~n5898 ;
  assign y6279 = n13305 ;
  assign y6280 = ~n13312 ;
  assign y6281 = ~n13315 ;
  assign y6282 = ~n13316 ;
  assign y6283 = n13318 ;
  assign y6284 = ~n13319 ;
  assign y6285 = n13320 ;
  assign y6286 = ~n13322 ;
  assign y6287 = ~1'b0 ;
  assign y6288 = ~1'b0 ;
  assign y6289 = ~1'b0 ;
  assign y6290 = ~1'b0 ;
  assign y6291 = n13325 ;
  assign y6292 = n13331 ;
  assign y6293 = ~n13335 ;
  assign y6294 = ~1'b0 ;
  assign y6295 = n13339 ;
  assign y6296 = n13345 ;
  assign y6297 = n13351 ;
  assign y6298 = ~1'b0 ;
  assign y6299 = ~n13352 ;
  assign y6300 = ~n13355 ;
  assign y6301 = ~n13359 ;
  assign y6302 = ~1'b0 ;
  assign y6303 = n13365 ;
  assign y6304 = ~1'b0 ;
  assign y6305 = n13366 ;
  assign y6306 = n13368 ;
  assign y6307 = ~n13375 ;
  assign y6308 = n13378 ;
  assign y6309 = n13379 ;
  assign y6310 = ~n13380 ;
  assign y6311 = ~n13381 ;
  assign y6312 = ~1'b0 ;
  assign y6313 = ~1'b0 ;
  assign y6314 = n13385 ;
  assign y6315 = ~1'b0 ;
  assign y6316 = ~n13391 ;
  assign y6317 = ~n13394 ;
  assign y6318 = ~n13399 ;
  assign y6319 = ~n13402 ;
  assign y6320 = ~1'b0 ;
  assign y6321 = n13404 ;
  assign y6322 = ~1'b0 ;
  assign y6323 = ~n13405 ;
  assign y6324 = n13409 ;
  assign y6325 = n13410 ;
  assign y6326 = n13412 ;
  assign y6327 = ~n13417 ;
  assign y6328 = ~n13423 ;
  assign y6329 = n13431 ;
  assign y6330 = ~n13440 ;
  assign y6331 = n5690 ;
  assign y6332 = ~n13443 ;
  assign y6333 = n13444 ;
  assign y6334 = ~n13452 ;
  assign y6335 = ~n13454 ;
  assign y6336 = ~1'b0 ;
  assign y6337 = ~1'b0 ;
  assign y6338 = ~1'b0 ;
  assign y6339 = n13459 ;
  assign y6340 = n13461 ;
  assign y6341 = ~1'b0 ;
  assign y6342 = ~n13462 ;
  assign y6343 = ~n8899 ;
  assign y6344 = ~1'b0 ;
  assign y6345 = ~n13463 ;
  assign y6346 = ~1'b0 ;
  assign y6347 = ~1'b0 ;
  assign y6348 = ~1'b0 ;
  assign y6349 = ~1'b0 ;
  assign y6350 = n13465 ;
  assign y6351 = ~1'b0 ;
  assign y6352 = ~1'b0 ;
  assign y6353 = n13468 ;
  assign y6354 = 1'b0 ;
  assign y6355 = ~1'b0 ;
  assign y6356 = n13470 ;
  assign y6357 = ~n13474 ;
  assign y6358 = ~n13476 ;
  assign y6359 = ~1'b0 ;
  assign y6360 = ~n13481 ;
  assign y6361 = ~n13485 ;
  assign y6362 = n13487 ;
  assign y6363 = n13491 ;
  assign y6364 = ~n9204 ;
  assign y6365 = ~1'b0 ;
  assign y6366 = n13494 ;
  assign y6367 = n13496 ;
  assign y6368 = n13502 ;
  assign y6369 = ~n13503 ;
  assign y6370 = ~n13504 ;
  assign y6371 = ~1'b0 ;
  assign y6372 = ~n13506 ;
  assign y6373 = ~1'b0 ;
  assign y6374 = n13510 ;
  assign y6375 = ~1'b0 ;
  assign y6376 = n13511 ;
  assign y6377 = ~1'b0 ;
  assign y6378 = n13520 ;
  assign y6379 = ~1'b0 ;
  assign y6380 = ~n13521 ;
  assign y6381 = ~1'b0 ;
  assign y6382 = ~n13523 ;
  assign y6383 = n13524 ;
  assign y6384 = n13525 ;
  assign y6385 = n13527 ;
  assign y6386 = ~1'b0 ;
  assign y6387 = n13528 ;
  assign y6388 = ~1'b0 ;
  assign y6389 = n13529 ;
  assign y6390 = ~n13531 ;
  assign y6391 = ~1'b0 ;
  assign y6392 = n858 ;
  assign y6393 = ~n13532 ;
  assign y6394 = ~1'b0 ;
  assign y6395 = ~n13533 ;
  assign y6396 = ~n13534 ;
  assign y6397 = n13537 ;
  assign y6398 = n13538 ;
  assign y6399 = n13539 ;
  assign y6400 = ~n13541 ;
  assign y6401 = ~n5058 ;
  assign y6402 = ~1'b0 ;
  assign y6403 = n13544 ;
  assign y6404 = ~n13545 ;
  assign y6405 = ~1'b0 ;
  assign y6406 = n13547 ;
  assign y6407 = ~n13550 ;
  assign y6408 = n13555 ;
  assign y6409 = ~1'b0 ;
  assign y6410 = ~1'b0 ;
  assign y6411 = n8607 ;
  assign y6412 = n13558 ;
  assign y6413 = ~1'b0 ;
  assign y6414 = ~1'b0 ;
  assign y6415 = n13567 ;
  assign y6416 = n13569 ;
  assign y6417 = ~n13571 ;
  assign y6418 = ~n13576 ;
  assign y6419 = ~1'b0 ;
  assign y6420 = ~1'b0 ;
  assign y6421 = ~n13578 ;
  assign y6422 = n13585 ;
  assign y6423 = n13592 ;
  assign y6424 = ~n13594 ;
  assign y6425 = ~1'b0 ;
  assign y6426 = ~n13598 ;
  assign y6427 = ~n13601 ;
  assign y6428 = ~n7855 ;
  assign y6429 = n5815 ;
  assign y6430 = ~1'b0 ;
  assign y6431 = ~n13603 ;
  assign y6432 = ~1'b0 ;
  assign y6433 = ~n13604 ;
  assign y6434 = ~1'b0 ;
  assign y6435 = ~1'b0 ;
  assign y6436 = ~n13606 ;
  assign y6437 = n13608 ;
  assign y6438 = n13610 ;
  assign y6439 = ~n13611 ;
  assign y6440 = n13615 ;
  assign y6441 = ~1'b0 ;
  assign y6442 = n13616 ;
  assign y6443 = 1'b0 ;
  assign y6444 = ~n13618 ;
  assign y6445 = ~1'b0 ;
  assign y6446 = ~n13628 ;
  assign y6447 = n13633 ;
  assign y6448 = n13635 ;
  assign y6449 = n13638 ;
  assign y6450 = n13640 ;
  assign y6451 = ~n13647 ;
  assign y6452 = ~n13650 ;
  assign y6453 = ~1'b0 ;
  assign y6454 = ~1'b0 ;
  assign y6455 = ~1'b0 ;
  assign y6456 = ~n13654 ;
  assign y6457 = n13658 ;
  assign y6458 = ~n13661 ;
  assign y6459 = ~1'b0 ;
  assign y6460 = ~1'b0 ;
  assign y6461 = ~n3706 ;
  assign y6462 = ~n13671 ;
  assign y6463 = ~n13673 ;
  assign y6464 = ~n13678 ;
  assign y6465 = ~1'b0 ;
  assign y6466 = ~1'b0 ;
  assign y6467 = ~n13682 ;
  assign y6468 = ~1'b0 ;
  assign y6469 = n13683 ;
  assign y6470 = ~n13685 ;
  assign y6471 = ~n13688 ;
  assign y6472 = n13690 ;
  assign y6473 = n13692 ;
  assign y6474 = ~n13697 ;
  assign y6475 = ~n13700 ;
  assign y6476 = ~n13701 ;
  assign y6477 = ~n13705 ;
  assign y6478 = ~n13706 ;
  assign y6479 = ~n13713 ;
  assign y6480 = n13718 ;
  assign y6481 = n13719 ;
  assign y6482 = ~n13720 ;
  assign y6483 = n13727 ;
  assign y6484 = n13730 ;
  assign y6485 = ~1'b0 ;
  assign y6486 = n13732 ;
  assign y6487 = n13738 ;
  assign y6488 = ~1'b0 ;
  assign y6489 = n13743 ;
  assign y6490 = ~n13745 ;
  assign y6491 = n5237 ;
  assign y6492 = ~1'b0 ;
  assign y6493 = ~1'b0 ;
  assign y6494 = ~1'b0 ;
  assign y6495 = ~n13756 ;
  assign y6496 = ~n13760 ;
  assign y6497 = ~1'b0 ;
  assign y6498 = ~1'b0 ;
  assign y6499 = ~n13762 ;
  assign y6500 = ~1'b0 ;
  assign y6501 = ~1'b0 ;
  assign y6502 = ~1'b0 ;
  assign y6503 = 1'b0 ;
  assign y6504 = n13763 ;
  assign y6505 = ~1'b0 ;
  assign y6506 = ~n13765 ;
  assign y6507 = n13766 ;
  assign y6508 = ~1'b0 ;
  assign y6509 = ~1'b0 ;
  assign y6510 = ~n13767 ;
  assign y6511 = ~n13768 ;
  assign y6512 = ~1'b0 ;
  assign y6513 = ~n13769 ;
  assign y6514 = ~1'b0 ;
  assign y6515 = ~n6879 ;
  assign y6516 = n3349 ;
  assign y6517 = n13777 ;
  assign y6518 = n13778 ;
  assign y6519 = ~1'b0 ;
  assign y6520 = ~1'b0 ;
  assign y6521 = n13780 ;
  assign y6522 = ~1'b0 ;
  assign y6523 = ~1'b0 ;
  assign y6524 = ~1'b0 ;
  assign y6525 = ~1'b0 ;
  assign y6526 = n13781 ;
  assign y6527 = n13782 ;
  assign y6528 = ~1'b0 ;
  assign y6529 = ~1'b0 ;
  assign y6530 = ~1'b0 ;
  assign y6531 = n13783 ;
  assign y6532 = n13787 ;
  assign y6533 = ~n13790 ;
  assign y6534 = ~1'b0 ;
  assign y6535 = n13793 ;
  assign y6536 = ~1'b0 ;
  assign y6537 = ~1'b0 ;
  assign y6538 = n4296 ;
  assign y6539 = ~1'b0 ;
  assign y6540 = ~n13796 ;
  assign y6541 = ~n13800 ;
  assign y6542 = ~1'b0 ;
  assign y6543 = n2387 ;
  assign y6544 = n13801 ;
  assign y6545 = ~n13802 ;
  assign y6546 = ~1'b0 ;
  assign y6547 = n4343 ;
  assign y6548 = n13805 ;
  assign y6549 = n13806 ;
  assign y6550 = n13807 ;
  assign y6551 = 1'b0 ;
  assign y6552 = ~n13808 ;
  assign y6553 = ~n13810 ;
  assign y6554 = ~1'b0 ;
  assign y6555 = ~n13812 ;
  assign y6556 = n13817 ;
  assign y6557 = ~n13607 ;
  assign y6558 = ~n13818 ;
  assign y6559 = ~n13823 ;
  assign y6560 = n13830 ;
  assign y6561 = ~1'b0 ;
  assign y6562 = n13834 ;
  assign y6563 = n13835 ;
  assign y6564 = ~n13836 ;
  assign y6565 = ~n13842 ;
  assign y6566 = ~n13844 ;
  assign y6567 = ~1'b0 ;
  assign y6568 = ~1'b0 ;
  assign y6569 = ~n13848 ;
  assign y6570 = ~1'b0 ;
  assign y6571 = ~n13849 ;
  assign y6572 = n13853 ;
  assign y6573 = ~n13855 ;
  assign y6574 = ~n13857 ;
  assign y6575 = n13860 ;
  assign y6576 = ~n13862 ;
  assign y6577 = ~n13863 ;
  assign y6578 = ~n13867 ;
  assign y6579 = ~1'b0 ;
  assign y6580 = n13869 ;
  assign y6581 = n13870 ;
  assign y6582 = ~n13875 ;
  assign y6583 = n13877 ;
  assign y6584 = 1'b0 ;
  assign y6585 = ~1'b0 ;
  assign y6586 = ~1'b0 ;
  assign y6587 = ~n13880 ;
  assign y6588 = ~1'b0 ;
  assign y6589 = ~n13883 ;
  assign y6590 = ~n13889 ;
  assign y6591 = n13892 ;
  assign y6592 = ~1'b0 ;
  assign y6593 = n13896 ;
  assign y6594 = ~1'b0 ;
  assign y6595 = n13897 ;
  assign y6596 = ~1'b0 ;
  assign y6597 = n13900 ;
  assign y6598 = ~1'b0 ;
  assign y6599 = n13903 ;
  assign y6600 = ~n2881 ;
  assign y6601 = n13906 ;
  assign y6602 = ~1'b0 ;
  assign y6603 = n13911 ;
  assign y6604 = ~1'b0 ;
  assign y6605 = ~1'b0 ;
  assign y6606 = ~1'b0 ;
  assign y6607 = n13912 ;
  assign y6608 = ~1'b0 ;
  assign y6609 = ~n13913 ;
  assign y6610 = ~1'b0 ;
  assign y6611 = ~n13919 ;
  assign y6612 = ~1'b0 ;
  assign y6613 = ~n13922 ;
  assign y6614 = n13923 ;
  assign y6615 = n13926 ;
  assign y6616 = n13931 ;
  assign y6617 = ~1'b0 ;
  assign y6618 = ~n13932 ;
  assign y6619 = ~n13936 ;
  assign y6620 = n13942 ;
  assign y6621 = n13946 ;
  assign y6622 = n13947 ;
  assign y6623 = ~n13951 ;
  assign y6624 = ~1'b0 ;
  assign y6625 = ~n13952 ;
  assign y6626 = n13954 ;
  assign y6627 = ~n13955 ;
  assign y6628 = ~1'b0 ;
  assign y6629 = ~n13957 ;
  assign y6630 = n13960 ;
  assign y6631 = ~1'b0 ;
  assign y6632 = ~n13964 ;
  assign y6633 = n13965 ;
  assign y6634 = n13966 ;
  assign y6635 = ~n13969 ;
  assign y6636 = ~1'b0 ;
  assign y6637 = n13973 ;
  assign y6638 = ~1'b0 ;
  assign y6639 = n13974 ;
  assign y6640 = ~1'b0 ;
  assign y6641 = ~n10111 ;
  assign y6642 = n13975 ;
  assign y6643 = ~1'b0 ;
  assign y6644 = ~n13979 ;
  assign y6645 = n13982 ;
  assign y6646 = ~1'b0 ;
  assign y6647 = n13985 ;
  assign y6648 = n13990 ;
  assign y6649 = ~n13992 ;
  assign y6650 = ~1'b0 ;
  assign y6651 = ~n13995 ;
  assign y6652 = ~1'b0 ;
  assign y6653 = ~1'b0 ;
  assign y6654 = ~n13999 ;
  assign y6655 = ~1'b0 ;
  assign y6656 = ~n14002 ;
  assign y6657 = ~n14003 ;
  assign y6658 = ~n14004 ;
  assign y6659 = n14005 ;
  assign y6660 = ~n14012 ;
  assign y6661 = ~n14014 ;
  assign y6662 = ~n14019 ;
  assign y6663 = ~1'b0 ;
  assign y6664 = ~n14020 ;
  assign y6665 = ~1'b0 ;
  assign y6666 = n14021 ;
  assign y6667 = ~n14022 ;
  assign y6668 = ~1'b0 ;
  assign y6669 = 1'b0 ;
  assign y6670 = ~n14023 ;
  assign y6671 = ~n14032 ;
  assign y6672 = ~n14036 ;
  assign y6673 = n14037 ;
  assign y6674 = ~n14044 ;
  assign y6675 = ~1'b0 ;
  assign y6676 = n14045 ;
  assign y6677 = ~1'b0 ;
  assign y6678 = ~1'b0 ;
  assign y6679 = ~1'b0 ;
  assign y6680 = ~n14048 ;
  assign y6681 = n14049 ;
  assign y6682 = ~n14052 ;
  assign y6683 = n14059 ;
  assign y6684 = n10552 ;
  assign y6685 = n14060 ;
  assign y6686 = n14062 ;
  assign y6687 = ~n10290 ;
  assign y6688 = ~n14063 ;
  assign y6689 = 1'b0 ;
  assign y6690 = ~n14064 ;
  assign y6691 = ~1'b0 ;
  assign y6692 = ~n14070 ;
  assign y6693 = ~n14073 ;
  assign y6694 = ~1'b0 ;
  assign y6695 = ~1'b0 ;
  assign y6696 = ~1'b0 ;
  assign y6697 = ~n14074 ;
  assign y6698 = n14076 ;
  assign y6699 = ~1'b0 ;
  assign y6700 = n14081 ;
  assign y6701 = ~n14083 ;
  assign y6702 = n10724 ;
  assign y6703 = ~1'b0 ;
  assign y6704 = n14084 ;
  assign y6705 = ~n14086 ;
  assign y6706 = n14088 ;
  assign y6707 = n14092 ;
  assign y6708 = n6163 ;
  assign y6709 = ~1'b0 ;
  assign y6710 = ~1'b0 ;
  assign y6711 = ~n14096 ;
  assign y6712 = ~1'b0 ;
  assign y6713 = n14097 ;
  assign y6714 = ~n14098 ;
  assign y6715 = ~1'b0 ;
  assign y6716 = ~1'b0 ;
  assign y6717 = n14104 ;
  assign y6718 = ~1'b0 ;
  assign y6719 = ~n14105 ;
  assign y6720 = n14115 ;
  assign y6721 = ~n14118 ;
  assign y6722 = ~1'b0 ;
  assign y6723 = n14122 ;
  assign y6724 = n7796 ;
  assign y6725 = ~n14124 ;
  assign y6726 = ~n14125 ;
  assign y6727 = n14126 ;
  assign y6728 = n14132 ;
  assign y6729 = ~n14133 ;
  assign y6730 = ~1'b0 ;
  assign y6731 = ~1'b0 ;
  assign y6732 = ~n14138 ;
  assign y6733 = n14139 ;
  assign y6734 = ~n6257 ;
  assign y6735 = ~1'b0 ;
  assign y6736 = n14140 ;
  assign y6737 = ~n4553 ;
  assign y6738 = ~n14142 ;
  assign y6739 = ~1'b0 ;
  assign y6740 = ~n14143 ;
  assign y6741 = ~1'b0 ;
  assign y6742 = n5785 ;
  assign y6743 = n14148 ;
  assign y6744 = ~1'b0 ;
  assign y6745 = ~n14152 ;
  assign y6746 = ~1'b0 ;
  assign y6747 = n14153 ;
  assign y6748 = n14155 ;
  assign y6749 = ~n14156 ;
  assign y6750 = ~n14158 ;
  assign y6751 = ~1'b0 ;
  assign y6752 = ~n14162 ;
  assign y6753 = ~1'b0 ;
  assign y6754 = ~n14164 ;
  assign y6755 = ~1'b0 ;
  assign y6756 = n14166 ;
  assign y6757 = n14168 ;
  assign y6758 = ~1'b0 ;
  assign y6759 = ~1'b0 ;
  assign y6760 = n14170 ;
  assign y6761 = ~n14174 ;
  assign y6762 = ~1'b0 ;
  assign y6763 = n14175 ;
  assign y6764 = ~n14177 ;
  assign y6765 = ~n14178 ;
  assign y6766 = n14179 ;
  assign y6767 = ~1'b0 ;
  assign y6768 = ~1'b0 ;
  assign y6769 = ~1'b0 ;
  assign y6770 = 1'b0 ;
  assign y6771 = n14181 ;
  assign y6772 = ~n14186 ;
  assign y6773 = ~1'b0 ;
  assign y6774 = n14187 ;
  assign y6775 = ~n14191 ;
  assign y6776 = ~1'b0 ;
  assign y6777 = ~1'b0 ;
  assign y6778 = ~1'b0 ;
  assign y6779 = n14192 ;
  assign y6780 = ~1'b0 ;
  assign y6781 = ~n14194 ;
  assign y6782 = ~n14198 ;
  assign y6783 = ~1'b0 ;
  assign y6784 = n14199 ;
  assign y6785 = ~1'b0 ;
  assign y6786 = n14201 ;
  assign y6787 = n14202 ;
  assign y6788 = n14203 ;
  assign y6789 = n14204 ;
  assign y6790 = ~1'b0 ;
  assign y6791 = n14212 ;
  assign y6792 = ~n14213 ;
  assign y6793 = ~n12621 ;
  assign y6794 = ~n14216 ;
  assign y6795 = ~n14220 ;
  assign y6796 = n14227 ;
  assign y6797 = ~1'b0 ;
  assign y6798 = ~1'b0 ;
  assign y6799 = ~1'b0 ;
  assign y6800 = n14228 ;
  assign y6801 = ~n14231 ;
  assign y6802 = ~n14232 ;
  assign y6803 = ~n14239 ;
  assign y6804 = ~1'b0 ;
  assign y6805 = ~n14244 ;
  assign y6806 = n14246 ;
  assign y6807 = ~n14247 ;
  assign y6808 = ~n14252 ;
  assign y6809 = n1153 ;
  assign y6810 = ~1'b0 ;
  assign y6811 = n14253 ;
  assign y6812 = n14254 ;
  assign y6813 = n14258 ;
  assign y6814 = ~n14261 ;
  assign y6815 = ~1'b0 ;
  assign y6816 = ~n14267 ;
  assign y6817 = ~1'b0 ;
  assign y6818 = ~n14269 ;
  assign y6819 = ~1'b0 ;
  assign y6820 = ~n14270 ;
  assign y6821 = ~1'b0 ;
  assign y6822 = ~1'b0 ;
  assign y6823 = ~1'b0 ;
  assign y6824 = ~1'b0 ;
  assign y6825 = ~1'b0 ;
  assign y6826 = ~1'b0 ;
  assign y6827 = ~n14271 ;
  assign y6828 = ~n14272 ;
  assign y6829 = ~n14277 ;
  assign y6830 = ~n14283 ;
  assign y6831 = n14287 ;
  assign y6832 = n14288 ;
  assign y6833 = ~n14291 ;
  assign y6834 = ~1'b0 ;
  assign y6835 = ~n14292 ;
  assign y6836 = n14294 ;
  assign y6837 = n14295 ;
  assign y6838 = ~n14297 ;
  assign y6839 = ~1'b0 ;
  assign y6840 = n13026 ;
  assign y6841 = ~n14301 ;
  assign y6842 = ~1'b0 ;
  assign y6843 = ~1'b0 ;
  assign y6844 = n14302 ;
  assign y6845 = ~n7334 ;
  assign y6846 = ~n14303 ;
  assign y6847 = ~1'b0 ;
  assign y6848 = ~n14307 ;
  assign y6849 = n14308 ;
  assign y6850 = n14310 ;
  assign y6851 = ~1'b0 ;
  assign y6852 = ~n14313 ;
  assign y6853 = n14318 ;
  assign y6854 = n14321 ;
  assign y6855 = ~n4685 ;
  assign y6856 = 1'b0 ;
  assign y6857 = ~1'b0 ;
  assign y6858 = ~1'b0 ;
  assign y6859 = ~n14324 ;
  assign y6860 = ~n14325 ;
  assign y6861 = n14326 ;
  assign y6862 = ~n14327 ;
  assign y6863 = ~1'b0 ;
  assign y6864 = ~1'b0 ;
  assign y6865 = n14330 ;
  assign y6866 = ~n14331 ;
  assign y6867 = ~n14336 ;
  assign y6868 = ~1'b0 ;
  assign y6869 = n14337 ;
  assign y6870 = ~n14339 ;
  assign y6871 = ~1'b0 ;
  assign y6872 = ~1'b0 ;
  assign y6873 = ~n14342 ;
  assign y6874 = ~1'b0 ;
  assign y6875 = n14347 ;
  assign y6876 = ~1'b0 ;
  assign y6877 = n11204 ;
  assign y6878 = n14351 ;
  assign y6879 = ~1'b0 ;
  assign y6880 = ~n14352 ;
  assign y6881 = ~n14355 ;
  assign y6882 = ~n14357 ;
  assign y6883 = n14358 ;
  assign y6884 = n14361 ;
  assign y6885 = ~n14366 ;
  assign y6886 = ~n14371 ;
  assign y6887 = ~n14373 ;
  assign y6888 = n14374 ;
  assign y6889 = n14376 ;
  assign y6890 = ~1'b0 ;
  assign y6891 = ~n2953 ;
  assign y6892 = n14377 ;
  assign y6893 = 1'b0 ;
  assign y6894 = ~1'b0 ;
  assign y6895 = n14387 ;
  assign y6896 = n14396 ;
  assign y6897 = ~1'b0 ;
  assign y6898 = ~n14399 ;
  assign y6899 = ~1'b0 ;
  assign y6900 = ~1'b0 ;
  assign y6901 = n14404 ;
  assign y6902 = ~1'b0 ;
  assign y6903 = n14405 ;
  assign y6904 = ~n14406 ;
  assign y6905 = n14408 ;
  assign y6906 = ~n14410 ;
  assign y6907 = n14415 ;
  assign y6908 = n14417 ;
  assign y6909 = ~n14419 ;
  assign y6910 = n14424 ;
  assign y6911 = ~1'b0 ;
  assign y6912 = 1'b0 ;
  assign y6913 = n14428 ;
  assign y6914 = ~n14430 ;
  assign y6915 = ~n14431 ;
  assign y6916 = ~n14444 ;
  assign y6917 = n14445 ;
  assign y6918 = ~1'b0 ;
  assign y6919 = ~n14447 ;
  assign y6920 = ~1'b0 ;
  assign y6921 = ~1'b0 ;
  assign y6922 = n14449 ;
  assign y6923 = ~1'b0 ;
  assign y6924 = ~n14453 ;
  assign y6925 = ~n14456 ;
  assign y6926 = ~1'b0 ;
  assign y6927 = ~n11655 ;
  assign y6928 = n14459 ;
  assign y6929 = ~n14460 ;
  assign y6930 = ~n14464 ;
  assign y6931 = ~1'b0 ;
  assign y6932 = ~n14469 ;
  assign y6933 = n14473 ;
  assign y6934 = ~n14475 ;
  assign y6935 = ~1'b0 ;
  assign y6936 = n14479 ;
  assign y6937 = ~1'b0 ;
  assign y6938 = ~n14480 ;
  assign y6939 = ~n5371 ;
  assign y6940 = ~1'b0 ;
  assign y6941 = ~n14481 ;
  assign y6942 = ~n4001 ;
  assign y6943 = 1'b0 ;
  assign y6944 = ~1'b0 ;
  assign y6945 = ~n14483 ;
  assign y6946 = ~n14484 ;
  assign y6947 = ~1'b0 ;
  assign y6948 = ~1'b0 ;
  assign y6949 = n14487 ;
  assign y6950 = ~1'b0 ;
  assign y6951 = n5539 ;
  assign y6952 = ~1'b0 ;
  assign y6953 = ~n14490 ;
  assign y6954 = ~n14493 ;
  assign y6955 = ~1'b0 ;
  assign y6956 = ~n14494 ;
  assign y6957 = n1447 ;
  assign y6958 = ~n14497 ;
  assign y6959 = n14500 ;
  assign y6960 = ~n14501 ;
  assign y6961 = ~1'b0 ;
  assign y6962 = ~1'b0 ;
  assign y6963 = ~1'b0 ;
  assign y6964 = ~1'b0 ;
  assign y6965 = ~1'b0 ;
  assign y6966 = ~n14505 ;
  assign y6967 = n14510 ;
  assign y6968 = ~1'b0 ;
  assign y6969 = n14511 ;
  assign y6970 = n14513 ;
  assign y6971 = ~n14518 ;
  assign y6972 = ~1'b0 ;
  assign y6973 = ~n12096 ;
  assign y6974 = ~1'b0 ;
  assign y6975 = ~n14519 ;
  assign y6976 = n14522 ;
  assign y6977 = ~1'b0 ;
  assign y6978 = n14523 ;
  assign y6979 = n14525 ;
  assign y6980 = ~n14529 ;
  assign y6981 = ~1'b0 ;
  assign y6982 = ~n14532 ;
  assign y6983 = ~n14534 ;
  assign y6984 = n1856 ;
  assign y6985 = n14535 ;
  assign y6986 = n14536 ;
  assign y6987 = ~n8785 ;
  assign y6988 = 1'b0 ;
  assign y6989 = ~n11369 ;
  assign y6990 = n6842 ;
  assign y6991 = ~n14537 ;
  assign y6992 = ~n14539 ;
  assign y6993 = ~n14543 ;
  assign y6994 = ~1'b0 ;
  assign y6995 = n14544 ;
  assign y6996 = n14549 ;
  assign y6997 = ~n14551 ;
  assign y6998 = n14555 ;
  assign y6999 = ~1'b0 ;
  assign y7000 = ~n14556 ;
  assign y7001 = ~n14557 ;
  assign y7002 = ~n14576 ;
  assign y7003 = ~1'b0 ;
  assign y7004 = ~1'b0 ;
  assign y7005 = ~n14588 ;
  assign y7006 = ~1'b0 ;
  assign y7007 = ~n14593 ;
  assign y7008 = n14598 ;
  assign y7009 = n14606 ;
  assign y7010 = ~1'b0 ;
  assign y7011 = ~1'b0 ;
  assign y7012 = n14607 ;
  assign y7013 = n14609 ;
  assign y7014 = ~1'b0 ;
  assign y7015 = ~n14612 ;
  assign y7016 = ~n14613 ;
  assign y7017 = n14616 ;
  assign y7018 = ~1'b0 ;
  assign y7019 = n14617 ;
  assign y7020 = ~1'b0 ;
  assign y7021 = n14618 ;
  assign y7022 = n14620 ;
  assign y7023 = ~n14626 ;
  assign y7024 = ~n14628 ;
  assign y7025 = n14631 ;
  assign y7026 = ~1'b0 ;
  assign y7027 = ~n14632 ;
  assign y7028 = n14635 ;
  assign y7029 = ~n14642 ;
  assign y7030 = n14644 ;
  assign y7031 = ~1'b0 ;
  assign y7032 = n14647 ;
  assign y7033 = ~n14649 ;
  assign y7034 = ~n14651 ;
  assign y7035 = n14655 ;
  assign y7036 = n14656 ;
  assign y7037 = ~n14660 ;
  assign y7038 = n14661 ;
  assign y7039 = n14664 ;
  assign y7040 = n14673 ;
  assign y7041 = n14675 ;
  assign y7042 = n11127 ;
  assign y7043 = ~n14679 ;
  assign y7044 = ~1'b0 ;
  assign y7045 = ~n14682 ;
  assign y7046 = ~n14687 ;
  assign y7047 = ~1'b0 ;
  assign y7048 = ~1'b0 ;
  assign y7049 = ~1'b0 ;
  assign y7050 = ~n4968 ;
  assign y7051 = n14688 ;
  assign y7052 = ~1'b0 ;
  assign y7053 = n1862 ;
  assign y7054 = ~1'b0 ;
  assign y7055 = n14692 ;
  assign y7056 = ~1'b0 ;
  assign y7057 = n14695 ;
  assign y7058 = ~1'b0 ;
  assign y7059 = n14696 ;
  assign y7060 = ~1'b0 ;
  assign y7061 = ~1'b0 ;
  assign y7062 = n14697 ;
  assign y7063 = n14698 ;
  assign y7064 = ~n14699 ;
  assign y7065 = n14706 ;
  assign y7066 = n14708 ;
  assign y7067 = ~1'b0 ;
  assign y7068 = ~1'b0 ;
  assign y7069 = ~1'b0 ;
  assign y7070 = n14711 ;
  assign y7071 = ~n14719 ;
  assign y7072 = n14720 ;
  assign y7073 = ~n14722 ;
  assign y7074 = ~1'b0 ;
  assign y7075 = ~n14732 ;
  assign y7076 = ~n14735 ;
  assign y7077 = ~n14740 ;
  assign y7078 = n14741 ;
  assign y7079 = n14744 ;
  assign y7080 = ~1'b0 ;
  assign y7081 = 1'b0 ;
  assign y7082 = ~n14745 ;
  assign y7083 = n14749 ;
  assign y7084 = n14750 ;
  assign y7085 = ~n14752 ;
  assign y7086 = n14760 ;
  assign y7087 = ~n14763 ;
  assign y7088 = ~n14770 ;
  assign y7089 = n14771 ;
  assign y7090 = n14772 ;
  assign y7091 = n14774 ;
  assign y7092 = n14784 ;
  assign y7093 = ~n14785 ;
  assign y7094 = n14796 ;
  assign y7095 = ~n14799 ;
  assign y7096 = ~n14801 ;
  assign y7097 = 1'b0 ;
  assign y7098 = ~n14807 ;
  assign y7099 = ~n14808 ;
  assign y7100 = n14814 ;
  assign y7101 = ~1'b0 ;
  assign y7102 = n14818 ;
  assign y7103 = n14820 ;
  assign y7104 = n14823 ;
  assign y7105 = n7972 ;
  assign y7106 = ~n14827 ;
  assign y7107 = n14836 ;
  assign y7108 = ~n14839 ;
  assign y7109 = ~n14847 ;
  assign y7110 = ~n14852 ;
  assign y7111 = ~1'b0 ;
  assign y7112 = n11605 ;
  assign y7113 = n14854 ;
  assign y7114 = n14855 ;
  assign y7115 = ~n14857 ;
  assign y7116 = ~n14859 ;
  assign y7117 = ~n14861 ;
  assign y7118 = n14864 ;
  assign y7119 = n14866 ;
  assign y7120 = ~1'b0 ;
  assign y7121 = ~1'b0 ;
  assign y7122 = ~1'b0 ;
  assign y7123 = ~n14870 ;
  assign y7124 = 1'b0 ;
  assign y7125 = ~n14872 ;
  assign y7126 = ~n14874 ;
  assign y7127 = n14875 ;
  assign y7128 = n14877 ;
  assign y7129 = ~1'b0 ;
  assign y7130 = ~n14885 ;
  assign y7131 = ~n14886 ;
  assign y7132 = ~1'b0 ;
  assign y7133 = n14889 ;
  assign y7134 = ~1'b0 ;
  assign y7135 = ~n14891 ;
  assign y7136 = ~n9850 ;
  assign y7137 = ~1'b0 ;
  assign y7138 = n14892 ;
  assign y7139 = ~n1633 ;
  assign y7140 = ~1'b0 ;
  assign y7141 = ~n14897 ;
  assign y7142 = ~1'b0 ;
  assign y7143 = n14898 ;
  assign y7144 = ~1'b0 ;
  assign y7145 = ~1'b0 ;
  assign y7146 = n14900 ;
  assign y7147 = ~1'b0 ;
  assign y7148 = ~n14902 ;
  assign y7149 = ~n14906 ;
  assign y7150 = ~1'b0 ;
  assign y7151 = x9 ;
  assign y7152 = ~1'b0 ;
  assign y7153 = n14909 ;
  assign y7154 = ~n14911 ;
  assign y7155 = ~n14913 ;
  assign y7156 = ~n14916 ;
  assign y7157 = n14918 ;
  assign y7158 = ~n14921 ;
  assign y7159 = ~1'b0 ;
  assign y7160 = ~1'b0 ;
  assign y7161 = n14922 ;
  assign y7162 = ~n14927 ;
  assign y7163 = ~n14932 ;
  assign y7164 = ~1'b0 ;
  assign y7165 = n14933 ;
  assign y7166 = ~n14935 ;
  assign y7167 = ~1'b0 ;
  assign y7168 = n14941 ;
  assign y7169 = ~n14946 ;
  assign y7170 = ~n14948 ;
  assign y7171 = n11492 ;
  assign y7172 = ~n14950 ;
  assign y7173 = ~n14954 ;
  assign y7174 = ~n14956 ;
  assign y7175 = ~n14958 ;
  assign y7176 = ~n14963 ;
  assign y7177 = ~n13672 ;
  assign y7178 = n14965 ;
  assign y7179 = ~n2394 ;
  assign y7180 = n14970 ;
  assign y7181 = ~1'b0 ;
  assign y7182 = n14977 ;
  assign y7183 = ~n14978 ;
  assign y7184 = ~1'b0 ;
  assign y7185 = ~n14981 ;
  assign y7186 = n14988 ;
  assign y7187 = ~n14991 ;
  assign y7188 = n14992 ;
  assign y7189 = ~1'b0 ;
  assign y7190 = ~1'b0 ;
  assign y7191 = ~n14993 ;
  assign y7192 = ~n14996 ;
  assign y7193 = ~n14997 ;
  assign y7194 = 1'b0 ;
  assign y7195 = ~n15003 ;
  assign y7196 = ~n15006 ;
  assign y7197 = ~n15014 ;
  assign y7198 = n15017 ;
  assign y7199 = ~n15019 ;
  assign y7200 = n15020 ;
  assign y7201 = n15024 ;
  assign y7202 = ~n15026 ;
  assign y7203 = n15027 ;
  assign y7204 = n15031 ;
  assign y7205 = n15034 ;
  assign y7206 = ~n15035 ;
  assign y7207 = ~n15037 ;
  assign y7208 = ~n15038 ;
  assign y7209 = ~1'b0 ;
  assign y7210 = n15039 ;
  assign y7211 = ~1'b0 ;
  assign y7212 = ~n15044 ;
  assign y7213 = n15046 ;
  assign y7214 = ~1'b0 ;
  assign y7215 = n15048 ;
  assign y7216 = n15049 ;
  assign y7217 = ~n15051 ;
  assign y7218 = n15053 ;
  assign y7219 = n15057 ;
  assign y7220 = ~1'b0 ;
  assign y7221 = ~n15063 ;
  assign y7222 = ~1'b0 ;
  assign y7223 = n15067 ;
  assign y7224 = n15068 ;
  assign y7225 = ~n15073 ;
  assign y7226 = ~1'b0 ;
  assign y7227 = ~n15074 ;
  assign y7228 = ~n15076 ;
  assign y7229 = ~n15079 ;
  assign y7230 = n15082 ;
  assign y7231 = ~n15084 ;
  assign y7232 = n15085 ;
  assign y7233 = n15089 ;
  assign y7234 = ~n15090 ;
  assign y7235 = n15095 ;
  assign y7236 = ~n15100 ;
  assign y7237 = n15101 ;
  assign y7238 = n15106 ;
  assign y7239 = n15109 ;
  assign y7240 = ~n15111 ;
  assign y7241 = ~n15112 ;
  assign y7242 = ~1'b0 ;
  assign y7243 = ~1'b0 ;
  assign y7244 = ~n15113 ;
  assign y7245 = ~n15115 ;
  assign y7246 = ~n15124 ;
  assign y7247 = ~1'b0 ;
  assign y7248 = ~n15126 ;
  assign y7249 = ~1'b0 ;
  assign y7250 = ~n15133 ;
  assign y7251 = ~n15135 ;
  assign y7252 = ~n15137 ;
  assign y7253 = n15139 ;
  assign y7254 = n15140 ;
  assign y7255 = n15141 ;
  assign y7256 = n15143 ;
  assign y7257 = ~n15151 ;
  assign y7258 = ~n15153 ;
  assign y7259 = ~1'b0 ;
  assign y7260 = ~n13800 ;
  assign y7261 = ~n15154 ;
  assign y7262 = ~n15155 ;
  assign y7263 = ~n15158 ;
  assign y7264 = ~n15162 ;
  assign y7265 = ~n15163 ;
  assign y7266 = n15166 ;
  assign y7267 = ~n15169 ;
  assign y7268 = n15171 ;
  assign y7269 = n15173 ;
  assign y7270 = ~n15176 ;
  assign y7271 = n15177 ;
  assign y7272 = n15181 ;
  assign y7273 = 1'b0 ;
  assign y7274 = n15183 ;
  assign y7275 = n15185 ;
  assign y7276 = ~1'b0 ;
  assign y7277 = ~1'b0 ;
  assign y7278 = n15188 ;
  assign y7279 = n15192 ;
  assign y7280 = n2819 ;
  assign y7281 = n15197 ;
  assign y7282 = n15201 ;
  assign y7283 = ~1'b0 ;
  assign y7284 = ~1'b0 ;
  assign y7285 = ~n15202 ;
  assign y7286 = ~n15209 ;
  assign y7287 = ~1'b0 ;
  assign y7288 = 1'b0 ;
  assign y7289 = n15214 ;
  assign y7290 = ~1'b0 ;
  assign y7291 = n15215 ;
  assign y7292 = ~n15216 ;
  assign y7293 = ~n15219 ;
  assign y7294 = ~n15220 ;
  assign y7295 = ~n15221 ;
  assign y7296 = n15224 ;
  assign y7297 = ~n15227 ;
  assign y7298 = ~1'b0 ;
  assign y7299 = ~n15228 ;
  assign y7300 = n11701 ;
  assign y7301 = ~1'b0 ;
  assign y7302 = n15232 ;
  assign y7303 = n15239 ;
  assign y7304 = n6730 ;
  assign y7305 = ~n15241 ;
  assign y7306 = ~1'b0 ;
  assign y7307 = ~1'b0 ;
  assign y7308 = n15245 ;
  assign y7309 = ~1'b0 ;
  assign y7310 = ~1'b0 ;
  assign y7311 = ~1'b0 ;
  assign y7312 = ~n15247 ;
  assign y7313 = ~n15251 ;
  assign y7314 = n15253 ;
  assign y7315 = n15255 ;
  assign y7316 = ~n15256 ;
  assign y7317 = n15257 ;
  assign y7318 = ~n15258 ;
  assign y7319 = ~n15263 ;
  assign y7320 = n15264 ;
  assign y7321 = ~1'b0 ;
  assign y7322 = ~n15266 ;
  assign y7323 = n15269 ;
  assign y7324 = ~1'b0 ;
  assign y7325 = n15271 ;
  assign y7326 = n15273 ;
  assign y7327 = ~1'b0 ;
  assign y7328 = ~1'b0 ;
  assign y7329 = n15276 ;
  assign y7330 = ~1'b0 ;
  assign y7331 = ~n15281 ;
  assign y7332 = ~n15283 ;
  assign y7333 = ~1'b0 ;
  assign y7334 = n15285 ;
  assign y7335 = n15286 ;
  assign y7336 = ~1'b0 ;
  assign y7337 = ~1'b0 ;
  assign y7338 = ~n15288 ;
  assign y7339 = n15292 ;
  assign y7340 = n15294 ;
  assign y7341 = ~n15297 ;
  assign y7342 = ~n15298 ;
  assign y7343 = ~n15301 ;
  assign y7344 = n15304 ;
  assign y7345 = ~n15307 ;
  assign y7346 = n15314 ;
  assign y7347 = ~1'b0 ;
  assign y7348 = 1'b0 ;
  assign y7349 = ~1'b0 ;
  assign y7350 = n15316 ;
  assign y7351 = n15320 ;
  assign y7352 = ~1'b0 ;
  assign y7353 = ~n15322 ;
  assign y7354 = n1402 ;
  assign y7355 = ~1'b0 ;
  assign y7356 = ~n15325 ;
  assign y7357 = ~n15328 ;
  assign y7358 = n15331 ;
  assign y7359 = ~1'b0 ;
  assign y7360 = ~1'b0 ;
  assign y7361 = ~n15332 ;
  assign y7362 = ~1'b0 ;
  assign y7363 = ~1'b0 ;
  assign y7364 = n15333 ;
  assign y7365 = ~1'b0 ;
  assign y7366 = ~1'b0 ;
  assign y7367 = n6629 ;
  assign y7368 = ~n15334 ;
  assign y7369 = ~n15335 ;
  assign y7370 = n15336 ;
  assign y7371 = ~1'b0 ;
  assign y7372 = ~1'b0 ;
  assign y7373 = ~n15342 ;
  assign y7374 = n15343 ;
  assign y7375 = n6857 ;
  assign y7376 = n15346 ;
  assign y7377 = ~1'b0 ;
  assign y7378 = 1'b0 ;
  assign y7379 = n15348 ;
  assign y7380 = ~1'b0 ;
  assign y7381 = ~n15349 ;
  assign y7382 = ~n15353 ;
  assign y7383 = ~1'b0 ;
  assign y7384 = ~1'b0 ;
  assign y7385 = ~1'b0 ;
  assign y7386 = n15354 ;
  assign y7387 = n15356 ;
  assign y7388 = n15360 ;
  assign y7389 = ~1'b0 ;
  assign y7390 = ~1'b0 ;
  assign y7391 = ~n3900 ;
  assign y7392 = n15365 ;
  assign y7393 = ~n15370 ;
  assign y7394 = ~n15372 ;
  assign y7395 = ~n15373 ;
  assign y7396 = ~1'b0 ;
  assign y7397 = ~n15375 ;
  assign y7398 = ~1'b0 ;
  assign y7399 = ~n15377 ;
  assign y7400 = ~1'b0 ;
  assign y7401 = ~n15378 ;
  assign y7402 = ~n15381 ;
  assign y7403 = n15383 ;
  assign y7404 = ~n15385 ;
  assign y7405 = n10731 ;
  assign y7406 = ~n15387 ;
  assign y7407 = ~n15390 ;
  assign y7408 = n13502 ;
  assign y7409 = n15394 ;
  assign y7410 = ~1'b0 ;
  assign y7411 = ~1'b0 ;
  assign y7412 = ~n15395 ;
  assign y7413 = n15399 ;
  assign y7414 = ~1'b0 ;
  assign y7415 = ~1'b0 ;
  assign y7416 = ~n15402 ;
  assign y7417 = ~1'b0 ;
  assign y7418 = ~n15408 ;
  assign y7419 = n15410 ;
  assign y7420 = ~1'b0 ;
  assign y7421 = ~1'b0 ;
  assign y7422 = ~n15414 ;
  assign y7423 = ~1'b0 ;
  assign y7424 = n15417 ;
  assign y7425 = ~1'b0 ;
  assign y7426 = n15420 ;
  assign y7427 = ~1'b0 ;
  assign y7428 = ~n15423 ;
  assign y7429 = ~n15425 ;
  assign y7430 = ~n15428 ;
  assign y7431 = n9872 ;
  assign y7432 = n15430 ;
  assign y7433 = n1428 ;
  assign y7434 = ~1'b0 ;
  assign y7435 = ~1'b0 ;
  assign y7436 = ~n15432 ;
  assign y7437 = n15433 ;
  assign y7438 = ~1'b0 ;
  assign y7439 = ~1'b0 ;
  assign y7440 = ~n15436 ;
  assign y7441 = ~1'b0 ;
  assign y7442 = ~1'b0 ;
  assign y7443 = n15438 ;
  assign y7444 = ~1'b0 ;
  assign y7445 = n15439 ;
  assign y7446 = ~n15441 ;
  assign y7447 = ~n15443 ;
  assign y7448 = ~n9627 ;
  assign y7449 = n15452 ;
  assign y7450 = n15455 ;
  assign y7451 = ~n15461 ;
  assign y7452 = n15464 ;
  assign y7453 = ~1'b0 ;
  assign y7454 = ~n15477 ;
  assign y7455 = ~n15483 ;
  assign y7456 = n15484 ;
  assign y7457 = ~1'b0 ;
  assign y7458 = ~n15485 ;
  assign y7459 = n15487 ;
  assign y7460 = n15492 ;
  assign y7461 = 1'b0 ;
  assign y7462 = n15495 ;
  assign y7463 = ~n15498 ;
  assign y7464 = n15501 ;
  assign y7465 = ~n15502 ;
  assign y7466 = ~n15506 ;
  assign y7467 = ~n15510 ;
  assign y7468 = n15512 ;
  assign y7469 = ~1'b0 ;
  assign y7470 = n15514 ;
  assign y7471 = n15516 ;
  assign y7472 = ~1'b0 ;
  assign y7473 = ~n15520 ;
  assign y7474 = ~n15521 ;
  assign y7475 = ~n15524 ;
  assign y7476 = n15526 ;
  assign y7477 = ~1'b0 ;
  assign y7478 = n15532 ;
  assign y7479 = n15534 ;
  assign y7480 = n15535 ;
  assign y7481 = n15537 ;
  assign y7482 = ~n15538 ;
  assign y7483 = ~n15539 ;
  assign y7484 = ~n15540 ;
  assign y7485 = n15545 ;
  assign y7486 = n15551 ;
  assign y7487 = ~n15555 ;
  assign y7488 = ~1'b0 ;
  assign y7489 = ~1'b0 ;
  assign y7490 = ~1'b0 ;
  assign y7491 = ~1'b0 ;
  assign y7492 = n3397 ;
  assign y7493 = ~n15559 ;
  assign y7494 = ~1'b0 ;
  assign y7495 = n15561 ;
  assign y7496 = n15563 ;
  assign y7497 = ~1'b0 ;
  assign y7498 = ~n15568 ;
  assign y7499 = ~n15570 ;
  assign y7500 = ~n15571 ;
  assign y7501 = ~n15573 ;
  assign y7502 = n15574 ;
  assign y7503 = ~1'b0 ;
  assign y7504 = n15577 ;
  assign y7505 = ~n15578 ;
  assign y7506 = 1'b0 ;
  assign y7507 = ~1'b0 ;
  assign y7508 = ~n15582 ;
  assign y7509 = ~1'b0 ;
  assign y7510 = ~n10057 ;
  assign y7511 = ~1'b0 ;
  assign y7512 = n15593 ;
  assign y7513 = ~1'b0 ;
  assign y7514 = ~n15596 ;
  assign y7515 = n15603 ;
  assign y7516 = ~n15611 ;
  assign y7517 = n15615 ;
  assign y7518 = ~n15616 ;
  assign y7519 = n15617 ;
  assign y7520 = ~1'b0 ;
  assign y7521 = n15619 ;
  assign y7522 = ~1'b0 ;
  assign y7523 = ~1'b0 ;
  assign y7524 = n3457 ;
  assign y7525 = ~n15624 ;
  assign y7526 = ~1'b0 ;
  assign y7527 = ~1'b0 ;
  assign y7528 = n15627 ;
  assign y7529 = n15629 ;
  assign y7530 = ~n15630 ;
  assign y7531 = ~n15633 ;
  assign y7532 = ~n15637 ;
  assign y7533 = ~1'b0 ;
  assign y7534 = ~1'b0 ;
  assign y7535 = ~1'b0 ;
  assign y7536 = n15639 ;
  assign y7537 = 1'b0 ;
  assign y7538 = ~n15640 ;
  assign y7539 = ~1'b0 ;
  assign y7540 = ~1'b0 ;
  assign y7541 = n15641 ;
  assign y7542 = 1'b0 ;
  assign y7543 = n15653 ;
  assign y7544 = ~x39 ;
  assign y7545 = n15658 ;
  assign y7546 = n15659 ;
  assign y7547 = ~n15662 ;
  assign y7548 = ~n15666 ;
  assign y7549 = n11497 ;
  assign y7550 = n15671 ;
  assign y7551 = n15672 ;
  assign y7552 = ~1'b0 ;
  assign y7553 = ~n5925 ;
  assign y7554 = ~n15678 ;
  assign y7555 = ~n15683 ;
  assign y7556 = ~1'b0 ;
  assign y7557 = n15684 ;
  assign y7558 = ~1'b0 ;
  assign y7559 = ~1'b0 ;
  assign y7560 = ~1'b0 ;
  assign y7561 = n15686 ;
  assign y7562 = ~1'b0 ;
  assign y7563 = ~n15687 ;
  assign y7564 = ~1'b0 ;
  assign y7565 = ~1'b0 ;
  assign y7566 = ~1'b0 ;
  assign y7567 = ~1'b0 ;
  assign y7568 = n15688 ;
  assign y7569 = ~n15691 ;
  assign y7570 = n15694 ;
  assign y7571 = ~1'b0 ;
  assign y7572 = ~1'b0 ;
  assign y7573 = n15697 ;
  assign y7574 = n15698 ;
  assign y7575 = ~n15700 ;
  assign y7576 = ~n3152 ;
  assign y7577 = n15701 ;
  assign y7578 = n15708 ;
  assign y7579 = ~1'b0 ;
  assign y7580 = n15709 ;
  assign y7581 = n15714 ;
  assign y7582 = n15715 ;
  assign y7583 = ~n15716 ;
  assign y7584 = ~n15718 ;
  assign y7585 = ~1'b0 ;
  assign y7586 = n15722 ;
  assign y7587 = ~1'b0 ;
  assign y7588 = ~1'b0 ;
  assign y7589 = ~1'b0 ;
  assign y7590 = ~n15729 ;
  assign y7591 = n15730 ;
  assign y7592 = ~1'b0 ;
  assign y7593 = n663 ;
  assign y7594 = ~1'b0 ;
  assign y7595 = ~1'b0 ;
  assign y7596 = n15732 ;
  assign y7597 = ~n15735 ;
  assign y7598 = ~1'b0 ;
  assign y7599 = ~n15743 ;
  assign y7600 = n15749 ;
  assign y7601 = ~1'b0 ;
  assign y7602 = ~n15750 ;
  assign y7603 = ~n15754 ;
  assign y7604 = n15756 ;
  assign y7605 = ~1'b0 ;
  assign y7606 = ~n15758 ;
  assign y7607 = ~n15761 ;
  assign y7608 = ~1'b0 ;
  assign y7609 = ~n15763 ;
  assign y7610 = ~1'b0 ;
  assign y7611 = n15765 ;
  assign y7612 = ~n15766 ;
  assign y7613 = n15772 ;
  assign y7614 = n15774 ;
  assign y7615 = ~1'b0 ;
  assign y7616 = ~1'b0 ;
  assign y7617 = n15787 ;
  assign y7618 = ~n15792 ;
  assign y7619 = n15793 ;
  assign y7620 = ~1'b0 ;
  assign y7621 = ~n5579 ;
  assign y7622 = ~1'b0 ;
  assign y7623 = ~1'b0 ;
  assign y7624 = ~n15797 ;
  assign y7625 = ~1'b0 ;
  assign y7626 = ~1'b0 ;
  assign y7627 = ~1'b0 ;
  assign y7628 = ~1'b0 ;
  assign y7629 = ~1'b0 ;
  assign y7630 = n15799 ;
  assign y7631 = ~1'b0 ;
  assign y7632 = ~n15803 ;
  assign y7633 = n15811 ;
  assign y7634 = n15812 ;
  assign y7635 = n15814 ;
  assign y7636 = n15818 ;
  assign y7637 = ~1'b0 ;
  assign y7638 = ~n15820 ;
  assign y7639 = n15825 ;
  assign y7640 = 1'b0 ;
  assign y7641 = ~1'b0 ;
  assign y7642 = ~n15826 ;
  assign y7643 = ~1'b0 ;
  assign y7644 = ~n15830 ;
  assign y7645 = ~n15832 ;
  assign y7646 = ~1'b0 ;
  assign y7647 = ~1'b0 ;
  assign y7648 = ~n15837 ;
  assign y7649 = ~n6805 ;
  assign y7650 = n15839 ;
  assign y7651 = ~n15841 ;
  assign y7652 = n15842 ;
  assign y7653 = n15843 ;
  assign y7654 = ~n15849 ;
  assign y7655 = ~1'b0 ;
  assign y7656 = ~1'b0 ;
  assign y7657 = n15857 ;
  assign y7658 = ~1'b0 ;
  assign y7659 = ~n10529 ;
  assign y7660 = n15858 ;
  assign y7661 = n15865 ;
  assign y7662 = ~1'b0 ;
  assign y7663 = ~1'b0 ;
  assign y7664 = n15867 ;
  assign y7665 = ~1'b0 ;
  assign y7666 = ~n15872 ;
  assign y7667 = 1'b0 ;
  assign y7668 = ~n15874 ;
  assign y7669 = n12338 ;
  assign y7670 = ~n9753 ;
  assign y7671 = n15875 ;
  assign y7672 = ~1'b0 ;
  assign y7673 = ~1'b0 ;
  assign y7674 = ~n15878 ;
  assign y7675 = ~n15880 ;
  assign y7676 = ~n15881 ;
  assign y7677 = n15882 ;
  assign y7678 = ~n15883 ;
  assign y7679 = ~n15887 ;
  assign y7680 = ~n15891 ;
  assign y7681 = n15892 ;
  assign y7682 = n15893 ;
  assign y7683 = n15894 ;
  assign y7684 = ~n15909 ;
  assign y7685 = ~n15911 ;
  assign y7686 = ~n14533 ;
  assign y7687 = ~1'b0 ;
  assign y7688 = ~n15914 ;
  assign y7689 = ~n15916 ;
  assign y7690 = ~n15921 ;
  assign y7691 = n15923 ;
  assign y7692 = n15924 ;
  assign y7693 = ~n15926 ;
  assign y7694 = ~1'b0 ;
  assign y7695 = ~n15927 ;
  assign y7696 = ~1'b0 ;
  assign y7697 = n15931 ;
  assign y7698 = n15943 ;
  assign y7699 = ~n15945 ;
  assign y7700 = ~n15950 ;
  assign y7701 = ~n15953 ;
  assign y7702 = ~1'b0 ;
  assign y7703 = ~n15954 ;
  assign y7704 = ~n15955 ;
  assign y7705 = n15956 ;
  assign y7706 = n15957 ;
  assign y7707 = n15958 ;
  assign y7708 = ~1'b0 ;
  assign y7709 = n15960 ;
  assign y7710 = ~n15964 ;
  assign y7711 = ~1'b0 ;
  assign y7712 = ~n15967 ;
  assign y7713 = n6979 ;
  assign y7714 = ~1'b0 ;
  assign y7715 = n15970 ;
  assign y7716 = n15973 ;
  assign y7717 = n15975 ;
  assign y7718 = 1'b0 ;
  assign y7719 = ~n15981 ;
  assign y7720 = ~1'b0 ;
  assign y7721 = n15983 ;
  assign y7722 = ~1'b0 ;
  assign y7723 = ~1'b0 ;
  assign y7724 = n15992 ;
  assign y7725 = n1008 ;
  assign y7726 = n15993 ;
  assign y7727 = n15998 ;
  assign y7728 = ~n15347 ;
  assign y7729 = ~n15999 ;
  assign y7730 = n16001 ;
  assign y7731 = n16006 ;
  assign y7732 = ~n16014 ;
  assign y7733 = n16015 ;
  assign y7734 = ~n16016 ;
  assign y7735 = ~n16017 ;
  assign y7736 = ~1'b0 ;
  assign y7737 = ~1'b0 ;
  assign y7738 = n16018 ;
  assign y7739 = 1'b0 ;
  assign y7740 = ~n2263 ;
  assign y7741 = ~n16033 ;
  assign y7742 = ~n15557 ;
  assign y7743 = ~n16037 ;
  assign y7744 = ~n16045 ;
  assign y7745 = ~n16047 ;
  assign y7746 = n16026 ;
  assign y7747 = n16049 ;
  assign y7748 = n16057 ;
  assign y7749 = n16062 ;
  assign y7750 = ~1'b0 ;
  assign y7751 = n16070 ;
  assign y7752 = ~1'b0 ;
  assign y7753 = ~n16071 ;
  assign y7754 = ~n16077 ;
  assign y7755 = n16078 ;
  assign y7756 = ~n13239 ;
  assign y7757 = ~n16079 ;
  assign y7758 = ~n16082 ;
  assign y7759 = ~n15809 ;
  assign y7760 = ~n16090 ;
  assign y7761 = ~n16093 ;
  assign y7762 = ~n16096 ;
  assign y7763 = ~1'b0 ;
  assign y7764 = n16098 ;
  assign y7765 = n16101 ;
  assign y7766 = ~n16102 ;
  assign y7767 = n10721 ;
  assign y7768 = ~1'b0 ;
  assign y7769 = n16106 ;
  assign y7770 = ~1'b0 ;
  assign y7771 = ~1'b0 ;
  assign y7772 = n16109 ;
  assign y7773 = n16112 ;
  assign y7774 = n16116 ;
  assign y7775 = n16122 ;
  assign y7776 = ~1'b0 ;
  assign y7777 = ~n16125 ;
  assign y7778 = n16126 ;
  assign y7779 = ~1'b0 ;
  assign y7780 = n16131 ;
  assign y7781 = ~n16132 ;
  assign y7782 = ~n16134 ;
  assign y7783 = n16138 ;
  assign y7784 = n12854 ;
  assign y7785 = ~1'b0 ;
  assign y7786 = ~1'b0 ;
  assign y7787 = n1042 ;
  assign y7788 = n15880 ;
  assign y7789 = ~1'b0 ;
  assign y7790 = n16139 ;
  assign y7791 = n16141 ;
  assign y7792 = ~1'b0 ;
  assign y7793 = ~n16142 ;
  assign y7794 = n16146 ;
  assign y7795 = ~n16148 ;
  assign y7796 = ~n16149 ;
  assign y7797 = ~n16152 ;
  assign y7798 = ~n16154 ;
  assign y7799 = ~1'b0 ;
  assign y7800 = n16156 ;
  assign y7801 = ~1'b0 ;
  assign y7802 = ~1'b0 ;
  assign y7803 = ~1'b0 ;
  assign y7804 = n16158 ;
  assign y7805 = ~1'b0 ;
  assign y7806 = ~n16160 ;
  assign y7807 = ~1'b0 ;
  assign y7808 = n16162 ;
  assign y7809 = n16164 ;
  assign y7810 = ~1'b0 ;
  assign y7811 = 1'b0 ;
  assign y7812 = 1'b0 ;
  assign y7813 = ~1'b0 ;
  assign y7814 = ~1'b0 ;
  assign y7815 = n16165 ;
  assign y7816 = ~n16167 ;
  assign y7817 = n16168 ;
  assign y7818 = ~n16170 ;
  assign y7819 = ~n16171 ;
  assign y7820 = n16172 ;
  assign y7821 = 1'b0 ;
  assign y7822 = ~n16178 ;
  assign y7823 = ~1'b0 ;
  assign y7824 = n16180 ;
  assign y7825 = ~n16181 ;
  assign y7826 = n16183 ;
  assign y7827 = ~n16184 ;
  assign y7828 = ~n16185 ;
  assign y7829 = ~n16187 ;
  assign y7830 = n16196 ;
  assign y7831 = n16198 ;
  assign y7832 = n16200 ;
  assign y7833 = n16208 ;
  assign y7834 = ~1'b0 ;
  assign y7835 = ~1'b0 ;
  assign y7836 = ~1'b0 ;
  assign y7837 = n16209 ;
  assign y7838 = ~n16213 ;
  assign y7839 = n16215 ;
  assign y7840 = ~n16216 ;
  assign y7841 = ~n16223 ;
  assign y7842 = ~1'b0 ;
  assign y7843 = ~n16228 ;
  assign y7844 = ~n16230 ;
  assign y7845 = ~n16233 ;
  assign y7846 = ~1'b0 ;
  assign y7847 = ~1'b0 ;
  assign y7848 = n16236 ;
  assign y7849 = ~n16241 ;
  assign y7850 = ~n16244 ;
  assign y7851 = n16247 ;
  assign y7852 = ~1'b0 ;
  assign y7853 = n16248 ;
  assign y7854 = ~n16252 ;
  assign y7855 = n4309 ;
  assign y7856 = ~n13725 ;
  assign y7857 = ~n16254 ;
  assign y7858 = n16260 ;
  assign y7859 = ~n16266 ;
  assign y7860 = ~n16269 ;
  assign y7861 = ~1'b0 ;
  assign y7862 = ~1'b0 ;
  assign y7863 = ~1'b0 ;
  assign y7864 = ~n16275 ;
  assign y7865 = ~1'b0 ;
  assign y7866 = ~1'b0 ;
  assign y7867 = ~1'b0 ;
  assign y7868 = n16276 ;
  assign y7869 = ~1'b0 ;
  assign y7870 = ~n16277 ;
  assign y7871 = ~n16280 ;
  assign y7872 = ~n16281 ;
  assign y7873 = n16283 ;
  assign y7874 = n16284 ;
  assign y7875 = n16286 ;
  assign y7876 = n16295 ;
  assign y7877 = ~1'b0 ;
  assign y7878 = n16297 ;
  assign y7879 = ~1'b0 ;
  assign y7880 = n16299 ;
  assign y7881 = ~1'b0 ;
  assign y7882 = 1'b0 ;
  assign y7883 = ~n16300 ;
  assign y7884 = ~n16301 ;
  assign y7885 = ~1'b0 ;
  assign y7886 = ~1'b0 ;
  assign y7887 = n16304 ;
  assign y7888 = n16305 ;
  assign y7889 = ~1'b0 ;
  assign y7890 = n16308 ;
  assign y7891 = ~1'b0 ;
  assign y7892 = n16309 ;
  assign y7893 = ~1'b0 ;
  assign y7894 = ~n16311 ;
  assign y7895 = ~n16313 ;
  assign y7896 = ~n16319 ;
  assign y7897 = ~n16320 ;
  assign y7898 = ~n16321 ;
  assign y7899 = n16322 ;
  assign y7900 = n16324 ;
  assign y7901 = ~1'b0 ;
  assign y7902 = n16326 ;
  assign y7903 = ~1'b0 ;
  assign y7904 = ~1'b0 ;
  assign y7905 = ~n16327 ;
  assign y7906 = n16329 ;
  assign y7907 = ~n7359 ;
  assign y7908 = n16332 ;
  assign y7909 = ~1'b0 ;
  assign y7910 = n16334 ;
  assign y7911 = ~1'b0 ;
  assign y7912 = n16341 ;
  assign y7913 = n16342 ;
  assign y7914 = ~n16343 ;
  assign y7915 = n7241 ;
  assign y7916 = ~1'b0 ;
  assign y7917 = ~n16344 ;
  assign y7918 = ~n16355 ;
  assign y7919 = ~1'b0 ;
  assign y7920 = n16356 ;
  assign y7921 = ~n16361 ;
  assign y7922 = ~n16362 ;
  assign y7923 = n16366 ;
  assign y7924 = ~n14647 ;
  assign y7925 = n16368 ;
  assign y7926 = ~n6818 ;
  assign y7927 = ~n16371 ;
  assign y7928 = ~n16372 ;
  assign y7929 = 1'b0 ;
  assign y7930 = ~1'b0 ;
  assign y7931 = ~n16373 ;
  assign y7932 = n16375 ;
  assign y7933 = ~n16379 ;
  assign y7934 = ~1'b0 ;
  assign y7935 = ~n16380 ;
  assign y7936 = n16386 ;
  assign y7937 = ~n16388 ;
  assign y7938 = ~1'b0 ;
  assign y7939 = ~n16390 ;
  assign y7940 = ~1'b0 ;
  assign y7941 = ~n16393 ;
  assign y7942 = n16395 ;
  assign y7943 = ~1'b0 ;
  assign y7944 = ~1'b0 ;
  assign y7945 = ~n16401 ;
  assign y7946 = ~1'b0 ;
  assign y7947 = ~n11863 ;
  assign y7948 = 1'b0 ;
  assign y7949 = n16403 ;
  assign y7950 = ~n11002 ;
  assign y7951 = n16404 ;
  assign y7952 = 1'b0 ;
  assign y7953 = n16407 ;
  assign y7954 = n16412 ;
  assign y7955 = ~1'b0 ;
  assign y7956 = n16416 ;
  assign y7957 = n16419 ;
  assign y7958 = ~1'b0 ;
  assign y7959 = ~1'b0 ;
  assign y7960 = ~1'b0 ;
  assign y7961 = n16420 ;
  assign y7962 = ~n16421 ;
  assign y7963 = n16423 ;
  assign y7964 = n16425 ;
  assign y7965 = ~n9028 ;
  assign y7966 = n16430 ;
  assign y7967 = n14905 ;
  assign y7968 = ~1'b0 ;
  assign y7969 = n16435 ;
  assign y7970 = ~n16436 ;
  assign y7971 = ~n16440 ;
  assign y7972 = n16442 ;
  assign y7973 = n16445 ;
  assign y7974 = ~1'b0 ;
  assign y7975 = ~1'b0 ;
  assign y7976 = n16447 ;
  assign y7977 = ~n16450 ;
  assign y7978 = n16453 ;
  assign y7979 = ~1'b0 ;
  assign y7980 = ~n16455 ;
  assign y7981 = ~1'b0 ;
  assign y7982 = n16456 ;
  assign y7983 = ~n16457 ;
  assign y7984 = n16460 ;
  assign y7985 = ~1'b0 ;
  assign y7986 = ~n16463 ;
  assign y7987 = ~n16466 ;
  assign y7988 = n14794 ;
  assign y7989 = n16474 ;
  assign y7990 = ~1'b0 ;
  assign y7991 = n16475 ;
  assign y7992 = n16477 ;
  assign y7993 = ~n16478 ;
  assign y7994 = ~1'b0 ;
  assign y7995 = ~n16479 ;
  assign y7996 = ~n16486 ;
  assign y7997 = n16490 ;
  assign y7998 = ~1'b0 ;
  assign y7999 = ~1'b0 ;
  assign y8000 = ~1'b0 ;
  assign y8001 = ~n16492 ;
  assign y8002 = n16493 ;
  assign y8003 = n16494 ;
  assign y8004 = ~1'b0 ;
  assign y8005 = ~n4723 ;
  assign y8006 = ~1'b0 ;
  assign y8007 = 1'b0 ;
  assign y8008 = ~n16497 ;
  assign y8009 = n16500 ;
  assign y8010 = n16505 ;
  assign y8011 = n16509 ;
  assign y8012 = n16511 ;
  assign y8013 = ~n16517 ;
  assign y8014 = n16522 ;
  assign y8015 = ~1'b0 ;
  assign y8016 = n16525 ;
  assign y8017 = ~n16528 ;
  assign y8018 = n6179 ;
  assign y8019 = ~n16531 ;
  assign y8020 = ~1'b0 ;
  assign y8021 = n16537 ;
  assign y8022 = ~n16539 ;
  assign y8023 = n14109 ;
  assign y8024 = ~n16540 ;
  assign y8025 = ~n16542 ;
  assign y8026 = n16549 ;
  assign y8027 = ~n16564 ;
  assign y8028 = n16567 ;
  assign y8029 = ~n16568 ;
  assign y8030 = ~n16573 ;
  assign y8031 = ~n16578 ;
  assign y8032 = ~n8545 ;
  assign y8033 = ~1'b0 ;
  assign y8034 = n16584 ;
  assign y8035 = ~n16586 ;
  assign y8036 = ~n16588 ;
  assign y8037 = ~n16590 ;
  assign y8038 = ~1'b0 ;
  assign y8039 = ~n16592 ;
  assign y8040 = ~n16593 ;
  assign y8041 = ~n16595 ;
  assign y8042 = n16597 ;
  assign y8043 = n16600 ;
  assign y8044 = ~1'b0 ;
  assign y8045 = 1'b0 ;
  assign y8046 = n16604 ;
  assign y8047 = n16608 ;
  assign y8048 = n16609 ;
  assign y8049 = ~1'b0 ;
  assign y8050 = n16610 ;
  assign y8051 = n16613 ;
  assign y8052 = ~1'b0 ;
  assign y8053 = ~1'b0 ;
  assign y8054 = ~1'b0 ;
  assign y8055 = ~n16614 ;
  assign y8056 = ~n16615 ;
  assign y8057 = ~n16618 ;
  assign y8058 = ~n16621 ;
  assign y8059 = ~1'b0 ;
  assign y8060 = ~1'b0 ;
  assign y8061 = n16622 ;
  assign y8062 = n16623 ;
  assign y8063 = ~n16627 ;
  assign y8064 = ~n16630 ;
  assign y8065 = ~n16632 ;
  assign y8066 = ~n16634 ;
  assign y8067 = n16637 ;
  assign y8068 = n16638 ;
  assign y8069 = n16642 ;
  assign y8070 = ~n16645 ;
  assign y8071 = ~n16653 ;
  assign y8072 = n16655 ;
  assign y8073 = ~n16661 ;
  assign y8074 = ~1'b0 ;
  assign y8075 = ~n16662 ;
  assign y8076 = ~n16664 ;
  assign y8077 = ~n16669 ;
  assign y8078 = n16670 ;
  assign y8079 = ~1'b0 ;
  assign y8080 = ~n16672 ;
  assign y8081 = ~1'b0 ;
  assign y8082 = ~n16673 ;
  assign y8083 = n16678 ;
  assign y8084 = ~n16681 ;
  assign y8085 = n16683 ;
  assign y8086 = ~n886 ;
  assign y8087 = ~1'b0 ;
  assign y8088 = ~1'b0 ;
  assign y8089 = ~n16685 ;
  assign y8090 = n16688 ;
  assign y8091 = ~1'b0 ;
  assign y8092 = ~1'b0 ;
  assign y8093 = n16691 ;
  assign y8094 = ~1'b0 ;
  assign y8095 = n16693 ;
  assign y8096 = ~1'b0 ;
  assign y8097 = ~n3286 ;
  assign y8098 = ~n16695 ;
  assign y8099 = ~n16699 ;
  assign y8100 = n16700 ;
  assign y8101 = ~1'b0 ;
  assign y8102 = n16705 ;
  assign y8103 = ~n16707 ;
  assign y8104 = n16708 ;
  assign y8105 = ~n16716 ;
  assign y8106 = ~n16718 ;
  assign y8107 = n425 ;
  assign y8108 = n16719 ;
  assign y8109 = ~1'b0 ;
  assign y8110 = 1'b0 ;
  assign y8111 = n3189 ;
  assign y8112 = ~1'b0 ;
  assign y8113 = n16723 ;
  assign y8114 = ~n16724 ;
  assign y8115 = ~n16727 ;
  assign y8116 = n16739 ;
  assign y8117 = ~n16740 ;
  assign y8118 = 1'b0 ;
  assign y8119 = ~n16743 ;
  assign y8120 = ~1'b0 ;
  assign y8121 = ~1'b0 ;
  assign y8122 = ~n16747 ;
  assign y8123 = ~n16749 ;
  assign y8124 = ~1'b0 ;
  assign y8125 = n16751 ;
  assign y8126 = n16759 ;
  assign y8127 = n16760 ;
  assign y8128 = n16767 ;
  assign y8129 = ~n16770 ;
  assign y8130 = ~n16777 ;
  assign y8131 = ~1'b0 ;
  assign y8132 = 1'b0 ;
  assign y8133 = ~n16779 ;
  assign y8134 = ~1'b0 ;
  assign y8135 = ~n16780 ;
  assign y8136 = ~1'b0 ;
  assign y8137 = ~n16783 ;
  assign y8138 = ~n16784 ;
  assign y8139 = ~1'b0 ;
  assign y8140 = ~n16790 ;
  assign y8141 = n16791 ;
  assign y8142 = ~n16792 ;
  assign y8143 = ~1'b0 ;
  assign y8144 = n16795 ;
  assign y8145 = ~n16797 ;
  assign y8146 = ~n16800 ;
  assign y8147 = ~n16803 ;
  assign y8148 = n16809 ;
  assign y8149 = 1'b0 ;
  assign y8150 = ~n16810 ;
  assign y8151 = ~1'b0 ;
  assign y8152 = ~1'b0 ;
  assign y8153 = ~1'b0 ;
  assign y8154 = n16812 ;
  assign y8155 = n15932 ;
  assign y8156 = ~1'b0 ;
  assign y8157 = ~n16813 ;
  assign y8158 = n16817 ;
  assign y8159 = ~n16819 ;
  assign y8160 = ~n16820 ;
  assign y8161 = ~1'b0 ;
  assign y8162 = ~1'b0 ;
  assign y8163 = ~1'b0 ;
  assign y8164 = ~1'b0 ;
  assign y8165 = ~1'b0 ;
  assign y8166 = n5704 ;
  assign y8167 = n16824 ;
  assign y8168 = n16826 ;
  assign y8169 = n16830 ;
  assign y8170 = ~n16832 ;
  assign y8171 = n16836 ;
  assign y8172 = n16837 ;
  assign y8173 = n16838 ;
  assign y8174 = 1'b0 ;
  assign y8175 = n10738 ;
  assign y8176 = ~1'b0 ;
  assign y8177 = ~n16842 ;
  assign y8178 = 1'b0 ;
  assign y8179 = ~n6965 ;
  assign y8180 = n16848 ;
  assign y8181 = n16855 ;
  assign y8182 = ~n16858 ;
  assign y8183 = n16864 ;
  assign y8184 = ~1'b0 ;
  assign y8185 = ~1'b0 ;
  assign y8186 = ~n16865 ;
  assign y8187 = n16866 ;
  assign y8188 = ~1'b0 ;
  assign y8189 = ~n16868 ;
  assign y8190 = ~1'b0 ;
  assign y8191 = n16870 ;
  assign y8192 = n1692 ;
  assign y8193 = ~n16873 ;
  assign y8194 = ~n16874 ;
  assign y8195 = ~1'b0 ;
  assign y8196 = ~1'b0 ;
  assign y8197 = n16875 ;
  assign y8198 = n16878 ;
  assign y8199 = ~1'b0 ;
  assign y8200 = n9053 ;
  assign y8201 = n16884 ;
  assign y8202 = ~1'b0 ;
  assign y8203 = n16886 ;
  assign y8204 = n16887 ;
  assign y8205 = ~n16888 ;
  assign y8206 = ~1'b0 ;
  assign y8207 = n16893 ;
  assign y8208 = n16895 ;
  assign y8209 = ~n16897 ;
  assign y8210 = ~n16900 ;
  assign y8211 = n16905 ;
  assign y8212 = ~n16907 ;
  assign y8213 = ~n3513 ;
  assign y8214 = ~n16911 ;
  assign y8215 = ~n16912 ;
  assign y8216 = ~1'b0 ;
  assign y8217 = n16913 ;
  assign y8218 = ~n16919 ;
  assign y8219 = ~1'b0 ;
  assign y8220 = ~n16921 ;
  assign y8221 = n16927 ;
  assign y8222 = ~n16929 ;
  assign y8223 = n4953 ;
  assign y8224 = ~1'b0 ;
  assign y8225 = n16930 ;
  assign y8226 = ~n16935 ;
  assign y8227 = ~n16936 ;
  assign y8228 = ~1'b0 ;
  assign y8229 = ~n16937 ;
  assign y8230 = n16938 ;
  assign y8231 = ~n16939 ;
  assign y8232 = ~n16940 ;
  assign y8233 = n16947 ;
  assign y8234 = n16949 ;
  assign y8235 = ~1'b0 ;
  assign y8236 = ~1'b0 ;
  assign y8237 = n16950 ;
  assign y8238 = n16952 ;
  assign y8239 = ~n16953 ;
  assign y8240 = ~1'b0 ;
  assign y8241 = n16956 ;
  assign y8242 = ~1'b0 ;
  assign y8243 = ~n16958 ;
  assign y8244 = n16960 ;
  assign y8245 = ~1'b0 ;
  assign y8246 = n16961 ;
  assign y8247 = ~n16962 ;
  assign y8248 = ~n16964 ;
  assign y8249 = ~n16965 ;
  assign y8250 = n16966 ;
  assign y8251 = n16968 ;
  assign y8252 = ~n16969 ;
  assign y8253 = ~n16970 ;
  assign y8254 = ~1'b0 ;
  assign y8255 = n16974 ;
  assign y8256 = ~1'b0 ;
  assign y8257 = n16976 ;
  assign y8258 = n16978 ;
  assign y8259 = n16983 ;
  assign y8260 = ~1'b0 ;
  assign y8261 = n16987 ;
  assign y8262 = n16988 ;
  assign y8263 = ~1'b0 ;
  assign y8264 = ~1'b0 ;
  assign y8265 = ~1'b0 ;
  assign y8266 = ~1'b0 ;
  assign y8267 = ~1'b0 ;
  assign y8268 = n16991 ;
  assign y8269 = ~n16992 ;
  assign y8270 = ~1'b0 ;
  assign y8271 = ~n16998 ;
  assign y8272 = ~1'b0 ;
  assign y8273 = ~1'b0 ;
  assign y8274 = ~1'b0 ;
  assign y8275 = ~1'b0 ;
  assign y8276 = ~n16999 ;
  assign y8277 = ~n17005 ;
  assign y8278 = ~1'b0 ;
  assign y8279 = n17010 ;
  assign y8280 = ~1'b0 ;
  assign y8281 = n17017 ;
  assign y8282 = n17018 ;
  assign y8283 = n17019 ;
  assign y8284 = n17023 ;
  assign y8285 = ~n17025 ;
  assign y8286 = ~1'b0 ;
  assign y8287 = ~n17031 ;
  assign y8288 = n913 ;
  assign y8289 = n17039 ;
  assign y8290 = 1'b0 ;
  assign y8291 = ~n17043 ;
  assign y8292 = ~n17047 ;
  assign y8293 = ~1'b0 ;
  assign y8294 = n17049 ;
  assign y8295 = n5034 ;
  assign y8296 = ~1'b0 ;
  assign y8297 = n17055 ;
  assign y8298 = ~n17058 ;
  assign y8299 = ~n17070 ;
  assign y8300 = ~n17074 ;
  assign y8301 = ~n17077 ;
  assign y8302 = n17079 ;
  assign y8303 = n9801 ;
  assign y8304 = ~n2366 ;
  assign y8305 = n17080 ;
  assign y8306 = ~n17082 ;
  assign y8307 = ~n17084 ;
  assign y8308 = ~n17086 ;
  assign y8309 = n17087 ;
  assign y8310 = ~1'b0 ;
  assign y8311 = n17093 ;
  assign y8312 = ~1'b0 ;
  assign y8313 = ~n17095 ;
  assign y8314 = ~1'b0 ;
  assign y8315 = ~n17098 ;
  assign y8316 = ~1'b0 ;
  assign y8317 = ~1'b0 ;
  assign y8318 = ~1'b0 ;
  assign y8319 = ~n17102 ;
  assign y8320 = ~n17103 ;
  assign y8321 = ~n17112 ;
  assign y8322 = n17116 ;
  assign y8323 = ~n17118 ;
  assign y8324 = ~1'b0 ;
  assign y8325 = ~1'b0 ;
  assign y8326 = ~1'b0 ;
  assign y8327 = ~n17120 ;
  assign y8328 = ~n17121 ;
  assign y8329 = ~n17122 ;
  assign y8330 = ~1'b0 ;
  assign y8331 = ~1'b0 ;
  assign y8332 = ~n14437 ;
  assign y8333 = ~1'b0 ;
  assign y8334 = ~n17124 ;
  assign y8335 = ~1'b0 ;
  assign y8336 = ~n2297 ;
  assign y8337 = n17129 ;
  assign y8338 = ~1'b0 ;
  assign y8339 = ~n17137 ;
  assign y8340 = ~1'b0 ;
  assign y8341 = ~n293 ;
  assign y8342 = ~n17140 ;
  assign y8343 = n17143 ;
  assign y8344 = n17146 ;
  assign y8345 = ~n17148 ;
  assign y8346 = ~1'b0 ;
  assign y8347 = n17152 ;
  assign y8348 = ~n17153 ;
  assign y8349 = ~n17162 ;
  assign y8350 = n17164 ;
  assign y8351 = ~1'b0 ;
  assign y8352 = n17165 ;
  assign y8353 = ~n17167 ;
  assign y8354 = ~1'b0 ;
  assign y8355 = ~n17168 ;
  assign y8356 = ~n17170 ;
  assign y8357 = n17171 ;
  assign y8358 = ~1'b0 ;
  assign y8359 = ~1'b0 ;
  assign y8360 = ~n17175 ;
  assign y8361 = ~1'b0 ;
  assign y8362 = ~n17181 ;
  assign y8363 = n17184 ;
  assign y8364 = ~n17190 ;
  assign y8365 = ~n17193 ;
  assign y8366 = ~n17195 ;
  assign y8367 = ~1'b0 ;
  assign y8368 = n17196 ;
  assign y8369 = ~n17201 ;
  assign y8370 = n17202 ;
  assign y8371 = n17216 ;
  assign y8372 = ~1'b0 ;
  assign y8373 = n17222 ;
  assign y8374 = ~1'b0 ;
  assign y8375 = ~n17223 ;
  assign y8376 = ~1'b0 ;
  assign y8377 = n17224 ;
  assign y8378 = n17231 ;
  assign y8379 = n17232 ;
  assign y8380 = ~n17235 ;
  assign y8381 = n17242 ;
  assign y8382 = ~n17243 ;
  assign y8383 = ~1'b0 ;
  assign y8384 = ~n17244 ;
  assign y8385 = ~n17251 ;
  assign y8386 = ~n17253 ;
  assign y8387 = n17254 ;
  assign y8388 = ~1'b0 ;
  assign y8389 = n17257 ;
  assign y8390 = n17261 ;
  assign y8391 = n17264 ;
  assign y8392 = ~1'b0 ;
  assign y8393 = n17266 ;
  assign y8394 = ~n17269 ;
  assign y8395 = ~1'b0 ;
  assign y8396 = n16146 ;
  assign y8397 = ~n17271 ;
  assign y8398 = ~1'b0 ;
  assign y8399 = ~1'b0 ;
  assign y8400 = ~n17275 ;
  assign y8401 = n17277 ;
  assign y8402 = ~n17278 ;
  assign y8403 = ~n17280 ;
  assign y8404 = n17283 ;
  assign y8405 = n17287 ;
  assign y8406 = ~n17289 ;
  assign y8407 = n17296 ;
  assign y8408 = ~1'b0 ;
  assign y8409 = ~n17299 ;
  assign y8410 = n17300 ;
  assign y8411 = n17301 ;
  assign y8412 = 1'b0 ;
  assign y8413 = ~1'b0 ;
  assign y8414 = ~1'b0 ;
  assign y8415 = n17302 ;
  assign y8416 = n12963 ;
  assign y8417 = n17304 ;
  assign y8418 = ~1'b0 ;
  assign y8419 = ~1'b0 ;
  assign y8420 = n17310 ;
  assign y8421 = ~1'b0 ;
  assign y8422 = n17316 ;
  assign y8423 = ~n17317 ;
  assign y8424 = n17319 ;
  assign y8425 = n17323 ;
  assign y8426 = ~1'b0 ;
  assign y8427 = n17324 ;
  assign y8428 = ~n17330 ;
  assign y8429 = ~1'b0 ;
  assign y8430 = ~n17331 ;
  assign y8431 = ~1'b0 ;
  assign y8432 = n17332 ;
  assign y8433 = ~n17333 ;
  assign y8434 = ~n17334 ;
  assign y8435 = n17339 ;
  assign y8436 = n7524 ;
  assign y8437 = ~n17340 ;
  assign y8438 = ~1'b0 ;
  assign y8439 = ~1'b0 ;
  assign y8440 = ~n17345 ;
  assign y8441 = n17347 ;
  assign y8442 = ~n17349 ;
  assign y8443 = n17350 ;
  assign y8444 = n17353 ;
  assign y8445 = ~1'b0 ;
  assign y8446 = ~n17358 ;
  assign y8447 = ~n17360 ;
  assign y8448 = ~n17361 ;
  assign y8449 = ~n17369 ;
  assign y8450 = ~1'b0 ;
  assign y8451 = n17370 ;
  assign y8452 = ~n17380 ;
  assign y8453 = n17383 ;
  assign y8454 = ~n17384 ;
  assign y8455 = ~1'b0 ;
  assign y8456 = ~n17390 ;
  assign y8457 = ~1'b0 ;
  assign y8458 = ~n17393 ;
  assign y8459 = ~n17396 ;
  assign y8460 = 1'b0 ;
  assign y8461 = ~n17397 ;
  assign y8462 = ~1'b0 ;
  assign y8463 = n1998 ;
  assign y8464 = ~n17399 ;
  assign y8465 = ~1'b0 ;
  assign y8466 = ~n17402 ;
  assign y8467 = ~n17403 ;
  assign y8468 = ~n17408 ;
  assign y8469 = ~1'b0 ;
  assign y8470 = n15779 ;
  assign y8471 = ~1'b0 ;
  assign y8472 = n17411 ;
  assign y8473 = n17412 ;
  assign y8474 = n17414 ;
  assign y8475 = n15391 ;
  assign y8476 = ~n17419 ;
  assign y8477 = n17421 ;
  assign y8478 = ~n17423 ;
  assign y8479 = ~n17427 ;
  assign y8480 = ~1'b0 ;
  assign y8481 = n17428 ;
  assign y8482 = n17429 ;
  assign y8483 = ~1'b0 ;
  assign y8484 = ~n17431 ;
  assign y8485 = n17433 ;
  assign y8486 = ~n17434 ;
  assign y8487 = n13231 ;
  assign y8488 = ~1'b0 ;
  assign y8489 = ~1'b0 ;
  assign y8490 = ~n17435 ;
  assign y8491 = ~1'b0 ;
  assign y8492 = ~1'b0 ;
  assign y8493 = ~n17439 ;
  assign y8494 = n17442 ;
  assign y8495 = ~n2372 ;
  assign y8496 = ~1'b0 ;
  assign y8497 = 1'b0 ;
  assign y8498 = ~n17443 ;
  assign y8499 = n17446 ;
  assign y8500 = ~n4428 ;
  assign y8501 = ~n17453 ;
  assign y8502 = n3855 ;
  assign y8503 = ~1'b0 ;
  assign y8504 = ~1'b0 ;
  assign y8505 = ~1'b0 ;
  assign y8506 = ~1'b0 ;
  assign y8507 = ~n17454 ;
  assign y8508 = n17459 ;
  assign y8509 = n17460 ;
  assign y8510 = n17465 ;
  assign y8511 = ~1'b0 ;
  assign y8512 = ~n17467 ;
  assign y8513 = ~n17468 ;
  assign y8514 = n17474 ;
  assign y8515 = ~n17482 ;
  assign y8516 = n13474 ;
  assign y8517 = ~n17483 ;
  assign y8518 = ~n17484 ;
  assign y8519 = ~1'b0 ;
  assign y8520 = n17490 ;
  assign y8521 = n17494 ;
  assign y8522 = n17496 ;
  assign y8523 = n17497 ;
  assign y8524 = ~1'b0 ;
  assign y8525 = ~n17500 ;
  assign y8526 = n17501 ;
  assign y8527 = ~n8381 ;
  assign y8528 = ~1'b0 ;
  assign y8529 = ~1'b0 ;
  assign y8530 = ~n17507 ;
  assign y8531 = ~n17511 ;
  assign y8532 = ~1'b0 ;
  assign y8533 = ~1'b0 ;
  assign y8534 = n17515 ;
  assign y8535 = ~1'b0 ;
  assign y8536 = n17521 ;
  assign y8537 = n17522 ;
  assign y8538 = ~n14014 ;
  assign y8539 = ~n17524 ;
  assign y8540 = ~n17528 ;
  assign y8541 = ~n17536 ;
  assign y8542 = ~n17537 ;
  assign y8543 = ~1'b0 ;
  assign y8544 = ~n17538 ;
  assign y8545 = ~n17540 ;
  assign y8546 = ~n17541 ;
  assign y8547 = n17545 ;
  assign y8548 = ~n1021 ;
  assign y8549 = ~n17550 ;
  assign y8550 = n17551 ;
  assign y8551 = ~1'b0 ;
  assign y8552 = ~n17553 ;
  assign y8553 = ~n17555 ;
  assign y8554 = n17556 ;
  assign y8555 = n17557 ;
  assign y8556 = ~1'b0 ;
  assign y8557 = ~1'b0 ;
  assign y8558 = ~1'b0 ;
  assign y8559 = 1'b0 ;
  assign y8560 = ~n17558 ;
  assign y8561 = ~1'b0 ;
  assign y8562 = ~1'b0 ;
  assign y8563 = ~n17560 ;
  assign y8564 = ~n13300 ;
  assign y8565 = n17565 ;
  assign y8566 = n17566 ;
  assign y8567 = ~1'b0 ;
  assign y8568 = ~n17567 ;
  assign y8569 = ~1'b0 ;
  assign y8570 = n17568 ;
  assign y8571 = n17570 ;
  assign y8572 = n17571 ;
  assign y8573 = n17573 ;
  assign y8574 = ~1'b0 ;
  assign y8575 = 1'b0 ;
  assign y8576 = ~n17574 ;
  assign y8577 = ~1'b0 ;
  assign y8578 = n17575 ;
  assign y8579 = ~n17576 ;
  assign y8580 = n17578 ;
  assign y8581 = ~1'b0 ;
  assign y8582 = n17582 ;
  assign y8583 = n17583 ;
  assign y8584 = ~1'b0 ;
  assign y8585 = ~1'b0 ;
  assign y8586 = ~1'b0 ;
  assign y8587 = ~1'b0 ;
  assign y8588 = ~n17587 ;
  assign y8589 = ~n17588 ;
  assign y8590 = ~n10299 ;
  assign y8591 = ~n17590 ;
  assign y8592 = n17599 ;
  assign y8593 = ~1'b0 ;
  assign y8594 = n17602 ;
  assign y8595 = ~n17605 ;
  assign y8596 = ~1'b0 ;
  assign y8597 = ~1'b0 ;
  assign y8598 = n17610 ;
  assign y8599 = ~n17611 ;
  assign y8600 = ~n17612 ;
  assign y8601 = ~1'b0 ;
  assign y8602 = n17613 ;
  assign y8603 = n17616 ;
  assign y8604 = ~n17628 ;
  assign y8605 = ~1'b0 ;
  assign y8606 = n17635 ;
  assign y8607 = n17637 ;
  assign y8608 = ~n17639 ;
  assign y8609 = ~n17642 ;
  assign y8610 = ~n17643 ;
  assign y8611 = ~n17645 ;
  assign y8612 = ~n17646 ;
  assign y8613 = ~1'b0 ;
  assign y8614 = n17655 ;
  assign y8615 = ~n17663 ;
  assign y8616 = ~1'b0 ;
  assign y8617 = ~n17668 ;
  assign y8618 = n17673 ;
  assign y8619 = n17685 ;
  assign y8620 = n17687 ;
  assign y8621 = n17692 ;
  assign y8622 = n17697 ;
  assign y8623 = ~1'b0 ;
  assign y8624 = ~n17699 ;
  assign y8625 = n17701 ;
  assign y8626 = ~n17703 ;
  assign y8627 = ~n17709 ;
  assign y8628 = ~n17710 ;
  assign y8629 = ~n9226 ;
  assign y8630 = ~1'b0 ;
  assign y8631 = ~1'b0 ;
  assign y8632 = ~n14389 ;
  assign y8633 = n17713 ;
  assign y8634 = ~n17716 ;
  assign y8635 = ~n17718 ;
  assign y8636 = ~1'b0 ;
  assign y8637 = ~n17719 ;
  assign y8638 = ~n14470 ;
  assign y8639 = n11983 ;
  assign y8640 = ~n17722 ;
  assign y8641 = ~n17723 ;
  assign y8642 = ~n10420 ;
  assign y8643 = ~n17725 ;
  assign y8644 = ~n17726 ;
  assign y8645 = ~n17732 ;
  assign y8646 = ~1'b0 ;
  assign y8647 = ~n17733 ;
  assign y8648 = n17737 ;
  assign y8649 = n17738 ;
  assign y8650 = n17739 ;
  assign y8651 = ~1'b0 ;
  assign y8652 = ~n17745 ;
  assign y8653 = 1'b0 ;
  assign y8654 = n17748 ;
  assign y8655 = ~n17750 ;
  assign y8656 = ~n17751 ;
  assign y8657 = n17755 ;
  assign y8658 = ~1'b0 ;
  assign y8659 = ~n17758 ;
  assign y8660 = n17761 ;
  assign y8661 = 1'b0 ;
  assign y8662 = n17764 ;
  assign y8663 = ~n17766 ;
  assign y8664 = 1'b0 ;
  assign y8665 = ~1'b0 ;
  assign y8666 = n17768 ;
  assign y8667 = n17771 ;
  assign y8668 = ~1'b0 ;
  assign y8669 = ~1'b0 ;
  assign y8670 = ~1'b0 ;
  assign y8671 = n17772 ;
  assign y8672 = ~n17773 ;
  assign y8673 = n17775 ;
  assign y8674 = n17777 ;
  assign y8675 = ~1'b0 ;
  assign y8676 = n8121 ;
  assign y8677 = ~1'b0 ;
  assign y8678 = ~n17778 ;
  assign y8679 = ~1'b0 ;
  assign y8680 = ~n17783 ;
  assign y8681 = ~n17785 ;
  assign y8682 = ~1'b0 ;
  assign y8683 = ~n17788 ;
  assign y8684 = ~1'b0 ;
  assign y8685 = ~1'b0 ;
  assign y8686 = n15459 ;
  assign y8687 = n17790 ;
  assign y8688 = ~n17791 ;
  assign y8689 = n17793 ;
  assign y8690 = n17797 ;
  assign y8691 = ~n17804 ;
  assign y8692 = n17806 ;
  assign y8693 = n17809 ;
  assign y8694 = n17812 ;
  assign y8695 = n17813 ;
  assign y8696 = n17814 ;
  assign y8697 = ~1'b0 ;
  assign y8698 = ~n17817 ;
  assign y8699 = ~n17820 ;
  assign y8700 = n17821 ;
  assign y8701 = ~n17823 ;
  assign y8702 = ~n17824 ;
  assign y8703 = ~n17825 ;
  assign y8704 = ~n17826 ;
  assign y8705 = ~1'b0 ;
  assign y8706 = ~1'b0 ;
  assign y8707 = ~1'b0 ;
  assign y8708 = n14313 ;
  assign y8709 = n17827 ;
  assign y8710 = ~n17828 ;
  assign y8711 = n17832 ;
  assign y8712 = ~n17836 ;
  assign y8713 = n17840 ;
  assign y8714 = n17843 ;
  assign y8715 = ~1'b0 ;
  assign y8716 = n17844 ;
  assign y8717 = 1'b0 ;
  assign y8718 = ~n17846 ;
  assign y8719 = ~n17847 ;
  assign y8720 = ~1'b0 ;
  assign y8721 = n17850 ;
  assign y8722 = n17856 ;
  assign y8723 = ~n17863 ;
  assign y8724 = ~1'b0 ;
  assign y8725 = n17865 ;
  assign y8726 = 1'b0 ;
  assign y8727 = ~n17866 ;
  assign y8728 = n17868 ;
  assign y8729 = n17869 ;
  assign y8730 = ~n17872 ;
  assign y8731 = n17873 ;
  assign y8732 = n17875 ;
  assign y8733 = ~n17876 ;
  assign y8734 = n17879 ;
  assign y8735 = n17881 ;
  assign y8736 = ~n17884 ;
  assign y8737 = n17885 ;
  assign y8738 = n17886 ;
  assign y8739 = ~1'b0 ;
  assign y8740 = ~n17887 ;
  assign y8741 = ~n17888 ;
  assign y8742 = n17890 ;
  assign y8743 = n17896 ;
  assign y8744 = ~1'b0 ;
  assign y8745 = ~1'b0 ;
  assign y8746 = n17901 ;
  assign y8747 = ~1'b0 ;
  assign y8748 = n17902 ;
  assign y8749 = ~n17906 ;
  assign y8750 = ~1'b0 ;
  assign y8751 = ~1'b0 ;
  assign y8752 = n17907 ;
  assign y8753 = ~n17908 ;
  assign y8754 = n17251 ;
  assign y8755 = ~1'b0 ;
  assign y8756 = ~n17910 ;
  assign y8757 = n17912 ;
  assign y8758 = 1'b0 ;
  assign y8759 = ~n17914 ;
  assign y8760 = ~n17916 ;
  assign y8761 = ~1'b0 ;
  assign y8762 = ~n17921 ;
  assign y8763 = ~1'b0 ;
  assign y8764 = ~1'b0 ;
  assign y8765 = ~1'b0 ;
  assign y8766 = ~n17923 ;
  assign y8767 = ~x115 ;
  assign y8768 = ~1'b0 ;
  assign y8769 = ~n17925 ;
  assign y8770 = ~1'b0 ;
  assign y8771 = ~n2644 ;
  assign y8772 = ~n17926 ;
  assign y8773 = ~1'b0 ;
  assign y8774 = n17932 ;
  assign y8775 = ~1'b0 ;
  assign y8776 = ~1'b0 ;
  assign y8777 = ~n17935 ;
  assign y8778 = ~n17936 ;
  assign y8779 = ~1'b0 ;
  assign y8780 = ~n17939 ;
  assign y8781 = ~n17942 ;
  assign y8782 = n17944 ;
  assign y8783 = n17946 ;
  assign y8784 = ~1'b0 ;
  assign y8785 = n17950 ;
  assign y8786 = ~1'b0 ;
  assign y8787 = n17951 ;
  assign y8788 = ~n17952 ;
  assign y8789 = n17953 ;
  assign y8790 = ~n17956 ;
  assign y8791 = ~n17963 ;
  assign y8792 = n11506 ;
  assign y8793 = n17964 ;
  assign y8794 = ~n17972 ;
  assign y8795 = ~n17976 ;
  assign y8796 = ~n17979 ;
  assign y8797 = ~n17981 ;
  assign y8798 = ~1'b0 ;
  assign y8799 = n17985 ;
  assign y8800 = n17986 ;
  assign y8801 = ~n17991 ;
  assign y8802 = ~n10731 ;
  assign y8803 = ~n9200 ;
  assign y8804 = ~n7263 ;
  assign y8805 = ~n17992 ;
  assign y8806 = ~n17993 ;
  assign y8807 = ~1'b0 ;
  assign y8808 = n17996 ;
  assign y8809 = n18000 ;
  assign y8810 = ~n18005 ;
  assign y8811 = ~n18009 ;
  assign y8812 = n18013 ;
  assign y8813 = n18014 ;
  assign y8814 = n18017 ;
  assign y8815 = ~n18020 ;
  assign y8816 = n18022 ;
  assign y8817 = ~1'b0 ;
  assign y8818 = ~n18023 ;
  assign y8819 = n18028 ;
  assign y8820 = ~n18033 ;
  assign y8821 = n18035 ;
  assign y8822 = n18037 ;
  assign y8823 = n18039 ;
  assign y8824 = ~n18040 ;
  assign y8825 = n18041 ;
  assign y8826 = ~n18048 ;
  assign y8827 = ~n18050 ;
  assign y8828 = ~n18052 ;
  assign y8829 = ~n18053 ;
  assign y8830 = ~1'b0 ;
  assign y8831 = ~1'b0 ;
  assign y8832 = n18054 ;
  assign y8833 = ~n18055 ;
  assign y8834 = ~1'b0 ;
  assign y8835 = 1'b0 ;
  assign y8836 = n18057 ;
  assign y8837 = ~1'b0 ;
  assign y8838 = ~n18064 ;
  assign y8839 = ~1'b0 ;
  assign y8840 = ~1'b0 ;
  assign y8841 = n18065 ;
  assign y8842 = n18070 ;
  assign y8843 = ~1'b0 ;
  assign y8844 = ~n18071 ;
  assign y8845 = ~n18072 ;
  assign y8846 = ~1'b0 ;
  assign y8847 = ~1'b0 ;
  assign y8848 = n18076 ;
  assign y8849 = ~1'b0 ;
  assign y8850 = ~1'b0 ;
  assign y8851 = n18078 ;
  assign y8852 = n18079 ;
  assign y8853 = ~1'b0 ;
  assign y8854 = 1'b0 ;
  assign y8855 = ~n18083 ;
  assign y8856 = ~1'b0 ;
  assign y8857 = ~n18089 ;
  assign y8858 = n18099 ;
  assign y8859 = ~1'b0 ;
  assign y8860 = ~n18106 ;
  assign y8861 = ~n18107 ;
  assign y8862 = ~n18110 ;
  assign y8863 = n18112 ;
  assign y8864 = ~n18118 ;
  assign y8865 = n18124 ;
  assign y8866 = ~1'b0 ;
  assign y8867 = ~n18137 ;
  assign y8868 = n18138 ;
  assign y8869 = ~1'b0 ;
  assign y8870 = n18142 ;
  assign y8871 = ~1'b0 ;
  assign y8872 = n18145 ;
  assign y8873 = ~n18152 ;
  assign y8874 = ~1'b0 ;
  assign y8875 = ~1'b0 ;
  assign y8876 = ~n18155 ;
  assign y8877 = n18157 ;
  assign y8878 = ~1'b0 ;
  assign y8879 = n18158 ;
  assign y8880 = ~n18160 ;
  assign y8881 = n18162 ;
  assign y8882 = ~n18163 ;
  assign y8883 = n18166 ;
  assign y8884 = ~1'b0 ;
  assign y8885 = ~n18169 ;
  assign y8886 = n18171 ;
  assign y8887 = ~n18174 ;
  assign y8888 = ~n18183 ;
  assign y8889 = ~n18184 ;
  assign y8890 = ~1'b0 ;
  assign y8891 = ~n18186 ;
  assign y8892 = ~1'b0 ;
  assign y8893 = ~n18188 ;
  assign y8894 = n18192 ;
  assign y8895 = n18196 ;
  assign y8896 = ~n18198 ;
  assign y8897 = ~n18204 ;
  assign y8898 = n18205 ;
  assign y8899 = ~1'b0 ;
  assign y8900 = n18209 ;
  assign y8901 = n18211 ;
  assign y8902 = ~n18218 ;
  assign y8903 = n18219 ;
  assign y8904 = ~1'b0 ;
  assign y8905 = ~n18223 ;
  assign y8906 = ~n1125 ;
  assign y8907 = ~1'b0 ;
  assign y8908 = ~1'b0 ;
  assign y8909 = n18228 ;
  assign y8910 = ~n18231 ;
  assign y8911 = n18232 ;
  assign y8912 = n18233 ;
  assign y8913 = ~n18237 ;
  assign y8914 = ~n18239 ;
  assign y8915 = ~n18242 ;
  assign y8916 = n2875 ;
  assign y8917 = n18243 ;
  assign y8918 = ~n2225 ;
  assign y8919 = ~n18244 ;
  assign y8920 = ~n18246 ;
  assign y8921 = ~1'b0 ;
  assign y8922 = ~n18250 ;
  assign y8923 = ~1'b0 ;
  assign y8924 = n18253 ;
  assign y8925 = ~n18254 ;
  assign y8926 = n18257 ;
  assign y8927 = n18261 ;
  assign y8928 = n18263 ;
  assign y8929 = ~1'b0 ;
  assign y8930 = ~n18266 ;
  assign y8931 = ~n18267 ;
  assign y8932 = n18276 ;
  assign y8933 = ~n18277 ;
  assign y8934 = n18284 ;
  assign y8935 = ~n18287 ;
  assign y8936 = ~n18290 ;
  assign y8937 = ~n18293 ;
  assign y8938 = n18295 ;
  assign y8939 = n18296 ;
  assign y8940 = ~1'b0 ;
  assign y8941 = ~1'b0 ;
  assign y8942 = ~n1051 ;
  assign y8943 = ~n18302 ;
  assign y8944 = n18303 ;
  assign y8945 = n18309 ;
  assign y8946 = n18312 ;
  assign y8947 = ~1'b0 ;
  assign y8948 = ~n18313 ;
  assign y8949 = n18315 ;
  assign y8950 = 1'b0 ;
  assign y8951 = ~n18317 ;
  assign y8952 = n18318 ;
  assign y8953 = n18319 ;
  assign y8954 = n18321 ;
  assign y8955 = ~1'b0 ;
  assign y8956 = ~1'b0 ;
  assign y8957 = 1'b0 ;
  assign y8958 = ~n18323 ;
  assign y8959 = n18324 ;
  assign y8960 = ~1'b0 ;
  assign y8961 = ~n18325 ;
  assign y8962 = n18330 ;
  assign y8963 = ~1'b0 ;
  assign y8964 = ~n18331 ;
  assign y8965 = ~n18340 ;
  assign y8966 = ~1'b0 ;
  assign y8967 = n1648 ;
  assign y8968 = n18341 ;
  assign y8969 = n18345 ;
  assign y8970 = ~1'b0 ;
  assign y8971 = ~n18348 ;
  assign y8972 = n2570 ;
  assign y8973 = ~1'b0 ;
  assign y8974 = ~1'b0 ;
  assign y8975 = 1'b0 ;
  assign y8976 = n18350 ;
  assign y8977 = n18354 ;
  assign y8978 = ~1'b0 ;
  assign y8979 = ~n18356 ;
  assign y8980 = n18357 ;
  assign y8981 = ~n18360 ;
  assign y8982 = n18365 ;
  assign y8983 = ~n18367 ;
  assign y8984 = ~n5806 ;
  assign y8985 = n18369 ;
  assign y8986 = ~n18378 ;
  assign y8987 = n18380 ;
  assign y8988 = ~n18384 ;
  assign y8989 = ~n18386 ;
  assign y8990 = n18390 ;
  assign y8991 = ~1'b0 ;
  assign y8992 = ~n18396 ;
  assign y8993 = n18397 ;
  assign y8994 = ~n18399 ;
  assign y8995 = ~n18400 ;
  assign y8996 = ~1'b0 ;
  assign y8997 = ~1'b0 ;
  assign y8998 = ~n18401 ;
  assign y8999 = n18402 ;
  assign y9000 = 1'b0 ;
  assign y9001 = ~1'b0 ;
  assign y9002 = 1'b0 ;
  assign y9003 = ~1'b0 ;
  assign y9004 = ~1'b0 ;
  assign y9005 = ~n18406 ;
  assign y9006 = ~1'b0 ;
  assign y9007 = ~1'b0 ;
  assign y9008 = n18408 ;
  assign y9009 = n18411 ;
  assign y9010 = n18414 ;
  assign y9011 = ~n18415 ;
  assign y9012 = ~1'b0 ;
  assign y9013 = ~1'b0 ;
  assign y9014 = n18416 ;
  assign y9015 = ~1'b0 ;
  assign y9016 = ~1'b0 ;
  assign y9017 = n18419 ;
  assign y9018 = n18422 ;
  assign y9019 = n18423 ;
  assign y9020 = n18428 ;
  assign y9021 = n18430 ;
  assign y9022 = 1'b0 ;
  assign y9023 = ~1'b0 ;
  assign y9024 = ~n18432 ;
  assign y9025 = ~1'b0 ;
  assign y9026 = n18433 ;
  assign y9027 = n18447 ;
  assign y9028 = n18449 ;
  assign y9029 = n18453 ;
  assign y9030 = n18458 ;
  assign y9031 = ~n18459 ;
  assign y9032 = ~1'b0 ;
  assign y9033 = n18462 ;
  assign y9034 = ~1'b0 ;
  assign y9035 = ~1'b0 ;
  assign y9036 = ~1'b0 ;
  assign y9037 = ~1'b0 ;
  assign y9038 = ~n18465 ;
  assign y9039 = ~1'b0 ;
  assign y9040 = n18472 ;
  assign y9041 = ~n18474 ;
  assign y9042 = ~1'b0 ;
  assign y9043 = n18475 ;
  assign y9044 = ~n18481 ;
  assign y9045 = n18482 ;
  assign y9046 = ~n18486 ;
  assign y9047 = ~n18491 ;
  assign y9048 = ~1'b0 ;
  assign y9049 = ~n18493 ;
  assign y9050 = n18495 ;
  assign y9051 = n2297 ;
  assign y9052 = ~1'b0 ;
  assign y9053 = 1'b0 ;
  assign y9054 = ~n18500 ;
  assign y9055 = n11121 ;
  assign y9056 = ~1'b0 ;
  assign y9057 = ~1'b0 ;
  assign y9058 = n18509 ;
  assign y9059 = ~n18511 ;
  assign y9060 = ~n18514 ;
  assign y9061 = ~1'b0 ;
  assign y9062 = ~1'b0 ;
  assign y9063 = ~1'b0 ;
  assign y9064 = ~1'b0 ;
  assign y9065 = ~1'b0 ;
  assign y9066 = n18515 ;
  assign y9067 = ~n4222 ;
  assign y9068 = n18520 ;
  assign y9069 = ~1'b0 ;
  assign y9070 = n18453 ;
  assign y9071 = ~1'b0 ;
  assign y9072 = ~n18521 ;
  assign y9073 = ~n18530 ;
  assign y9074 = ~n18533 ;
  assign y9075 = n18534 ;
  assign y9076 = ~n18535 ;
  assign y9077 = ~n18536 ;
  assign y9078 = ~1'b0 ;
  assign y9079 = ~n18538 ;
  assign y9080 = ~n18550 ;
  assign y9081 = ~1'b0 ;
  assign y9082 = ~1'b0 ;
  assign y9083 = n18552 ;
  assign y9084 = ~n18555 ;
  assign y9085 = n18558 ;
  assign y9086 = n18572 ;
  assign y9087 = ~n18576 ;
  assign y9088 = n18582 ;
  assign y9089 = ~1'b0 ;
  assign y9090 = ~1'b0 ;
  assign y9091 = n18584 ;
  assign y9092 = ~n18587 ;
  assign y9093 = ~n18588 ;
  assign y9094 = ~n18592 ;
  assign y9095 = ~n18595 ;
  assign y9096 = n8236 ;
  assign y9097 = n6881 ;
  assign y9098 = ~n18599 ;
  assign y9099 = ~n18604 ;
  assign y9100 = ~1'b0 ;
  assign y9101 = ~n18606 ;
  assign y9102 = n18610 ;
  assign y9103 = n18620 ;
  assign y9104 = ~n18626 ;
  assign y9105 = n18629 ;
  assign y9106 = n18635 ;
  assign y9107 = n18638 ;
  assign y9108 = n18643 ;
  assign y9109 = n18645 ;
  assign y9110 = ~1'b0 ;
  assign y9111 = ~1'b0 ;
  assign y9112 = ~1'b0 ;
  assign y9113 = ~1'b0 ;
  assign y9114 = ~n18649 ;
  assign y9115 = n18652 ;
  assign y9116 = n18656 ;
  assign y9117 = ~n18658 ;
  assign y9118 = n18659 ;
  assign y9119 = n18666 ;
  assign y9120 = n18668 ;
  assign y9121 = ~1'b0 ;
  assign y9122 = ~n18670 ;
  assign y9123 = ~1'b0 ;
  assign y9124 = n18671 ;
  assign y9125 = ~n18675 ;
  assign y9126 = ~1'b0 ;
  assign y9127 = ~1'b0 ;
  assign y9128 = n18677 ;
  assign y9129 = ~n18680 ;
  assign y9130 = n18682 ;
  assign y9131 = ~1'b0 ;
  assign y9132 = ~n18688 ;
  assign y9133 = n18698 ;
  assign y9134 = n18702 ;
  assign y9135 = ~n18704 ;
  assign y9136 = n18712 ;
  assign y9137 = n5293 ;
  assign y9138 = n18715 ;
  assign y9139 = ~n18720 ;
  assign y9140 = n18722 ;
  assign y9141 = n18727 ;
  assign y9142 = 1'b0 ;
  assign y9143 = ~n7825 ;
  assign y9144 = ~1'b0 ;
  assign y9145 = n3494 ;
  assign y9146 = ~1'b0 ;
  assign y9147 = ~n18730 ;
  assign y9148 = ~n18731 ;
  assign y9149 = ~n18735 ;
  assign y9150 = n18737 ;
  assign y9151 = ~n18738 ;
  assign y9152 = ~n18739 ;
  assign y9153 = n18740 ;
  assign y9154 = n18744 ;
  assign y9155 = ~n18747 ;
  assign y9156 = 1'b0 ;
  assign y9157 = ~1'b0 ;
  assign y9158 = ~n18750 ;
  assign y9159 = ~n18751 ;
  assign y9160 = ~1'b0 ;
  assign y9161 = ~1'b0 ;
  assign y9162 = ~1'b0 ;
  assign y9163 = n18756 ;
  assign y9164 = ~n18757 ;
  assign y9165 = n18763 ;
  assign y9166 = ~1'b0 ;
  assign y9167 = n6582 ;
  assign y9168 = ~1'b0 ;
  assign y9169 = n18770 ;
  assign y9170 = n18773 ;
  assign y9171 = ~n18781 ;
  assign y9172 = ~n18782 ;
  assign y9173 = ~1'b0 ;
  assign y9174 = n18783 ;
  assign y9175 = ~1'b0 ;
  assign y9176 = n18785 ;
  assign y9177 = n18789 ;
  assign y9178 = n18792 ;
  assign y9179 = n18796 ;
  assign y9180 = n18798 ;
  assign y9181 = n18800 ;
  assign y9182 = ~1'b0 ;
  assign y9183 = ~1'b0 ;
  assign y9184 = n5165 ;
  assign y9185 = ~n18801 ;
  assign y9186 = ~n18804 ;
  assign y9187 = ~n18000 ;
  assign y9188 = ~n18805 ;
  assign y9189 = ~n18807 ;
  assign y9190 = n18808 ;
  assign y9191 = n18810 ;
  assign y9192 = n18813 ;
  assign y9193 = n18815 ;
  assign y9194 = n18816 ;
  assign y9195 = ~n18817 ;
  assign y9196 = ~n11650 ;
  assign y9197 = n18819 ;
  assign y9198 = ~n18824 ;
  assign y9199 = n18830 ;
  assign y9200 = n18832 ;
  assign y9201 = n18839 ;
  assign y9202 = n18846 ;
  assign y9203 = n18847 ;
  assign y9204 = n18848 ;
  assign y9205 = ~n18854 ;
  assign y9206 = ~1'b0 ;
  assign y9207 = ~n18858 ;
  assign y9208 = n18859 ;
  assign y9209 = n18865 ;
  assign y9210 = ~n18866 ;
  assign y9211 = n18869 ;
  assign y9212 = ~n18871 ;
  assign y9213 = n18873 ;
  assign y9214 = ~1'b0 ;
  assign y9215 = n18876 ;
  assign y9216 = ~1'b0 ;
  assign y9217 = ~n18877 ;
  assign y9218 = ~n8322 ;
  assign y9219 = n18879 ;
  assign y9220 = ~n18882 ;
  assign y9221 = n18884 ;
  assign y9222 = ~n18886 ;
  assign y9223 = ~1'b0 ;
  assign y9224 = ~1'b0 ;
  assign y9225 = n18887 ;
  assign y9226 = n18888 ;
  assign y9227 = n15341 ;
  assign y9228 = n18891 ;
  assign y9229 = ~1'b0 ;
  assign y9230 = ~n18895 ;
  assign y9231 = n18898 ;
  assign y9232 = n18902 ;
  assign y9233 = ~n18908 ;
  assign y9234 = n18909 ;
  assign y9235 = ~1'b0 ;
  assign y9236 = ~1'b0 ;
  assign y9237 = ~1'b0 ;
  assign y9238 = ~1'b0 ;
  assign y9239 = n18913 ;
  assign y9240 = ~n18918 ;
  assign y9241 = ~n860 ;
  assign y9242 = ~n18921 ;
  assign y9243 = ~n18927 ;
  assign y9244 = ~1'b0 ;
  assign y9245 = ~n1185 ;
  assign y9246 = ~n18930 ;
  assign y9247 = 1'b0 ;
  assign y9248 = ~1'b0 ;
  assign y9249 = ~1'b0 ;
  assign y9250 = n18932 ;
  assign y9251 = ~n18934 ;
  assign y9252 = ~1'b0 ;
  assign y9253 = ~1'b0 ;
  assign y9254 = ~n18939 ;
  assign y9255 = ~n18941 ;
  assign y9256 = ~n18944 ;
  assign y9257 = ~n18950 ;
  assign y9258 = ~1'b0 ;
  assign y9259 = n18952 ;
  assign y9260 = ~n18954 ;
  assign y9261 = ~n18957 ;
  assign y9262 = n18961 ;
  assign y9263 = n18962 ;
  assign y9264 = n18964 ;
  assign y9265 = ~n18966 ;
  assign y9266 = n18969 ;
  assign y9267 = ~n18970 ;
  assign y9268 = ~n18971 ;
  assign y9269 = n18974 ;
  assign y9270 = n19002 ;
  assign y9271 = ~1'b0 ;
  assign y9272 = ~1'b0 ;
  assign y9273 = ~n19007 ;
  assign y9274 = ~n19008 ;
  assign y9275 = ~1'b0 ;
  assign y9276 = ~n19010 ;
  assign y9277 = ~n19011 ;
  assign y9278 = n19012 ;
  assign y9279 = ~1'b0 ;
  assign y9280 = ~n19013 ;
  assign y9281 = n19014 ;
  assign y9282 = ~1'b0 ;
  assign y9283 = n19017 ;
  assign y9284 = ~n19018 ;
  assign y9285 = n19021 ;
  assign y9286 = ~1'b0 ;
  assign y9287 = ~n19024 ;
  assign y9288 = ~1'b0 ;
  assign y9289 = ~1'b0 ;
  assign y9290 = n19028 ;
  assign y9291 = n19031 ;
  assign y9292 = n19035 ;
  assign y9293 = n19040 ;
  assign y9294 = n19041 ;
  assign y9295 = ~1'b0 ;
  assign y9296 = ~n19042 ;
  assign y9297 = n1626 ;
  assign y9298 = ~1'b0 ;
  assign y9299 = ~1'b0 ;
  assign y9300 = ~n19049 ;
  assign y9301 = ~1'b0 ;
  assign y9302 = ~1'b0 ;
  assign y9303 = ~1'b0 ;
  assign y9304 = n19050 ;
  assign y9305 = n19052 ;
  assign y9306 = ~n19054 ;
  assign y9307 = ~n19057 ;
  assign y9308 = ~n19061 ;
  assign y9309 = ~n19065 ;
  assign y9310 = ~n19071 ;
  assign y9311 = ~n19073 ;
  assign y9312 = ~n5608 ;
  assign y9313 = n19074 ;
  assign y9314 = n19077 ;
  assign y9315 = n19078 ;
  assign y9316 = ~n19080 ;
  assign y9317 = ~1'b0 ;
  assign y9318 = 1'b0 ;
  assign y9319 = ~1'b0 ;
  assign y9320 = ~1'b0 ;
  assign y9321 = ~1'b0 ;
  assign y9322 = ~n19085 ;
  assign y9323 = ~1'b0 ;
  assign y9324 = n19086 ;
  assign y9325 = n19087 ;
  assign y9326 = n6718 ;
  assign y9327 = ~n19090 ;
  assign y9328 = 1'b0 ;
  assign y9329 = n19093 ;
  assign y9330 = ~n19095 ;
  assign y9331 = n19096 ;
  assign y9332 = ~1'b0 ;
  assign y9333 = ~1'b0 ;
  assign y9334 = n19108 ;
  assign y9335 = ~1'b0 ;
  assign y9336 = n19109 ;
  assign y9337 = ~n19110 ;
  assign y9338 = n19111 ;
  assign y9339 = n19115 ;
  assign y9340 = ~n19117 ;
  assign y9341 = ~n19119 ;
  assign y9342 = ~n19120 ;
  assign y9343 = n19121 ;
  assign y9344 = n19122 ;
  assign y9345 = 1'b0 ;
  assign y9346 = n19123 ;
  assign y9347 = ~n19126 ;
  assign y9348 = ~1'b0 ;
  assign y9349 = n19130 ;
  assign y9350 = n19131 ;
  assign y9351 = n19133 ;
  assign y9352 = ~1'b0 ;
  assign y9353 = n671 ;
  assign y9354 = n19135 ;
  assign y9355 = ~1'b0 ;
  assign y9356 = ~n19136 ;
  assign y9357 = ~n3494 ;
  assign y9358 = n12754 ;
  assign y9359 = ~n19141 ;
  assign y9360 = n19142 ;
  assign y9361 = ~n14497 ;
  assign y9362 = ~1'b0 ;
  assign y9363 = ~1'b0 ;
  assign y9364 = n19143 ;
  assign y9365 = n19148 ;
  assign y9366 = n19150 ;
  assign y9367 = ~n19153 ;
  assign y9368 = n19154 ;
  assign y9369 = ~1'b0 ;
  assign y9370 = ~n19155 ;
  assign y9371 = ~1'b0 ;
  assign y9372 = n19160 ;
  assign y9373 = 1'b0 ;
  assign y9374 = n19164 ;
  assign y9375 = ~n19165 ;
  assign y9376 = ~1'b0 ;
  assign y9377 = ~1'b0 ;
  assign y9378 = ~n19167 ;
  assign y9379 = ~n19169 ;
  assign y9380 = ~n19170 ;
  assign y9381 = n19171 ;
  assign y9382 = n19173 ;
  assign y9383 = ~1'b0 ;
  assign y9384 = ~n9635 ;
  assign y9385 = ~1'b0 ;
  assign y9386 = ~n19177 ;
  assign y9387 = ~1'b0 ;
  assign y9388 = ~1'b0 ;
  assign y9389 = ~n19178 ;
  assign y9390 = ~1'b0 ;
  assign y9391 = ~n19179 ;
  assign y9392 = ~1'b0 ;
  assign y9393 = n19181 ;
  assign y9394 = n19182 ;
  assign y9395 = ~n19183 ;
  assign y9396 = ~n19185 ;
  assign y9397 = n19189 ;
  assign y9398 = ~n19191 ;
  assign y9399 = n19193 ;
  assign y9400 = n19196 ;
  assign y9401 = n19197 ;
  assign y9402 = ~n14885 ;
  assign y9403 = n19198 ;
  assign y9404 = ~n19204 ;
  assign y9405 = ~n19208 ;
  assign y9406 = n19209 ;
  assign y9407 = ~1'b0 ;
  assign y9408 = n19217 ;
  assign y9409 = ~n19219 ;
  assign y9410 = ~1'b0 ;
  assign y9411 = n19223 ;
  assign y9412 = ~n19225 ;
  assign y9413 = n19227 ;
  assign y9414 = ~n19228 ;
  assign y9415 = ~n18499 ;
  assign y9416 = n19233 ;
  assign y9417 = n5975 ;
  assign y9418 = n19236 ;
  assign y9419 = ~n19242 ;
  assign y9420 = ~n19244 ;
  assign y9421 = ~1'b0 ;
  assign y9422 = n17438 ;
  assign y9423 = n19245 ;
  assign y9424 = ~1'b0 ;
  assign y9425 = ~1'b0 ;
  assign y9426 = ~1'b0 ;
  assign y9427 = n19246 ;
  assign y9428 = n19248 ;
  assign y9429 = ~1'b0 ;
  assign y9430 = ~n19252 ;
  assign y9431 = n19253 ;
  assign y9432 = ~n19254 ;
  assign y9433 = ~1'b0 ;
  assign y9434 = n19257 ;
  assign y9435 = ~1'b0 ;
  assign y9436 = ~1'b0 ;
  assign y9437 = ~1'b0 ;
  assign y9438 = n19259 ;
  assign y9439 = n19263 ;
  assign y9440 = n19265 ;
  assign y9441 = n19269 ;
  assign y9442 = n4222 ;
  assign y9443 = ~n19270 ;
  assign y9444 = ~1'b0 ;
  assign y9445 = ~n19271 ;
  assign y9446 = ~n19278 ;
  assign y9447 = ~n19281 ;
  assign y9448 = ~1'b0 ;
  assign y9449 = ~n671 ;
  assign y9450 = n19286 ;
  assign y9451 = ~1'b0 ;
  assign y9452 = n19287 ;
  assign y9453 = ~1'b0 ;
  assign y9454 = ~1'b0 ;
  assign y9455 = ~1'b0 ;
  assign y9456 = ~n19288 ;
  assign y9457 = n19292 ;
  assign y9458 = ~1'b0 ;
  assign y9459 = ~1'b0 ;
  assign y9460 = ~n8690 ;
  assign y9461 = n19294 ;
  assign y9462 = ~1'b0 ;
  assign y9463 = ~1'b0 ;
  assign y9464 = n19295 ;
  assign y9465 = n19303 ;
  assign y9466 = ~n19304 ;
  assign y9467 = 1'b0 ;
  assign y9468 = ~n19314 ;
  assign y9469 = ~1'b0 ;
  assign y9470 = ~1'b0 ;
  assign y9471 = ~1'b0 ;
  assign y9472 = ~1'b0 ;
  assign y9473 = n19318 ;
  assign y9474 = ~n19322 ;
  assign y9475 = ~n19323 ;
  assign y9476 = ~n19326 ;
  assign y9477 = ~n19327 ;
  assign y9478 = n19330 ;
  assign y9479 = ~n19331 ;
  assign y9480 = ~n19332 ;
  assign y9481 = ~1'b0 ;
  assign y9482 = ~n19333 ;
  assign y9483 = ~1'b0 ;
  assign y9484 = ~n17223 ;
  assign y9485 = ~n19340 ;
  assign y9486 = n19347 ;
  assign y9487 = ~n19354 ;
  assign y9488 = n19362 ;
  assign y9489 = n19364 ;
  assign y9490 = n19366 ;
  assign y9491 = ~1'b0 ;
  assign y9492 = n18557 ;
  assign y9493 = n19369 ;
  assign y9494 = ~1'b0 ;
  assign y9495 = n10329 ;
  assign y9496 = ~n19371 ;
  assign y9497 = ~1'b0 ;
  assign y9498 = 1'b0 ;
  assign y9499 = 1'b0 ;
  assign y9500 = ~1'b0 ;
  assign y9501 = ~1'b0 ;
  assign y9502 = ~1'b0 ;
  assign y9503 = n19380 ;
  assign y9504 = ~1'b0 ;
  assign y9505 = n19385 ;
  assign y9506 = 1'b0 ;
  assign y9507 = ~1'b0 ;
  assign y9508 = n19389 ;
  assign y9509 = n19392 ;
  assign y9510 = ~n19397 ;
  assign y9511 = ~n19401 ;
  assign y9512 = ~n19402 ;
  assign y9513 = n19408 ;
  assign y9514 = ~n4637 ;
  assign y9515 = n19409 ;
  assign y9516 = ~n19412 ;
  assign y9517 = ~n19419 ;
  assign y9518 = ~n19420 ;
  assign y9519 = 1'b0 ;
  assign y9520 = ~n19425 ;
  assign y9521 = ~n19427 ;
  assign y9522 = ~n19428 ;
  assign y9523 = n19432 ;
  assign y9524 = n7958 ;
  assign y9525 = ~1'b0 ;
  assign y9526 = 1'b0 ;
  assign y9527 = n19433 ;
  assign y9528 = n19441 ;
  assign y9529 = 1'b0 ;
  assign y9530 = ~n19447 ;
  assign y9531 = ~1'b0 ;
  assign y9532 = ~1'b0 ;
  assign y9533 = n19450 ;
  assign y9534 = ~1'b0 ;
  assign y9535 = n19451 ;
  assign y9536 = ~1'b0 ;
  assign y9537 = n19453 ;
  assign y9538 = n19458 ;
  assign y9539 = ~n19459 ;
  assign y9540 = ~1'b0 ;
  assign y9541 = n19462 ;
  assign y9542 = n19463 ;
  assign y9543 = ~1'b0 ;
  assign y9544 = ~1'b0 ;
  assign y9545 = n19464 ;
  assign y9546 = ~n19479 ;
  assign y9547 = ~1'b0 ;
  assign y9548 = n19485 ;
  assign y9549 = n19492 ;
  assign y9550 = n19494 ;
  assign y9551 = n19502 ;
  assign y9552 = ~1'b0 ;
  assign y9553 = ~n14394 ;
  assign y9554 = n19507 ;
  assign y9555 = n19517 ;
  assign y9556 = ~n19519 ;
  assign y9557 = ~1'b0 ;
  assign y9558 = n19523 ;
  assign y9559 = ~n19527 ;
  assign y9560 = ~n19532 ;
  assign y9561 = n19533 ;
  assign y9562 = ~n19534 ;
  assign y9563 = ~n19538 ;
  assign y9564 = n19543 ;
  assign y9565 = n19545 ;
  assign y9566 = ~1'b0 ;
  assign y9567 = ~1'b0 ;
  assign y9568 = n19547 ;
  assign y9569 = ~n19548 ;
  assign y9570 = n19549 ;
  assign y9571 = n19553 ;
  assign y9572 = n19557 ;
  assign y9573 = ~n9758 ;
  assign y9574 = n19558 ;
  assign y9575 = n19559 ;
  assign y9576 = ~n3693 ;
  assign y9577 = ~1'b0 ;
  assign y9578 = ~1'b0 ;
  assign y9579 = ~1'b0 ;
  assign y9580 = ~n19568 ;
  assign y9581 = ~n19569 ;
  assign y9582 = n19571 ;
  assign y9583 = 1'b0 ;
  assign y9584 = ~n19572 ;
  assign y9585 = ~1'b0 ;
  assign y9586 = ~n19573 ;
  assign y9587 = n19575 ;
  assign y9588 = n5686 ;
  assign y9589 = n19578 ;
  assign y9590 = ~n19323 ;
  assign y9591 = ~n6357 ;
  assign y9592 = ~n19581 ;
  assign y9593 = n19585 ;
  assign y9594 = ~1'b0 ;
  assign y9595 = ~n19587 ;
  assign y9596 = n19594 ;
  assign y9597 = ~n19599 ;
  assign y9598 = ~n19600 ;
  assign y9599 = ~1'b0 ;
  assign y9600 = ~1'b0 ;
  assign y9601 = ~1'b0 ;
  assign y9602 = ~1'b0 ;
  assign y9603 = ~n19603 ;
  assign y9604 = 1'b0 ;
  assign y9605 = ~n19604 ;
  assign y9606 = ~n19605 ;
  assign y9607 = ~1'b0 ;
  assign y9608 = n19606 ;
  assign y9609 = n19612 ;
  assign y9610 = ~n19613 ;
  assign y9611 = n19617 ;
  assign y9612 = n19618 ;
  assign y9613 = n19623 ;
  assign y9614 = n19625 ;
  assign y9615 = n19626 ;
  assign y9616 = ~1'b0 ;
  assign y9617 = ~1'b0 ;
  assign y9618 = ~n19630 ;
  assign y9619 = ~n19631 ;
  assign y9620 = ~n19633 ;
  assign y9621 = ~n19634 ;
  assign y9622 = n1292 ;
  assign y9623 = ~1'b0 ;
  assign y9624 = ~1'b0 ;
  assign y9625 = ~n19636 ;
  assign y9626 = ~n19642 ;
  assign y9627 = n19644 ;
  assign y9628 = n19645 ;
  assign y9629 = ~1'b0 ;
  assign y9630 = ~n19646 ;
  assign y9631 = n19651 ;
  assign y9632 = n19653 ;
  assign y9633 = n19657 ;
  assign y9634 = ~n19658 ;
  assign y9635 = n19659 ;
  assign y9636 = n19660 ;
  assign y9637 = ~1'b0 ;
  assign y9638 = ~n19662 ;
  assign y9639 = ~n19663 ;
  assign y9640 = n19666 ;
  assign y9641 = ~n19670 ;
  assign y9642 = ~n19675 ;
  assign y9643 = n19679 ;
  assign y9644 = ~n19685 ;
  assign y9645 = ~1'b0 ;
  assign y9646 = ~n19686 ;
  assign y9647 = ~n19693 ;
  assign y9648 = ~n19694 ;
  assign y9649 = ~n19696 ;
  assign y9650 = ~1'b0 ;
  assign y9651 = ~1'b0 ;
  assign y9652 = ~1'b0 ;
  assign y9653 = n19698 ;
  assign y9654 = 1'b0 ;
  assign y9655 = ~1'b0 ;
  assign y9656 = ~n19702 ;
  assign y9657 = ~n19709 ;
  assign y9658 = n19710 ;
  assign y9659 = ~1'b0 ;
  assign y9660 = 1'b0 ;
  assign y9661 = ~n19711 ;
  assign y9662 = n19712 ;
  assign y9663 = n19715 ;
  assign y9664 = n19721 ;
  assign y9665 = n19725 ;
  assign y9666 = n19727 ;
  assign y9667 = n19728 ;
  assign y9668 = ~n19729 ;
  assign y9669 = ~n19732 ;
  assign y9670 = ~1'b0 ;
  assign y9671 = n19735 ;
  assign y9672 = n19736 ;
  assign y9673 = ~n19738 ;
  assign y9674 = ~n19740 ;
  assign y9675 = n19742 ;
  assign y9676 = ~n19743 ;
  assign y9677 = ~n19745 ;
  assign y9678 = ~1'b0 ;
  assign y9679 = ~n19747 ;
  assign y9680 = ~n19749 ;
  assign y9681 = ~n19751 ;
  assign y9682 = ~n9708 ;
  assign y9683 = ~n19754 ;
  assign y9684 = ~n19761 ;
  assign y9685 = n19763 ;
  assign y9686 = n19769 ;
  assign y9687 = ~n9865 ;
  assign y9688 = ~1'b0 ;
  assign y9689 = ~n19770 ;
  assign y9690 = ~n19772 ;
  assign y9691 = ~1'b0 ;
  assign y9692 = n19774 ;
  assign y9693 = ~n19016 ;
  assign y9694 = n451 ;
  assign y9695 = ~n19776 ;
  assign y9696 = ~n19782 ;
  assign y9697 = ~n19784 ;
  assign y9698 = ~1'b0 ;
  assign y9699 = n19789 ;
  assign y9700 = n19790 ;
  assign y9701 = n19793 ;
  assign y9702 = n19796 ;
  assign y9703 = ~1'b0 ;
  assign y9704 = ~1'b0 ;
  assign y9705 = n19802 ;
  assign y9706 = n12274 ;
  assign y9707 = ~n19803 ;
  assign y9708 = n19805 ;
  assign y9709 = ~1'b0 ;
  assign y9710 = ~1'b0 ;
  assign y9711 = ~n19807 ;
  assign y9712 = ~1'b0 ;
  assign y9713 = 1'b0 ;
  assign y9714 = n19809 ;
  assign y9715 = ~1'b0 ;
  assign y9716 = ~1'b0 ;
  assign y9717 = ~1'b0 ;
  assign y9718 = n19811 ;
  assign y9719 = n19812 ;
  assign y9720 = ~1'b0 ;
  assign y9721 = ~1'b0 ;
  assign y9722 = n19817 ;
  assign y9723 = ~n19818 ;
  assign y9724 = ~1'b0 ;
  assign y9725 = n19821 ;
  assign y9726 = ~n19834 ;
  assign y9727 = ~n19836 ;
  assign y9728 = ~n19837 ;
  assign y9729 = 1'b0 ;
  assign y9730 = ~n19839 ;
  assign y9731 = ~n19858 ;
  assign y9732 = ~n19860 ;
  assign y9733 = n19861 ;
  assign y9734 = ~1'b0 ;
  assign y9735 = ~1'b0 ;
  assign y9736 = ~n19863 ;
  assign y9737 = ~n19865 ;
  assign y9738 = n19867 ;
  assign y9739 = ~n19869 ;
  assign y9740 = ~1'b0 ;
  assign y9741 = ~n19871 ;
  assign y9742 = n19872 ;
  assign y9743 = n19873 ;
  assign y9744 = ~n19877 ;
  assign y9745 = n1387 ;
  assign y9746 = ~1'b0 ;
  assign y9747 = n17747 ;
  assign y9748 = ~n19878 ;
  assign y9749 = ~n19880 ;
  assign y9750 = ~x147 ;
  assign y9751 = ~n19883 ;
  assign y9752 = ~n19892 ;
  assign y9753 = ~1'b0 ;
  assign y9754 = n19895 ;
  assign y9755 = ~n19898 ;
  assign y9756 = ~n4013 ;
  assign y9757 = 1'b0 ;
  assign y9758 = ~1'b0 ;
  assign y9759 = ~1'b0 ;
  assign y9760 = ~1'b0 ;
  assign y9761 = ~n19900 ;
  assign y9762 = n19901 ;
  assign y9763 = ~1'b0 ;
  assign y9764 = n19903 ;
  assign y9765 = ~1'b0 ;
  assign y9766 = n19905 ;
  assign y9767 = ~n19908 ;
  assign y9768 = ~n19909 ;
  assign y9769 = ~n19910 ;
  assign y9770 = n19911 ;
  assign y9771 = n19914 ;
  assign y9772 = ~n19917 ;
  assign y9773 = n19919 ;
  assign y9774 = ~1'b0 ;
  assign y9775 = ~n19921 ;
  assign y9776 = ~n19923 ;
  assign y9777 = 1'b0 ;
  assign y9778 = n16859 ;
  assign y9779 = ~n19926 ;
  assign y9780 = ~n19927 ;
  assign y9781 = n19928 ;
  assign y9782 = n2192 ;
  assign y9783 = ~n6524 ;
  assign y9784 = n19929 ;
  assign y9785 = n19930 ;
  assign y9786 = n19932 ;
  assign y9787 = 1'b0 ;
  assign y9788 = ~n19934 ;
  assign y9789 = n19939 ;
  assign y9790 = ~1'b0 ;
  assign y9791 = ~n19941 ;
  assign y9792 = ~1'b0 ;
  assign y9793 = ~1'b0 ;
  assign y9794 = ~n19943 ;
  assign y9795 = ~1'b0 ;
  assign y9796 = n13620 ;
  assign y9797 = n19944 ;
  assign y9798 = ~1'b0 ;
  assign y9799 = n19947 ;
  assign y9800 = ~n19948 ;
  assign y9801 = n19950 ;
  assign y9802 = ~n19953 ;
  assign y9803 = n19954 ;
  assign y9804 = ~n19955 ;
  assign y9805 = ~1'b0 ;
  assign y9806 = ~n19956 ;
  assign y9807 = ~1'b0 ;
  assign y9808 = n19960 ;
  assign y9809 = n19961 ;
  assign y9810 = ~n19967 ;
  assign y9811 = ~n19969 ;
  assign y9812 = ~n19971 ;
  assign y9813 = ~n19973 ;
  assign y9814 = ~1'b0 ;
  assign y9815 = n19977 ;
  assign y9816 = 1'b0 ;
  assign y9817 = ~n19980 ;
  assign y9818 = 1'b0 ;
  assign y9819 = n19982 ;
  assign y9820 = ~n19984 ;
  assign y9821 = ~1'b0 ;
  assign y9822 = ~1'b0 ;
  assign y9823 = n19985 ;
  assign y9824 = n19987 ;
  assign y9825 = ~n19992 ;
  assign y9826 = ~1'b0 ;
  assign y9827 = ~1'b0 ;
  assign y9828 = ~n19996 ;
  assign y9829 = ~n19998 ;
  assign y9830 = n20001 ;
  assign y9831 = ~1'b0 ;
  assign y9832 = ~n20008 ;
  assign y9833 = ~n20017 ;
  assign y9834 = ~n20019 ;
  assign y9835 = ~n20020 ;
  assign y9836 = 1'b0 ;
  assign y9837 = ~1'b0 ;
  assign y9838 = ~1'b0 ;
  assign y9839 = n20021 ;
  assign y9840 = ~1'b0 ;
  assign y9841 = ~n20024 ;
  assign y9842 = ~n20026 ;
  assign y9843 = n20028 ;
  assign y9844 = n20030 ;
  assign y9845 = ~n20032 ;
  assign y9846 = ~n8529 ;
  assign y9847 = ~1'b0 ;
  assign y9848 = ~n20033 ;
  assign y9849 = ~n20034 ;
  assign y9850 = n14150 ;
  assign y9851 = n20037 ;
  assign y9852 = ~n20038 ;
  assign y9853 = ~1'b0 ;
  assign y9854 = ~1'b0 ;
  assign y9855 = ~n20043 ;
  assign y9856 = n20044 ;
  assign y9857 = ~1'b0 ;
  assign y9858 = ~1'b0 ;
  assign y9859 = ~n20052 ;
  assign y9860 = ~n20055 ;
  assign y9861 = ~n20058 ;
  assign y9862 = ~n20060 ;
  assign y9863 = ~1'b0 ;
  assign y9864 = n19104 ;
  assign y9865 = ~n8087 ;
  assign y9866 = n20064 ;
  assign y9867 = n20069 ;
  assign y9868 = ~n20071 ;
  assign y9869 = ~1'b0 ;
  assign y9870 = ~1'b0 ;
  assign y9871 = ~1'b0 ;
  assign y9872 = n20083 ;
  assign y9873 = n8980 ;
  assign y9874 = ~1'b0 ;
  assign y9875 = n20086 ;
  assign y9876 = ~n20088 ;
  assign y9877 = n20090 ;
  assign y9878 = ~n20093 ;
  assign y9879 = ~n20094 ;
  assign y9880 = n20095 ;
  assign y9881 = ~1'b0 ;
  assign y9882 = ~1'b0 ;
  assign y9883 = ~n20098 ;
  assign y9884 = ~n20100 ;
  assign y9885 = ~1'b0 ;
  assign y9886 = ~1'b0 ;
  assign y9887 = n20106 ;
  assign y9888 = ~n20107 ;
  assign y9889 = n20110 ;
  assign y9890 = ~1'b0 ;
  assign y9891 = ~n20115 ;
  assign y9892 = ~n6522 ;
  assign y9893 = n20116 ;
  assign y9894 = ~1'b0 ;
  assign y9895 = ~1'b0 ;
  assign y9896 = ~1'b0 ;
  assign y9897 = ~1'b0 ;
  assign y9898 = ~n20119 ;
  assign y9899 = ~n20121 ;
  assign y9900 = ~n20126 ;
  assign y9901 = n20128 ;
  assign y9902 = n20129 ;
  assign y9903 = ~n20130 ;
  assign y9904 = n20131 ;
  assign y9905 = n20134 ;
  assign y9906 = ~1'b0 ;
  assign y9907 = ~n20136 ;
  assign y9908 = ~n20138 ;
  assign y9909 = n20140 ;
  assign y9910 = ~n20141 ;
  assign y9911 = n20143 ;
  assign y9912 = ~1'b0 ;
  assign y9913 = ~1'b0 ;
  assign y9914 = n20151 ;
  assign y9915 = ~n10666 ;
  assign y9916 = ~n20154 ;
  assign y9917 = ~n20159 ;
  assign y9918 = n20166 ;
  assign y9919 = n10981 ;
  assign y9920 = n20169 ;
  assign y9921 = ~n20170 ;
  assign y9922 = ~n20172 ;
  assign y9923 = ~n20177 ;
  assign y9924 = ~n20179 ;
  assign y9925 = ~n5091 ;
  assign y9926 = ~1'b0 ;
  assign y9927 = ~n20180 ;
  assign y9928 = ~n20182 ;
  assign y9929 = n20184 ;
  assign y9930 = n20186 ;
  assign y9931 = ~n20187 ;
  assign y9932 = n20188 ;
  assign y9933 = ~n20190 ;
  assign y9934 = ~1'b0 ;
  assign y9935 = ~1'b0 ;
  assign y9936 = 1'b0 ;
  assign y9937 = n20193 ;
  assign y9938 = n20197 ;
  assign y9939 = n20198 ;
  assign y9940 = ~n20200 ;
  assign y9941 = n11871 ;
  assign y9942 = ~n20202 ;
  assign y9943 = n20203 ;
  assign y9944 = ~n20210 ;
  assign y9945 = ~n20211 ;
  assign y9946 = ~1'b0 ;
  assign y9947 = ~n10911 ;
  assign y9948 = ~n20216 ;
  assign y9949 = n20217 ;
  assign y9950 = ~n20221 ;
  assign y9951 = n20222 ;
  assign y9952 = ~1'b0 ;
  assign y9953 = ~n4031 ;
  assign y9954 = ~n20223 ;
  assign y9955 = ~n20227 ;
  assign y9956 = ~1'b0 ;
  assign y9957 = ~n20231 ;
  assign y9958 = ~1'b0 ;
  assign y9959 = n20243 ;
  assign y9960 = ~n20245 ;
  assign y9961 = ~n20247 ;
  assign y9962 = ~1'b0 ;
  assign y9963 = ~1'b0 ;
  assign y9964 = ~1'b0 ;
  assign y9965 = n20249 ;
  assign y9966 = ~n19769 ;
  assign y9967 = ~1'b0 ;
  assign y9968 = ~n20250 ;
  assign y9969 = ~1'b0 ;
  assign y9970 = ~n20251 ;
  assign y9971 = ~1'b0 ;
  assign y9972 = ~1'b0 ;
  assign y9973 = n20252 ;
  assign y9974 = ~1'b0 ;
  assign y9975 = ~n20253 ;
  assign y9976 = 1'b0 ;
  assign y9977 = n20260 ;
  assign y9978 = n20262 ;
  assign y9979 = ~n10129 ;
  assign y9980 = ~n20264 ;
  assign y9981 = n20265 ;
  assign y9982 = n20269 ;
  assign y9983 = n20270 ;
  assign y9984 = n20271 ;
  assign y9985 = n16980 ;
  assign y9986 = n20273 ;
  assign y9987 = ~n15689 ;
  assign y9988 = n20275 ;
  assign y9989 = n20278 ;
  assign y9990 = ~n20281 ;
  assign y9991 = ~n20283 ;
  assign y9992 = ~n20292 ;
  assign y9993 = n20295 ;
  assign y9994 = n20302 ;
  assign y9995 = ~n20306 ;
  assign y9996 = n20308 ;
  assign y9997 = ~1'b0 ;
  assign y9998 = n20310 ;
  assign y9999 = n20312 ;
  assign y10000 = n20317 ;
  assign y10001 = ~n20322 ;
  assign y10002 = n20324 ;
  assign y10003 = ~n20326 ;
  assign y10004 = ~n20332 ;
  assign y10005 = ~1'b0 ;
  assign y10006 = ~n20333 ;
  assign y10007 = n20336 ;
  assign y10008 = n20337 ;
  assign y10009 = n20338 ;
  assign y10010 = ~1'b0 ;
  assign y10011 = ~1'b0 ;
  assign y10012 = ~1'b0 ;
  assign y10013 = ~n20339 ;
  assign y10014 = n20340 ;
  assign y10015 = ~n20341 ;
  assign y10016 = ~1'b0 ;
  assign y10017 = ~n20342 ;
  assign y10018 = n20346 ;
  assign y10019 = ~1'b0 ;
  assign y10020 = ~1'b0 ;
  assign y10021 = ~n20349 ;
  assign y10022 = n20350 ;
  assign y10023 = ~1'b0 ;
  assign y10024 = ~1'b0 ;
  assign y10025 = n20351 ;
  assign y10026 = ~1'b0 ;
  assign y10027 = ~n18630 ;
  assign y10028 = ~1'b0 ;
  assign y10029 = ~1'b0 ;
  assign y10030 = ~1'b0 ;
  assign y10031 = ~n20356 ;
  assign y10032 = n20358 ;
  assign y10033 = n20370 ;
  assign y10034 = n20372 ;
  assign y10035 = ~1'b0 ;
  assign y10036 = n20374 ;
  assign y10037 = n20376 ;
  assign y10038 = n20377 ;
  assign y10039 = n20378 ;
  assign y10040 = ~n20380 ;
  assign y10041 = n20381 ;
  assign y10042 = ~1'b0 ;
  assign y10043 = 1'b0 ;
  assign y10044 = ~n20383 ;
  assign y10045 = 1'b0 ;
  assign y10046 = ~n3703 ;
  assign y10047 = n20384 ;
  assign y10048 = ~n20387 ;
  assign y10049 = n20388 ;
  assign y10050 = ~1'b0 ;
  assign y10051 = ~n20392 ;
  assign y10052 = ~1'b0 ;
  assign y10053 = n20394 ;
  assign y10054 = ~n20395 ;
  assign y10055 = ~1'b0 ;
  assign y10056 = 1'b0 ;
  assign y10057 = ~n20396 ;
  assign y10058 = ~1'b0 ;
  assign y10059 = n20404 ;
  assign y10060 = n20405 ;
  assign y10061 = ~n4132 ;
  assign y10062 = n20408 ;
  assign y10063 = ~n20411 ;
  assign y10064 = ~n20413 ;
  assign y10065 = ~1'b0 ;
  assign y10066 = ~n20421 ;
  assign y10067 = n20423 ;
  assign y10068 = 1'b0 ;
  assign y10069 = n20427 ;
  assign y10070 = n20431 ;
  assign y10071 = ~1'b0 ;
  assign y10072 = ~n20434 ;
  assign y10073 = n20437 ;
  assign y10074 = n20439 ;
  assign y10075 = ~n20440 ;
  assign y10076 = ~n20443 ;
  assign y10077 = ~n20446 ;
  assign y10078 = ~n20448 ;
  assign y10079 = n20449 ;
  assign y10080 = ~1'b0 ;
  assign y10081 = ~n20451 ;
  assign y10082 = ~n20453 ;
  assign y10083 = ~n20459 ;
  assign y10084 = n20462 ;
  assign y10085 = ~1'b0 ;
  assign y10086 = ~1'b0 ;
  assign y10087 = ~1'b0 ;
  assign y10088 = n20463 ;
  assign y10089 = ~n20464 ;
  assign y10090 = ~1'b0 ;
  assign y10091 = n20465 ;
  assign y10092 = ~n20466 ;
  assign y10093 = n20468 ;
  assign y10094 = ~n3325 ;
  assign y10095 = ~n20470 ;
  assign y10096 = n20476 ;
  assign y10097 = n20477 ;
  assign y10098 = ~n20483 ;
  assign y10099 = n20486 ;
  assign y10100 = ~1'b0 ;
  assign y10101 = ~1'b0 ;
  assign y10102 = n20487 ;
  assign y10103 = ~n20492 ;
  assign y10104 = ~n20495 ;
  assign y10105 = n20500 ;
  assign y10106 = ~n20501 ;
  assign y10107 = n20502 ;
  assign y10108 = ~n20504 ;
  assign y10109 = ~n20511 ;
  assign y10110 = ~1'b0 ;
  assign y10111 = n20512 ;
  assign y10112 = ~n20514 ;
  assign y10113 = ~1'b0 ;
  assign y10114 = ~n20515 ;
  assign y10115 = n10963 ;
  assign y10116 = n20519 ;
  assign y10117 = ~1'b0 ;
  assign y10118 = ~n20522 ;
  assign y10119 = ~n20523 ;
  assign y10120 = ~n20529 ;
  assign y10121 = ~n10498 ;
  assign y10122 = n20530 ;
  assign y10123 = ~n20538 ;
  assign y10124 = ~n9993 ;
  assign y10125 = n20544 ;
  assign y10126 = n20545 ;
  assign y10127 = ~n20548 ;
  assign y10128 = ~1'b0 ;
  assign y10129 = ~1'b0 ;
  assign y10130 = ~1'b0 ;
  assign y10131 = ~1'b0 ;
  assign y10132 = ~n20551 ;
  assign y10133 = n20556 ;
  assign y10134 = ~1'b0 ;
  assign y10135 = n20560 ;
  assign y10136 = n20561 ;
  assign y10137 = ~1'b0 ;
  assign y10138 = n20564 ;
  assign y10139 = n20568 ;
  assign y10140 = ~n20569 ;
  assign y10141 = n20570 ;
  assign y10142 = ~1'b0 ;
  assign y10143 = n20571 ;
  assign y10144 = ~n306 ;
  assign y10145 = ~n12224 ;
  assign y10146 = n20575 ;
  assign y10147 = n20578 ;
  assign y10148 = ~n20579 ;
  assign y10149 = n20583 ;
  assign y10150 = ~1'b0 ;
  assign y10151 = ~n671 ;
  assign y10152 = ~n20586 ;
  assign y10153 = ~1'b0 ;
  assign y10154 = n20590 ;
  assign y10155 = ~n20594 ;
  assign y10156 = ~n20596 ;
  assign y10157 = n20601 ;
  assign y10158 = ~1'b0 ;
  assign y10159 = ~1'b0 ;
  assign y10160 = n20603 ;
  assign y10161 = ~n20605 ;
  assign y10162 = ~1'b0 ;
  assign y10163 = ~n20606 ;
  assign y10164 = ~n12517 ;
  assign y10165 = ~1'b0 ;
  assign y10166 = ~n20611 ;
  assign y10167 = ~1'b0 ;
  assign y10168 = ~n20616 ;
  assign y10169 = n20617 ;
  assign y10170 = n20623 ;
  assign y10171 = n20626 ;
  assign y10172 = 1'b0 ;
  assign y10173 = n20635 ;
  assign y10174 = ~n20639 ;
  assign y10175 = n20642 ;
  assign y10176 = n8838 ;
  assign y10177 = ~n20645 ;
  assign y10178 = ~n20646 ;
  assign y10179 = n20649 ;
  assign y10180 = n20651 ;
  assign y10181 = ~n20652 ;
  assign y10182 = ~1'b0 ;
  assign y10183 = 1'b0 ;
  assign y10184 = ~1'b0 ;
  assign y10185 = ~1'b0 ;
  assign y10186 = ~1'b0 ;
  assign y10187 = ~1'b0 ;
  assign y10188 = ~1'b0 ;
  assign y10189 = n1146 ;
  assign y10190 = ~1'b0 ;
  assign y10191 = ~1'b0 ;
  assign y10192 = ~n8225 ;
  assign y10193 = n20655 ;
  assign y10194 = n20661 ;
  assign y10195 = n20666 ;
  assign y10196 = ~n20667 ;
  assign y10197 = n20669 ;
  assign y10198 = ~n13847 ;
  assign y10199 = n20670 ;
  assign y10200 = ~1'b0 ;
  assign y10201 = ~1'b0 ;
  assign y10202 = ~n20672 ;
  assign y10203 = ~1'b0 ;
  assign y10204 = ~1'b0 ;
  assign y10205 = ~1'b0 ;
  assign y10206 = ~n20678 ;
  assign y10207 = ~n20679 ;
  assign y10208 = n20680 ;
  assign y10209 = ~n20681 ;
  assign y10210 = n20684 ;
  assign y10211 = ~n20690 ;
  assign y10212 = n20691 ;
  assign y10213 = 1'b0 ;
  assign y10214 = ~n20692 ;
  assign y10215 = ~n20695 ;
  assign y10216 = ~n20698 ;
  assign y10217 = ~1'b0 ;
  assign y10218 = 1'b0 ;
  assign y10219 = n20700 ;
  assign y10220 = n20707 ;
  assign y10221 = ~1'b0 ;
  assign y10222 = n20710 ;
  assign y10223 = n20712 ;
  assign y10224 = n20714 ;
  assign y10225 = ~1'b0 ;
  assign y10226 = ~n20715 ;
  assign y10227 = n20721 ;
  assign y10228 = n19283 ;
  assign y10229 = n20726 ;
  assign y10230 = ~n20727 ;
  assign y10231 = n20728 ;
  assign y10232 = ~n20731 ;
  assign y10233 = ~n20739 ;
  assign y10234 = n20741 ;
  assign y10235 = ~n20745 ;
  assign y10236 = ~n20750 ;
  assign y10237 = ~n20753 ;
  assign y10238 = ~n20755 ;
  assign y10239 = ~1'b0 ;
  assign y10240 = ~1'b0 ;
  assign y10241 = ~1'b0 ;
  assign y10242 = ~1'b0 ;
  assign y10243 = n20757 ;
  assign y10244 = n20761 ;
  assign y10245 = n20762 ;
  assign y10246 = n17765 ;
  assign y10247 = n20767 ;
  assign y10248 = ~1'b0 ;
  assign y10249 = ~1'b0 ;
  assign y10250 = n20771 ;
  assign y10251 = ~1'b0 ;
  assign y10252 = ~n20774 ;
  assign y10253 = ~1'b0 ;
  assign y10254 = ~1'b0 ;
  assign y10255 = ~n20778 ;
  assign y10256 = ~n20779 ;
  assign y10257 = n20784 ;
  assign y10258 = n8633 ;
  assign y10259 = ~n20788 ;
  assign y10260 = n20789 ;
  assign y10261 = ~1'b0 ;
  assign y10262 = ~n20792 ;
  assign y10263 = ~n20794 ;
  assign y10264 = ~n20795 ;
  assign y10265 = ~1'b0 ;
  assign y10266 = ~n20326 ;
  assign y10267 = n20797 ;
  assign y10268 = ~n1492 ;
  assign y10269 = ~n20802 ;
  assign y10270 = ~1'b0 ;
  assign y10271 = ~1'b0 ;
  assign y10272 = n20803 ;
  assign y10273 = n20805 ;
  assign y10274 = ~n16804 ;
  assign y10275 = ~1'b0 ;
  assign y10276 = n20806 ;
  assign y10277 = ~n20807 ;
  assign y10278 = ~n20810 ;
  assign y10279 = ~n20811 ;
  assign y10280 = n20815 ;
  assign y10281 = n20816 ;
  assign y10282 = ~1'b0 ;
  assign y10283 = n20822 ;
  assign y10284 = ~n20824 ;
  assign y10285 = ~1'b0 ;
  assign y10286 = ~n20826 ;
  assign y10287 = n20827 ;
  assign y10288 = ~n20834 ;
  assign y10289 = ~n20836 ;
  assign y10290 = n20840 ;
  assign y10291 = n4218 ;
  assign y10292 = ~1'b0 ;
  assign y10293 = ~n20842 ;
  assign y10294 = n20843 ;
  assign y10295 = ~n20846 ;
  assign y10296 = ~n20847 ;
  assign y10297 = ~n20849 ;
  assign y10298 = ~n1244 ;
  assign y10299 = n20855 ;
  assign y10300 = ~n20857 ;
  assign y10301 = n20858 ;
  assign y10302 = ~n20861 ;
  assign y10303 = ~n20863 ;
  assign y10304 = ~1'b0 ;
  assign y10305 = n20864 ;
  assign y10306 = n20316 ;
  assign y10307 = ~1'b0 ;
  assign y10308 = ~n20867 ;
  assign y10309 = ~n20868 ;
  assign y10310 = n20869 ;
  assign y10311 = ~n20870 ;
  assign y10312 = n20872 ;
  assign y10313 = ~n16982 ;
  assign y10314 = ~n20874 ;
  assign y10315 = n20877 ;
  assign y10316 = ~n20886 ;
  assign y10317 = ~n20892 ;
  assign y10318 = ~1'b0 ;
  assign y10319 = ~1'b0 ;
  assign y10320 = ~n7749 ;
  assign y10321 = ~n20894 ;
  assign y10322 = ~1'b0 ;
  assign y10323 = ~n20898 ;
  assign y10324 = n20899 ;
  assign y10325 = n20900 ;
  assign y10326 = ~1'b0 ;
  assign y10327 = ~n20903 ;
  assign y10328 = n20904 ;
  assign y10329 = ~n20905 ;
  assign y10330 = ~1'b0 ;
  assign y10331 = ~n20906 ;
  assign y10332 = ~n20912 ;
  assign y10333 = ~n20923 ;
  assign y10334 = ~n20924 ;
  assign y10335 = ~1'b0 ;
  assign y10336 = n20929 ;
  assign y10337 = n688 ;
  assign y10338 = n20931 ;
  assign y10339 = n20940 ;
  assign y10340 = n20942 ;
  assign y10341 = ~n20834 ;
  assign y10342 = ~1'b0 ;
  assign y10343 = ~n20943 ;
  assign y10344 = ~1'b0 ;
  assign y10345 = n20949 ;
  assign y10346 = ~1'b0 ;
  assign y10347 = n20953 ;
  assign y10348 = n18062 ;
  assign y10349 = n20954 ;
  assign y10350 = ~1'b0 ;
  assign y10351 = n20955 ;
  assign y10352 = n20958 ;
  assign y10353 = ~n20961 ;
  assign y10354 = n20963 ;
  assign y10355 = n20965 ;
  assign y10356 = n20967 ;
  assign y10357 = ~n20968 ;
  assign y10358 = ~1'b0 ;
  assign y10359 = ~n20969 ;
  assign y10360 = ~n20971 ;
  assign y10361 = n20972 ;
  assign y10362 = n20975 ;
  assign y10363 = ~n20979 ;
  assign y10364 = ~n2141 ;
  assign y10365 = ~n20983 ;
  assign y10366 = n20984 ;
  assign y10367 = ~n20986 ;
  assign y10368 = n20988 ;
  assign y10369 = ~n20989 ;
  assign y10370 = n20991 ;
  assign y10371 = ~1'b0 ;
  assign y10372 = ~n20992 ;
  assign y10373 = n20994 ;
  assign y10374 = ~n20995 ;
  assign y10375 = ~1'b0 ;
  assign y10376 = ~n20996 ;
  assign y10377 = n21000 ;
  assign y10378 = n21003 ;
  assign y10379 = ~n21008 ;
  assign y10380 = ~n21010 ;
  assign y10381 = ~n21011 ;
  assign y10382 = n3054 ;
  assign y10383 = ~n21013 ;
  assign y10384 = ~n21016 ;
  assign y10385 = n21020 ;
  assign y10386 = n21024 ;
  assign y10387 = ~1'b0 ;
  assign y10388 = ~n21025 ;
  assign y10389 = ~1'b0 ;
  assign y10390 = n21029 ;
  assign y10391 = n21033 ;
  assign y10392 = n21034 ;
  assign y10393 = ~n21035 ;
  assign y10394 = n21037 ;
  assign y10395 = ~1'b0 ;
  assign y10396 = ~1'b0 ;
  assign y10397 = ~1'b0 ;
  assign y10398 = ~1'b0 ;
  assign y10399 = ~1'b0 ;
  assign y10400 = ~n21039 ;
  assign y10401 = ~n21044 ;
  assign y10402 = ~n7298 ;
  assign y10403 = ~n21046 ;
  assign y10404 = ~n21051 ;
  assign y10405 = ~1'b0 ;
  assign y10406 = ~n3380 ;
  assign y10407 = ~n21058 ;
  assign y10408 = ~1'b0 ;
  assign y10409 = ~1'b0 ;
  assign y10410 = ~n21059 ;
  assign y10411 = n21060 ;
  assign y10412 = ~1'b0 ;
  assign y10413 = n21062 ;
  assign y10414 = ~1'b0 ;
  assign y10415 = n21064 ;
  assign y10416 = ~n21068 ;
  assign y10417 = n21071 ;
  assign y10418 = x112 ;
  assign y10419 = ~1'b0 ;
  assign y10420 = n21074 ;
  assign y10421 = ~n21076 ;
  assign y10422 = ~1'b0 ;
  assign y10423 = ~1'b0 ;
  assign y10424 = ~n9684 ;
  assign y10425 = n21077 ;
  assign y10426 = n21078 ;
  assign y10427 = ~1'b0 ;
  assign y10428 = 1'b0 ;
  assign y10429 = ~n21080 ;
  assign y10430 = ~n21081 ;
  assign y10431 = n4673 ;
  assign y10432 = ~n21083 ;
  assign y10433 = ~n21085 ;
  assign y10434 = ~1'b0 ;
  assign y10435 = ~1'b0 ;
  assign y10436 = ~n21086 ;
  assign y10437 = n21089 ;
  assign y10438 = ~n21093 ;
  assign y10439 = ~1'b0 ;
  assign y10440 = ~1'b0 ;
  assign y10441 = ~1'b0 ;
  assign y10442 = ~n21098 ;
  assign y10443 = ~n21099 ;
  assign y10444 = n21101 ;
  assign y10445 = n21104 ;
  assign y10446 = ~n21106 ;
  assign y10447 = ~1'b0 ;
  assign y10448 = n14777 ;
  assign y10449 = ~n21108 ;
  assign y10450 = n21109 ;
  assign y10451 = ~n21112 ;
  assign y10452 = ~1'b0 ;
  assign y10453 = ~1'b0 ;
  assign y10454 = ~n21115 ;
  assign y10455 = n21116 ;
  assign y10456 = ~n21118 ;
  assign y10457 = ~n21120 ;
  assign y10458 = ~n21124 ;
  assign y10459 = ~n21128 ;
  assign y10460 = ~1'b0 ;
  assign y10461 = ~1'b0 ;
  assign y10462 = ~n21130 ;
  assign y10463 = ~n21135 ;
  assign y10464 = ~n21138 ;
  assign y10465 = ~1'b0 ;
  assign y10466 = n21139 ;
  assign y10467 = ~n21141 ;
  assign y10468 = ~1'b0 ;
  assign y10469 = ~n21143 ;
  assign y10470 = ~1'b0 ;
  assign y10471 = n21146 ;
  assign y10472 = ~n21147 ;
  assign y10473 = ~n21149 ;
  assign y10474 = ~1'b0 ;
  assign y10475 = ~n21153 ;
  assign y10476 = n21154 ;
  assign y10477 = ~1'b0 ;
  assign y10478 = ~n21155 ;
  assign y10479 = n21159 ;
  assign y10480 = ~n21160 ;
  assign y10481 = ~n12372 ;
  assign y10482 = ~1'b0 ;
  assign y10483 = n21166 ;
  assign y10484 = n21167 ;
  assign y10485 = n21168 ;
  assign y10486 = n21173 ;
  assign y10487 = n21174 ;
  assign y10488 = ~1'b0 ;
  assign y10489 = ~1'b0 ;
  assign y10490 = ~1'b0 ;
  assign y10491 = ~n21176 ;
  assign y10492 = ~1'b0 ;
  assign y10493 = n21177 ;
  assign y10494 = ~n6817 ;
  assign y10495 = n21178 ;
  assign y10496 = ~n21183 ;
  assign y10497 = ~n21185 ;
  assign y10498 = n21192 ;
  assign y10499 = ~1'b0 ;
  assign y10500 = n21196 ;
  assign y10501 = ~n21200 ;
  assign y10502 = ~n21201 ;
  assign y10503 = n21204 ;
  assign y10504 = ~1'b0 ;
  assign y10505 = n21207 ;
  assign y10506 = ~n21209 ;
  assign y10507 = n21212 ;
  assign y10508 = ~n21213 ;
  assign y10509 = n21215 ;
  assign y10510 = n21216 ;
  assign y10511 = n21220 ;
  assign y10512 = 1'b0 ;
  assign y10513 = ~1'b0 ;
  assign y10514 = n1129 ;
  assign y10515 = ~n21222 ;
  assign y10516 = ~n21224 ;
  assign y10517 = n21228 ;
  assign y10518 = n21230 ;
  assign y10519 = ~1'b0 ;
  assign y10520 = n21231 ;
  assign y10521 = ~n21232 ;
  assign y10522 = ~n21233 ;
  assign y10523 = ~1'b0 ;
  assign y10524 = ~1'b0 ;
  assign y10525 = ~1'b0 ;
  assign y10526 = n21235 ;
  assign y10527 = ~n21238 ;
  assign y10528 = n21240 ;
  assign y10529 = ~1'b0 ;
  assign y10530 = ~n21244 ;
  assign y10531 = ~1'b0 ;
  assign y10532 = n19797 ;
  assign y10533 = ~1'b0 ;
  assign y10534 = ~n21250 ;
  assign y10535 = ~n21251 ;
  assign y10536 = ~n4083 ;
  assign y10537 = ~n11541 ;
  assign y10538 = ~1'b0 ;
  assign y10539 = ~1'b0 ;
  assign y10540 = ~n21253 ;
  assign y10541 = ~1'b0 ;
  assign y10542 = ~n21257 ;
  assign y10543 = n21258 ;
  assign y10544 = n21259 ;
  assign y10545 = ~n21261 ;
  assign y10546 = n21263 ;
  assign y10547 = ~1'b0 ;
  assign y10548 = n11956 ;
  assign y10549 = n21264 ;
  assign y10550 = ~1'b0 ;
  assign y10551 = ~1'b0 ;
  assign y10552 = n21265 ;
  assign y10553 = n21271 ;
  assign y10554 = n21272 ;
  assign y10555 = n21273 ;
  assign y10556 = ~n21274 ;
  assign y10557 = n21280 ;
  assign y10558 = n21283 ;
  assign y10559 = ~n21285 ;
  assign y10560 = ~n21287 ;
  assign y10561 = ~n21292 ;
  assign y10562 = ~n21294 ;
  assign y10563 = ~n21295 ;
  assign y10564 = ~1'b0 ;
  assign y10565 = ~1'b0 ;
  assign y10566 = ~1'b0 ;
  assign y10567 = ~1'b0 ;
  assign y10568 = ~n21297 ;
  assign y10569 = 1'b0 ;
  assign y10570 = ~n14873 ;
  assign y10571 = ~n21299 ;
  assign y10572 = ~1'b0 ;
  assign y10573 = n21302 ;
  assign y10574 = ~1'b0 ;
  assign y10575 = ~n21303 ;
  assign y10576 = n21305 ;
  assign y10577 = n21307 ;
  assign y10578 = ~n21308 ;
  assign y10579 = n6414 ;
  assign y10580 = ~1'b0 ;
  assign y10581 = ~n21310 ;
  assign y10582 = n21317 ;
  assign y10583 = ~n21319 ;
  assign y10584 = ~n21325 ;
  assign y10585 = n21329 ;
  assign y10586 = ~n21332 ;
  assign y10587 = n21333 ;
  assign y10588 = ~n21336 ;
  assign y10589 = n21338 ;
  assign y10590 = n21340 ;
  assign y10591 = ~1'b0 ;
  assign y10592 = ~1'b0 ;
  assign y10593 = ~n21342 ;
  assign y10594 = ~n21346 ;
  assign y10595 = ~n21348 ;
  assign y10596 = ~n21349 ;
  assign y10597 = ~n21350 ;
  assign y10598 = n21351 ;
  assign y10599 = ~n21352 ;
  assign y10600 = n21357 ;
  assign y10601 = n21360 ;
  assign y10602 = ~1'b0 ;
  assign y10603 = ~n21368 ;
  assign y10604 = n21370 ;
  assign y10605 = n21371 ;
  assign y10606 = ~1'b0 ;
  assign y10607 = n21373 ;
  assign y10608 = ~1'b0 ;
  assign y10609 = ~n21375 ;
  assign y10610 = ~n21384 ;
  assign y10611 = ~1'b0 ;
  assign y10612 = ~n21386 ;
  assign y10613 = n21395 ;
  assign y10614 = ~1'b0 ;
  assign y10615 = n21396 ;
  assign y10616 = ~n14989 ;
  assign y10617 = ~n21398 ;
  assign y10618 = ~1'b0 ;
  assign y10619 = 1'b0 ;
  assign y10620 = ~1'b0 ;
  assign y10621 = 1'b0 ;
  assign y10622 = ~1'b0 ;
  assign y10623 = ~n21400 ;
  assign y10624 = n21401 ;
  assign y10625 = ~n21402 ;
  assign y10626 = ~n21409 ;
  assign y10627 = n21416 ;
  assign y10628 = ~n4711 ;
  assign y10629 = ~n21418 ;
  assign y10630 = ~n21419 ;
  assign y10631 = n21420 ;
  assign y10632 = n21421 ;
  assign y10633 = n10470 ;
  assign y10634 = n21422 ;
  assign y10635 = ~1'b0 ;
  assign y10636 = ~n21424 ;
  assign y10637 = n21430 ;
  assign y10638 = n21439 ;
  assign y10639 = ~n21444 ;
  assign y10640 = n21445 ;
  assign y10641 = n21447 ;
  assign y10642 = ~n21450 ;
  assign y10643 = n21455 ;
  assign y10644 = n21457 ;
  assign y10645 = ~1'b0 ;
  assign y10646 = ~n21459 ;
  assign y10647 = ~n21460 ;
  assign y10648 = ~1'b0 ;
  assign y10649 = ~n21462 ;
  assign y10650 = n21470 ;
  assign y10651 = ~n21473 ;
  assign y10652 = ~1'b0 ;
  assign y10653 = ~1'b0 ;
  assign y10654 = n21475 ;
  assign y10655 = ~1'b0 ;
  assign y10656 = ~n21477 ;
  assign y10657 = ~1'b0 ;
  assign y10658 = ~n21478 ;
  assign y10659 = ~1'b0 ;
  assign y10660 = ~n21480 ;
  assign y10661 = n21486 ;
  assign y10662 = ~1'b0 ;
  assign y10663 = ~1'b0 ;
  assign y10664 = n21488 ;
  assign y10665 = n21489 ;
  assign y10666 = ~1'b0 ;
  assign y10667 = ~1'b0 ;
  assign y10668 = ~1'b0 ;
  assign y10669 = ~n21495 ;
  assign y10670 = n21499 ;
  assign y10671 = ~1'b0 ;
  assign y10672 = n21500 ;
  assign y10673 = ~n21501 ;
  assign y10674 = n21503 ;
  assign y10675 = ~1'b0 ;
  assign y10676 = n21504 ;
  assign y10677 = n6204 ;
  assign y10678 = ~1'b0 ;
  assign y10679 = n21506 ;
  assign y10680 = ~1'b0 ;
  assign y10681 = ~1'b0 ;
  assign y10682 = ~1'b0 ;
  assign y10683 = ~n21513 ;
  assign y10684 = ~n21515 ;
  assign y10685 = ~n10961 ;
  assign y10686 = ~1'b0 ;
  assign y10687 = ~n21520 ;
  assign y10688 = n21524 ;
  assign y10689 = n21532 ;
  assign y10690 = n21533 ;
  assign y10691 = ~1'b0 ;
  assign y10692 = n21539 ;
  assign y10693 = n17456 ;
  assign y10694 = ~n21541 ;
  assign y10695 = ~1'b0 ;
  assign y10696 = ~n21545 ;
  assign y10697 = ~1'b0 ;
  assign y10698 = n21546 ;
  assign y10699 = ~1'b0 ;
  assign y10700 = ~1'b0 ;
  assign y10701 = n21551 ;
  assign y10702 = n21552 ;
  assign y10703 = ~n21553 ;
  assign y10704 = ~n21558 ;
  assign y10705 = n21562 ;
  assign y10706 = ~1'b0 ;
  assign y10707 = ~n12329 ;
  assign y10708 = ~n21563 ;
  assign y10709 = n21571 ;
  assign y10710 = n21574 ;
  assign y10711 = ~n6945 ;
  assign y10712 = n21576 ;
  assign y10713 = ~1'b0 ;
  assign y10714 = n18100 ;
  assign y10715 = ~1'b0 ;
  assign y10716 = ~1'b0 ;
  assign y10717 = 1'b0 ;
  assign y10718 = n19971 ;
  assign y10719 = ~n21579 ;
  assign y10720 = n21581 ;
  assign y10721 = n21583 ;
  assign y10722 = n21588 ;
  assign y10723 = ~n21592 ;
  assign y10724 = ~n21593 ;
  assign y10725 = n21596 ;
  assign y10726 = n21599 ;
  assign y10727 = ~n21608 ;
  assign y10728 = 1'b0 ;
  assign y10729 = ~n21610 ;
  assign y10730 = ~n21611 ;
  assign y10731 = ~n21613 ;
  assign y10732 = ~n21616 ;
  assign y10733 = ~1'b0 ;
  assign y10734 = ~1'b0 ;
  assign y10735 = ~x115 ;
  assign y10736 = n21617 ;
  assign y10737 = ~1'b0 ;
  assign y10738 = ~n21618 ;
  assign y10739 = ~1'b0 ;
  assign y10740 = ~n21620 ;
  assign y10741 = ~1'b0 ;
  assign y10742 = ~n21623 ;
  assign y10743 = ~n21625 ;
  assign y10744 = ~n21628 ;
  assign y10745 = ~1'b0 ;
  assign y10746 = ~n21631 ;
  assign y10747 = ~n4927 ;
  assign y10748 = ~1'b0 ;
  assign y10749 = ~n21634 ;
  assign y10750 = ~n21635 ;
  assign y10751 = n21639 ;
  assign y10752 = n21641 ;
  assign y10753 = ~n21645 ;
  assign y10754 = n21646 ;
  assign y10755 = ~n21651 ;
  assign y10756 = n21653 ;
  assign y10757 = ~n21655 ;
  assign y10758 = ~n21657 ;
  assign y10759 = n21658 ;
  assign y10760 = ~n21661 ;
  assign y10761 = ~1'b0 ;
  assign y10762 = ~n21663 ;
  assign y10763 = ~1'b0 ;
  assign y10764 = ~n21671 ;
  assign y10765 = ~n21673 ;
  assign y10766 = n21675 ;
  assign y10767 = 1'b0 ;
  assign y10768 = n21676 ;
  assign y10769 = ~1'b0 ;
  assign y10770 = ~n21682 ;
  assign y10771 = ~1'b0 ;
  assign y10772 = n21683 ;
  assign y10773 = ~n21684 ;
  assign y10774 = ~1'b0 ;
  assign y10775 = ~n21689 ;
  assign y10776 = ~1'b0 ;
  assign y10777 = n21694 ;
  assign y10778 = ~n21698 ;
  assign y10779 = ~n21699 ;
  assign y10780 = ~n21703 ;
  assign y10781 = n21705 ;
  assign y10782 = n21707 ;
  assign y10783 = ~1'b0 ;
  assign y10784 = n21710 ;
  assign y10785 = ~n21716 ;
  assign y10786 = ~1'b0 ;
  assign y10787 = ~n21718 ;
  assign y10788 = ~n21719 ;
  assign y10789 = n21721 ;
  assign y10790 = ~n21724 ;
  assign y10791 = ~n21728 ;
  assign y10792 = ~1'b0 ;
  assign y10793 = ~n21732 ;
  assign y10794 = n10516 ;
  assign y10795 = ~n9164 ;
  assign y10796 = n21736 ;
  assign y10797 = ~n21740 ;
  assign y10798 = n21741 ;
  assign y10799 = n21744 ;
  assign y10800 = ~n21751 ;
  assign y10801 = ~1'b0 ;
  assign y10802 = ~n15537 ;
  assign y10803 = ~n21753 ;
  assign y10804 = ~n21754 ;
  assign y10805 = ~n21755 ;
  assign y10806 = ~n21758 ;
  assign y10807 = ~n21761 ;
  assign y10808 = 1'b0 ;
  assign y10809 = ~1'b0 ;
  assign y10810 = ~n21763 ;
  assign y10811 = ~n21764 ;
  assign y10812 = ~1'b0 ;
  assign y10813 = ~n1379 ;
  assign y10814 = ~1'b0 ;
  assign y10815 = ~1'b0 ;
  assign y10816 = ~1'b0 ;
  assign y10817 = ~n8722 ;
  assign y10818 = ~1'b0 ;
  assign y10819 = ~n21770 ;
  assign y10820 = n21771 ;
  assign y10821 = ~1'b0 ;
  assign y10822 = ~n21772 ;
  assign y10823 = ~1'b0 ;
  assign y10824 = ~1'b0 ;
  assign y10825 = ~1'b0 ;
  assign y10826 = n21779 ;
  assign y10827 = n21782 ;
  assign y10828 = n21783 ;
  assign y10829 = n21786 ;
  assign y10830 = ~n21790 ;
  assign y10831 = ~1'b0 ;
  assign y10832 = ~n21792 ;
  assign y10833 = n21795 ;
  assign y10834 = n21796 ;
  assign y10835 = ~n3985 ;
  assign y10836 = ~n543 ;
  assign y10837 = ~n21797 ;
  assign y10838 = ~1'b0 ;
  assign y10839 = ~n21798 ;
  assign y10840 = ~n21804 ;
  assign y10841 = n20047 ;
  assign y10842 = ~1'b0 ;
  assign y10843 = n21805 ;
  assign y10844 = ~n6618 ;
  assign y10845 = n20152 ;
  assign y10846 = ~n21806 ;
  assign y10847 = n21810 ;
  assign y10848 = ~n21812 ;
  assign y10849 = ~n21813 ;
  assign y10850 = ~n21822 ;
  assign y10851 = n21826 ;
  assign y10852 = n21831 ;
  assign y10853 = ~1'b0 ;
  assign y10854 = ~n21833 ;
  assign y10855 = n21837 ;
  assign y10856 = ~n21838 ;
  assign y10857 = ~n21839 ;
  assign y10858 = ~n21844 ;
  assign y10859 = ~n21845 ;
  assign y10860 = ~1'b0 ;
  assign y10861 = ~1'b0 ;
  assign y10862 = n21847 ;
  assign y10863 = ~n21848 ;
  assign y10864 = ~n21851 ;
  assign y10865 = n21852 ;
  assign y10866 = ~n21856 ;
  assign y10867 = ~n21860 ;
  assign y10868 = ~n21861 ;
  assign y10869 = ~n21868 ;
  assign y10870 = n21869 ;
  assign y10871 = n21870 ;
  assign y10872 = n21875 ;
  assign y10873 = x123 ;
  assign y10874 = ~1'b0 ;
  assign y10875 = n21876 ;
  assign y10876 = ~1'b0 ;
  assign y10877 = ~1'b0 ;
  assign y10878 = ~n9814 ;
  assign y10879 = n21877 ;
  assign y10880 = ~1'b0 ;
  assign y10881 = ~n21304 ;
  assign y10882 = ~1'b0 ;
  assign y10883 = n21878 ;
  assign y10884 = ~n21880 ;
  assign y10885 = ~1'b0 ;
  assign y10886 = ~1'b0 ;
  assign y10887 = ~n21883 ;
  assign y10888 = ~n21884 ;
  assign y10889 = n4481 ;
  assign y10890 = n21888 ;
  assign y10891 = ~n21897 ;
  assign y10892 = n21898 ;
  assign y10893 = ~1'b0 ;
  assign y10894 = ~n21899 ;
  assign y10895 = ~n21903 ;
  assign y10896 = x251 ;
  assign y10897 = n21905 ;
  assign y10898 = ~1'b0 ;
  assign y10899 = ~1'b0 ;
  assign y10900 = ~n7996 ;
  assign y10901 = 1'b0 ;
  assign y10902 = n21907 ;
  assign y10903 = ~n21910 ;
  assign y10904 = ~n21912 ;
  assign y10905 = n21913 ;
  assign y10906 = ~n21914 ;
  assign y10907 = n17730 ;
  assign y10908 = ~n21921 ;
  assign y10909 = ~n21922 ;
  assign y10910 = ~n21924 ;
  assign y10911 = ~n21935 ;
  assign y10912 = ~n21937 ;
  assign y10913 = ~n21938 ;
  assign y10914 = ~1'b0 ;
  assign y10915 = ~1'b0 ;
  assign y10916 = ~1'b0 ;
  assign y10917 = ~n21939 ;
  assign y10918 = ~n21940 ;
  assign y10919 = ~1'b0 ;
  assign y10920 = ~n21948 ;
  assign y10921 = ~n21949 ;
  assign y10922 = ~1'b0 ;
  assign y10923 = ~n21950 ;
  assign y10924 = ~1'b0 ;
  assign y10925 = ~1'b0 ;
  assign y10926 = ~n21960 ;
  assign y10927 = n21962 ;
  assign y10928 = ~n21965 ;
  assign y10929 = n2701 ;
  assign y10930 = ~n21966 ;
  assign y10931 = ~n21969 ;
  assign y10932 = ~1'b0 ;
  assign y10933 = ~1'b0 ;
  assign y10934 = ~n21970 ;
  assign y10935 = n21971 ;
  assign y10936 = ~n21974 ;
  assign y10937 = ~n21977 ;
  assign y10938 = ~n21978 ;
  assign y10939 = ~n12305 ;
  assign y10940 = n17626 ;
  assign y10941 = ~n21980 ;
  assign y10942 = n21981 ;
  assign y10943 = ~n21985 ;
  assign y10944 = ~1'b0 ;
  assign y10945 = n21986 ;
  assign y10946 = ~n9336 ;
  assign y10947 = ~1'b0 ;
  assign y10948 = ~1'b0 ;
  assign y10949 = n1748 ;
  assign y10950 = ~n21988 ;
  assign y10951 = 1'b0 ;
  assign y10952 = n21989 ;
  assign y10953 = n21991 ;
  assign y10954 = ~n21997 ;
  assign y10955 = ~n22003 ;
  assign y10956 = ~1'b0 ;
  assign y10957 = n22004 ;
  assign y10958 = n22005 ;
  assign y10959 = n22008 ;
  assign y10960 = n22009 ;
  assign y10961 = ~n22010 ;
  assign y10962 = ~n22012 ;
  assign y10963 = ~1'b0 ;
  assign y10964 = n22014 ;
  assign y10965 = n22018 ;
  assign y10966 = ~n22023 ;
  assign y10967 = ~1'b0 ;
  assign y10968 = ~n22024 ;
  assign y10969 = n22027 ;
  assign y10970 = ~1'b0 ;
  assign y10971 = ~1'b0 ;
  assign y10972 = n22028 ;
  assign y10973 = ~n22029 ;
  assign y10974 = ~n22030 ;
  assign y10975 = n22031 ;
  assign y10976 = ~n22037 ;
  assign y10977 = n22039 ;
  assign y10978 = ~n22043 ;
  assign y10979 = ~n22047 ;
  assign y10980 = n22049 ;
  assign y10981 = ~n22050 ;
  assign y10982 = ~n22057 ;
  assign y10983 = n22060 ;
  assign y10984 = ~n22068 ;
  assign y10985 = ~1'b0 ;
  assign y10986 = n13032 ;
  assign y10987 = ~n22069 ;
  assign y10988 = ~n22071 ;
  assign y10989 = ~1'b0 ;
  assign y10990 = ~n22072 ;
  assign y10991 = n22073 ;
  assign y10992 = n22075 ;
  assign y10993 = ~1'b0 ;
  assign y10994 = ~1'b0 ;
  assign y10995 = n22077 ;
  assign y10996 = n22079 ;
  assign y10997 = n22083 ;
  assign y10998 = n22088 ;
  assign y10999 = n22090 ;
  assign y11000 = n22092 ;
  assign y11001 = n22094 ;
  assign y11002 = ~n22095 ;
  assign y11003 = ~1'b0 ;
  assign y11004 = ~1'b0 ;
  assign y11005 = ~n22097 ;
  assign y11006 = ~1'b0 ;
  assign y11007 = ~1'b0 ;
  assign y11008 = ~1'b0 ;
  assign y11009 = ~n22104 ;
  assign y11010 = n1307 ;
  assign y11011 = ~n14236 ;
  assign y11012 = ~n22109 ;
  assign y11013 = n4843 ;
  assign y11014 = ~n22111 ;
  assign y11015 = ~1'b0 ;
  assign y11016 = ~1'b0 ;
  assign y11017 = ~n22114 ;
  assign y11018 = n22119 ;
  assign y11019 = ~1'b0 ;
  assign y11020 = n22121 ;
  assign y11021 = ~1'b0 ;
  assign y11022 = n15498 ;
  assign y11023 = n8827 ;
  assign y11024 = ~1'b0 ;
  assign y11025 = ~1'b0 ;
  assign y11026 = n22122 ;
  assign y11027 = n22124 ;
  assign y11028 = ~1'b0 ;
  assign y11029 = ~1'b0 ;
  assign y11030 = n22126 ;
  assign y11031 = ~1'b0 ;
  assign y11032 = ~n22128 ;
  assign y11033 = ~1'b0 ;
  assign y11034 = ~1'b0 ;
  assign y11035 = ~n22131 ;
  assign y11036 = ~n22133 ;
  assign y11037 = n20888 ;
  assign y11038 = n22137 ;
  assign y11039 = n22138 ;
  assign y11040 = ~1'b0 ;
  assign y11041 = n22140 ;
  assign y11042 = ~n2264 ;
  assign y11043 = ~n22141 ;
  assign y11044 = n22142 ;
  assign y11045 = ~1'b0 ;
  assign y11046 = ~n22150 ;
  assign y11047 = n22151 ;
  assign y11048 = ~1'b0 ;
  assign y11049 = n10676 ;
  assign y11050 = ~1'b0 ;
  assign y11051 = ~1'b0 ;
  assign y11052 = ~n22152 ;
  assign y11053 = ~1'b0 ;
  assign y11054 = n22161 ;
  assign y11055 = ~1'b0 ;
  assign y11056 = ~n22165 ;
  assign y11057 = ~n22167 ;
  assign y11058 = n22168 ;
  assign y11059 = ~n12581 ;
  assign y11060 = n22171 ;
  assign y11061 = n22172 ;
  assign y11062 = n1749 ;
  assign y11063 = n22174 ;
  assign y11064 = n22180 ;
  assign y11065 = n15979 ;
  assign y11066 = ~n22181 ;
  assign y11067 = n22186 ;
  assign y11068 = n22188 ;
  assign y11069 = ~1'b0 ;
  assign y11070 = ~1'b0 ;
  assign y11071 = ~n22191 ;
  assign y11072 = ~n22194 ;
  assign y11073 = n22196 ;
  assign y11074 = ~n22198 ;
  assign y11075 = ~n22203 ;
  assign y11076 = ~1'b0 ;
  assign y11077 = ~n22206 ;
  assign y11078 = ~1'b0 ;
  assign y11079 = ~1'b0 ;
  assign y11080 = ~n22208 ;
  assign y11081 = n22210 ;
  assign y11082 = n22211 ;
  assign y11083 = ~n1708 ;
  assign y11084 = ~n22215 ;
  assign y11085 = ~n22220 ;
  assign y11086 = ~n22221 ;
  assign y11087 = ~n22223 ;
  assign y11088 = n16739 ;
  assign y11089 = ~n22226 ;
  assign y11090 = ~n22230 ;
  assign y11091 = ~n22233 ;
  assign y11092 = n22238 ;
  assign y11093 = ~n22239 ;
  assign y11094 = ~n22242 ;
  assign y11095 = ~1'b0 ;
  assign y11096 = ~1'b0 ;
  assign y11097 = ~n22251 ;
  assign y11098 = n22254 ;
  assign y11099 = ~n22258 ;
  assign y11100 = ~1'b0 ;
  assign y11101 = ~n22260 ;
  assign y11102 = ~1'b0 ;
  assign y11103 = n20673 ;
  assign y11104 = n22267 ;
  assign y11105 = ~1'b0 ;
  assign y11106 = ~1'b0 ;
  assign y11107 = n22268 ;
  assign y11108 = ~1'b0 ;
  assign y11109 = ~n18551 ;
  assign y11110 = ~1'b0 ;
  assign y11111 = ~n22270 ;
  assign y11112 = ~1'b0 ;
  assign y11113 = n22274 ;
  assign y11114 = ~1'b0 ;
  assign y11115 = n1628 ;
  assign y11116 = n22279 ;
  assign y11117 = ~n1926 ;
  assign y11118 = ~1'b0 ;
  assign y11119 = n22282 ;
  assign y11120 = n22283 ;
  assign y11121 = ~1'b0 ;
  assign y11122 = ~n16252 ;
  assign y11123 = n22285 ;
  assign y11124 = ~1'b0 ;
  assign y11125 = ~1'b0 ;
  assign y11126 = n22288 ;
  assign y11127 = n22290 ;
  assign y11128 = n22294 ;
  assign y11129 = ~n22298 ;
  assign y11130 = n1815 ;
  assign y11131 = ~n22301 ;
  assign y11132 = ~1'b0 ;
  assign y11133 = ~1'b0 ;
  assign y11134 = n22303 ;
  assign y11135 = ~n22305 ;
  assign y11136 = n22308 ;
  assign y11137 = ~n22309 ;
  assign y11138 = ~1'b0 ;
  assign y11139 = ~n22314 ;
  assign y11140 = n9241 ;
  assign y11141 = n22320 ;
  assign y11142 = 1'b0 ;
  assign y11143 = ~n22323 ;
  assign y11144 = n22326 ;
  assign y11145 = n22327 ;
  assign y11146 = ~n22328 ;
  assign y11147 = ~n22329 ;
  assign y11148 = ~1'b0 ;
  assign y11149 = ~n22331 ;
  assign y11150 = ~n22333 ;
  assign y11151 = ~1'b0 ;
  assign y11152 = ~n22335 ;
  assign y11153 = n22341 ;
  assign y11154 = n22346 ;
  assign y11155 = ~n22351 ;
  assign y11156 = ~1'b0 ;
  assign y11157 = ~n22354 ;
  assign y11158 = n22355 ;
  assign y11159 = ~n22359 ;
  assign y11160 = ~1'b0 ;
  assign y11161 = n22360 ;
  assign y11162 = ~1'b0 ;
  assign y11163 = ~1'b0 ;
  assign y11164 = ~n22362 ;
  assign y11165 = n20776 ;
  assign y11166 = ~n22363 ;
  assign y11167 = n22367 ;
  assign y11168 = n22369 ;
  assign y11169 = n22371 ;
  assign y11170 = ~1'b0 ;
  assign y11171 = ~n22372 ;
  assign y11172 = ~1'b0 ;
  assign y11173 = ~1'b0 ;
  assign y11174 = ~1'b0 ;
  assign y11175 = ~n22374 ;
  assign y11176 = ~1'b0 ;
  assign y11177 = ~n22375 ;
  assign y11178 = ~n22376 ;
  assign y11179 = ~n22379 ;
  assign y11180 = n22383 ;
  assign y11181 = ~n22385 ;
  assign y11182 = ~1'b0 ;
  assign y11183 = ~n583 ;
  assign y11184 = ~n22387 ;
  assign y11185 = ~1'b0 ;
  assign y11186 = n22388 ;
  assign y11187 = ~1'b0 ;
  assign y11188 = ~n22390 ;
  assign y11189 = ~n22393 ;
  assign y11190 = ~n22394 ;
  assign y11191 = ~n22401 ;
  assign y11192 = ~1'b0 ;
  assign y11193 = 1'b0 ;
  assign y11194 = n22404 ;
  assign y11195 = n22405 ;
  assign y11196 = ~n22408 ;
  assign y11197 = ~n20566 ;
  assign y11198 = ~1'b0 ;
  assign y11199 = n22409 ;
  assign y11200 = n22414 ;
  assign y11201 = ~n22416 ;
  assign y11202 = ~n22421 ;
  assign y11203 = n22427 ;
  assign y11204 = n10405 ;
  assign y11205 = ~n22428 ;
  assign y11206 = n22430 ;
  assign y11207 = ~1'b0 ;
  assign y11208 = ~n22438 ;
  assign y11209 = ~n10781 ;
  assign y11210 = ~1'b0 ;
  assign y11211 = ~1'b0 ;
  assign y11212 = ~n22441 ;
  assign y11213 = ~n22443 ;
  assign y11214 = ~1'b0 ;
  assign y11215 = n4325 ;
  assign y11216 = n22447 ;
  assign y11217 = ~1'b0 ;
  assign y11218 = ~1'b0 ;
  assign y11219 = n3894 ;
  assign y11220 = n22449 ;
  assign y11221 = ~1'b0 ;
  assign y11222 = n22451 ;
  assign y11223 = n22461 ;
  assign y11224 = ~n22462 ;
  assign y11225 = ~1'b0 ;
  assign y11226 = n22463 ;
  assign y11227 = n22464 ;
  assign y11228 = n22466 ;
  assign y11229 = n22468 ;
  assign y11230 = n22471 ;
  assign y11231 = n22482 ;
  assign y11232 = ~1'b0 ;
  assign y11233 = ~1'b0 ;
  assign y11234 = ~n13083 ;
  assign y11235 = ~1'b0 ;
  assign y11236 = ~n22486 ;
  assign y11237 = n22489 ;
  assign y11238 = n22491 ;
  assign y11239 = ~n22492 ;
  assign y11240 = ~n22494 ;
  assign y11241 = ~n22495 ;
  assign y11242 = ~n22496 ;
  assign y11243 = ~1'b0 ;
  assign y11244 = ~n22497 ;
  assign y11245 = ~n22498 ;
  assign y11246 = ~1'b0 ;
  assign y11247 = n22501 ;
  assign y11248 = ~n22504 ;
  assign y11249 = n22506 ;
  assign y11250 = ~1'b0 ;
  assign y11251 = ~n22507 ;
  assign y11252 = n22517 ;
  assign y11253 = n22519 ;
  assign y11254 = n22522 ;
  assign y11255 = n22525 ;
  assign y11256 = n22526 ;
  assign y11257 = n22528 ;
  assign y11258 = ~n22529 ;
  assign y11259 = n22536 ;
  assign y11260 = n22545 ;
  assign y11261 = n22549 ;
  assign y11262 = ~1'b0 ;
  assign y11263 = n22552 ;
  assign y11264 = ~1'b0 ;
  assign y11265 = ~n22554 ;
  assign y11266 = n22559 ;
  assign y11267 = ~n22560 ;
  assign y11268 = ~n22562 ;
  assign y11269 = ~n22564 ;
  assign y11270 = ~n22565 ;
  assign y11271 = n22567 ;
  assign y11272 = n22571 ;
  assign y11273 = ~n22574 ;
  assign y11274 = ~n22576 ;
  assign y11275 = ~1'b0 ;
  assign y11276 = ~1'b0 ;
  assign y11277 = ~1'b0 ;
  assign y11278 = ~n22578 ;
  assign y11279 = ~n22584 ;
  assign y11280 = ~n3134 ;
  assign y11281 = n22586 ;
  assign y11282 = n22589 ;
  assign y11283 = ~n22591 ;
  assign y11284 = 1'b0 ;
  assign y11285 = n14752 ;
  assign y11286 = ~n22594 ;
  assign y11287 = ~1'b0 ;
  assign y11288 = ~n22597 ;
  assign y11289 = n22598 ;
  assign y11290 = ~n22599 ;
  assign y11291 = n22601 ;
  assign y11292 = ~1'b0 ;
  assign y11293 = ~1'b0 ;
  assign y11294 = ~n22603 ;
  assign y11295 = n22605 ;
  assign y11296 = ~n22607 ;
  assign y11297 = ~n22612 ;
  assign y11298 = ~1'b0 ;
  assign y11299 = ~1'b0 ;
  assign y11300 = ~n22615 ;
  assign y11301 = 1'b0 ;
  assign y11302 = n22616 ;
  assign y11303 = ~1'b0 ;
  assign y11304 = ~1'b0 ;
  assign y11305 = ~1'b0 ;
  assign y11306 = ~n22618 ;
  assign y11307 = n22624 ;
  assign y11308 = ~n22625 ;
  assign y11309 = ~1'b0 ;
  assign y11310 = 1'b0 ;
  assign y11311 = ~1'b0 ;
  assign y11312 = n22628 ;
  assign y11313 = ~n22632 ;
  assign y11314 = ~n22639 ;
  assign y11315 = ~1'b0 ;
  assign y11316 = ~1'b0 ;
  assign y11317 = ~n22642 ;
  assign y11318 = n22647 ;
  assign y11319 = ~1'b0 ;
  assign y11320 = n22649 ;
  assign y11321 = n22650 ;
  assign y11322 = ~n22652 ;
  assign y11323 = ~n22655 ;
  assign y11324 = ~1'b0 ;
  assign y11325 = n22659 ;
  assign y11326 = n22660 ;
  assign y11327 = ~n22661 ;
  assign y11328 = n22662 ;
  assign y11329 = n22663 ;
  assign y11330 = ~1'b0 ;
  assign y11331 = 1'b0 ;
  assign y11332 = ~n21318 ;
  assign y11333 = ~n22666 ;
  assign y11334 = ~1'b0 ;
  assign y11335 = ~n22671 ;
  assign y11336 = ~n22674 ;
  assign y11337 = ~n22678 ;
  assign y11338 = n22682 ;
  assign y11339 = ~1'b0 ;
  assign y11340 = n22686 ;
  assign y11341 = ~n22688 ;
  assign y11342 = n22689 ;
  assign y11343 = ~n22690 ;
  assign y11344 = n15723 ;
  assign y11345 = ~n21096 ;
  assign y11346 = n22692 ;
  assign y11347 = ~1'b0 ;
  assign y11348 = n22695 ;
  assign y11349 = n22696 ;
  assign y11350 = ~1'b0 ;
  assign y11351 = ~n22697 ;
  assign y11352 = n22700 ;
  assign y11353 = ~n22703 ;
  assign y11354 = n22704 ;
  assign y11355 = n22712 ;
  assign y11356 = n22713 ;
  assign y11357 = n22715 ;
  assign y11358 = ~n22716 ;
  assign y11359 = ~n22717 ;
  assign y11360 = n7828 ;
  assign y11361 = n22719 ;
  assign y11362 = n22721 ;
  assign y11363 = n22723 ;
  assign y11364 = n22724 ;
  assign y11365 = ~n22728 ;
  assign y11366 = ~n22730 ;
  assign y11367 = 1'b0 ;
  assign y11368 = n22733 ;
  assign y11369 = ~1'b0 ;
  assign y11370 = ~1'b0 ;
  assign y11371 = ~n22735 ;
  assign y11372 = ~n22741 ;
  assign y11373 = n14259 ;
  assign y11374 = n22742 ;
  assign y11375 = n22745 ;
  assign y11376 = n4009 ;
  assign y11377 = ~n22747 ;
  assign y11378 = n22749 ;
  assign y11379 = n22752 ;
  assign y11380 = ~n22761 ;
  assign y11381 = ~n22762 ;
  assign y11382 = ~n22766 ;
  assign y11383 = ~n22768 ;
  assign y11384 = n417 ;
  assign y11385 = ~1'b0 ;
  assign y11386 = ~1'b0 ;
  assign y11387 = n22771 ;
  assign y11388 = ~1'b0 ;
  assign y11389 = n22772 ;
  assign y11390 = n6754 ;
  assign y11391 = ~1'b0 ;
  assign y11392 = ~1'b0 ;
  assign y11393 = n22774 ;
  assign y11394 = n22778 ;
  assign y11395 = n22780 ;
  assign y11396 = n22781 ;
  assign y11397 = ~n22782 ;
  assign y11398 = 1'b0 ;
  assign y11399 = ~1'b0 ;
  assign y11400 = ~n22789 ;
  assign y11401 = ~n22790 ;
  assign y11402 = ~n22791 ;
  assign y11403 = ~n22794 ;
  assign y11404 = n22796 ;
  assign y11405 = ~1'b0 ;
  assign y11406 = n22799 ;
  assign y11407 = ~n22803 ;
  assign y11408 = ~1'b0 ;
  assign y11409 = n22806 ;
  assign y11410 = n22808 ;
  assign y11411 = n22811 ;
  assign y11412 = n22815 ;
  assign y11413 = ~1'b0 ;
  assign y11414 = ~1'b0 ;
  assign y11415 = ~1'b0 ;
  assign y11416 = ~1'b0 ;
  assign y11417 = ~n22822 ;
  assign y11418 = ~1'b0 ;
  assign y11419 = ~n22825 ;
  assign y11420 = n22827 ;
  assign y11421 = 1'b0 ;
  assign y11422 = n22835 ;
  assign y11423 = n22836 ;
  assign y11424 = ~1'b0 ;
  assign y11425 = n22839 ;
  assign y11426 = ~1'b0 ;
  assign y11427 = ~1'b0 ;
  assign y11428 = n22841 ;
  assign y11429 = ~1'b0 ;
  assign y11430 = ~n22843 ;
  assign y11431 = n22846 ;
  assign y11432 = ~1'b0 ;
  assign y11433 = ~1'b0 ;
  assign y11434 = n22849 ;
  assign y11435 = ~n22850 ;
  assign y11436 = ~n6785 ;
  assign y11437 = ~1'b0 ;
  assign y11438 = ~n22852 ;
  assign y11439 = ~n22855 ;
  assign y11440 = n22859 ;
  assign y11441 = ~n22860 ;
  assign y11442 = n22861 ;
  assign y11443 = ~n22864 ;
  assign y11444 = n22865 ;
  assign y11445 = n22866 ;
  assign y11446 = ~1'b0 ;
  assign y11447 = 1'b0 ;
  assign y11448 = ~n21068 ;
  assign y11449 = ~n22868 ;
  assign y11450 = ~1'b0 ;
  assign y11451 = ~1'b0 ;
  assign y11452 = n22869 ;
  assign y11453 = n22871 ;
  assign y11454 = ~n22872 ;
  assign y11455 = ~n22876 ;
  assign y11456 = n22877 ;
  assign y11457 = n22885 ;
  assign y11458 = ~n22892 ;
  assign y11459 = ~1'b0 ;
  assign y11460 = ~1'b0 ;
  assign y11461 = ~1'b0 ;
  assign y11462 = ~n22894 ;
  assign y11463 = ~1'b0 ;
  assign y11464 = n22895 ;
  assign y11465 = n22896 ;
  assign y11466 = n22897 ;
  assign y11467 = ~1'b0 ;
  assign y11468 = ~1'b0 ;
  assign y11469 = ~n22898 ;
  assign y11470 = ~n22900 ;
  assign y11471 = ~1'b0 ;
  assign y11472 = n22903 ;
  assign y11473 = ~n22904 ;
  assign y11474 = n22912 ;
  assign y11475 = ~n22915 ;
  assign y11476 = ~n22917 ;
  assign y11477 = ~1'b0 ;
  assign y11478 = ~1'b0 ;
  assign y11479 = n22918 ;
  assign y11480 = ~n22919 ;
  assign y11481 = ~1'b0 ;
  assign y11482 = ~1'b0 ;
  assign y11483 = ~n22923 ;
  assign y11484 = ~1'b0 ;
  assign y11485 = ~n22925 ;
  assign y11486 = n22928 ;
  assign y11487 = ~n22940 ;
  assign y11488 = 1'b0 ;
  assign y11489 = ~n10690 ;
  assign y11490 = ~n22951 ;
  assign y11491 = ~n22952 ;
  assign y11492 = ~n22953 ;
  assign y11493 = ~n22957 ;
  assign y11494 = ~n22959 ;
  assign y11495 = ~n22967 ;
  assign y11496 = ~1'b0 ;
  assign y11497 = n22968 ;
  assign y11498 = n13097 ;
  assign y11499 = n22972 ;
  assign y11500 = n22979 ;
  assign y11501 = n22980 ;
  assign y11502 = n22981 ;
  assign y11503 = ~1'b0 ;
  assign y11504 = ~n22983 ;
  assign y11505 = ~n22984 ;
  assign y11506 = ~1'b0 ;
  assign y11507 = ~n22985 ;
  assign y11508 = ~n22987 ;
  assign y11509 = ~1'b0 ;
  assign y11510 = ~1'b0 ;
  assign y11511 = ~1'b0 ;
  assign y11512 = ~n22989 ;
  assign y11513 = n22991 ;
  assign y11514 = n22992 ;
  assign y11515 = ~1'b0 ;
  assign y11516 = ~1'b0 ;
  assign y11517 = ~n22996 ;
  assign y11518 = ~n18472 ;
  assign y11519 = ~n22483 ;
  assign y11520 = ~n22999 ;
  assign y11521 = ~1'b0 ;
  assign y11522 = n23001 ;
  assign y11523 = ~n23008 ;
  assign y11524 = n23013 ;
  assign y11525 = n23015 ;
  assign y11526 = ~n23020 ;
  assign y11527 = ~n23021 ;
  assign y11528 = ~n23022 ;
  assign y11529 = ~n23023 ;
  assign y11530 = ~n23027 ;
  assign y11531 = n23029 ;
  assign y11532 = ~n23032 ;
  assign y11533 = n23033 ;
  assign y11534 = n23037 ;
  assign y11535 = n692 ;
  assign y11536 = n23041 ;
  assign y11537 = ~n14666 ;
  assign y11538 = ~n23044 ;
  assign y11539 = ~n23046 ;
  assign y11540 = ~1'b0 ;
  assign y11541 = ~n18282 ;
  assign y11542 = n2950 ;
  assign y11543 = ~n23052 ;
  assign y11544 = n23055 ;
  assign y11545 = n23056 ;
  assign y11546 = ~n23057 ;
  assign y11547 = n23062 ;
  assign y11548 = ~1'b0 ;
  assign y11549 = n23063 ;
  assign y11550 = ~n23066 ;
  assign y11551 = n23070 ;
  assign y11552 = n21588 ;
  assign y11553 = ~n23072 ;
  assign y11554 = ~n23075 ;
  assign y11555 = ~n23076 ;
  assign y11556 = ~n23080 ;
  assign y11557 = ~n23082 ;
  assign y11558 = ~1'b0 ;
  assign y11559 = ~1'b0 ;
  assign y11560 = 1'b0 ;
  assign y11561 = ~1'b0 ;
  assign y11562 = ~n23087 ;
  assign y11563 = ~n23089 ;
  assign y11564 = ~1'b0 ;
  assign y11565 = ~1'b0 ;
  assign y11566 = ~n23090 ;
  assign y11567 = n23092 ;
  assign y11568 = ~n23093 ;
  assign y11569 = n23094 ;
  assign y11570 = n23095 ;
  assign y11571 = ~n23096 ;
  assign y11572 = n23100 ;
  assign y11573 = ~1'b0 ;
  assign y11574 = n23103 ;
  assign y11575 = n7018 ;
  assign y11576 = n23107 ;
  assign y11577 = n23113 ;
  assign y11578 = ~n23114 ;
  assign y11579 = ~1'b0 ;
  assign y11580 = ~1'b0 ;
  assign y11581 = ~1'b0 ;
  assign y11582 = n23115 ;
  assign y11583 = ~n23116 ;
  assign y11584 = ~n23118 ;
  assign y11585 = ~n23120 ;
  assign y11586 = ~1'b0 ;
  assign y11587 = n23121 ;
  assign y11588 = ~n23122 ;
  assign y11589 = ~n23129 ;
  assign y11590 = ~n23136 ;
  assign y11591 = ~1'b0 ;
  assign y11592 = ~n23141 ;
  assign y11593 = ~n23142 ;
  assign y11594 = ~n23143 ;
  assign y11595 = n23150 ;
  assign y11596 = n23152 ;
  assign y11597 = ~n23153 ;
  assign y11598 = n10944 ;
  assign y11599 = ~n23154 ;
  assign y11600 = ~n23155 ;
  assign y11601 = ~n23157 ;
  assign y11602 = n23159 ;
  assign y11603 = ~n23163 ;
  assign y11604 = ~n23164 ;
  assign y11605 = ~n23165 ;
  assign y11606 = ~n23166 ;
  assign y11607 = n23167 ;
  assign y11608 = ~n23172 ;
  assign y11609 = n23178 ;
  assign y11610 = ~n23181 ;
  assign y11611 = ~1'b0 ;
  assign y11612 = n23182 ;
  assign y11613 = n23188 ;
  assign y11614 = n23189 ;
  assign y11615 = n23190 ;
  assign y11616 = ~n23192 ;
  assign y11617 = n23194 ;
  assign y11618 = ~n23197 ;
  assign y11619 = ~n23200 ;
  assign y11620 = ~n23204 ;
  assign y11621 = ~n23206 ;
  assign y11622 = ~1'b0 ;
  assign y11623 = ~1'b0 ;
  assign y11624 = ~1'b0 ;
  assign y11625 = ~n23210 ;
  assign y11626 = ~1'b0 ;
  assign y11627 = ~n23212 ;
  assign y11628 = ~n23216 ;
  assign y11629 = ~1'b0 ;
  assign y11630 = n23217 ;
  assign y11631 = n23223 ;
  assign y11632 = ~n23226 ;
  assign y11633 = ~n23228 ;
  assign y11634 = n23236 ;
  assign y11635 = ~1'b0 ;
  assign y11636 = n19227 ;
  assign y11637 = ~n23239 ;
  assign y11638 = ~1'b0 ;
  assign y11639 = n23240 ;
  assign y11640 = ~1'b0 ;
  assign y11641 = ~n23241 ;
  assign y11642 = ~1'b0 ;
  assign y11643 = ~n23243 ;
  assign y11644 = n23245 ;
  assign y11645 = n23248 ;
  assign y11646 = n23250 ;
  assign y11647 = n23252 ;
  assign y11648 = ~n19292 ;
  assign y11649 = ~n23259 ;
  assign y11650 = ~n23261 ;
  assign y11651 = ~1'b0 ;
  assign y11652 = n23264 ;
  assign y11653 = ~n23265 ;
  assign y11654 = n23267 ;
  assign y11655 = ~n23268 ;
  assign y11656 = ~1'b0 ;
  assign y11657 = ~1'b0 ;
  assign y11658 = ~n14664 ;
  assign y11659 = n16519 ;
  assign y11660 = ~n23272 ;
  assign y11661 = ~1'b0 ;
  assign y11662 = ~n23273 ;
  assign y11663 = ~1'b0 ;
  assign y11664 = ~1'b0 ;
  assign y11665 = n23275 ;
  assign y11666 = n23277 ;
  assign y11667 = n23279 ;
  assign y11668 = ~1'b0 ;
  assign y11669 = ~1'b0 ;
  assign y11670 = ~1'b0 ;
  assign y11671 = ~n23281 ;
  assign y11672 = ~n23283 ;
  assign y11673 = ~1'b0 ;
  assign y11674 = ~n23287 ;
  assign y11675 = 1'b0 ;
  assign y11676 = n23290 ;
  assign y11677 = ~1'b0 ;
  assign y11678 = n23299 ;
  assign y11679 = n23301 ;
  assign y11680 = n23302 ;
  assign y11681 = ~1'b0 ;
  assign y11682 = n19370 ;
  assign y11683 = ~n23303 ;
  assign y11684 = n23305 ;
  assign y11685 = n23306 ;
  assign y11686 = n23307 ;
  assign y11687 = ~1'b0 ;
  assign y11688 = ~1'b0 ;
  assign y11689 = n23309 ;
  assign y11690 = ~n23311 ;
  assign y11691 = ~1'b0 ;
  assign y11692 = ~n23312 ;
  assign y11693 = ~1'b0 ;
  assign y11694 = ~1'b0 ;
  assign y11695 = n23314 ;
  assign y11696 = ~1'b0 ;
  assign y11697 = ~1'b0 ;
  assign y11698 = ~1'b0 ;
  assign y11699 = n23316 ;
  assign y11700 = ~1'b0 ;
  assign y11701 = n16609 ;
  assign y11702 = n23319 ;
  assign y11703 = n23322 ;
  assign y11704 = n23324 ;
  assign y11705 = ~1'b0 ;
  assign y11706 = ~n23330 ;
  assign y11707 = n23331 ;
  assign y11708 = ~n23332 ;
  assign y11709 = n23337 ;
  assign y11710 = n23338 ;
  assign y11711 = n23339 ;
  assign y11712 = ~n23340 ;
  assign y11713 = ~n23341 ;
  assign y11714 = n23350 ;
  assign y11715 = ~1'b0 ;
  assign y11716 = ~n23353 ;
  assign y11717 = ~n23356 ;
  assign y11718 = ~n537 ;
  assign y11719 = n23359 ;
  assign y11720 = n23361 ;
  assign y11721 = n23364 ;
  assign y11722 = ~n7998 ;
  assign y11723 = ~n23365 ;
  assign y11724 = ~n23366 ;
  assign y11725 = n23367 ;
  assign y11726 = ~1'b0 ;
  assign y11727 = ~n23370 ;
  assign y11728 = ~n23374 ;
  assign y11729 = ~n23377 ;
  assign y11730 = ~n23378 ;
  assign y11731 = n23380 ;
  assign y11732 = ~1'b0 ;
  assign y11733 = ~1'b0 ;
  assign y11734 = ~n23381 ;
  assign y11735 = n23383 ;
  assign y11736 = ~n23384 ;
  assign y11737 = n23388 ;
  assign y11738 = n23392 ;
  assign y11739 = ~n23393 ;
  assign y11740 = ~n23395 ;
  assign y11741 = ~n23398 ;
  assign y11742 = ~n23404 ;
  assign y11743 = ~1'b0 ;
  assign y11744 = n23408 ;
  assign y11745 = ~n23411 ;
  assign y11746 = ~1'b0 ;
  assign y11747 = n23413 ;
  assign y11748 = ~1'b0 ;
  assign y11749 = ~1'b0 ;
  assign y11750 = ~n23416 ;
  assign y11751 = ~1'b0 ;
  assign y11752 = ~1'b0 ;
  assign y11753 = n6113 ;
  assign y11754 = ~1'b0 ;
  assign y11755 = ~n23418 ;
  assign y11756 = ~n23419 ;
  assign y11757 = n23421 ;
  assign y11758 = n13620 ;
  assign y11759 = ~n23423 ;
  assign y11760 = ~1'b0 ;
  assign y11761 = ~n23425 ;
  assign y11762 = ~n23426 ;
  assign y11763 = n23428 ;
  assign y11764 = ~n23432 ;
  assign y11765 = ~n4010 ;
  assign y11766 = ~n23435 ;
  assign y11767 = 1'b0 ;
  assign y11768 = ~n23438 ;
  assign y11769 = n23441 ;
  assign y11770 = n23442 ;
  assign y11771 = ~n1966 ;
  assign y11772 = n23444 ;
  assign y11773 = ~n23449 ;
  assign y11774 = n23451 ;
  assign y11775 = n23452 ;
  assign y11776 = n23456 ;
  assign y11777 = n19503 ;
  assign y11778 = ~n23459 ;
  assign y11779 = ~n23461 ;
  assign y11780 = ~1'b0 ;
  assign y11781 = ~n23465 ;
  assign y11782 = ~n23466 ;
  assign y11783 = ~1'b0 ;
  assign y11784 = n23467 ;
  assign y11785 = ~n23470 ;
  assign y11786 = n23471 ;
  assign y11787 = n23472 ;
  assign y11788 = ~n23476 ;
  assign y11789 = ~n23477 ;
  assign y11790 = ~1'b0 ;
  assign y11791 = n23487 ;
  assign y11792 = n23488 ;
  assign y11793 = n23491 ;
  assign y11794 = 1'b0 ;
  assign y11795 = n23493 ;
  assign y11796 = ~n23495 ;
  assign y11797 = ~n23496 ;
  assign y11798 = ~1'b0 ;
  assign y11799 = ~1'b0 ;
  assign y11800 = ~1'b0 ;
  assign y11801 = ~1'b0 ;
  assign y11802 = ~1'b0 ;
  assign y11803 = n23498 ;
  assign y11804 = n23502 ;
  assign y11805 = ~1'b0 ;
  assign y11806 = n23507 ;
  assign y11807 = n23508 ;
  assign y11808 = n23515 ;
  assign y11809 = ~1'b0 ;
  assign y11810 = ~n23519 ;
  assign y11811 = ~n23520 ;
  assign y11812 = n23521 ;
  assign y11813 = ~1'b0 ;
  assign y11814 = ~1'b0 ;
  assign y11815 = ~1'b0 ;
  assign y11816 = 1'b0 ;
  assign y11817 = n23528 ;
  assign y11818 = ~n23529 ;
  assign y11819 = ~1'b0 ;
  assign y11820 = ~n13714 ;
  assign y11821 = ~1'b0 ;
  assign y11822 = ~1'b0 ;
  assign y11823 = ~n23531 ;
  assign y11824 = n23532 ;
  assign y11825 = ~1'b0 ;
  assign y11826 = n23534 ;
  assign y11827 = ~1'b0 ;
  assign y11828 = n14752 ;
  assign y11829 = ~n23536 ;
  assign y11830 = ~n23540 ;
  assign y11831 = n17275 ;
  assign y11832 = n23543 ;
  assign y11833 = ~n23545 ;
  assign y11834 = ~n23546 ;
  assign y11835 = ~1'b0 ;
  assign y11836 = ~n6602 ;
  assign y11837 = ~1'b0 ;
  assign y11838 = ~1'b0 ;
  assign y11839 = ~n23547 ;
  assign y11840 = ~n23549 ;
  assign y11841 = ~1'b0 ;
  assign y11842 = ~n14143 ;
  assign y11843 = ~1'b0 ;
  assign y11844 = ~n23551 ;
  assign y11845 = ~1'b0 ;
  assign y11846 = ~n23553 ;
  assign y11847 = ~1'b0 ;
  assign y11848 = ~1'b0 ;
  assign y11849 = ~n23556 ;
  assign y11850 = ~n23561 ;
  assign y11851 = ~n14698 ;
  assign y11852 = ~n23569 ;
  assign y11853 = ~n23571 ;
  assign y11854 = ~1'b0 ;
  assign y11855 = ~n23577 ;
  assign y11856 = ~n469 ;
  assign y11857 = n2049 ;
  assign y11858 = n23581 ;
  assign y11859 = ~1'b0 ;
  assign y11860 = n23583 ;
  assign y11861 = ~1'b0 ;
  assign y11862 = ~n23587 ;
  assign y11863 = ~1'b0 ;
  assign y11864 = n23588 ;
  assign y11865 = ~1'b0 ;
  assign y11866 = ~n23589 ;
  assign y11867 = ~1'b0 ;
  assign y11868 = ~1'b0 ;
  assign y11869 = n23592 ;
  assign y11870 = n23594 ;
  assign y11871 = ~n23598 ;
  assign y11872 = ~n23601 ;
  assign y11873 = n23602 ;
  assign y11874 = n23604 ;
  assign y11875 = ~1'b0 ;
  assign y11876 = 1'b0 ;
  assign y11877 = ~n23605 ;
  assign y11878 = ~n23609 ;
  assign y11879 = ~n23610 ;
  assign y11880 = ~1'b0 ;
  assign y11881 = ~1'b0 ;
  assign y11882 = n23613 ;
  assign y11883 = ~1'b0 ;
  assign y11884 = ~n1917 ;
  assign y11885 = ~n23617 ;
  assign y11886 = n23621 ;
  assign y11887 = 1'b0 ;
  assign y11888 = ~n23623 ;
  assign y11889 = ~n23635 ;
  assign y11890 = n23640 ;
  assign y11891 = n23641 ;
  assign y11892 = ~1'b0 ;
  assign y11893 = ~n23647 ;
  assign y11894 = ~1'b0 ;
  assign y11895 = ~1'b0 ;
  assign y11896 = 1'b0 ;
  assign y11897 = n15015 ;
  assign y11898 = ~n23649 ;
  assign y11899 = ~n23651 ;
  assign y11900 = ~1'b0 ;
  assign y11901 = ~n23652 ;
  assign y11902 = n23655 ;
  assign y11903 = ~1'b0 ;
  assign y11904 = ~n23657 ;
  assign y11905 = n23658 ;
  assign y11906 = ~n23660 ;
  assign y11907 = n23663 ;
  assign y11908 = ~1'b0 ;
  assign y11909 = ~1'b0 ;
  assign y11910 = n23664 ;
  assign y11911 = ~n23665 ;
  assign y11912 = ~1'b0 ;
  assign y11913 = ~n23671 ;
  assign y11914 = ~1'b0 ;
  assign y11915 = ~1'b0 ;
  assign y11916 = ~n23673 ;
  assign y11917 = n23674 ;
  assign y11918 = ~1'b0 ;
  assign y11919 = ~1'b0 ;
  assign y11920 = n9907 ;
  assign y11921 = ~1'b0 ;
  assign y11922 = n23679 ;
  assign y11923 = ~n23683 ;
  assign y11924 = ~1'b0 ;
  assign y11925 = ~1'b0 ;
  assign y11926 = ~n23684 ;
  assign y11927 = n23690 ;
  assign y11928 = ~1'b0 ;
  assign y11929 = ~n23694 ;
  assign y11930 = ~1'b0 ;
  assign y11931 = ~n23695 ;
  assign y11932 = ~n23698 ;
  assign y11933 = ~1'b0 ;
  assign y11934 = n23702 ;
  assign y11935 = ~1'b0 ;
  assign y11936 = n23706 ;
  assign y11937 = ~1'b0 ;
  assign y11938 = ~n23709 ;
  assign y11939 = ~n23713 ;
  assign y11940 = 1'b0 ;
  assign y11941 = n23715 ;
  assign y11942 = ~1'b0 ;
  assign y11943 = ~1'b0 ;
  assign y11944 = ~n23716 ;
  assign y11945 = n23722 ;
  assign y11946 = ~n23725 ;
  assign y11947 = ~n23729 ;
  assign y11948 = n23731 ;
  assign y11949 = ~1'b0 ;
  assign y11950 = n23732 ;
  assign y11951 = ~n23739 ;
  assign y11952 = ~1'b0 ;
  assign y11953 = ~1'b0 ;
  assign y11954 = ~n23741 ;
  assign y11955 = n23742 ;
  assign y11956 = ~1'b0 ;
  assign y11957 = n23743 ;
  assign y11958 = ~1'b0 ;
  assign y11959 = ~n23745 ;
  assign y11960 = n23746 ;
  assign y11961 = ~n23747 ;
  assign y11962 = n23748 ;
  assign y11963 = ~1'b0 ;
  assign y11964 = n23749 ;
  assign y11965 = ~1'b0 ;
  assign y11966 = n23750 ;
  assign y11967 = ~1'b0 ;
  assign y11968 = ~1'b0 ;
  assign y11969 = ~n23752 ;
  assign y11970 = ~1'b0 ;
  assign y11971 = ~1'b0 ;
  assign y11972 = ~1'b0 ;
  assign y11973 = ~n23753 ;
  assign y11974 = ~n23755 ;
  assign y11975 = ~1'b0 ;
  assign y11976 = n23759 ;
  assign y11977 = ~1'b0 ;
  assign y11978 = ~1'b0 ;
  assign y11979 = n23768 ;
  assign y11980 = ~n23772 ;
  assign y11981 = ~n23773 ;
  assign y11982 = ~n23775 ;
  assign y11983 = ~n23777 ;
  assign y11984 = n23784 ;
  assign y11985 = n23787 ;
  assign y11986 = ~1'b0 ;
  assign y11987 = ~n23793 ;
  assign y11988 = ~n23794 ;
  assign y11989 = ~1'b0 ;
  assign y11990 = ~1'b0 ;
  assign y11991 = ~1'b0 ;
  assign y11992 = ~n11633 ;
  assign y11993 = n23796 ;
  assign y11994 = ~1'b0 ;
  assign y11995 = ~n23798 ;
  assign y11996 = ~1'b0 ;
  assign y11997 = ~1'b0 ;
  assign y11998 = ~n23800 ;
  assign y11999 = ~n20450 ;
  assign y12000 = ~n23803 ;
  assign y12001 = ~n23807 ;
  assign y12002 = n23808 ;
  assign y12003 = ~n23810 ;
  assign y12004 = ~n23813 ;
  assign y12005 = ~n23816 ;
  assign y12006 = ~n23827 ;
  assign y12007 = n23828 ;
  assign y12008 = ~1'b0 ;
  assign y12009 = n23832 ;
  assign y12010 = n23835 ;
  assign y12011 = 1'b0 ;
  assign y12012 = n23837 ;
  assign y12013 = n23839 ;
  assign y12014 = ~1'b0 ;
  assign y12015 = ~n23842 ;
  assign y12016 = ~1'b0 ;
  assign y12017 = n23848 ;
  assign y12018 = n23849 ;
  assign y12019 = n23850 ;
  assign y12020 = ~1'b0 ;
  assign y12021 = n23854 ;
  assign y12022 = ~n23858 ;
  assign y12023 = ~n23862 ;
  assign y12024 = ~1'b0 ;
  assign y12025 = ~1'b0 ;
  assign y12026 = ~n23871 ;
  assign y12027 = n23879 ;
  assign y12028 = x116 ;
  assign y12029 = ~1'b0 ;
  assign y12030 = ~n23880 ;
  assign y12031 = n23881 ;
  assign y12032 = ~n23886 ;
  assign y12033 = n23888 ;
  assign y12034 = ~1'b0 ;
  assign y12035 = ~n23889 ;
  assign y12036 = ~n23890 ;
  assign y12037 = n23893 ;
  assign y12038 = n23895 ;
  assign y12039 = ~1'b0 ;
  assign y12040 = ~n23896 ;
  assign y12041 = n13354 ;
  assign y12042 = n23905 ;
  assign y12043 = ~1'b0 ;
  assign y12044 = ~n23909 ;
  assign y12045 = n23911 ;
  assign y12046 = ~1'b0 ;
  assign y12047 = n23933 ;
  assign y12048 = ~1'b0 ;
  assign y12049 = n23934 ;
  assign y12050 = ~1'b0 ;
  assign y12051 = ~n23936 ;
  assign y12052 = ~1'b0 ;
  assign y12053 = ~n23937 ;
  assign y12054 = ~1'b0 ;
  assign y12055 = ~n23938 ;
  assign y12056 = ~n23939 ;
  assign y12057 = n23940 ;
  assign y12058 = ~1'b0 ;
  assign y12059 = n23942 ;
  assign y12060 = ~1'b0 ;
  assign y12061 = n23946 ;
  assign y12062 = ~n23947 ;
  assign y12063 = ~1'b0 ;
  assign y12064 = ~n23949 ;
  assign y12065 = n23959 ;
  assign y12066 = ~n23961 ;
  assign y12067 = ~n23962 ;
  assign y12068 = n23965 ;
  assign y12069 = ~1'b0 ;
  assign y12070 = n23968 ;
  assign y12071 = n23970 ;
  assign y12072 = n23972 ;
  assign y12073 = ~n23974 ;
  assign y12074 = n23977 ;
  assign y12075 = ~n23978 ;
  assign y12076 = n23979 ;
  assign y12077 = n23980 ;
  assign y12078 = ~n23982 ;
  assign y12079 = ~n23985 ;
  assign y12080 = ~n23987 ;
  assign y12081 = n23989 ;
  assign y12082 = ~n5746 ;
  assign y12083 = ~1'b0 ;
  assign y12084 = n23992 ;
  assign y12085 = ~1'b0 ;
  assign y12086 = ~1'b0 ;
  assign y12087 = n23995 ;
  assign y12088 = n23997 ;
  assign y12089 = ~n24002 ;
  assign y12090 = ~1'b0 ;
  assign y12091 = n24004 ;
  assign y12092 = ~1'b0 ;
  assign y12093 = n24005 ;
  assign y12094 = ~1'b0 ;
  assign y12095 = ~1'b0 ;
  assign y12096 = n24007 ;
  assign y12097 = ~1'b0 ;
  assign y12098 = n23184 ;
  assign y12099 = ~1'b0 ;
  assign y12100 = ~n24009 ;
  assign y12101 = ~n24015 ;
  assign y12102 = ~n24017 ;
  assign y12103 = n24018 ;
  assign y12104 = n6565 ;
  assign y12105 = ~n24022 ;
  assign y12106 = ~n24024 ;
  assign y12107 = ~1'b0 ;
  assign y12108 = n24025 ;
  assign y12109 = ~n24026 ;
  assign y12110 = n24027 ;
  assign y12111 = n24028 ;
  assign y12112 = ~1'b0 ;
  assign y12113 = ~n24034 ;
  assign y12114 = n24036 ;
  assign y12115 = n24039 ;
  assign y12116 = n24040 ;
  assign y12117 = n24047 ;
  assign y12118 = n24048 ;
  assign y12119 = n24050 ;
  assign y12120 = ~1'b0 ;
  assign y12121 = n24051 ;
  assign y12122 = ~n24055 ;
  assign y12123 = ~n24058 ;
  assign y12124 = n24059 ;
  assign y12125 = ~n24062 ;
  assign y12126 = ~1'b0 ;
  assign y12127 = ~n24063 ;
  assign y12128 = ~n24065 ;
  assign y12129 = ~n24067 ;
  assign y12130 = ~n24069 ;
  assign y12131 = n24072 ;
  assign y12132 = ~1'b0 ;
  assign y12133 = ~1'b0 ;
  assign y12134 = ~1'b0 ;
  assign y12135 = ~n24074 ;
  assign y12136 = ~1'b0 ;
  assign y12137 = ~1'b0 ;
  assign y12138 = ~1'b0 ;
  assign y12139 = n24076 ;
  assign y12140 = ~1'b0 ;
  assign y12141 = ~n24082 ;
  assign y12142 = n24083 ;
  assign y12143 = ~n24086 ;
  assign y12144 = ~1'b0 ;
  assign y12145 = ~1'b0 ;
  assign y12146 = n24087 ;
  assign y12147 = ~n3036 ;
  assign y12148 = ~n24089 ;
  assign y12149 = ~n24093 ;
  assign y12150 = ~n24094 ;
  assign y12151 = n24095 ;
  assign y12152 = n24101 ;
  assign y12153 = ~1'b0 ;
  assign y12154 = n24102 ;
  assign y12155 = ~1'b0 ;
  assign y12156 = ~n24103 ;
  assign y12157 = ~1'b0 ;
  assign y12158 = n24105 ;
  assign y12159 = ~1'b0 ;
  assign y12160 = ~n24107 ;
  assign y12161 = ~n16252 ;
  assign y12162 = n24121 ;
  assign y12163 = ~n24124 ;
  assign y12164 = ~1'b0 ;
  assign y12165 = ~1'b0 ;
  assign y12166 = n24125 ;
  assign y12167 = ~n24126 ;
  assign y12168 = ~n10174 ;
  assign y12169 = ~n24129 ;
  assign y12170 = ~n3189 ;
  assign y12171 = n24130 ;
  assign y12172 = 1'b0 ;
  assign y12173 = ~1'b0 ;
  assign y12174 = ~1'b0 ;
  assign y12175 = ~1'b0 ;
  assign y12176 = ~n24133 ;
  assign y12177 = ~n1859 ;
  assign y12178 = n24135 ;
  assign y12179 = n24138 ;
  assign y12180 = ~n24142 ;
  assign y12181 = n24143 ;
  assign y12182 = ~1'b0 ;
  assign y12183 = ~n24145 ;
  assign y12184 = ~1'b0 ;
  assign y12185 = ~n24148 ;
  assign y12186 = ~1'b0 ;
  assign y12187 = ~n24150 ;
  assign y12188 = ~n24152 ;
  assign y12189 = ~n24158 ;
  assign y12190 = ~n24161 ;
  assign y12191 = ~1'b0 ;
  assign y12192 = ~1'b0 ;
  assign y12193 = n14949 ;
  assign y12194 = ~n24164 ;
  assign y12195 = ~n24165 ;
  assign y12196 = ~n24166 ;
  assign y12197 = n24173 ;
  assign y12198 = ~n24175 ;
  assign y12199 = ~n645 ;
  assign y12200 = n24178 ;
  assign y12201 = ~1'b0 ;
  assign y12202 = ~1'b0 ;
  assign y12203 = n24180 ;
  assign y12204 = n3823 ;
  assign y12205 = ~1'b0 ;
  assign y12206 = n24184 ;
  assign y12207 = 1'b0 ;
  assign y12208 = ~n24186 ;
  assign y12209 = ~1'b0 ;
  assign y12210 = ~1'b0 ;
  assign y12211 = n24187 ;
  assign y12212 = n24190 ;
  assign y12213 = ~1'b0 ;
  assign y12214 = ~n24191 ;
  assign y12215 = ~1'b0 ;
  assign y12216 = ~n24196 ;
  assign y12217 = ~n7029 ;
  assign y12218 = n24201 ;
  assign y12219 = ~1'b0 ;
  assign y12220 = ~n24204 ;
  assign y12221 = ~1'b0 ;
  assign y12222 = n24206 ;
  assign y12223 = ~n24209 ;
  assign y12224 = n24211 ;
  assign y12225 = ~n24212 ;
  assign y12226 = ~n24217 ;
  assign y12227 = n24220 ;
  assign y12228 = n24224 ;
  assign y12229 = ~n24226 ;
  assign y12230 = ~n9290 ;
  assign y12231 = n24235 ;
  assign y12232 = ~1'b0 ;
  assign y12233 = ~n24239 ;
  assign y12234 = n24243 ;
  assign y12235 = ~1'b0 ;
  assign y12236 = n3400 ;
  assign y12237 = 1'b0 ;
  assign y12238 = n24244 ;
  assign y12239 = ~1'b0 ;
  assign y12240 = ~1'b0 ;
  assign y12241 = ~1'b0 ;
  assign y12242 = ~n24245 ;
  assign y12243 = ~n24249 ;
  assign y12244 = ~1'b0 ;
  assign y12245 = 1'b0 ;
  assign y12246 = ~n24252 ;
  assign y12247 = n24256 ;
  assign y12248 = ~1'b0 ;
  assign y12249 = ~n24259 ;
  assign y12250 = ~n24260 ;
  assign y12251 = ~n24264 ;
  assign y12252 = n9782 ;
  assign y12253 = n24265 ;
  assign y12254 = ~1'b0 ;
  assign y12255 = ~n24269 ;
  assign y12256 = ~n19704 ;
  assign y12257 = n24271 ;
  assign y12258 = ~n24273 ;
  assign y12259 = ~1'b0 ;
  assign y12260 = n24277 ;
  assign y12261 = n24278 ;
  assign y12262 = n24283 ;
  assign y12263 = n24287 ;
  assign y12264 = ~1'b0 ;
  assign y12265 = n24288 ;
  assign y12266 = n19148 ;
  assign y12267 = n24289 ;
  assign y12268 = n24291 ;
  assign y12269 = ~1'b0 ;
  assign y12270 = n24294 ;
  assign y12271 = ~n24295 ;
  assign y12272 = n24299 ;
  assign y12273 = ~n24300 ;
  assign y12274 = ~n24302 ;
  assign y12275 = n24303 ;
  assign y12276 = n24305 ;
  assign y12277 = ~1'b0 ;
  assign y12278 = n24309 ;
  assign y12279 = ~n24310 ;
  assign y12280 = ~n24315 ;
  assign y12281 = n24319 ;
  assign y12282 = ~1'b0 ;
  assign y12283 = ~1'b0 ;
  assign y12284 = ~n23891 ;
  assign y12285 = n24320 ;
  assign y12286 = ~n24321 ;
  assign y12287 = ~1'b0 ;
  assign y12288 = ~n24326 ;
  assign y12289 = ~1'b0 ;
  assign y12290 = ~n874 ;
  assign y12291 = n24328 ;
  assign y12292 = n24329 ;
  assign y12293 = ~n24335 ;
  assign y12294 = ~1'b0 ;
  assign y12295 = ~1'b0 ;
  assign y12296 = ~n24337 ;
  assign y12297 = n24338 ;
  assign y12298 = n24340 ;
  assign y12299 = ~n24342 ;
  assign y12300 = n24346 ;
  assign y12301 = ~n24351 ;
  assign y12302 = ~n24354 ;
  assign y12303 = ~n24357 ;
  assign y12304 = n24358 ;
  assign y12305 = ~1'b0 ;
  assign y12306 = ~1'b0 ;
  assign y12307 = ~n24360 ;
  assign y12308 = ~1'b0 ;
  assign y12309 = ~1'b0 ;
  assign y12310 = ~1'b0 ;
  assign y12311 = ~n24363 ;
  assign y12312 = ~n16177 ;
  assign y12313 = ~n24366 ;
  assign y12314 = ~n24368 ;
  assign y12315 = ~1'b0 ;
  assign y12316 = ~n24369 ;
  assign y12317 = ~n24370 ;
  assign y12318 = n24371 ;
  assign y12319 = n24372 ;
  assign y12320 = ~1'b0 ;
  assign y12321 = n24373 ;
  assign y12322 = ~n23396 ;
  assign y12323 = n24376 ;
  assign y12324 = n24377 ;
  assign y12325 = ~1'b0 ;
  assign y12326 = ~1'b0 ;
  assign y12327 = n24379 ;
  assign y12328 = x35 ;
  assign y12329 = n24380 ;
  assign y12330 = n24381 ;
  assign y12331 = ~n24383 ;
  assign y12332 = ~n20172 ;
  assign y12333 = n24384 ;
  assign y12334 = ~1'b0 ;
  assign y12335 = ~1'b0 ;
  assign y12336 = ~1'b0 ;
  assign y12337 = ~n7925 ;
  assign y12338 = ~n24385 ;
  assign y12339 = n24388 ;
  assign y12340 = ~1'b0 ;
  assign y12341 = ~1'b0 ;
  assign y12342 = n24389 ;
  assign y12343 = n24390 ;
  assign y12344 = ~1'b0 ;
  assign y12345 = ~1'b0 ;
  assign y12346 = n24391 ;
  assign y12347 = ~n24392 ;
  assign y12348 = n24395 ;
  assign y12349 = ~n24397 ;
  assign y12350 = ~n24400 ;
  assign y12351 = ~n1265 ;
  assign y12352 = ~n24405 ;
  assign y12353 = n24407 ;
  assign y12354 = n17507 ;
  assign y12355 = n24408 ;
  assign y12356 = ~1'b0 ;
  assign y12357 = ~n24411 ;
  assign y12358 = ~n24422 ;
  assign y12359 = ~n24426 ;
  assign y12360 = ~n24432 ;
  assign y12361 = ~1'b0 ;
  assign y12362 = ~1'b0 ;
  assign y12363 = ~n24434 ;
  assign y12364 = ~n24435 ;
  assign y12365 = n24442 ;
  assign y12366 = ~1'b0 ;
  assign y12367 = ~n24445 ;
  assign y12368 = n24446 ;
  assign y12369 = n24447 ;
  assign y12370 = n24448 ;
  assign y12371 = ~1'b0 ;
  assign y12372 = n24450 ;
  assign y12373 = ~n24454 ;
  assign y12374 = ~1'b0 ;
  assign y12375 = n24459 ;
  assign y12376 = n24463 ;
  assign y12377 = ~1'b0 ;
  assign y12378 = ~1'b0 ;
  assign y12379 = n24466 ;
  assign y12380 = n24470 ;
  assign y12381 = ~1'b0 ;
  assign y12382 = ~1'b0 ;
  assign y12383 = n24471 ;
  assign y12384 = n24479 ;
  assign y12385 = 1'b0 ;
  assign y12386 = ~n24481 ;
  assign y12387 = ~n24485 ;
  assign y12388 = ~n24488 ;
  assign y12389 = n24489 ;
  assign y12390 = n24492 ;
  assign y12391 = n24494 ;
  assign y12392 = ~n24496 ;
  assign y12393 = ~n24497 ;
  assign y12394 = n24499 ;
  assign y12395 = n24500 ;
  assign y12396 = n24507 ;
  assign y12397 = ~1'b0 ;
  assign y12398 = n24508 ;
  assign y12399 = n24510 ;
  assign y12400 = ~1'b0 ;
  assign y12401 = ~1'b0 ;
  assign y12402 = ~1'b0 ;
  assign y12403 = ~1'b0 ;
  assign y12404 = n24511 ;
  assign y12405 = ~1'b0 ;
  assign y12406 = n24518 ;
  assign y12407 = n24520 ;
  assign y12408 = ~n24522 ;
  assign y12409 = ~n24529 ;
  assign y12410 = n24530 ;
  assign y12411 = ~1'b0 ;
  assign y12412 = ~1'b0 ;
  assign y12413 = n24532 ;
  assign y12414 = n24533 ;
  assign y12415 = ~n24535 ;
  assign y12416 = n24539 ;
  assign y12417 = ~1'b0 ;
  assign y12418 = n24541 ;
  assign y12419 = ~n24543 ;
  assign y12420 = ~n24548 ;
  assign y12421 = ~n24551 ;
  assign y12422 = ~1'b0 ;
  assign y12423 = n24553 ;
  assign y12424 = n24554 ;
  assign y12425 = ~1'b0 ;
  assign y12426 = ~1'b0 ;
  assign y12427 = n24555 ;
  assign y12428 = ~n814 ;
  assign y12429 = 1'b0 ;
  assign y12430 = 1'b0 ;
  assign y12431 = ~1'b0 ;
  assign y12432 = n24560 ;
  assign y12433 = ~1'b0 ;
  assign y12434 = n24562 ;
  assign y12435 = ~1'b0 ;
  assign y12436 = n24564 ;
  assign y12437 = n24565 ;
  assign y12438 = ~n24566 ;
  assign y12439 = n24569 ;
  assign y12440 = n24570 ;
  assign y12441 = ~1'b0 ;
  assign y12442 = n24575 ;
  assign y12443 = ~n24579 ;
  assign y12444 = ~1'b0 ;
  assign y12445 = ~1'b0 ;
  assign y12446 = ~1'b0 ;
  assign y12447 = n24582 ;
  assign y12448 = n24586 ;
  assign y12449 = ~n24588 ;
  assign y12450 = ~n24589 ;
  assign y12451 = ~n24591 ;
  assign y12452 = ~1'b0 ;
  assign y12453 = ~1'b0 ;
  assign y12454 = ~1'b0 ;
  assign y12455 = n24594 ;
  assign y12456 = n24597 ;
  assign y12457 = ~n24599 ;
  assign y12458 = ~n24605 ;
  assign y12459 = ~1'b0 ;
  assign y12460 = ~n24607 ;
  assign y12461 = ~1'b0 ;
  assign y12462 = ~1'b0 ;
  assign y12463 = ~n24613 ;
  assign y12464 = n24618 ;
  assign y12465 = n24619 ;
  assign y12466 = n24622 ;
  assign y12467 = n24623 ;
  assign y12468 = ~1'b0 ;
  assign y12469 = n24628 ;
  assign y12470 = ~n24630 ;
  assign y12471 = n24632 ;
  assign y12472 = n13173 ;
  assign y12473 = ~n24637 ;
  assign y12474 = ~n24638 ;
  assign y12475 = n24639 ;
  assign y12476 = n24640 ;
  assign y12477 = ~n24642 ;
  assign y12478 = 1'b0 ;
  assign y12479 = ~1'b0 ;
  assign y12480 = ~1'b0 ;
  assign y12481 = ~n24650 ;
  assign y12482 = ~n24651 ;
  assign y12483 = ~n24652 ;
  assign y12484 = ~n24653 ;
  assign y12485 = n19068 ;
  assign y12486 = n24655 ;
  assign y12487 = n24659 ;
  assign y12488 = ~n24661 ;
  assign y12489 = ~1'b0 ;
  assign y12490 = n24668 ;
  assign y12491 = ~1'b0 ;
  assign y12492 = ~1'b0 ;
  assign y12493 = ~n24672 ;
  assign y12494 = ~1'b0 ;
  assign y12495 = n24673 ;
  assign y12496 = n24674 ;
  assign y12497 = ~1'b0 ;
  assign y12498 = ~n24676 ;
  assign y12499 = ~n24677 ;
  assign y12500 = n24683 ;
  assign y12501 = ~n24684 ;
  assign y12502 = n8449 ;
  assign y12503 = ~n24685 ;
  assign y12504 = n24686 ;
  assign y12505 = n24688 ;
  assign y12506 = 1'b0 ;
  assign y12507 = n24690 ;
  assign y12508 = ~n24695 ;
  assign y12509 = ~n24696 ;
  assign y12510 = ~n24697 ;
  assign y12511 = n24699 ;
  assign y12512 = ~1'b0 ;
  assign y12513 = ~1'b0 ;
  assign y12514 = ~n24700 ;
  assign y12515 = ~n24701 ;
  assign y12516 = n4328 ;
  assign y12517 = ~n24703 ;
  assign y12518 = ~n24704 ;
  assign y12519 = ~n24707 ;
  assign y12520 = ~1'b0 ;
  assign y12521 = n24708 ;
  assign y12522 = ~n24709 ;
  assign y12523 = ~n24710 ;
  assign y12524 = ~1'b0 ;
  assign y12525 = ~n24712 ;
  assign y12526 = ~n24717 ;
  assign y12527 = ~n24718 ;
  assign y12528 = ~1'b0 ;
  assign y12529 = n24720 ;
  assign y12530 = n19344 ;
  assign y12531 = ~n24722 ;
  assign y12532 = ~n24723 ;
  assign y12533 = n24728 ;
  assign y12534 = ~1'b0 ;
  assign y12535 = ~1'b0 ;
  assign y12536 = n24729 ;
  assign y12537 = ~n4910 ;
  assign y12538 = n24730 ;
  assign y12539 = n24732 ;
  assign y12540 = ~n24740 ;
  assign y12541 = ~n24743 ;
  assign y12542 = ~1'b0 ;
  assign y12543 = ~1'b0 ;
  assign y12544 = ~1'b0 ;
  assign y12545 = n24746 ;
  assign y12546 = n24747 ;
  assign y12547 = n24748 ;
  assign y12548 = n24749 ;
  assign y12549 = n24753 ;
  assign y12550 = ~n24758 ;
  assign y12551 = ~1'b0 ;
  assign y12552 = ~n24760 ;
  assign y12553 = ~n24762 ;
  assign y12554 = ~1'b0 ;
  assign y12555 = ~n24769 ;
  assign y12556 = n24772 ;
  assign y12557 = ~n24778 ;
  assign y12558 = n24779 ;
  assign y12559 = n24780 ;
  assign y12560 = ~n24781 ;
  assign y12561 = ~n24782 ;
  assign y12562 = ~n21179 ;
  assign y12563 = n24783 ;
  assign y12564 = 1'b0 ;
  assign y12565 = n24784 ;
  assign y12566 = ~n24796 ;
  assign y12567 = ~1'b0 ;
  assign y12568 = ~n7586 ;
  assign y12569 = n24798 ;
  assign y12570 = ~1'b0 ;
  assign y12571 = ~n24799 ;
  assign y12572 = 1'b0 ;
  assign y12573 = ~n24800 ;
  assign y12574 = n24802 ;
  assign y12575 = ~n24803 ;
  assign y12576 = n24804 ;
  assign y12577 = n24807 ;
  assign y12578 = ~n24810 ;
  assign y12579 = ~1'b0 ;
  assign y12580 = ~n24811 ;
  assign y12581 = n24814 ;
  assign y12582 = n24818 ;
  assign y12583 = ~1'b0 ;
  assign y12584 = ~1'b0 ;
  assign y12585 = ~n24819 ;
  assign y12586 = ~1'b0 ;
  assign y12587 = ~n24821 ;
  assign y12588 = ~1'b0 ;
  assign y12589 = ~1'b0 ;
  assign y12590 = ~n24826 ;
  assign y12591 = ~n6177 ;
  assign y12592 = n24829 ;
  assign y12593 = ~1'b0 ;
  assign y12594 = ~n24833 ;
  assign y12595 = n24834 ;
  assign y12596 = ~1'b0 ;
  assign y12597 = ~n24837 ;
  assign y12598 = n24845 ;
  assign y12599 = n24846 ;
  assign y12600 = ~n24849 ;
  assign y12601 = n24852 ;
  assign y12602 = 1'b0 ;
  assign y12603 = n24853 ;
  assign y12604 = n5210 ;
  assign y12605 = ~1'b0 ;
  assign y12606 = ~1'b0 ;
  assign y12607 = ~1'b0 ;
  assign y12608 = n24854 ;
  assign y12609 = ~n24855 ;
  assign y12610 = n24856 ;
  assign y12611 = n24859 ;
  assign y12612 = n11234 ;
  assign y12613 = ~1'b0 ;
  assign y12614 = ~1'b0 ;
  assign y12615 = ~n24860 ;
  assign y12616 = ~1'b0 ;
  assign y12617 = n24864 ;
  assign y12618 = ~n24869 ;
  assign y12619 = ~n24873 ;
  assign y12620 = ~1'b0 ;
  assign y12621 = ~1'b0 ;
  assign y12622 = n24874 ;
  assign y12623 = n2014 ;
  assign y12624 = ~1'b0 ;
  assign y12625 = n24883 ;
  assign y12626 = n24889 ;
  assign y12627 = n24893 ;
  assign y12628 = ~n14080 ;
  assign y12629 = ~n24895 ;
  assign y12630 = ~1'b0 ;
  assign y12631 = ~1'b0 ;
  assign y12632 = ~1'b0 ;
  assign y12633 = ~1'b0 ;
  assign y12634 = ~1'b0 ;
  assign y12635 = ~n24897 ;
  assign y12636 = ~1'b0 ;
  assign y12637 = ~1'b0 ;
  assign y12638 = ~n24898 ;
  assign y12639 = ~1'b0 ;
  assign y12640 = ~n24900 ;
  assign y12641 = ~1'b0 ;
  assign y12642 = ~n24905 ;
  assign y12643 = n24906 ;
  assign y12644 = ~n24910 ;
  assign y12645 = ~n24912 ;
  assign y12646 = ~n7809 ;
  assign y12647 = ~1'b0 ;
  assign y12648 = n24913 ;
  assign y12649 = n1261 ;
  assign y12650 = ~n12754 ;
  assign y12651 = ~n24914 ;
  assign y12652 = n24919 ;
  assign y12653 = n24922 ;
  assign y12654 = n24925 ;
  assign y12655 = ~n24926 ;
  assign y12656 = n24927 ;
  assign y12657 = n24928 ;
  assign y12658 = n24933 ;
  assign y12659 = n24938 ;
  assign y12660 = n24939 ;
  assign y12661 = n24942 ;
  assign y12662 = n24944 ;
  assign y12663 = ~n24945 ;
  assign y12664 = ~1'b0 ;
  assign y12665 = ~1'b0 ;
  assign y12666 = n24948 ;
  assign y12667 = ~n24952 ;
  assign y12668 = ~1'b0 ;
  assign y12669 = ~1'b0 ;
  assign y12670 = ~n24955 ;
  assign y12671 = n24958 ;
  assign y12672 = ~n24962 ;
  assign y12673 = ~n14017 ;
  assign y12674 = ~n8816 ;
  assign y12675 = ~n24972 ;
  assign y12676 = ~n24974 ;
  assign y12677 = ~1'b0 ;
  assign y12678 = ~1'b0 ;
  assign y12679 = n24978 ;
  assign y12680 = ~n23305 ;
  assign y12681 = n24980 ;
  assign y12682 = n24983 ;
  assign y12683 = n24989 ;
  assign y12684 = ~1'b0 ;
  assign y12685 = ~1'b0 ;
  assign y12686 = ~1'b0 ;
  assign y12687 = n24991 ;
  assign y12688 = n24993 ;
  assign y12689 = n24995 ;
  assign y12690 = ~1'b0 ;
  assign y12691 = ~n25001 ;
  assign y12692 = n25004 ;
  assign y12693 = 1'b0 ;
  assign y12694 = ~n25006 ;
  assign y12695 = ~n25008 ;
  assign y12696 = ~n25019 ;
  assign y12697 = ~1'b0 ;
  assign y12698 = ~n25021 ;
  assign y12699 = ~n25022 ;
  assign y12700 = ~n25026 ;
  assign y12701 = ~1'b0 ;
  assign y12702 = ~1'b0 ;
  assign y12703 = ~n25027 ;
  assign y12704 = ~1'b0 ;
  assign y12705 = ~n25031 ;
  assign y12706 = n25033 ;
  assign y12707 = ~n18465 ;
  assign y12708 = ~n25038 ;
  assign y12709 = ~n25041 ;
  assign y12710 = ~1'b0 ;
  assign y12711 = n25043 ;
  assign y12712 = ~1'b0 ;
  assign y12713 = ~n25044 ;
  assign y12714 = ~n25046 ;
  assign y12715 = n25049 ;
  assign y12716 = ~1'b0 ;
  assign y12717 = n6533 ;
  assign y12718 = ~1'b0 ;
  assign y12719 = ~n25059 ;
  assign y12720 = n25061 ;
  assign y12721 = ~n25062 ;
  assign y12722 = ~1'b0 ;
  assign y12723 = ~n25063 ;
  assign y12724 = ~n25064 ;
  assign y12725 = ~1'b0 ;
  assign y12726 = n25066 ;
  assign y12727 = ~n25068 ;
  assign y12728 = ~n25080 ;
  assign y12729 = ~1'b0 ;
  assign y12730 = ~n4269 ;
  assign y12731 = n5792 ;
  assign y12732 = ~n25082 ;
  assign y12733 = ~1'b0 ;
  assign y12734 = n25084 ;
  assign y12735 = ~n11277 ;
  assign y12736 = ~1'b0 ;
  assign y12737 = n25086 ;
  assign y12738 = ~n25091 ;
  assign y12739 = n25092 ;
  assign y12740 = ~n25093 ;
  assign y12741 = ~n25096 ;
  assign y12742 = ~n25098 ;
  assign y12743 = ~n25100 ;
  assign y12744 = n25105 ;
  assign y12745 = ~1'b0 ;
  assign y12746 = ~n25112 ;
  assign y12747 = ~n25113 ;
  assign y12748 = ~1'b0 ;
  assign y12749 = ~n25116 ;
  assign y12750 = ~n25119 ;
  assign y12751 = 1'b0 ;
  assign y12752 = n25121 ;
  assign y12753 = ~n10349 ;
  assign y12754 = n25126 ;
  assign y12755 = n25128 ;
  assign y12756 = ~1'b0 ;
  assign y12757 = ~n25136 ;
  assign y12758 = n25142 ;
  assign y12759 = ~1'b0 ;
  assign y12760 = ~n25143 ;
  assign y12761 = ~1'b0 ;
  assign y12762 = ~n25144 ;
  assign y12763 = n25147 ;
  assign y12764 = ~n25149 ;
  assign y12765 = ~n10000 ;
  assign y12766 = ~n25152 ;
  assign y12767 = ~n25156 ;
  assign y12768 = ~n7271 ;
  assign y12769 = n25157 ;
  assign y12770 = n25159 ;
  assign y12771 = n25160 ;
  assign y12772 = n25162 ;
  assign y12773 = ~n25163 ;
  assign y12774 = ~1'b0 ;
  assign y12775 = n25164 ;
  assign y12776 = n3942 ;
  assign y12777 = n25166 ;
  assign y12778 = ~1'b0 ;
  assign y12779 = ~n25170 ;
  assign y12780 = ~n25172 ;
  assign y12781 = n25173 ;
  assign y12782 = ~n25179 ;
  assign y12783 = n25181 ;
  assign y12784 = n25182 ;
  assign y12785 = n25185 ;
  assign y12786 = n25193 ;
  assign y12787 = n23475 ;
  assign y12788 = n25196 ;
  assign y12789 = ~n25198 ;
  assign y12790 = ~n11440 ;
  assign y12791 = ~1'b0 ;
  assign y12792 = ~n25202 ;
  assign y12793 = ~1'b0 ;
  assign y12794 = ~1'b0 ;
  assign y12795 = n25204 ;
  assign y12796 = n25206 ;
  assign y12797 = ~1'b0 ;
  assign y12798 = n25207 ;
  assign y12799 = n25209 ;
  assign y12800 = ~n25210 ;
  assign y12801 = ~n25212 ;
  assign y12802 = ~n25214 ;
  assign y12803 = ~n25215 ;
  assign y12804 = ~1'b0 ;
  assign y12805 = n25217 ;
  assign y12806 = ~1'b0 ;
  assign y12807 = n25220 ;
  assign y12808 = ~n13162 ;
  assign y12809 = ~1'b0 ;
  assign y12810 = ~1'b0 ;
  assign y12811 = ~n25223 ;
  assign y12812 = ~n25225 ;
  assign y12813 = n3411 ;
  assign y12814 = ~n25228 ;
  assign y12815 = n25230 ;
  assign y12816 = ~n25237 ;
  assign y12817 = ~n7623 ;
  assign y12818 = ~1'b0 ;
  assign y12819 = 1'b0 ;
  assign y12820 = ~1'b0 ;
  assign y12821 = n25238 ;
  assign y12822 = ~1'b0 ;
  assign y12823 = n25243 ;
  assign y12824 = n25246 ;
  assign y12825 = n25247 ;
  assign y12826 = ~1'b0 ;
  assign y12827 = ~1'b0 ;
  assign y12828 = n25249 ;
  assign y12829 = ~n25252 ;
  assign y12830 = ~n3378 ;
  assign y12831 = n25254 ;
  assign y12832 = ~1'b0 ;
  assign y12833 = ~n25258 ;
  assign y12834 = n25261 ;
  assign y12835 = ~n25263 ;
  assign y12836 = ~n25264 ;
  assign y12837 = ~1'b0 ;
  assign y12838 = ~1'b0 ;
  assign y12839 = ~n9622 ;
  assign y12840 = n25266 ;
  assign y12841 = 1'b0 ;
  assign y12842 = n25270 ;
  assign y12843 = ~n25271 ;
  assign y12844 = n25279 ;
  assign y12845 = n25282 ;
  assign y12846 = ~n25283 ;
  assign y12847 = ~n25285 ;
  assign y12848 = ~n25286 ;
  assign y12849 = ~n25288 ;
  assign y12850 = n25289 ;
  assign y12851 = n18222 ;
  assign y12852 = ~n25299 ;
  assign y12853 = ~n2320 ;
  assign y12854 = n25301 ;
  assign y12855 = n25304 ;
  assign y12856 = ~n5442 ;
  assign y12857 = ~1'b0 ;
  assign y12858 = n25305 ;
  assign y12859 = n25307 ;
  assign y12860 = ~1'b0 ;
  assign y12861 = n25308 ;
  assign y12862 = n25315 ;
  assign y12863 = n25321 ;
  assign y12864 = n25325 ;
  assign y12865 = ~n25326 ;
  assign y12866 = ~1'b0 ;
  assign y12867 = ~n25329 ;
  assign y12868 = n25333 ;
  assign y12869 = ~n25334 ;
  assign y12870 = ~1'b0 ;
  assign y12871 = 1'b0 ;
  assign y12872 = ~n25335 ;
  assign y12873 = ~n12812 ;
  assign y12874 = ~1'b0 ;
  assign y12875 = ~1'b0 ;
  assign y12876 = ~n13628 ;
  assign y12877 = ~1'b0 ;
  assign y12878 = ~n25337 ;
  assign y12879 = ~n25347 ;
  assign y12880 = n23842 ;
  assign y12881 = n25349 ;
  assign y12882 = ~1'b0 ;
  assign y12883 = ~1'b0 ;
  assign y12884 = ~n25353 ;
  assign y12885 = ~n25355 ;
  assign y12886 = ~1'b0 ;
  assign y12887 = ~1'b0 ;
  assign y12888 = ~n25359 ;
  assign y12889 = ~n25363 ;
  assign y12890 = n25368 ;
  assign y12891 = n25373 ;
  assign y12892 = ~1'b0 ;
  assign y12893 = ~n25376 ;
  assign y12894 = ~n14845 ;
  assign y12895 = n25378 ;
  assign y12896 = ~n6521 ;
  assign y12897 = ~n25379 ;
  assign y12898 = n25381 ;
  assign y12899 = ~n25382 ;
  assign y12900 = n25383 ;
  assign y12901 = ~1'b0 ;
  assign y12902 = n25387 ;
  assign y12903 = ~1'b0 ;
  assign y12904 = 1'b0 ;
  assign y12905 = n25388 ;
  assign y12906 = ~n25391 ;
  assign y12907 = n25395 ;
  assign y12908 = n7222 ;
  assign y12909 = ~n25398 ;
  assign y12910 = n25404 ;
  assign y12911 = ~n25406 ;
  assign y12912 = ~1'b0 ;
  assign y12913 = n25408 ;
  assign y12914 = ~1'b0 ;
  assign y12915 = ~1'b0 ;
  assign y12916 = ~n25409 ;
  assign y12917 = ~n25412 ;
  assign y12918 = n25414 ;
  assign y12919 = ~1'b0 ;
  assign y12920 = n25415 ;
  assign y12921 = ~1'b0 ;
  assign y12922 = ~1'b0 ;
  assign y12923 = ~1'b0 ;
  assign y12924 = ~n25417 ;
  assign y12925 = ~1'b0 ;
  assign y12926 = ~n25419 ;
  assign y12927 = n25424 ;
  assign y12928 = ~n25428 ;
  assign y12929 = n25438 ;
  assign y12930 = n15059 ;
  assign y12931 = ~n25443 ;
  assign y12932 = n25446 ;
  assign y12933 = n25449 ;
  assign y12934 = 1'b0 ;
  assign y12935 = ~n25451 ;
  assign y12936 = ~1'b0 ;
  assign y12937 = ~n25457 ;
  assign y12938 = ~n25460 ;
  assign y12939 = ~n25461 ;
  assign y12940 = ~1'b0 ;
  assign y12941 = n25463 ;
  assign y12942 = ~1'b0 ;
  assign y12943 = n25464 ;
  assign y12944 = n25466 ;
  assign y12945 = n25471 ;
  assign y12946 = n25477 ;
  assign y12947 = ~1'b0 ;
  assign y12948 = ~1'b0 ;
  assign y12949 = ~n25479 ;
  assign y12950 = n25480 ;
  assign y12951 = ~1'b0 ;
  assign y12952 = ~n25484 ;
  assign y12953 = ~n13671 ;
  assign y12954 = n25485 ;
  assign y12955 = n25488 ;
  assign y12956 = n25489 ;
  assign y12957 = ~n25496 ;
  assign y12958 = ~1'b0 ;
  assign y12959 = n25498 ;
  assign y12960 = n25501 ;
  assign y12961 = ~1'b0 ;
  assign y12962 = ~n25503 ;
  assign y12963 = ~1'b0 ;
  assign y12964 = n25505 ;
  assign y12965 = ~1'b0 ;
  assign y12966 = ~n25506 ;
  assign y12967 = ~n25508 ;
  assign y12968 = ~n25514 ;
  assign y12969 = n25518 ;
  assign y12970 = n25522 ;
  assign y12971 = x177 ;
  assign y12972 = ~n12690 ;
  assign y12973 = ~n25529 ;
  assign y12974 = n25532 ;
  assign y12975 = ~n25541 ;
  assign y12976 = ~1'b0 ;
  assign y12977 = ~1'b0 ;
  assign y12978 = n25543 ;
  assign y12979 = ~n25547 ;
  assign y12980 = ~1'b0 ;
  assign y12981 = ~n25549 ;
  assign y12982 = ~n25553 ;
  assign y12983 = ~n25556 ;
  assign y12984 = n25558 ;
  assign y12985 = ~1'b0 ;
  assign y12986 = n25559 ;
  assign y12987 = ~n25572 ;
  assign y12988 = ~1'b0 ;
  assign y12989 = ~n25574 ;
  assign y12990 = ~n25581 ;
  assign y12991 = n25584 ;
  assign y12992 = n25587 ;
  assign y12993 = ~1'b0 ;
  assign y12994 = ~1'b0 ;
  assign y12995 = ~1'b0 ;
  assign y12996 = n25589 ;
  assign y12997 = ~1'b0 ;
  assign y12998 = ~n25590 ;
  assign y12999 = n25595 ;
  assign y13000 = n21356 ;
  assign y13001 = n25601 ;
  assign y13002 = n25602 ;
  assign y13003 = ~1'b0 ;
  assign y13004 = n25606 ;
  assign y13005 = ~1'b0 ;
  assign y13006 = n13370 ;
  assign y13007 = ~n25609 ;
  assign y13008 = n25611 ;
  assign y13009 = ~1'b0 ;
  assign y13010 = ~n25614 ;
  assign y13011 = ~n25621 ;
  assign y13012 = ~n25624 ;
  assign y13013 = ~1'b0 ;
  assign y13014 = ~1'b0 ;
  assign y13015 = n25625 ;
  assign y13016 = ~n25627 ;
  assign y13017 = n13521 ;
  assign y13018 = ~n25628 ;
  assign y13019 = n25629 ;
  assign y13020 = ~n25640 ;
  assign y13021 = ~1'b0 ;
  assign y13022 = n25641 ;
  assign y13023 = ~1'b0 ;
  assign y13024 = ~n2877 ;
  assign y13025 = n25642 ;
  assign y13026 = n25646 ;
  assign y13027 = ~n25655 ;
  assign y13028 = ~n25662 ;
  assign y13029 = n25663 ;
  assign y13030 = ~n25665 ;
  assign y13031 = n25667 ;
  assign y13032 = 1'b0 ;
  assign y13033 = ~n25669 ;
  assign y13034 = ~n25674 ;
  assign y13035 = ~n25679 ;
  assign y13036 = n25680 ;
  assign y13037 = ~1'b0 ;
  assign y13038 = ~1'b0 ;
  assign y13039 = ~1'b0 ;
  assign y13040 = ~1'b0 ;
  assign y13041 = n25686 ;
  assign y13042 = n25687 ;
  assign y13043 = ~1'b0 ;
  assign y13044 = ~1'b0 ;
  assign y13045 = ~n25690 ;
  assign y13046 = ~n25694 ;
  assign y13047 = ~n25697 ;
  assign y13048 = ~n25698 ;
  assign y13049 = ~1'b0 ;
  assign y13050 = n25701 ;
  assign y13051 = n25704 ;
  assign y13052 = ~n25706 ;
  assign y13053 = ~n25712 ;
  assign y13054 = ~n25717 ;
  assign y13055 = ~1'b0 ;
  assign y13056 = ~n25722 ;
  assign y13057 = n25726 ;
  assign y13058 = n25727 ;
  assign y13059 = ~1'b0 ;
  assign y13060 = n25730 ;
  assign y13061 = ~n1039 ;
  assign y13062 = ~1'b0 ;
  assign y13063 = ~n25735 ;
  assign y13064 = ~n25737 ;
  assign y13065 = ~1'b0 ;
  assign y13066 = n25741 ;
  assign y13067 = n25742 ;
  assign y13068 = ~1'b0 ;
  assign y13069 = n25743 ;
  assign y13070 = n7291 ;
  assign y13071 = ~n25745 ;
  assign y13072 = ~n25757 ;
  assign y13073 = ~n25758 ;
  assign y13074 = ~n25759 ;
  assign y13075 = n25762 ;
  assign y13076 = ~n25763 ;
  assign y13077 = n25764 ;
  assign y13078 = ~1'b0 ;
  assign y13079 = ~n9801 ;
  assign y13080 = 1'b0 ;
  assign y13081 = ~n25766 ;
  assign y13082 = ~1'b0 ;
  assign y13083 = ~n25767 ;
  assign y13084 = n24559 ;
  assign y13085 = n25773 ;
  assign y13086 = ~1'b0 ;
  assign y13087 = ~n25775 ;
  assign y13088 = ~1'b0 ;
  assign y13089 = n25778 ;
  assign y13090 = n25780 ;
  assign y13091 = ~1'b0 ;
  assign y13092 = 1'b0 ;
  assign y13093 = n25781 ;
  assign y13094 = ~1'b0 ;
  assign y13095 = ~n25782 ;
  assign y13096 = n25783 ;
  assign y13097 = n25784 ;
  assign y13098 = n25785 ;
  assign y13099 = ~n25788 ;
  assign y13100 = ~n25790 ;
  assign y13101 = ~1'b0 ;
  assign y13102 = n25793 ;
  assign y13103 = ~n25797 ;
  assign y13104 = n25798 ;
  assign y13105 = ~n25800 ;
  assign y13106 = n25804 ;
  assign y13107 = ~n1309 ;
  assign y13108 = ~1'b0 ;
  assign y13109 = ~n25805 ;
  assign y13110 = ~n24688 ;
  assign y13111 = ~n25807 ;
  assign y13112 = ~n25814 ;
  assign y13113 = ~1'b0 ;
  assign y13114 = n25815 ;
  assign y13115 = n6849 ;
  assign y13116 = n25816 ;
  assign y13117 = ~1'b0 ;
  assign y13118 = ~1'b0 ;
  assign y13119 = ~1'b0 ;
  assign y13120 = ~n25818 ;
  assign y13121 = n25821 ;
  assign y13122 = n25823 ;
  assign y13123 = n25824 ;
  assign y13124 = n867 ;
  assign y13125 = ~n25825 ;
  assign y13126 = ~n18042 ;
  assign y13127 = n25830 ;
  assign y13128 = ~1'b0 ;
  assign y13129 = ~n25833 ;
  assign y13130 = ~n25851 ;
  assign y13131 = ~n25852 ;
  assign y13132 = ~1'b0 ;
  assign y13133 = ~n25858 ;
  assign y13134 = ~n25861 ;
  assign y13135 = 1'b0 ;
  assign y13136 = ~n25865 ;
  assign y13137 = ~n9064 ;
  assign y13138 = n25868 ;
  assign y13139 = n25870 ;
  assign y13140 = n25872 ;
  assign y13141 = n25874 ;
  assign y13142 = ~n8216 ;
  assign y13143 = ~n25881 ;
  assign y13144 = ~n25883 ;
  assign y13145 = ~1'b0 ;
  assign y13146 = ~n5750 ;
  assign y13147 = ~n25884 ;
  assign y13148 = n25887 ;
  assign y13149 = 1'b0 ;
  assign y13150 = n25888 ;
  assign y13151 = ~1'b0 ;
  assign y13152 = n25890 ;
  assign y13153 = n25891 ;
  assign y13154 = n25892 ;
  assign y13155 = ~n14663 ;
  assign y13156 = n25898 ;
  assign y13157 = ~n25903 ;
  assign y13158 = ~1'b0 ;
  assign y13159 = ~n25904 ;
  assign y13160 = 1'b0 ;
  assign y13161 = ~n25907 ;
  assign y13162 = n25912 ;
  assign y13163 = ~n25915 ;
  assign y13164 = ~1'b0 ;
  assign y13165 = n6155 ;
  assign y13166 = n25917 ;
  assign y13167 = ~1'b0 ;
  assign y13168 = ~n25919 ;
  assign y13169 = n25923 ;
  assign y13170 = ~n21868 ;
  assign y13171 = ~n25924 ;
  assign y13172 = ~n25926 ;
  assign y13173 = n7532 ;
  assign y13174 = ~n11450 ;
  assign y13175 = ~1'b0 ;
  assign y13176 = n25929 ;
  assign y13177 = ~n25930 ;
  assign y13178 = ~n16615 ;
  assign y13179 = n25931 ;
  assign y13180 = ~1'b0 ;
  assign y13181 = n25933 ;
  assign y13182 = ~1'b0 ;
  assign y13183 = ~n25936 ;
  assign y13184 = ~n25941 ;
  assign y13185 = ~1'b0 ;
  assign y13186 = n25944 ;
  assign y13187 = n25946 ;
  assign y13188 = n25947 ;
  assign y13189 = ~n25948 ;
  assign y13190 = ~1'b0 ;
  assign y13191 = ~1'b0 ;
  assign y13192 = ~1'b0 ;
  assign y13193 = ~n25949 ;
  assign y13194 = n25950 ;
  assign y13195 = ~1'b0 ;
  assign y13196 = n25951 ;
  assign y13197 = n25952 ;
  assign y13198 = n25953 ;
  assign y13199 = ~1'b0 ;
  assign y13200 = ~n25955 ;
  assign y13201 = n25959 ;
  assign y13202 = ~n25961 ;
  assign y13203 = ~n25966 ;
  assign y13204 = ~n25967 ;
  assign y13205 = n25970 ;
  assign y13206 = ~n25980 ;
  assign y13207 = n25982 ;
  assign y13208 = n25983 ;
  assign y13209 = ~1'b0 ;
  assign y13210 = ~n25988 ;
  assign y13211 = ~1'b0 ;
  assign y13212 = ~n25991 ;
  assign y13213 = ~1'b0 ;
  assign y13214 = ~n25993 ;
  assign y13215 = ~n25996 ;
  assign y13216 = n26000 ;
  assign y13217 = ~n26003 ;
  assign y13218 = ~1'b0 ;
  assign y13219 = n26008 ;
  assign y13220 = ~1'b0 ;
  assign y13221 = ~n26010 ;
  assign y13222 = ~n26014 ;
  assign y13223 = ~n26016 ;
  assign y13224 = n394 ;
  assign y13225 = n26018 ;
  assign y13226 = n2961 ;
  assign y13227 = ~1'b0 ;
  assign y13228 = ~1'b0 ;
  assign y13229 = ~n26026 ;
  assign y13230 = n26028 ;
  assign y13231 = n26029 ;
  assign y13232 = ~1'b0 ;
  assign y13233 = n26030 ;
  assign y13234 = ~n11038 ;
  assign y13235 = ~n26032 ;
  assign y13236 = 1'b0 ;
  assign y13237 = ~1'b0 ;
  assign y13238 = ~1'b0 ;
  assign y13239 = ~1'b0 ;
  assign y13240 = n8861 ;
  assign y13241 = n26033 ;
  assign y13242 = ~n26034 ;
  assign y13243 = ~1'b0 ;
  assign y13244 = ~1'b0 ;
  assign y13245 = n26035 ;
  assign y13246 = ~n26039 ;
  assign y13247 = n26040 ;
  assign y13248 = ~n26044 ;
  assign y13249 = n26047 ;
  assign y13250 = ~n26048 ;
  assign y13251 = ~1'b0 ;
  assign y13252 = n26050 ;
  assign y13253 = n26065 ;
  assign y13254 = ~n26066 ;
  assign y13255 = n26067 ;
  assign y13256 = n26070 ;
  assign y13257 = ~n10832 ;
  assign y13258 = n26072 ;
  assign y13259 = n26073 ;
  assign y13260 = ~n26076 ;
  assign y13261 = ~n26077 ;
  assign y13262 = n26082 ;
  assign y13263 = n26083 ;
  assign y13264 = ~1'b0 ;
  assign y13265 = ~n26087 ;
  assign y13266 = ~n26090 ;
  assign y13267 = n26091 ;
  assign y13268 = n26096 ;
  assign y13269 = n26097 ;
  assign y13270 = ~1'b0 ;
  assign y13271 = ~1'b0 ;
  assign y13272 = ~1'b0 ;
  assign y13273 = 1'b0 ;
  assign y13274 = ~n26102 ;
  assign y13275 = n26108 ;
  assign y13276 = ~n26110 ;
  assign y13277 = ~n26114 ;
  assign y13278 = n26116 ;
  assign y13279 = n21358 ;
  assign y13280 = ~n26117 ;
  assign y13281 = ~n26124 ;
  assign y13282 = ~n26128 ;
  assign y13283 = n26130 ;
  assign y13284 = ~n26135 ;
  assign y13285 = ~1'b0 ;
  assign y13286 = n26136 ;
  assign y13287 = n26137 ;
  assign y13288 = ~1'b0 ;
  assign y13289 = n26139 ;
  assign y13290 = ~n26141 ;
  assign y13291 = ~n26142 ;
  assign y13292 = ~1'b0 ;
  assign y13293 = ~n26144 ;
  assign y13294 = n26147 ;
  assign y13295 = ~n26151 ;
  assign y13296 = ~1'b0 ;
  assign y13297 = ~n26154 ;
  assign y13298 = ~1'b0 ;
  assign y13299 = ~n26159 ;
  assign y13300 = ~1'b0 ;
  assign y13301 = ~1'b0 ;
  assign y13302 = n26160 ;
  assign y13303 = ~1'b0 ;
  assign y13304 = n26162 ;
  assign y13305 = ~n26164 ;
  assign y13306 = ~n26165 ;
  assign y13307 = ~1'b0 ;
  assign y13308 = ~n26169 ;
  assign y13309 = n26173 ;
  assign y13310 = n26175 ;
  assign y13311 = n26178 ;
  assign y13312 = n26179 ;
  assign y13313 = ~n26180 ;
  assign y13314 = n26184 ;
  assign y13315 = ~n22931 ;
  assign y13316 = n26187 ;
  assign y13317 = ~n26188 ;
  assign y13318 = ~1'b0 ;
  assign y13319 = ~n26191 ;
  assign y13320 = ~n16740 ;
  assign y13321 = ~n26193 ;
  assign y13322 = n26197 ;
  assign y13323 = ~n26199 ;
  assign y13324 = ~1'b0 ;
  assign y13325 = ~n26202 ;
  assign y13326 = n26205 ;
  assign y13327 = n26206 ;
  assign y13328 = ~1'b0 ;
  assign y13329 = ~1'b0 ;
  assign y13330 = ~1'b0 ;
  assign y13331 = n26208 ;
  assign y13332 = ~1'b0 ;
  assign y13333 = n24755 ;
  assign y13334 = n26212 ;
  assign y13335 = n26214 ;
  assign y13336 = n26216 ;
  assign y13337 = ~1'b0 ;
  assign y13338 = n26219 ;
  assign y13339 = ~1'b0 ;
  assign y13340 = n26225 ;
  assign y13341 = n26228 ;
  assign y13342 = ~1'b0 ;
  assign y13343 = ~n24695 ;
  assign y13344 = n26232 ;
  assign y13345 = ~1'b0 ;
  assign y13346 = n26233 ;
  assign y13347 = ~n26236 ;
  assign y13348 = 1'b0 ;
  assign y13349 = n26240 ;
  assign y13350 = n26242 ;
  assign y13351 = n26243 ;
  assign y13352 = ~n26245 ;
  assign y13353 = n26251 ;
  assign y13354 = ~n21520 ;
  assign y13355 = n26252 ;
  assign y13356 = ~1'b0 ;
  assign y13357 = ~1'b0 ;
  assign y13358 = n26254 ;
  assign y13359 = ~1'b0 ;
  assign y13360 = ~1'b0 ;
  assign y13361 = n26256 ;
  assign y13362 = 1'b0 ;
  assign y13363 = ~1'b0 ;
  assign y13364 = n26258 ;
  assign y13365 = 1'b0 ;
  assign y13366 = ~n26263 ;
  assign y13367 = ~n26264 ;
  assign y13368 = n26267 ;
  assign y13369 = ~1'b0 ;
  assign y13370 = ~n26272 ;
  assign y13371 = ~n26274 ;
  assign y13372 = n26279 ;
  assign y13373 = ~n26282 ;
  assign y13374 = n26284 ;
  assign y13375 = ~1'b0 ;
  assign y13376 = ~n15119 ;
  assign y13377 = ~n26288 ;
  assign y13378 = n26289 ;
  assign y13379 = n26291 ;
  assign y13380 = n26293 ;
  assign y13381 = ~n26294 ;
  assign y13382 = ~n26301 ;
  assign y13383 = n26302 ;
  assign y13384 = ~n26305 ;
  assign y13385 = ~n26306 ;
  assign y13386 = ~n26310 ;
  assign y13387 = n26315 ;
  assign y13388 = n26316 ;
  assign y13389 = ~1'b0 ;
  assign y13390 = ~n26318 ;
  assign y13391 = ~n6268 ;
  assign y13392 = n26321 ;
  assign y13393 = ~1'b0 ;
  assign y13394 = ~1'b0 ;
  assign y13395 = ~1'b0 ;
  assign y13396 = ~n26325 ;
  assign y13397 = ~n26328 ;
  assign y13398 = ~1'b0 ;
  assign y13399 = ~n26329 ;
  assign y13400 = ~n26330 ;
  assign y13401 = ~n26331 ;
  assign y13402 = ~n26332 ;
  assign y13403 = n26337 ;
  assign y13404 = 1'b0 ;
  assign y13405 = n26338 ;
  assign y13406 = ~n26346 ;
  assign y13407 = ~n26348 ;
  assign y13408 = ~n26350 ;
  assign y13409 = n26352 ;
  assign y13410 = ~1'b0 ;
  assign y13411 = ~n26356 ;
  assign y13412 = ~1'b0 ;
  assign y13413 = 1'b0 ;
  assign y13414 = n26365 ;
  assign y13415 = ~1'b0 ;
  assign y13416 = ~n14526 ;
  assign y13417 = ~n26368 ;
  assign y13418 = ~1'b0 ;
  assign y13419 = ~1'b0 ;
  assign y13420 = ~n26369 ;
  assign y13421 = ~n26370 ;
  assign y13422 = ~1'b0 ;
  assign y13423 = ~n26374 ;
  assign y13424 = ~1'b0 ;
  assign y13425 = ~n26375 ;
  assign y13426 = n26378 ;
  assign y13427 = n26380 ;
  assign y13428 = n26381 ;
  assign y13429 = ~1'b0 ;
  assign y13430 = n26385 ;
  assign y13431 = ~1'b0 ;
  assign y13432 = ~n26386 ;
  assign y13433 = ~n26390 ;
  assign y13434 = ~n26392 ;
  assign y13435 = n26393 ;
  assign y13436 = ~n26395 ;
  assign y13437 = n26402 ;
  assign y13438 = ~1'b0 ;
  assign y13439 = ~1'b0 ;
  assign y13440 = ~n26404 ;
  assign y13441 = ~n26406 ;
  assign y13442 = ~n26408 ;
  assign y13443 = ~1'b0 ;
  assign y13444 = n26411 ;
  assign y13445 = ~1'b0 ;
  assign y13446 = ~1'b0 ;
  assign y13447 = n26412 ;
  assign y13448 = ~n26415 ;
  assign y13449 = n26421 ;
  assign y13450 = n26425 ;
  assign y13451 = n26427 ;
  assign y13452 = n26429 ;
  assign y13453 = ~1'b0 ;
  assign y13454 = n17488 ;
  assign y13455 = ~1'b0 ;
  assign y13456 = n26431 ;
  assign y13457 = n26433 ;
  assign y13458 = ~n26434 ;
  assign y13459 = n26444 ;
  assign y13460 = ~n26445 ;
  assign y13461 = ~n26454 ;
  assign y13462 = ~n26458 ;
  assign y13463 = ~1'b0 ;
  assign y13464 = n26464 ;
  assign y13465 = n26465 ;
  assign y13466 = n26466 ;
  assign y13467 = ~n26469 ;
  assign y13468 = ~1'b0 ;
  assign y13469 = ~1'b0 ;
  assign y13470 = ~1'b0 ;
  assign y13471 = ~1'b0 ;
  assign y13472 = ~1'b0 ;
  assign y13473 = n26472 ;
  assign y13474 = ~n26473 ;
  assign y13475 = ~n1342 ;
  assign y13476 = ~1'b0 ;
  assign y13477 = n26476 ;
  assign y13478 = ~1'b0 ;
  assign y13479 = ~n26478 ;
  assign y13480 = ~n26487 ;
  assign y13481 = n26490 ;
  assign y13482 = ~1'b0 ;
  assign y13483 = ~n26491 ;
  assign y13484 = ~n26492 ;
  assign y13485 = ~n589 ;
  assign y13486 = ~n26494 ;
  assign y13487 = n26497 ;
  assign y13488 = n26499 ;
  assign y13489 = ~1'b0 ;
  assign y13490 = ~1'b0 ;
  assign y13491 = n26506 ;
  assign y13492 = ~1'b0 ;
  assign y13493 = ~n26507 ;
  assign y13494 = ~n26508 ;
  assign y13495 = n26509 ;
  assign y13496 = ~1'b0 ;
  assign y13497 = ~n26513 ;
  assign y13498 = n26517 ;
  assign y13499 = ~1'b0 ;
  assign y13500 = ~1'b0 ;
  assign y13501 = ~n26518 ;
  assign y13502 = ~n26523 ;
  assign y13503 = n26526 ;
  assign y13504 = ~n26527 ;
  assign y13505 = n26528 ;
  assign y13506 = ~n26529 ;
  assign y13507 = 1'b0 ;
  assign y13508 = ~1'b0 ;
  assign y13509 = n26531 ;
  assign y13510 = ~n19174 ;
  assign y13511 = n26537 ;
  assign y13512 = n21757 ;
  assign y13513 = ~1'b0 ;
  assign y13514 = ~1'b0 ;
  assign y13515 = ~n26545 ;
  assign y13516 = ~n26550 ;
  assign y13517 = ~n26551 ;
  assign y13518 = n26553 ;
  assign y13519 = n9114 ;
  assign y13520 = ~n26555 ;
  assign y13521 = ~n26556 ;
  assign y13522 = ~1'b0 ;
  assign y13523 = ~n26559 ;
  assign y13524 = n26564 ;
  assign y13525 = n26565 ;
  assign y13526 = ~1'b0 ;
  assign y13527 = n26567 ;
  assign y13528 = ~n26568 ;
  assign y13529 = n26569 ;
  assign y13530 = ~n26571 ;
  assign y13531 = ~n26575 ;
  assign y13532 = ~1'b0 ;
  assign y13533 = ~1'b0 ;
  assign y13534 = n26577 ;
  assign y13535 = n26579 ;
  assign y13536 = ~n26580 ;
  assign y13537 = n26581 ;
  assign y13538 = n26582 ;
  assign y13539 = ~1'b0 ;
  assign y13540 = n26584 ;
  assign y13541 = n26589 ;
  assign y13542 = ~1'b0 ;
  assign y13543 = n26592 ;
  assign y13544 = ~1'b0 ;
  assign y13545 = n26595 ;
  assign y13546 = ~n26601 ;
  assign y13547 = ~n26603 ;
  assign y13548 = n26607 ;
  assign y13549 = n26610 ;
  assign y13550 = n12281 ;
  assign y13551 = ~n26611 ;
  assign y13552 = ~1'b0 ;
  assign y13553 = ~n26612 ;
  assign y13554 = n2523 ;
  assign y13555 = ~n26615 ;
  assign y13556 = ~n26618 ;
  assign y13557 = n12940 ;
  assign y13558 = n26620 ;
  assign y13559 = n26621 ;
  assign y13560 = 1'b0 ;
  assign y13561 = n26623 ;
  assign y13562 = n26625 ;
  assign y13563 = ~1'b0 ;
  assign y13564 = n26627 ;
  assign y13565 = ~n26629 ;
  assign y13566 = ~n26631 ;
  assign y13567 = ~n26632 ;
  assign y13568 = ~1'b0 ;
  assign y13569 = ~1'b0 ;
  assign y13570 = ~n26633 ;
  assign y13571 = ~1'b0 ;
  assign y13572 = ~n26634 ;
  assign y13573 = ~n26637 ;
  assign y13574 = n26645 ;
  assign y13575 = ~n26646 ;
  assign y13576 = n26649 ;
  assign y13577 = ~1'b0 ;
  assign y13578 = n26651 ;
  assign y13579 = n26654 ;
  assign y13580 = n26659 ;
  assign y13581 = ~1'b0 ;
  assign y13582 = ~1'b0 ;
  assign y13583 = ~1'b0 ;
  assign y13584 = ~1'b0 ;
  assign y13585 = n26660 ;
  assign y13586 = n26662 ;
  assign y13587 = n26663 ;
  assign y13588 = ~1'b0 ;
  assign y13589 = ~1'b0 ;
  assign y13590 = ~n26667 ;
  assign y13591 = ~n4716 ;
  assign y13592 = ~1'b0 ;
  assign y13593 = ~1'b0 ;
  assign y13594 = n26669 ;
  assign y13595 = ~1'b0 ;
  assign y13596 = ~1'b0 ;
  assign y13597 = ~1'b0 ;
  assign y13598 = ~n26673 ;
  assign y13599 = n26674 ;
  assign y13600 = n26679 ;
  assign y13601 = ~1'b0 ;
  assign y13602 = n26684 ;
  assign y13603 = n26687 ;
  assign y13604 = ~n26688 ;
  assign y13605 = n26691 ;
  assign y13606 = ~n26692 ;
  assign y13607 = ~n26694 ;
  assign y13608 = ~1'b0 ;
  assign y13609 = ~1'b0 ;
  assign y13610 = ~n26697 ;
  assign y13611 = ~n26698 ;
  assign y13612 = ~n26703 ;
  assign y13613 = ~n26705 ;
  assign y13614 = ~n26706 ;
  assign y13615 = ~n26708 ;
  assign y13616 = n26710 ;
  assign y13617 = ~n26712 ;
  assign y13618 = n26714 ;
  assign y13619 = n26717 ;
  assign y13620 = n26721 ;
  assign y13621 = ~n1206 ;
  assign y13622 = ~1'b0 ;
  assign y13623 = ~n24418 ;
  assign y13624 = ~n8547 ;
  assign y13625 = n26722 ;
  assign y13626 = ~n26724 ;
  assign y13627 = ~n26725 ;
  assign y13628 = ~1'b0 ;
  assign y13629 = ~n26733 ;
  assign y13630 = n26735 ;
  assign y13631 = n26737 ;
  assign y13632 = ~n26739 ;
  assign y13633 = n26741 ;
  assign y13634 = ~1'b0 ;
  assign y13635 = ~1'b0 ;
  assign y13636 = ~n26749 ;
  assign y13637 = ~n26750 ;
  assign y13638 = ~n26763 ;
  assign y13639 = ~n26765 ;
  assign y13640 = ~1'b0 ;
  assign y13641 = n26767 ;
  assign y13642 = n26770 ;
  assign y13643 = ~n26773 ;
  assign y13644 = ~1'b0 ;
  assign y13645 = n26775 ;
  assign y13646 = ~n26776 ;
  assign y13647 = n26778 ;
  assign y13648 = n26780 ;
  assign y13649 = n26781 ;
  assign y13650 = ~1'b0 ;
  assign y13651 = ~n26782 ;
  assign y13652 = ~1'b0 ;
  assign y13653 = ~n26785 ;
  assign y13654 = n26786 ;
  assign y13655 = ~n26792 ;
  assign y13656 = ~n26793 ;
  assign y13657 = n6342 ;
  assign y13658 = ~1'b0 ;
  assign y13659 = ~n14479 ;
  assign y13660 = ~n26800 ;
  assign y13661 = n26808 ;
  assign y13662 = ~1'b0 ;
  assign y13663 = ~1'b0 ;
  assign y13664 = n26814 ;
  assign y13665 = ~n26816 ;
  assign y13666 = n9352 ;
  assign y13667 = ~1'b0 ;
  assign y13668 = ~1'b0 ;
  assign y13669 = n26817 ;
  assign y13670 = ~n26820 ;
  assign y13671 = n509 ;
  assign y13672 = ~1'b0 ;
  assign y13673 = n10327 ;
  assign y13674 = n26824 ;
  assign y13675 = n26825 ;
  assign y13676 = ~n19469 ;
  assign y13677 = ~n26827 ;
  assign y13678 = n26832 ;
  assign y13679 = n26838 ;
  assign y13680 = n26840 ;
  assign y13681 = n26843 ;
  assign y13682 = ~1'b0 ;
  assign y13683 = ~n19494 ;
  assign y13684 = ~1'b0 ;
  assign y13685 = ~1'b0 ;
  assign y13686 = n26844 ;
  assign y13687 = 1'b0 ;
  assign y13688 = ~1'b0 ;
  assign y13689 = ~1'b0 ;
  assign y13690 = ~n26846 ;
  assign y13691 = ~1'b0 ;
  assign y13692 = n26849 ;
  assign y13693 = n26853 ;
  assign y13694 = n6769 ;
  assign y13695 = n26854 ;
  assign y13696 = n26856 ;
  assign y13697 = ~1'b0 ;
  assign y13698 = ~1'b0 ;
  assign y13699 = ~1'b0 ;
  assign y13700 = ~n26861 ;
  assign y13701 = n26862 ;
  assign y13702 = n26863 ;
  assign y13703 = ~1'b0 ;
  assign y13704 = 1'b0 ;
  assign y13705 = 1'b0 ;
  assign y13706 = ~n26866 ;
  assign y13707 = x242 ;
  assign y13708 = n26870 ;
  assign y13709 = n26872 ;
  assign y13710 = ~1'b0 ;
  assign y13711 = ~1'b0 ;
  assign y13712 = ~1'b0 ;
  assign y13713 = ~n26873 ;
  assign y13714 = ~n26593 ;
  assign y13715 = n26877 ;
  assign y13716 = ~1'b0 ;
  assign y13717 = ~n26883 ;
  assign y13718 = n26884 ;
  assign y13719 = ~1'b0 ;
  assign y13720 = ~n26885 ;
  assign y13721 = ~n26887 ;
  assign y13722 = ~n26888 ;
  assign y13723 = ~1'b0 ;
  assign y13724 = ~n26890 ;
  assign y13725 = n26892 ;
  assign y13726 = ~n26893 ;
  assign y13727 = ~n26894 ;
  assign y13728 = n26902 ;
  assign y13729 = n26903 ;
  assign y13730 = ~n8941 ;
  assign y13731 = n26905 ;
  assign y13732 = n26908 ;
  assign y13733 = ~1'b0 ;
  assign y13734 = ~n26909 ;
  assign y13735 = ~n26910 ;
  assign y13736 = n26912 ;
  assign y13737 = n26913 ;
  assign y13738 = ~1'b0 ;
  assign y13739 = ~n26915 ;
  assign y13740 = ~n26919 ;
  assign y13741 = ~1'b0 ;
  assign y13742 = n26928 ;
  assign y13743 = ~1'b0 ;
  assign y13744 = ~n26933 ;
  assign y13745 = ~n26936 ;
  assign y13746 = ~n5054 ;
  assign y13747 = ~1'b0 ;
  assign y13748 = ~1'b0 ;
  assign y13749 = ~n26937 ;
  assign y13750 = n26938 ;
  assign y13751 = n26939 ;
  assign y13752 = n26941 ;
  assign y13753 = ~n26942 ;
  assign y13754 = ~n26944 ;
  assign y13755 = ~1'b0 ;
  assign y13756 = ~n26945 ;
  assign y13757 = n26947 ;
  assign y13758 = ~n25497 ;
  assign y13759 = n26948 ;
  assign y13760 = n26954 ;
  assign y13761 = ~1'b0 ;
  assign y13762 = n26956 ;
  assign y13763 = ~1'b0 ;
  assign y13764 = ~n26958 ;
  assign y13765 = ~n7491 ;
  assign y13766 = ~1'b0 ;
  assign y13767 = ~n26961 ;
  assign y13768 = ~1'b0 ;
  assign y13769 = n26963 ;
  assign y13770 = ~1'b0 ;
  assign y13771 = n12532 ;
  assign y13772 = ~1'b0 ;
  assign y13773 = ~n3996 ;
  assign y13774 = n26965 ;
  assign y13775 = ~n26966 ;
  assign y13776 = ~n26968 ;
  assign y13777 = ~1'b0 ;
  assign y13778 = ~1'b0 ;
  assign y13779 = n26969 ;
  assign y13780 = x159 ;
  assign y13781 = ~1'b0 ;
  assign y13782 = ~n26972 ;
  assign y13783 = ~1'b0 ;
  assign y13784 = ~1'b0 ;
  assign y13785 = ~n26977 ;
  assign y13786 = ~n26978 ;
  assign y13787 = ~1'b0 ;
  assign y13788 = ~n26981 ;
  assign y13789 = n18793 ;
  assign y13790 = ~n26984 ;
  assign y13791 = ~1'b0 ;
  assign y13792 = ~1'b0 ;
  assign y13793 = ~n26992 ;
  assign y13794 = n26996 ;
  assign y13795 = ~1'b0 ;
  assign y13796 = ~n26997 ;
  assign y13797 = n26999 ;
  assign y13798 = ~n27000 ;
  assign y13799 = ~n27001 ;
  assign y13800 = ~n27002 ;
  assign y13801 = n27006 ;
  assign y13802 = ~1'b0 ;
  assign y13803 = ~1'b0 ;
  assign y13804 = ~n27007 ;
  assign y13805 = ~1'b0 ;
  assign y13806 = ~n27008 ;
  assign y13807 = n27011 ;
  assign y13808 = n27012 ;
  assign y13809 = n27013 ;
  assign y13810 = ~1'b0 ;
  assign y13811 = n27015 ;
  assign y13812 = ~n27016 ;
  assign y13813 = ~n27018 ;
  assign y13814 = n27025 ;
  assign y13815 = ~1'b0 ;
  assign y13816 = n27027 ;
  assign y13817 = ~1'b0 ;
  assign y13818 = n27033 ;
  assign y13819 = ~1'b0 ;
  assign y13820 = ~n27035 ;
  assign y13821 = ~1'b0 ;
  assign y13822 = ~n27039 ;
  assign y13823 = ~n27042 ;
  assign y13824 = n27043 ;
  assign y13825 = n27044 ;
  assign y13826 = ~1'b0 ;
  assign y13827 = n27046 ;
  assign y13828 = ~1'b0 ;
  assign y13829 = n27050 ;
  assign y13830 = ~n27052 ;
  assign y13831 = ~n27053 ;
  assign y13832 = n27057 ;
  assign y13833 = n27059 ;
  assign y13834 = ~1'b0 ;
  assign y13835 = n27060 ;
  assign y13836 = ~1'b0 ;
  assign y13837 = n27062 ;
  assign y13838 = n27063 ;
  assign y13839 = ~1'b0 ;
  assign y13840 = ~1'b0 ;
  assign y13841 = ~n27064 ;
  assign y13842 = 1'b0 ;
  assign y13843 = ~1'b0 ;
  assign y13844 = n5836 ;
  assign y13845 = n27065 ;
  assign y13846 = n24078 ;
  assign y13847 = ~1'b0 ;
  assign y13848 = ~1'b0 ;
  assign y13849 = ~n27067 ;
  assign y13850 = n17337 ;
  assign y13851 = ~1'b0 ;
  assign y13852 = ~n27068 ;
  assign y13853 = ~1'b0 ;
  assign y13854 = ~n27074 ;
  assign y13855 = n27075 ;
  assign y13856 = n27079 ;
  assign y13857 = ~1'b0 ;
  assign y13858 = ~n27080 ;
  assign y13859 = n27082 ;
  assign y13860 = n27084 ;
  assign y13861 = n27086 ;
  assign y13862 = n27087 ;
  assign y13863 = ~1'b0 ;
  assign y13864 = ~n27089 ;
  assign y13865 = ~n27090 ;
  assign y13866 = ~n3846 ;
  assign y13867 = ~n27091 ;
  assign y13868 = n27092 ;
  assign y13869 = n27095 ;
  assign y13870 = ~n27097 ;
  assign y13871 = n27101 ;
  assign y13872 = n27103 ;
  assign y13873 = n27104 ;
  assign y13874 = ~n27106 ;
  assign y13875 = ~n27108 ;
  assign y13876 = ~1'b0 ;
  assign y13877 = ~1'b0 ;
  assign y13878 = ~n27109 ;
  assign y13879 = ~n27110 ;
  assign y13880 = ~n27115 ;
  assign y13881 = ~x242 ;
  assign y13882 = ~1'b0 ;
  assign y13883 = n27118 ;
  assign y13884 = n27125 ;
  assign y13885 = ~1'b0 ;
  assign y13886 = n14949 ;
  assign y13887 = n27126 ;
  assign y13888 = ~n4498 ;
  assign y13889 = n27127 ;
  assign y13890 = n27130 ;
  assign y13891 = ~n27132 ;
  assign y13892 = n27137 ;
  assign y13893 = ~1'b0 ;
  assign y13894 = n27138 ;
  assign y13895 = ~1'b0 ;
  assign y13896 = ~n27141 ;
  assign y13897 = ~1'b0 ;
  assign y13898 = ~n27142 ;
  assign y13899 = ~1'b0 ;
  assign y13900 = ~n27144 ;
  assign y13901 = n27145 ;
  assign y13902 = ~n27147 ;
  assign y13903 = 1'b0 ;
  assign y13904 = n27148 ;
  assign y13905 = ~n27153 ;
  assign y13906 = n27155 ;
  assign y13907 = ~n10354 ;
  assign y13908 = ~1'b0 ;
  assign y13909 = ~n27158 ;
  assign y13910 = n27168 ;
  assign y13911 = ~n27169 ;
  assign y13912 = ~1'b0 ;
  assign y13913 = n27170 ;
  assign y13914 = n27172 ;
  assign y13915 = n27173 ;
  assign y13916 = n27175 ;
  assign y13917 = n27177 ;
  assign y13918 = ~n27180 ;
  assign y13919 = 1'b0 ;
  assign y13920 = ~n27181 ;
  assign y13921 = ~n27182 ;
  assign y13922 = ~1'b0 ;
  assign y13923 = ~1'b0 ;
  assign y13924 = ~n8645 ;
  assign y13925 = ~1'b0 ;
  assign y13926 = ~n27184 ;
  assign y13927 = n27186 ;
  assign y13928 = ~1'b0 ;
  assign y13929 = ~n27187 ;
  assign y13930 = ~n27190 ;
  assign y13931 = ~1'b0 ;
  assign y13932 = n27191 ;
  assign y13933 = ~1'b0 ;
  assign y13934 = ~n27192 ;
  assign y13935 = n27194 ;
  assign y13936 = ~n27195 ;
  assign y13937 = n27199 ;
  assign y13938 = n1361 ;
  assign y13939 = n27203 ;
  assign y13940 = ~n27204 ;
  assign y13941 = n274 ;
  assign y13942 = ~1'b0 ;
  assign y13943 = n27209 ;
  assign y13944 = n27213 ;
  assign y13945 = n27214 ;
  assign y13946 = n27216 ;
  assign y13947 = ~n27217 ;
  assign y13948 = n27222 ;
  assign y13949 = ~n27223 ;
  assign y13950 = n27224 ;
  assign y13951 = ~1'b0 ;
  assign y13952 = ~1'b0 ;
  assign y13953 = n27225 ;
  assign y13954 = n27226 ;
  assign y13955 = n27227 ;
  assign y13956 = n27229 ;
  assign y13957 = ~n27232 ;
  assign y13958 = n27235 ;
  assign y13959 = n27239 ;
  assign y13960 = ~1'b0 ;
  assign y13961 = ~1'b0 ;
  assign y13962 = n27240 ;
  assign y13963 = ~1'b0 ;
  assign y13964 = ~n27245 ;
  assign y13965 = ~n27246 ;
  assign y13966 = ~1'b0 ;
  assign y13967 = 1'b0 ;
  assign y13968 = n27248 ;
  assign y13969 = n27251 ;
  assign y13970 = ~1'b0 ;
  assign y13971 = n21590 ;
  assign y13972 = n27257 ;
  assign y13973 = ~n27258 ;
  assign y13974 = ~n27259 ;
  assign y13975 = ~n27266 ;
  assign y13976 = ~1'b0 ;
  assign y13977 = n14094 ;
  assign y13978 = n27267 ;
  assign y13979 = n27268 ;
  assign y13980 = ~n27270 ;
  assign y13981 = ~n27271 ;
  assign y13982 = ~1'b0 ;
  assign y13983 = ~n27273 ;
  assign y13984 = n27275 ;
  assign y13985 = ~n27278 ;
  assign y13986 = ~n27279 ;
  assign y13987 = ~1'b0 ;
  assign y13988 = n27281 ;
  assign y13989 = ~1'b0 ;
  assign y13990 = ~1'b0 ;
  assign y13991 = ~1'b0 ;
  assign y13992 = ~1'b0 ;
  assign y13993 = ~n27282 ;
  assign y13994 = ~n27285 ;
  assign y13995 = ~n27287 ;
  assign y13996 = ~1'b0 ;
  assign y13997 = ~n27289 ;
  assign y13998 = ~n27292 ;
  assign y13999 = ~1'b0 ;
  assign y14000 = ~n27293 ;
  assign y14001 = ~1'b0 ;
  assign y14002 = n27295 ;
  assign y14003 = ~n27296 ;
  assign y14004 = ~1'b0 ;
  assign y14005 = ~n27297 ;
  assign y14006 = ~n27298 ;
  assign y14007 = n27306 ;
  assign y14008 = n27308 ;
  assign y14009 = ~1'b0 ;
  assign y14010 = ~1'b0 ;
  assign y14011 = ~n27311 ;
  assign y14012 = ~n27315 ;
  assign y14013 = ~n18356 ;
  assign y14014 = n13562 ;
  assign y14015 = ~n27318 ;
  assign y14016 = ~1'b0 ;
  assign y14017 = n27319 ;
  assign y14018 = n6177 ;
  assign y14019 = n27325 ;
  assign y14020 = ~n27330 ;
  assign y14021 = ~n2473 ;
  assign y14022 = n27333 ;
  assign y14023 = ~1'b0 ;
  assign y14024 = ~n27337 ;
  assign y14025 = ~1'b0 ;
  assign y14026 = ~1'b0 ;
  assign y14027 = x220 ;
  assign y14028 = ~n27338 ;
  assign y14029 = ~n27010 ;
  assign y14030 = n27340 ;
  assign y14031 = ~n27345 ;
  assign y14032 = n27348 ;
  assign y14033 = n27349 ;
  assign y14034 = 1'b0 ;
  assign y14035 = n27351 ;
  assign y14036 = ~n5582 ;
  assign y14037 = ~n27352 ;
  assign y14038 = ~n27355 ;
  assign y14039 = n27367 ;
  assign y14040 = ~1'b0 ;
  assign y14041 = ~n27376 ;
  assign y14042 = n5650 ;
  assign y14043 = n18310 ;
  assign y14044 = ~n27378 ;
  assign y14045 = ~n27380 ;
  assign y14046 = ~1'b0 ;
  assign y14047 = n27383 ;
  assign y14048 = ~1'b0 ;
  assign y14049 = 1'b0 ;
  assign y14050 = ~1'b0 ;
  assign y14051 = ~1'b0 ;
  assign y14052 = ~n27386 ;
  assign y14053 = n7449 ;
  assign y14054 = n27390 ;
  assign y14055 = ~1'b0 ;
  assign y14056 = ~1'b0 ;
  assign y14057 = n27391 ;
  assign y14058 = n27392 ;
  assign y14059 = ~n27396 ;
  assign y14060 = ~n27399 ;
  assign y14061 = ~n27400 ;
  assign y14062 = ~n27403 ;
  assign y14063 = ~1'b0 ;
  assign y14064 = ~1'b0 ;
  assign y14065 = ~1'b0 ;
  assign y14066 = n27410 ;
  assign y14067 = ~1'b0 ;
  assign y14068 = n8905 ;
  assign y14069 = n27411 ;
  assign y14070 = ~n27413 ;
  assign y14071 = n27415 ;
  assign y14072 = n3561 ;
  assign y14073 = n27429 ;
  assign y14074 = n27430 ;
  assign y14075 = n4562 ;
  assign y14076 = ~1'b0 ;
  assign y14077 = ~n27436 ;
  assign y14078 = ~n27440 ;
  assign y14079 = n27441 ;
  assign y14080 = ~n27446 ;
  assign y14081 = ~n27448 ;
  assign y14082 = ~1'b0 ;
  assign y14083 = ~n27457 ;
  assign y14084 = ~n27458 ;
  assign y14085 = ~n27459 ;
  assign y14086 = n11087 ;
  assign y14087 = n27461 ;
  assign y14088 = n27464 ;
  assign y14089 = n27466 ;
  assign y14090 = ~n27468 ;
  assign y14091 = ~n27473 ;
  assign y14092 = ~1'b0 ;
  assign y14093 = ~1'b0 ;
  assign y14094 = ~n27476 ;
  assign y14095 = ~n27478 ;
  assign y14096 = 1'b0 ;
  assign y14097 = ~1'b0 ;
  assign y14098 = n27479 ;
  assign y14099 = ~n27482 ;
  assign y14100 = ~1'b0 ;
  assign y14101 = ~1'b0 ;
  assign y14102 = n27486 ;
  assign y14103 = ~n27488 ;
  assign y14104 = ~n27490 ;
  assign y14105 = ~n27496 ;
  assign y14106 = ~n27497 ;
  assign y14107 = ~n27499 ;
  assign y14108 = ~n27500 ;
  assign y14109 = n27502 ;
  assign y14110 = ~1'b0 ;
  assign y14111 = ~n22982 ;
  assign y14112 = ~1'b0 ;
  assign y14113 = ~n27503 ;
  assign y14114 = ~1'b0 ;
  assign y14115 = ~n27505 ;
  assign y14116 = n27506 ;
  assign y14117 = n27507 ;
  assign y14118 = n27508 ;
  assign y14119 = ~1'b0 ;
  assign y14120 = ~n27510 ;
  assign y14121 = ~1'b0 ;
  assign y14122 = ~n27511 ;
  assign y14123 = ~n27513 ;
  assign y14124 = ~n6983 ;
  assign y14125 = n27514 ;
  assign y14126 = n27516 ;
  assign y14127 = n27519 ;
  assign y14128 = ~n27520 ;
  assign y14129 = n27523 ;
  assign y14130 = ~1'b0 ;
  assign y14131 = ~n27524 ;
  assign y14132 = n27526 ;
  assign y14133 = ~n27532 ;
  assign y14134 = ~n8008 ;
  assign y14135 = ~1'b0 ;
  assign y14136 = ~1'b0 ;
  assign y14137 = 1'b0 ;
  assign y14138 = ~1'b0 ;
  assign y14139 = ~n27534 ;
  assign y14140 = n27535 ;
  assign y14141 = ~1'b0 ;
  assign y14142 = n27538 ;
  assign y14143 = ~n27542 ;
  assign y14144 = ~n27543 ;
  assign y14145 = ~1'b0 ;
  assign y14146 = ~n27545 ;
  assign y14147 = ~1'b0 ;
  assign y14148 = ~1'b0 ;
  assign y14149 = ~n27547 ;
  assign y14150 = ~1'b0 ;
  assign y14151 = ~n27548 ;
  assign y14152 = 1'b0 ;
  assign y14153 = ~n27557 ;
  assign y14154 = ~n27558 ;
  assign y14155 = ~n27565 ;
  assign y14156 = ~n27567 ;
  assign y14157 = ~1'b0 ;
  assign y14158 = n27572 ;
  assign y14159 = ~1'b0 ;
  assign y14160 = n27574 ;
  assign y14161 = ~n794 ;
  assign y14162 = n27577 ;
  assign y14163 = ~n27578 ;
  assign y14164 = n27582 ;
  assign y14165 = ~n27590 ;
  assign y14166 = ~n27591 ;
  assign y14167 = ~n27592 ;
  assign y14168 = n27593 ;
  assign y14169 = ~1'b0 ;
  assign y14170 = n27595 ;
  assign y14171 = ~1'b0 ;
  assign y14172 = n27597 ;
  assign y14173 = ~n27598 ;
  assign y14174 = n27599 ;
  assign y14175 = ~n27600 ;
  assign y14176 = ~n27610 ;
  assign y14177 = ~n27618 ;
  assign y14178 = ~n27620 ;
  assign y14179 = 1'b0 ;
  assign y14180 = ~n27621 ;
  assign y14181 = ~n27623 ;
  assign y14182 = ~1'b0 ;
  assign y14183 = ~n27624 ;
  assign y14184 = ~n27625 ;
  assign y14185 = ~n27627 ;
  assign y14186 = ~1'b0 ;
  assign y14187 = ~1'b0 ;
  assign y14188 = n27630 ;
  assign y14189 = ~n27632 ;
  assign y14190 = ~1'b0 ;
  assign y14191 = ~n27635 ;
  assign y14192 = ~1'b0 ;
  assign y14193 = ~n27638 ;
  assign y14194 = ~1'b0 ;
  assign y14195 = ~1'b0 ;
  assign y14196 = ~n27642 ;
  assign y14197 = n27644 ;
  assign y14198 = ~n16333 ;
  assign y14199 = ~1'b0 ;
  assign y14200 = ~1'b0 ;
  assign y14201 = ~1'b0 ;
  assign y14202 = ~1'b0 ;
  assign y14203 = n27652 ;
  assign y14204 = ~1'b0 ;
  assign y14205 = ~n27655 ;
  assign y14206 = ~n27657 ;
  assign y14207 = ~1'b0 ;
  assign y14208 = ~1'b0 ;
  assign y14209 = ~1'b0 ;
  assign y14210 = ~n27658 ;
  assign y14211 = n27661 ;
  assign y14212 = n27664 ;
  assign y14213 = n2980 ;
  assign y14214 = ~n27667 ;
  assign y14215 = n27668 ;
  assign y14216 = ~1'b0 ;
  assign y14217 = n10164 ;
  assign y14218 = ~n27671 ;
  assign y14219 = ~1'b0 ;
  assign y14220 = ~1'b0 ;
  assign y14221 = ~n27677 ;
  assign y14222 = ~n27680 ;
  assign y14223 = ~1'b0 ;
  assign y14224 = ~n2697 ;
  assign y14225 = 1'b0 ;
  assign y14226 = n27684 ;
  assign y14227 = ~1'b0 ;
  assign y14228 = ~1'b0 ;
  assign y14229 = n8886 ;
  assign y14230 = ~1'b0 ;
  assign y14231 = ~n27694 ;
  assign y14232 = ~n27696 ;
  assign y14233 = n27703 ;
  assign y14234 = ~n27705 ;
  assign y14235 = n27711 ;
  assign y14236 = n27713 ;
  assign y14237 = ~n27717 ;
  assign y14238 = ~n27718 ;
  assign y14239 = ~n27725 ;
  assign y14240 = ~n27726 ;
  assign y14241 = n27728 ;
  assign y14242 = ~n27729 ;
  assign y14243 = ~n25024 ;
  assign y14244 = ~1'b0 ;
  assign y14245 = ~1'b0 ;
  assign y14246 = n970 ;
  assign y14247 = ~1'b0 ;
  assign y14248 = ~n27732 ;
  assign y14249 = ~1'b0 ;
  assign y14250 = ~n27734 ;
  assign y14251 = ~n27735 ;
  assign y14252 = ~n27736 ;
  assign y14253 = ~1'b0 ;
  assign y14254 = ~1'b0 ;
  assign y14255 = ~1'b0 ;
  assign y14256 = ~n27738 ;
  assign y14257 = ~1'b0 ;
  assign y14258 = ~n27741 ;
  assign y14259 = ~1'b0 ;
  assign y14260 = n27744 ;
  assign y14261 = n27746 ;
  assign y14262 = ~1'b0 ;
  assign y14263 = ~n27758 ;
  assign y14264 = ~1'b0 ;
  assign y14265 = ~n27760 ;
  assign y14266 = ~n27761 ;
  assign y14267 = ~n26498 ;
  assign y14268 = n6811 ;
  assign y14269 = ~1'b0 ;
  assign y14270 = ~1'b0 ;
  assign y14271 = ~n27764 ;
  assign y14272 = n27777 ;
  assign y14273 = n27779 ;
  assign y14274 = n27780 ;
  assign y14275 = n27784 ;
  assign y14276 = ~n27786 ;
  assign y14277 = n27787 ;
  assign y14278 = ~1'b0 ;
  assign y14279 = ~n4976 ;
  assign y14280 = ~1'b0 ;
  assign y14281 = ~n27789 ;
  assign y14282 = n4443 ;
  assign y14283 = ~n12384 ;
  assign y14284 = n27790 ;
  assign y14285 = ~n27792 ;
  assign y14286 = n27795 ;
  assign y14287 = n27797 ;
  assign y14288 = ~n27798 ;
  assign y14289 = ~n27803 ;
  assign y14290 = ~n27805 ;
  assign y14291 = ~n27806 ;
  assign y14292 = 1'b0 ;
  assign y14293 = ~n27807 ;
  assign y14294 = ~n27815 ;
  assign y14295 = ~1'b0 ;
  assign y14296 = ~1'b0 ;
  assign y14297 = n27819 ;
  assign y14298 = ~1'b0 ;
  assign y14299 = ~1'b0 ;
  assign y14300 = n14937 ;
  assign y14301 = ~1'b0 ;
  assign y14302 = ~1'b0 ;
  assign y14303 = ~1'b0 ;
  assign y14304 = ~1'b0 ;
  assign y14305 = ~n27822 ;
  assign y14306 = n27824 ;
  assign y14307 = n27827 ;
  assign y14308 = ~1'b0 ;
  assign y14309 = ~n27829 ;
  assign y14310 = ~n27833 ;
  assign y14311 = ~1'b0 ;
  assign y14312 = ~n27336 ;
  assign y14313 = ~n27836 ;
  assign y14314 = n27839 ;
  assign y14315 = n27845 ;
  assign y14316 = ~n27847 ;
  assign y14317 = ~n27848 ;
  assign y14318 = ~n27849 ;
  assign y14319 = 1'b0 ;
  assign y14320 = ~n27851 ;
  assign y14321 = 1'b0 ;
  assign y14322 = ~1'b0 ;
  assign y14323 = ~1'b0 ;
  assign y14324 = ~1'b0 ;
  assign y14325 = n27854 ;
  assign y14326 = ~1'b0 ;
  assign y14327 = ~1'b0 ;
  assign y14328 = ~1'b0 ;
  assign y14329 = n27858 ;
  assign y14330 = ~1'b0 ;
  assign y14331 = ~n27861 ;
  assign y14332 = ~1'b0 ;
  assign y14333 = ~1'b0 ;
  assign y14334 = n13747 ;
  assign y14335 = ~n27862 ;
  assign y14336 = n27043 ;
  assign y14337 = ~n27863 ;
  assign y14338 = n27864 ;
  assign y14339 = ~n9597 ;
  assign y14340 = ~n27865 ;
  assign y14341 = ~n26619 ;
  assign y14342 = ~n27868 ;
  assign y14343 = 1'b0 ;
  assign y14344 = n27869 ;
  assign y14345 = n27877 ;
  assign y14346 = ~1'b0 ;
  assign y14347 = ~n27879 ;
  assign y14348 = ~1'b0 ;
  assign y14349 = 1'b0 ;
  assign y14350 = n26935 ;
  assign y14351 = ~n27883 ;
  assign y14352 = ~1'b0 ;
  assign y14353 = ~n27885 ;
  assign y14354 = n27887 ;
  assign y14355 = n27891 ;
  assign y14356 = ~n27897 ;
  assign y14357 = ~n27905 ;
  assign y14358 = n27907 ;
  assign y14359 = ~n27909 ;
  assign y14360 = ~n27913 ;
  assign y14361 = ~n27914 ;
  assign y14362 = ~n27915 ;
  assign y14363 = n27916 ;
  assign y14364 = ~1'b0 ;
  assign y14365 = ~n27918 ;
  assign y14366 = n27919 ;
  assign y14367 = ~1'b0 ;
  assign y14368 = n22079 ;
  assign y14369 = ~n27921 ;
  assign y14370 = ~n27922 ;
  assign y14371 = n27924 ;
  assign y14372 = n27925 ;
  assign y14373 = ~n27927 ;
  assign y14374 = ~n27935 ;
  assign y14375 = n27937 ;
  assign y14376 = n27945 ;
  assign y14377 = ~1'b0 ;
  assign y14378 = ~1'b0 ;
  assign y14379 = ~n27946 ;
  assign y14380 = ~1'b0 ;
  assign y14381 = ~1'b0 ;
  assign y14382 = 1'b0 ;
  assign y14383 = ~1'b0 ;
  assign y14384 = ~n19650 ;
  assign y14385 = ~n27947 ;
  assign y14386 = ~1'b0 ;
  assign y14387 = ~1'b0 ;
  assign y14388 = n27951 ;
  assign y14389 = ~1'b0 ;
  assign y14390 = ~n27952 ;
  assign y14391 = n27953 ;
  assign y14392 = ~n2560 ;
  assign y14393 = ~1'b0 ;
  assign y14394 = ~1'b0 ;
  assign y14395 = ~1'b0 ;
  assign y14396 = ~n27956 ;
  assign y14397 = ~n14493 ;
  assign y14398 = n27960 ;
  assign y14399 = ~n27966 ;
  assign y14400 = ~1'b0 ;
  assign y14401 = n27967 ;
  assign y14402 = n27972 ;
  assign y14403 = ~n27974 ;
  assign y14404 = ~1'b0 ;
  assign y14405 = n6454 ;
  assign y14406 = ~n27976 ;
  assign y14407 = ~n27977 ;
  assign y14408 = ~1'b0 ;
  assign y14409 = ~n27981 ;
  assign y14410 = ~1'b0 ;
  assign y14411 = ~n27986 ;
  assign y14412 = n27987 ;
  assign y14413 = n27988 ;
  assign y14414 = ~n27989 ;
  assign y14415 = 1'b0 ;
  assign y14416 = ~n27991 ;
  assign y14417 = ~n27993 ;
  assign y14418 = n27998 ;
  assign y14419 = n27999 ;
  assign y14420 = n28000 ;
  assign y14421 = ~n11234 ;
  assign y14422 = ~n28002 ;
  assign y14423 = n28005 ;
  assign y14424 = ~n28006 ;
  assign y14425 = ~n28007 ;
  assign y14426 = n28008 ;
  assign y14427 = ~1'b0 ;
  assign y14428 = ~n28011 ;
  assign y14429 = ~1'b0 ;
  assign y14430 = n28012 ;
  assign y14431 = n28014 ;
  assign y14432 = ~1'b0 ;
  assign y14433 = n28015 ;
  assign y14434 = n18572 ;
  assign y14435 = ~n28019 ;
  assign y14436 = ~1'b0 ;
  assign y14437 = n28020 ;
  assign y14438 = ~n28021 ;
  assign y14439 = ~n28025 ;
  assign y14440 = ~1'b0 ;
  assign y14441 = ~n28027 ;
  assign y14442 = ~1'b0 ;
  assign y14443 = ~n25729 ;
  assign y14444 = n28028 ;
  assign y14445 = ~n3353 ;
  assign y14446 = n28037 ;
  assign y14447 = ~1'b0 ;
  assign y14448 = n28039 ;
  assign y14449 = ~n28045 ;
  assign y14450 = n28051 ;
  assign y14451 = n28054 ;
  assign y14452 = ~n28059 ;
  assign y14453 = n28064 ;
  assign y14454 = ~n28065 ;
  assign y14455 = ~n16934 ;
  assign y14456 = n28070 ;
  assign y14457 = n28076 ;
  assign y14458 = n28080 ;
  assign y14459 = n4844 ;
  assign y14460 = n28081 ;
  assign y14461 = ~n28082 ;
  assign y14462 = ~1'b0 ;
  assign y14463 = ~1'b0 ;
  assign y14464 = ~n28089 ;
  assign y14465 = ~n28097 ;
  assign y14466 = ~n28099 ;
  assign y14467 = ~n28103 ;
  assign y14468 = ~1'b0 ;
  assign y14469 = 1'b0 ;
  assign y14470 = ~1'b0 ;
  assign y14471 = n28105 ;
  assign y14472 = ~1'b0 ;
  assign y14473 = ~1'b0 ;
  assign y14474 = ~1'b0 ;
  assign y14475 = n28106 ;
  assign y14476 = ~1'b0 ;
  assign y14477 = n5626 ;
  assign y14478 = n28109 ;
  assign y14479 = ~n28110 ;
  assign y14480 = ~1'b0 ;
  assign y14481 = ~1'b0 ;
  assign y14482 = ~n28114 ;
  assign y14483 = n28116 ;
  assign y14484 = ~n28118 ;
  assign y14485 = n28120 ;
  assign y14486 = n28126 ;
  assign y14487 = ~1'b0 ;
  assign y14488 = ~1'b0 ;
  assign y14489 = n28127 ;
  assign y14490 = n12857 ;
  assign y14491 = n28130 ;
  assign y14492 = ~1'b0 ;
  assign y14493 = ~1'b0 ;
  assign y14494 = n28132 ;
  assign y14495 = ~n19464 ;
  assign y14496 = ~n28134 ;
  assign y14497 = ~n28136 ;
  assign y14498 = ~n5530 ;
  assign y14499 = ~1'b0 ;
  assign y14500 = n28140 ;
  assign y14501 = ~n28147 ;
  assign y14502 = ~n28149 ;
  assign y14503 = n28151 ;
  assign y14504 = ~n28152 ;
  assign y14505 = ~1'b0 ;
  assign y14506 = n28153 ;
  assign y14507 = ~n28155 ;
  assign y14508 = ~1'b0 ;
  assign y14509 = ~n28157 ;
  assign y14510 = ~1'b0 ;
  assign y14511 = ~n28158 ;
  assign y14512 = ~n28161 ;
  assign y14513 = ~n28167 ;
  assign y14514 = ~1'b0 ;
  assign y14515 = ~1'b0 ;
  assign y14516 = ~1'b0 ;
  assign y14517 = ~n28171 ;
  assign y14518 = ~n19013 ;
  assign y14519 = ~1'b0 ;
  assign y14520 = ~1'b0 ;
  assign y14521 = ~n28173 ;
  assign y14522 = ~n28174 ;
  assign y14523 = ~n24070 ;
  assign y14524 = ~n28178 ;
  assign y14525 = n28181 ;
  assign y14526 = n28185 ;
  assign y14527 = ~n28189 ;
  assign y14528 = ~1'b0 ;
  assign y14529 = ~1'b0 ;
  assign y14530 = ~1'b0 ;
  assign y14531 = ~n28191 ;
  assign y14532 = ~1'b0 ;
  assign y14533 = ~1'b0 ;
  assign y14534 = ~n28192 ;
  assign y14535 = ~n6274 ;
  assign y14536 = ~n28194 ;
  assign y14537 = n28196 ;
  assign y14538 = ~1'b0 ;
  assign y14539 = ~n28201 ;
  assign y14540 = n28207 ;
  assign y14541 = ~1'b0 ;
  assign y14542 = ~n28208 ;
  assign y14543 = n28210 ;
  assign y14544 = ~n28219 ;
  assign y14545 = 1'b0 ;
  assign y14546 = ~1'b0 ;
  assign y14547 = ~n28221 ;
  assign y14548 = ~1'b0 ;
  assign y14549 = n28223 ;
  assign y14550 = n28227 ;
  assign y14551 = n28231 ;
  assign y14552 = n28243 ;
  assign y14553 = ~n28244 ;
  assign y14554 = ~1'b0 ;
  assign y14555 = n23891 ;
  assign y14556 = ~n9048 ;
  assign y14557 = ~1'b0 ;
  assign y14558 = n28246 ;
  assign y14559 = ~1'b0 ;
  assign y14560 = ~n10484 ;
  assign y14561 = n28248 ;
  assign y14562 = ~1'b0 ;
  assign y14563 = 1'b0 ;
  assign y14564 = ~1'b0 ;
  assign y14565 = ~1'b0 ;
  assign y14566 = n28252 ;
  assign y14567 = n28253 ;
  assign y14568 = n25084 ;
  assign y14569 = ~n28256 ;
  assign y14570 = ~n28259 ;
  assign y14571 = ~n28261 ;
  assign y14572 = ~1'b0 ;
  assign y14573 = ~n28262 ;
  assign y14574 = ~1'b0 ;
  assign y14575 = ~n16612 ;
  assign y14576 = n28263 ;
  assign y14577 = ~1'b0 ;
  assign y14578 = x188 ;
  assign y14579 = n28266 ;
  assign y14580 = n10770 ;
  assign y14581 = ~n28270 ;
  assign y14582 = ~n28274 ;
  assign y14583 = ~1'b0 ;
  assign y14584 = n28275 ;
  assign y14585 = n2337 ;
  assign y14586 = n28276 ;
  assign y14587 = n28277 ;
  assign y14588 = n28278 ;
  assign y14589 = n28279 ;
  assign y14590 = 1'b0 ;
  assign y14591 = ~n28285 ;
  assign y14592 = ~n28286 ;
  assign y14593 = ~n28291 ;
  assign y14594 = ~n28292 ;
  assign y14595 = ~1'b0 ;
  assign y14596 = ~1'b0 ;
  assign y14597 = ~n28293 ;
  assign y14598 = n28295 ;
  assign y14599 = ~1'b0 ;
  assign y14600 = n28296 ;
  assign y14601 = ~1'b0 ;
  assign y14602 = ~1'b0 ;
  assign y14603 = 1'b0 ;
  assign y14604 = ~1'b0 ;
  assign y14605 = n28297 ;
  assign y14606 = ~n28303 ;
  assign y14607 = ~n28306 ;
  assign y14608 = ~1'b0 ;
  assign y14609 = ~n28314 ;
  assign y14610 = ~n3588 ;
  assign y14611 = ~1'b0 ;
  assign y14612 = ~n28315 ;
  assign y14613 = ~n28316 ;
  assign y14614 = n28317 ;
  assign y14615 = ~n28324 ;
  assign y14616 = n28326 ;
  assign y14617 = n28327 ;
  assign y14618 = ~n28328 ;
  assign y14619 = n28332 ;
  assign y14620 = ~1'b0 ;
  assign y14621 = n28337 ;
  assign y14622 = ~1'b0 ;
  assign y14623 = n28340 ;
  assign y14624 = n28350 ;
  assign y14625 = n22334 ;
  assign y14626 = ~n28352 ;
  assign y14627 = n28357 ;
  assign y14628 = ~n28360 ;
  assign y14629 = 1'b0 ;
  assign y14630 = ~1'b0 ;
  assign y14631 = ~1'b0 ;
  assign y14632 = n28367 ;
  assign y14633 = ~n28370 ;
  assign y14634 = ~1'b0 ;
  assign y14635 = n28372 ;
  assign y14636 = n28374 ;
  assign y14637 = ~1'b0 ;
  assign y14638 = n28375 ;
  assign y14639 = n28381 ;
  assign y14640 = ~n28382 ;
  assign y14641 = n28345 ;
  assign y14642 = ~1'b0 ;
  assign y14643 = ~1'b0 ;
  assign y14644 = ~n28385 ;
  assign y14645 = ~n28388 ;
  assign y14646 = ~n28394 ;
  assign y14647 = ~n28410 ;
  assign y14648 = ~1'b0 ;
  assign y14649 = ~n28412 ;
  assign y14650 = ~1'b0 ;
  assign y14651 = ~n28414 ;
  assign y14652 = ~1'b0 ;
  assign y14653 = n28417 ;
  assign y14654 = n8309 ;
  assign y14655 = n28419 ;
  assign y14656 = n28420 ;
  assign y14657 = n28421 ;
  assign y14658 = ~n28422 ;
  assign y14659 = ~n16621 ;
  assign y14660 = ~n28428 ;
  assign y14661 = n28430 ;
  assign y14662 = ~n28431 ;
  assign y14663 = n28433 ;
  assign y14664 = ~1'b0 ;
  assign y14665 = n28436 ;
  assign y14666 = ~1'b0 ;
  assign y14667 = ~n28437 ;
  assign y14668 = n28438 ;
  assign y14669 = n28439 ;
  assign y14670 = 1'b0 ;
  assign y14671 = n28441 ;
  assign y14672 = ~n28444 ;
  assign y14673 = ~1'b0 ;
  assign y14674 = ~n28448 ;
  assign y14675 = ~n28452 ;
  assign y14676 = ~n28455 ;
  assign y14677 = n28462 ;
  assign y14678 = ~1'b0 ;
  assign y14679 = ~n28463 ;
  assign y14680 = n28080 ;
  assign y14681 = n28467 ;
  assign y14682 = n28470 ;
  assign y14683 = ~n7704 ;
  assign y14684 = n28474 ;
  assign y14685 = ~1'b0 ;
  assign y14686 = ~n26517 ;
  assign y14687 = ~1'b0 ;
  assign y14688 = ~n28476 ;
  assign y14689 = ~n28477 ;
  assign y14690 = n28489 ;
  assign y14691 = ~n28490 ;
  assign y14692 = ~n28493 ;
  assign y14693 = n15745 ;
  assign y14694 = n28494 ;
  assign y14695 = n28497 ;
  assign y14696 = 1'b0 ;
  assign y14697 = 1'b0 ;
  assign y14698 = n28500 ;
  assign y14699 = ~n28501 ;
  assign y14700 = ~1'b0 ;
  assign y14701 = ~1'b0 ;
  assign y14702 = ~1'b0 ;
  assign y14703 = n28504 ;
  assign y14704 = ~n28505 ;
  assign y14705 = ~n28507 ;
  assign y14706 = n15792 ;
  assign y14707 = ~n28509 ;
  assign y14708 = n28510 ;
  assign y14709 = n28514 ;
  assign y14710 = ~1'b0 ;
  assign y14711 = ~n28518 ;
  assign y14712 = ~n28520 ;
  assign y14713 = ~n28522 ;
  assign y14714 = ~1'b0 ;
  assign y14715 = n28527 ;
  assign y14716 = ~1'b0 ;
  assign y14717 = ~n28532 ;
  assign y14718 = n28540 ;
  assign y14719 = ~n28542 ;
  assign y14720 = ~n28545 ;
  assign y14721 = ~1'b0 ;
  assign y14722 = ~1'b0 ;
  assign y14723 = ~n28547 ;
  assign y14724 = ~n28553 ;
  assign y14725 = ~1'b0 ;
  assign y14726 = ~1'b0 ;
  assign y14727 = ~n28554 ;
  assign y14728 = ~n28556 ;
  assign y14729 = n28566 ;
  assign y14730 = ~1'b0 ;
  assign y14731 = ~n28569 ;
  assign y14732 = ~n28572 ;
  assign y14733 = n28575 ;
  assign y14734 = n26257 ;
  assign y14735 = ~n28577 ;
  assign y14736 = ~1'b0 ;
  assign y14737 = n28581 ;
  assign y14738 = ~1'b0 ;
  assign y14739 = ~n28590 ;
  assign y14740 = n28591 ;
  assign y14741 = n28594 ;
  assign y14742 = n28596 ;
  assign y14743 = ~n28598 ;
  assign y14744 = n28600 ;
  assign y14745 = ~1'b0 ;
  assign y14746 = ~n28602 ;
  assign y14747 = ~n28607 ;
  assign y14748 = ~n28608 ;
  assign y14749 = ~1'b0 ;
  assign y14750 = ~n28609 ;
  assign y14751 = ~1'b0 ;
  assign y14752 = ~1'b0 ;
  assign y14753 = n5835 ;
  assign y14754 = ~n28614 ;
  assign y14755 = ~n28618 ;
  assign y14756 = n357 ;
  assign y14757 = n28621 ;
  assign y14758 = ~n28626 ;
  assign y14759 = n28629 ;
  assign y14760 = ~1'b0 ;
  assign y14761 = ~n28631 ;
  assign y14762 = ~1'b0 ;
  assign y14763 = n28632 ;
  assign y14764 = ~1'b0 ;
  assign y14765 = ~1'b0 ;
  assign y14766 = ~1'b0 ;
  assign y14767 = n28635 ;
  assign y14768 = ~1'b0 ;
  assign y14769 = n28637 ;
  assign y14770 = ~1'b0 ;
  assign y14771 = ~1'b0 ;
  assign y14772 = n28641 ;
  assign y14773 = ~1'b0 ;
  assign y14774 = n28647 ;
  assign y14775 = n28653 ;
  assign y14776 = n28654 ;
  assign y14777 = ~n28660 ;
  assign y14778 = ~n28666 ;
  assign y14779 = ~1'b0 ;
  assign y14780 = 1'b0 ;
  assign y14781 = n28667 ;
  assign y14782 = ~1'b0 ;
  assign y14783 = ~1'b0 ;
  assign y14784 = ~1'b0 ;
  assign y14785 = ~n1545 ;
  assign y14786 = n28668 ;
  assign y14787 = n28670 ;
  assign y14788 = n28683 ;
  assign y14789 = ~n28684 ;
  assign y14790 = ~1'b0 ;
  assign y14791 = ~n28685 ;
  assign y14792 = ~n28688 ;
  assign y14793 = n28692 ;
  assign y14794 = ~n28694 ;
  assign y14795 = ~n28695 ;
  assign y14796 = n28697 ;
  assign y14797 = n28700 ;
  assign y14798 = ~1'b0 ;
  assign y14799 = ~1'b0 ;
  assign y14800 = ~1'b0 ;
  assign y14801 = n28701 ;
  assign y14802 = ~n28704 ;
  assign y14803 = ~n28709 ;
  assign y14804 = ~1'b0 ;
  assign y14805 = n28716 ;
  assign y14806 = ~n28717 ;
  assign y14807 = ~n28719 ;
  assign y14808 = ~n28721 ;
  assign y14809 = ~1'b0 ;
  assign y14810 = ~1'b0 ;
  assign y14811 = ~n28723 ;
  assign y14812 = 1'b0 ;
  assign y14813 = n4824 ;
  assign y14814 = ~n28726 ;
  assign y14815 = ~1'b0 ;
  assign y14816 = ~1'b0 ;
  assign y14817 = ~n28727 ;
  assign y14818 = ~n28729 ;
  assign y14819 = n28730 ;
  assign y14820 = ~1'b0 ;
  assign y14821 = ~1'b0 ;
  assign y14822 = n15026 ;
  assign y14823 = ~n28733 ;
  assign y14824 = ~n28735 ;
  assign y14825 = ~1'b0 ;
  assign y14826 = n14360 ;
  assign y14827 = ~n28737 ;
  assign y14828 = n28738 ;
  assign y14829 = ~n6046 ;
  assign y14830 = n28740 ;
  assign y14831 = ~1'b0 ;
  assign y14832 = n28743 ;
  assign y14833 = ~1'b0 ;
  assign y14834 = 1'b0 ;
  assign y14835 = n28744 ;
  assign y14836 = n28747 ;
  assign y14837 = n28748 ;
  assign y14838 = ~n28754 ;
  assign y14839 = ~n28757 ;
  assign y14840 = ~n28759 ;
  assign y14841 = ~1'b0 ;
  assign y14842 = 1'b0 ;
  assign y14843 = n28762 ;
  assign y14844 = ~n28769 ;
  assign y14845 = 1'b0 ;
  assign y14846 = 1'b0 ;
  assign y14847 = ~1'b0 ;
  assign y14848 = ~1'b0 ;
  assign y14849 = n28771 ;
  assign y14850 = ~n28772 ;
  assign y14851 = ~1'b0 ;
  assign y14852 = ~n28773 ;
  assign y14853 = n28779 ;
  assign y14854 = n19886 ;
  assign y14855 = ~1'b0 ;
  assign y14856 = n28780 ;
  assign y14857 = ~1'b0 ;
  assign y14858 = ~n28783 ;
  assign y14859 = ~n28784 ;
  assign y14860 = ~1'b0 ;
  assign y14861 = ~1'b0 ;
  assign y14862 = n28785 ;
  assign y14863 = n28786 ;
  assign y14864 = ~1'b0 ;
  assign y14865 = ~n28787 ;
  assign y14866 = ~1'b0 ;
  assign y14867 = n28791 ;
  assign y14868 = ~1'b0 ;
  assign y14869 = n28792 ;
  assign y14870 = ~n28798 ;
  assign y14871 = ~1'b0 ;
  assign y14872 = ~n28799 ;
  assign y14873 = ~1'b0 ;
  assign y14874 = ~n28801 ;
  assign y14875 = ~1'b0 ;
  assign y14876 = ~n28806 ;
  assign y14877 = n28807 ;
  assign y14878 = n28818 ;
  assign y14879 = ~n28821 ;
  assign y14880 = n28822 ;
  assign y14881 = n28825 ;
  assign y14882 = ~1'b0 ;
  assign y14883 = ~1'b0 ;
  assign y14884 = ~1'b0 ;
  assign y14885 = n20464 ;
  assign y14886 = ~n28826 ;
  assign y14887 = n28827 ;
  assign y14888 = n28829 ;
  assign y14889 = ~1'b0 ;
  assign y14890 = n28833 ;
  assign y14891 = n28834 ;
  assign y14892 = ~n28836 ;
  assign y14893 = ~n8578 ;
  assign y14894 = ~1'b0 ;
  assign y14895 = ~1'b0 ;
  assign y14896 = ~n28839 ;
  assign y14897 = ~n19297 ;
  assign y14898 = ~1'b0 ;
  assign y14899 = n28840 ;
  assign y14900 = ~n28843 ;
  assign y14901 = 1'b0 ;
  assign y14902 = ~n28844 ;
  assign y14903 = n28845 ;
  assign y14904 = ~n28847 ;
  assign y14905 = n28848 ;
  assign y14906 = n28852 ;
  assign y14907 = ~1'b0 ;
  assign y14908 = 1'b0 ;
  assign y14909 = ~n28854 ;
  assign y14910 = n28858 ;
  assign y14911 = ~n28863 ;
  assign y14912 = ~1'b0 ;
  assign y14913 = ~1'b0 ;
  assign y14914 = n28864 ;
  assign y14915 = ~1'b0 ;
  assign y14916 = n28869 ;
  assign y14917 = ~n28870 ;
  assign y14918 = n28873 ;
  assign y14919 = ~n28876 ;
  assign y14920 = n28879 ;
  assign y14921 = ~n7877 ;
  assign y14922 = n28880 ;
  assign y14923 = ~1'b0 ;
  assign y14924 = n28882 ;
  assign y14925 = n28887 ;
  assign y14926 = ~n25646 ;
  assign y14927 = ~n28897 ;
  assign y14928 = ~1'b0 ;
  assign y14929 = ~n1295 ;
  assign y14930 = n28898 ;
  assign y14931 = ~1'b0 ;
  assign y14932 = n28902 ;
  assign y14933 = ~n28907 ;
  assign y14934 = ~1'b0 ;
  assign y14935 = 1'b0 ;
  assign y14936 = ~1'b0 ;
  assign y14937 = ~1'b0 ;
  assign y14938 = ~n28911 ;
  assign y14939 = n28912 ;
  assign y14940 = ~n28915 ;
  assign y14941 = ~n28917 ;
  assign y14942 = n16137 ;
  assign y14943 = n28918 ;
  assign y14944 = ~1'b0 ;
  assign y14945 = n28919 ;
  assign y14946 = ~n28920 ;
  assign y14947 = n28921 ;
  assign y14948 = n8974 ;
  assign y14949 = n28923 ;
  assign y14950 = n19491 ;
  assign y14951 = ~n28924 ;
  assign y14952 = ~1'b0 ;
  assign y14953 = ~n28927 ;
  assign y14954 = n28929 ;
  assign y14955 = ~n28931 ;
  assign y14956 = ~n28932 ;
  assign y14957 = n28933 ;
  assign y14958 = ~n28934 ;
  assign y14959 = ~n28935 ;
  assign y14960 = n28938 ;
  assign y14961 = ~1'b0 ;
  assign y14962 = n28939 ;
  assign y14963 = n28940 ;
  assign y14964 = ~1'b0 ;
  assign y14965 = ~1'b0 ;
  assign y14966 = 1'b0 ;
  assign y14967 = n28943 ;
  assign y14968 = n28944 ;
  assign y14969 = n28950 ;
  assign y14970 = ~1'b0 ;
  assign y14971 = n28952 ;
  assign y14972 = n28954 ;
  assign y14973 = ~1'b0 ;
  assign y14974 = n28955 ;
  assign y14975 = ~1'b0 ;
  assign y14976 = ~n28957 ;
  assign y14977 = ~1'b0 ;
  assign y14978 = n28958 ;
  assign y14979 = ~1'b0 ;
  assign y14980 = ~1'b0 ;
  assign y14981 = ~1'b0 ;
  assign y14982 = ~n28959 ;
  assign y14983 = ~n28964 ;
  assign y14984 = ~1'b0 ;
  assign y14985 = n28966 ;
  assign y14986 = ~n7222 ;
  assign y14987 = ~n28056 ;
  assign y14988 = n28967 ;
  assign y14989 = ~n28968 ;
  assign y14990 = 1'b0 ;
  assign y14991 = ~n28969 ;
  assign y14992 = ~1'b0 ;
  assign y14993 = ~1'b0 ;
  assign y14994 = n28972 ;
  assign y14995 = n28973 ;
  assign y14996 = n28978 ;
  assign y14997 = ~1'b0 ;
  assign y14998 = n28981 ;
  assign y14999 = ~1'b0 ;
  assign y15000 = ~n28984 ;
  assign y15001 = ~n28993 ;
  assign y15002 = ~n28995 ;
  assign y15003 = ~1'b0 ;
  assign y15004 = n28996 ;
  assign y15005 = n28997 ;
  assign y15006 = ~n29002 ;
  assign y15007 = n29005 ;
  assign y15008 = ~n29015 ;
  assign y15009 = ~n29018 ;
  assign y15010 = ~n29020 ;
  assign y15011 = n29021 ;
  assign y15012 = ~1'b0 ;
  assign y15013 = ~1'b0 ;
  assign y15014 = ~1'b0 ;
  assign y15015 = ~n29023 ;
  assign y15016 = 1'b0 ;
  assign y15017 = n29027 ;
  assign y15018 = ~1'b0 ;
  assign y15019 = ~n29029 ;
  assign y15020 = ~n29030 ;
  assign y15021 = n29034 ;
  assign y15022 = ~n29035 ;
  assign y15023 = ~1'b0 ;
  assign y15024 = n29036 ;
  assign y15025 = ~n29041 ;
  assign y15026 = ~n29044 ;
  assign y15027 = ~n29047 ;
  assign y15028 = ~1'b0 ;
  assign y15029 = ~1'b0 ;
  assign y15030 = n29051 ;
  assign y15031 = n29052 ;
  assign y15032 = ~n29057 ;
  assign y15033 = ~n29062 ;
  assign y15034 = ~n29064 ;
  assign y15035 = ~1'b0 ;
  assign y15036 = n29066 ;
  assign y15037 = n29069 ;
  assign y15038 = ~n29072 ;
  assign y15039 = n11699 ;
  assign y15040 = n29073 ;
  assign y15041 = n29074 ;
  assign y15042 = ~n29076 ;
  assign y15043 = ~1'b0 ;
  assign y15044 = ~1'b0 ;
  assign y15045 = ~1'b0 ;
  assign y15046 = ~1'b0 ;
  assign y15047 = ~n29078 ;
  assign y15048 = ~1'b0 ;
  assign y15049 = ~n29080 ;
  assign y15050 = ~n29085 ;
  assign y15051 = ~1'b0 ;
  assign y15052 = ~n29086 ;
  assign y15053 = ~1'b0 ;
  assign y15054 = ~1'b0 ;
  assign y15055 = n29093 ;
  assign y15056 = ~n29095 ;
  assign y15057 = n29101 ;
  assign y15058 = n29102 ;
  assign y15059 = ~1'b0 ;
  assign y15060 = ~1'b0 ;
  assign y15061 = n29104 ;
  assign y15062 = n29105 ;
  assign y15063 = n29107 ;
  assign y15064 = n29108 ;
  assign y15065 = n29109 ;
  assign y15066 = ~1'b0 ;
  assign y15067 = ~1'b0 ;
  assign y15068 = n29112 ;
  assign y15069 = n29114 ;
  assign y15070 = ~1'b0 ;
  assign y15071 = n29116 ;
  assign y15072 = 1'b0 ;
  assign y15073 = ~1'b0 ;
  assign y15074 = ~1'b0 ;
  assign y15075 = ~1'b0 ;
  assign y15076 = ~1'b0 ;
  assign y15077 = ~1'b0 ;
  assign y15078 = n29117 ;
  assign y15079 = ~1'b0 ;
  assign y15080 = ~1'b0 ;
  assign y15081 = ~1'b0 ;
  assign y15082 = ~1'b0 ;
  assign y15083 = n29118 ;
  assign y15084 = ~n29121 ;
  assign y15085 = ~1'b0 ;
  assign y15086 = ~1'b0 ;
  assign y15087 = n16495 ;
  assign y15088 = ~n29123 ;
  assign y15089 = ~n29125 ;
  assign y15090 = ~n29127 ;
  assign y15091 = ~1'b0 ;
  assign y15092 = ~n29132 ;
  assign y15093 = n29133 ;
  assign y15094 = ~n29136 ;
  assign y15095 = ~n29138 ;
  assign y15096 = ~n29140 ;
  assign y15097 = n29142 ;
  assign y15098 = ~n29144 ;
  assign y15099 = ~1'b0 ;
  assign y15100 = ~1'b0 ;
  assign y15101 = ~n29152 ;
  assign y15102 = n29155 ;
  assign y15103 = ~1'b0 ;
  assign y15104 = n29156 ;
  assign y15105 = ~n29157 ;
  assign y15106 = ~n29158 ;
  assign y15107 = n29161 ;
  assign y15108 = ~n29165 ;
  assign y15109 = n29166 ;
  assign y15110 = n29169 ;
  assign y15111 = ~n29173 ;
  assign y15112 = ~1'b0 ;
  assign y15113 = ~1'b0 ;
  assign y15114 = n29177 ;
  assign y15115 = ~n29178 ;
  assign y15116 = n29182 ;
  assign y15117 = ~n29184 ;
  assign y15118 = n29185 ;
  assign y15119 = n29187 ;
  assign y15120 = ~1'b0 ;
  assign y15121 = ~n29191 ;
  assign y15122 = ~1'b0 ;
  assign y15123 = n29194 ;
  assign y15124 = ~n29195 ;
  assign y15125 = ~1'b0 ;
  assign y15126 = n29197 ;
  assign y15127 = ~n29198 ;
  assign y15128 = ~n29204 ;
  assign y15129 = n29207 ;
  assign y15130 = n29211 ;
  assign y15131 = n20067 ;
  assign y15132 = ~1'b0 ;
  assign y15133 = n29213 ;
  assign y15134 = ~n6402 ;
  assign y15135 = n29214 ;
  assign y15136 = ~n29217 ;
  assign y15137 = ~1'b0 ;
  assign y15138 = ~n29223 ;
  assign y15139 = ~1'b0 ;
  assign y15140 = n2133 ;
  assign y15141 = n29225 ;
  assign y15142 = ~n29226 ;
  assign y15143 = ~n29230 ;
  assign y15144 = ~1'b0 ;
  assign y15145 = n29232 ;
  assign y15146 = n29235 ;
  assign y15147 = ~1'b0 ;
  assign y15148 = ~1'b0 ;
  assign y15149 = n29246 ;
  assign y15150 = ~n29247 ;
  assign y15151 = ~n29248 ;
  assign y15152 = ~n29251 ;
  assign y15153 = ~1'b0 ;
  assign y15154 = ~n29254 ;
  assign y15155 = n29255 ;
  assign y15156 = n29259 ;
  assign y15157 = n3435 ;
  assign y15158 = ~n7449 ;
  assign y15159 = n17441 ;
  assign y15160 = n29262 ;
  assign y15161 = ~n29263 ;
  assign y15162 = n29266 ;
  assign y15163 = ~n29271 ;
  assign y15164 = n29274 ;
  assign y15165 = ~1'b0 ;
  assign y15166 = n29276 ;
  assign y15167 = n29277 ;
  assign y15168 = ~1'b0 ;
  assign y15169 = ~1'b0 ;
  assign y15170 = n29280 ;
  assign y15171 = ~n10615 ;
  assign y15172 = 1'b0 ;
  assign y15173 = ~1'b0 ;
  assign y15174 = ~n29283 ;
  assign y15175 = n29286 ;
  assign y15176 = 1'b0 ;
  assign y15177 = ~1'b0 ;
  assign y15178 = ~n29288 ;
  assign y15179 = ~n29292 ;
  assign y15180 = n29294 ;
  assign y15181 = ~n23936 ;
  assign y15182 = ~n29297 ;
  assign y15183 = n29298 ;
  assign y15184 = ~1'b0 ;
  assign y15185 = ~n29301 ;
  assign y15186 = ~n29302 ;
  assign y15187 = ~n1891 ;
  assign y15188 = n29304 ;
  assign y15189 = n29305 ;
  assign y15190 = n29306 ;
  assign y15191 = ~1'b0 ;
  assign y15192 = ~1'b0 ;
  assign y15193 = n29307 ;
  assign y15194 = n29308 ;
  assign y15195 = n29310 ;
  assign y15196 = n29312 ;
  assign y15197 = n29320 ;
  assign y15198 = ~1'b0 ;
  assign y15199 = ~n29322 ;
  assign y15200 = n29325 ;
  assign y15201 = n29328 ;
  assign y15202 = n29329 ;
  assign y15203 = ~n29330 ;
  assign y15204 = ~n29333 ;
  assign y15205 = n29335 ;
  assign y15206 = ~1'b0 ;
  assign y15207 = ~n29336 ;
  assign y15208 = n29337 ;
  assign y15209 = n29338 ;
  assign y15210 = ~n29339 ;
  assign y15211 = 1'b0 ;
  assign y15212 = n29343 ;
  assign y15213 = n29345 ;
  assign y15214 = ~n29347 ;
  assign y15215 = n29348 ;
  assign y15216 = ~1'b0 ;
  assign y15217 = ~n29350 ;
  assign y15218 = n13960 ;
  assign y15219 = ~1'b0 ;
  assign y15220 = n29351 ;
  assign y15221 = ~1'b0 ;
  assign y15222 = n29353 ;
  assign y15223 = n29355 ;
  assign y15224 = ~n29356 ;
  assign y15225 = n29358 ;
  assign y15226 = n29360 ;
  assign y15227 = n13731 ;
  assign y15228 = ~n19824 ;
  assign y15229 = ~1'b0 ;
  assign y15230 = ~1'b0 ;
  assign y15231 = ~n29361 ;
  assign y15232 = n29376 ;
  assign y15233 = n29378 ;
  assign y15234 = ~n29379 ;
  assign y15235 = ~n29382 ;
  assign y15236 = ~1'b0 ;
  assign y15237 = ~n29387 ;
  assign y15238 = ~n6200 ;
  assign y15239 = ~1'b0 ;
  assign y15240 = ~n29389 ;
  assign y15241 = ~1'b0 ;
  assign y15242 = n29390 ;
  assign y15243 = n29391 ;
  assign y15244 = ~n20249 ;
  assign y15245 = ~1'b0 ;
  assign y15246 = ~1'b0 ;
  assign y15247 = n29394 ;
  assign y15248 = ~n29398 ;
  assign y15249 = n29401 ;
  assign y15250 = ~1'b0 ;
  assign y15251 = n29402 ;
  assign y15252 = n29405 ;
  assign y15253 = ~n29410 ;
  assign y15254 = n29411 ;
  assign y15255 = ~n29415 ;
  assign y15256 = n29418 ;
  assign y15257 = ~n29421 ;
  assign y15258 = ~n29422 ;
  assign y15259 = ~1'b0 ;
  assign y15260 = ~1'b0 ;
  assign y15261 = ~n29425 ;
  assign y15262 = n21107 ;
  assign y15263 = ~1'b0 ;
  assign y15264 = 1'b0 ;
  assign y15265 = n29426 ;
  assign y15266 = n29427 ;
  assign y15267 = ~n29438 ;
  assign y15268 = ~n29440 ;
  assign y15269 = ~n29442 ;
  assign y15270 = ~1'b0 ;
  assign y15271 = n29443 ;
  assign y15272 = ~1'b0 ;
  assign y15273 = ~1'b0 ;
  assign y15274 = ~n29446 ;
  assign y15275 = 1'b0 ;
  assign y15276 = n29449 ;
  assign y15277 = n28201 ;
  assign y15278 = n29452 ;
  assign y15279 = ~1'b0 ;
  assign y15280 = ~n29456 ;
  assign y15281 = ~n29457 ;
  assign y15282 = ~1'b0 ;
  assign y15283 = ~n29459 ;
  assign y15284 = n29461 ;
  assign y15285 = n29462 ;
  assign y15286 = ~1'b0 ;
  assign y15287 = ~1'b0 ;
  assign y15288 = ~n29463 ;
  assign y15289 = ~n29465 ;
  assign y15290 = ~n29467 ;
  assign y15291 = ~n29469 ;
  assign y15292 = ~n29476 ;
  assign y15293 = n29477 ;
  assign y15294 = ~n29481 ;
  assign y15295 = n29483 ;
  assign y15296 = ~n29485 ;
  assign y15297 = ~1'b0 ;
  assign y15298 = ~n29487 ;
  assign y15299 = ~1'b0 ;
  assign y15300 = n29489 ;
  assign y15301 = ~1'b0 ;
  assign y15302 = ~n29492 ;
  assign y15303 = ~n29496 ;
  assign y15304 = ~n29498 ;
  assign y15305 = ~n6970 ;
  assign y15306 = ~1'b0 ;
  assign y15307 = n29504 ;
  assign y15308 = n29507 ;
  assign y15309 = ~1'b0 ;
  assign y15310 = ~1'b0 ;
  assign y15311 = ~n29512 ;
  assign y15312 = ~1'b0 ;
  assign y15313 = n29513 ;
  assign y15314 = n13888 ;
  assign y15315 = n29515 ;
  assign y15316 = n29516 ;
  assign y15317 = ~1'b0 ;
  assign y15318 = ~n19364 ;
  assign y15319 = n29518 ;
  assign y15320 = ~1'b0 ;
  assign y15321 = ~n17911 ;
  assign y15322 = ~1'b0 ;
  assign y15323 = ~1'b0 ;
  assign y15324 = n29520 ;
  assign y15325 = n29522 ;
  assign y15326 = n26685 ;
  assign y15327 = ~1'b0 ;
  assign y15328 = ~1'b0 ;
  assign y15329 = n29524 ;
  assign y15330 = n29525 ;
  assign y15331 = n29527 ;
  assign y15332 = ~n29530 ;
  assign y15333 = n29531 ;
  assign y15334 = ~n15895 ;
  assign y15335 = ~1'b0 ;
  assign y15336 = ~1'b0 ;
  assign y15337 = n29533 ;
  assign y15338 = n29537 ;
  assign y15339 = ~1'b0 ;
  assign y15340 = n29540 ;
  assign y15341 = ~n29544 ;
  assign y15342 = ~1'b0 ;
  assign y15343 = ~n29545 ;
  assign y15344 = n29547 ;
  assign y15345 = ~1'b0 ;
  assign y15346 = ~1'b0 ;
  assign y15347 = n29548 ;
  assign y15348 = n29549 ;
  assign y15349 = ~n29553 ;
  assign y15350 = ~n29555 ;
  assign y15351 = ~1'b0 ;
  assign y15352 = ~n29557 ;
  assign y15353 = ~1'b0 ;
  assign y15354 = n29560 ;
  assign y15355 = ~n29561 ;
  assign y15356 = ~1'b0 ;
  assign y15357 = ~1'b0 ;
  assign y15358 = ~n29570 ;
  assign y15359 = ~n29576 ;
  assign y15360 = ~n29582 ;
  assign y15361 = ~1'b0 ;
  assign y15362 = ~n29584 ;
  assign y15363 = n29586 ;
  assign y15364 = n29591 ;
  assign y15365 = ~n24131 ;
  assign y15366 = ~1'b0 ;
  assign y15367 = n29592 ;
  assign y15368 = ~n29596 ;
  assign y15369 = ~n29598 ;
  assign y15370 = ~n29600 ;
  assign y15371 = ~n29607 ;
  assign y15372 = n29609 ;
  assign y15373 = n29610 ;
  assign y15374 = ~1'b0 ;
  assign y15375 = ~n29611 ;
  assign y15376 = ~n29612 ;
  assign y15377 = ~1'b0 ;
  assign y15378 = n29615 ;
  assign y15379 = ~1'b0 ;
  assign y15380 = ~n29618 ;
  assign y15381 = n29619 ;
  assign y15382 = ~n29620 ;
  assign y15383 = n10055 ;
  assign y15384 = ~n29626 ;
  assign y15385 = 1'b0 ;
  assign y15386 = n29629 ;
  assign y15387 = ~1'b0 ;
  assign y15388 = ~1'b0 ;
  assign y15389 = n7053 ;
  assign y15390 = n29630 ;
  assign y15391 = ~1'b0 ;
  assign y15392 = ~1'b0 ;
  assign y15393 = n12669 ;
  assign y15394 = ~1'b0 ;
  assign y15395 = ~n29633 ;
  assign y15396 = ~1'b0 ;
  assign y15397 = ~1'b0 ;
  assign y15398 = ~1'b0 ;
  assign y15399 = ~n29639 ;
  assign y15400 = ~1'b0 ;
  assign y15401 = ~n29641 ;
  assign y15402 = n20004 ;
  assign y15403 = ~n29642 ;
  assign y15404 = ~1'b0 ;
  assign y15405 = n29643 ;
  assign y15406 = ~1'b0 ;
  assign y15407 = ~n29645 ;
  assign y15408 = n29646 ;
  assign y15409 = n29648 ;
  assign y15410 = n29650 ;
  assign y15411 = ~n29653 ;
  assign y15412 = ~n29655 ;
  assign y15413 = ~n29657 ;
  assign y15414 = ~1'b0 ;
  assign y15415 = n23862 ;
  assign y15416 = n29658 ;
  assign y15417 = ~n29662 ;
  assign y15418 = ~n29663 ;
  assign y15419 = ~1'b0 ;
  assign y15420 = ~n29664 ;
  assign y15421 = ~1'b0 ;
  assign y15422 = n29665 ;
  assign y15423 = ~1'b0 ;
  assign y15424 = n29666 ;
  assign y15425 = n29668 ;
  assign y15426 = ~n29670 ;
  assign y15427 = 1'b0 ;
  assign y15428 = ~1'b0 ;
  assign y15429 = ~1'b0 ;
  assign y15430 = ~1'b0 ;
  assign y15431 = ~n29671 ;
  assign y15432 = ~n29678 ;
  assign y15433 = n29680 ;
  assign y15434 = ~n29681 ;
  assign y15435 = ~1'b0 ;
  assign y15436 = ~n29682 ;
  assign y15437 = n29684 ;
  assign y15438 = ~1'b0 ;
  assign y15439 = ~1'b0 ;
  assign y15440 = ~n29690 ;
  assign y15441 = ~n29691 ;
  assign y15442 = n29692 ;
  assign y15443 = ~n29694 ;
  assign y15444 = ~n29698 ;
  assign y15445 = ~1'b0 ;
  assign y15446 = ~n29700 ;
  assign y15447 = n14752 ;
  assign y15448 = n29702 ;
  assign y15449 = n29703 ;
  assign y15450 = ~1'b0 ;
  assign y15451 = ~1'b0 ;
  assign y15452 = ~1'b0 ;
  assign y15453 = ~n29704 ;
  assign y15454 = ~n29705 ;
  assign y15455 = ~n29707 ;
  assign y15456 = ~1'b0 ;
  assign y15457 = ~1'b0 ;
  assign y15458 = ~n29708 ;
  assign y15459 = ~n29710 ;
  assign y15460 = ~1'b0 ;
  assign y15461 = n3783 ;
  assign y15462 = n29711 ;
  assign y15463 = ~n29713 ;
  assign y15464 = n26892 ;
  assign y15465 = ~n17377 ;
  assign y15466 = ~n29717 ;
  assign y15467 = ~1'b0 ;
  assign y15468 = ~1'b0 ;
  assign y15469 = ~1'b0 ;
  assign y15470 = n29718 ;
  assign y15471 = n29720 ;
  assign y15472 = n29722 ;
  assign y15473 = n29723 ;
  assign y15474 = ~n29724 ;
  assign y15475 = ~1'b0 ;
  assign y15476 = ~1'b0 ;
  assign y15477 = ~1'b0 ;
  assign y15478 = ~n29725 ;
  assign y15479 = ~n29730 ;
  assign y15480 = ~n29736 ;
  assign y15481 = n29738 ;
  assign y15482 = ~n29740 ;
  assign y15483 = n29741 ;
  assign y15484 = ~n29742 ;
  assign y15485 = ~1'b0 ;
  assign y15486 = ~n29743 ;
  assign y15487 = ~1'b0 ;
  assign y15488 = n29744 ;
  assign y15489 = ~1'b0 ;
  assign y15490 = n29747 ;
  assign y15491 = ~n29748 ;
  assign y15492 = n29762 ;
  assign y15493 = ~1'b0 ;
  assign y15494 = ~n29763 ;
  assign y15495 = n29765 ;
  assign y15496 = ~1'b0 ;
  assign y15497 = ~n10144 ;
  assign y15498 = n29772 ;
  assign y15499 = ~n29776 ;
  assign y15500 = ~n29777 ;
  assign y15501 = ~1'b0 ;
  assign y15502 = 1'b0 ;
  assign y15503 = ~n29778 ;
  assign y15504 = n29779 ;
  assign y15505 = n29785 ;
  assign y15506 = ~n19124 ;
  assign y15507 = ~1'b0 ;
  assign y15508 = ~n29787 ;
  assign y15509 = ~n29790 ;
  assign y15510 = 1'b0 ;
  assign y15511 = ~n29794 ;
  assign y15512 = ~1'b0 ;
  assign y15513 = ~1'b0 ;
  assign y15514 = ~1'b0 ;
  assign y15515 = ~1'b0 ;
  assign y15516 = n29796 ;
  assign y15517 = ~1'b0 ;
  assign y15518 = ~n29797 ;
  assign y15519 = n29800 ;
  assign y15520 = ~n29802 ;
  assign y15521 = n29804 ;
  assign y15522 = ~n29806 ;
  assign y15523 = n29808 ;
  assign y15524 = ~1'b0 ;
  assign y15525 = ~n29809 ;
  assign y15526 = n29812 ;
  assign y15527 = ~n29813 ;
  assign y15528 = ~n29814 ;
  assign y15529 = ~n29815 ;
  assign y15530 = n29816 ;
  assign y15531 = ~1'b0 ;
  assign y15532 = ~n29819 ;
  assign y15533 = ~1'b0 ;
  assign y15534 = ~1'b0 ;
  assign y15535 = n29821 ;
  assign y15536 = n29827 ;
  assign y15537 = ~1'b0 ;
  assign y15538 = ~n29830 ;
  assign y15539 = n29831 ;
  assign y15540 = ~1'b0 ;
  assign y15541 = ~1'b0 ;
  assign y15542 = ~1'b0 ;
  assign y15543 = ~n29833 ;
  assign y15544 = n13312 ;
  assign y15545 = n29835 ;
  assign y15546 = ~n29841 ;
  assign y15547 = n29842 ;
  assign y15548 = n29843 ;
  assign y15549 = ~1'b0 ;
  assign y15550 = n29847 ;
  assign y15551 = ~n14831 ;
  assign y15552 = ~n29848 ;
  assign y15553 = n29852 ;
  assign y15554 = ~1'b0 ;
  assign y15555 = ~n25051 ;
  assign y15556 = ~n29855 ;
  assign y15557 = ~n4251 ;
  assign y15558 = ~1'b0 ;
  assign y15559 = ~n29860 ;
  assign y15560 = ~n29861 ;
  assign y15561 = ~n29862 ;
  assign y15562 = n29863 ;
  assign y15563 = n29866 ;
  assign y15564 = ~1'b0 ;
  assign y15565 = ~1'b0 ;
  assign y15566 = n29868 ;
  assign y15567 = ~n29870 ;
  assign y15568 = ~n29872 ;
  assign y15569 = ~n29873 ;
  assign y15570 = ~n7706 ;
  assign y15571 = ~1'b0 ;
  assign y15572 = ~n16028 ;
  assign y15573 = n29875 ;
  assign y15574 = n29876 ;
  assign y15575 = ~1'b0 ;
  assign y15576 = n29877 ;
  assign y15577 = n29883 ;
  assign y15578 = ~1'b0 ;
  assign y15579 = n29885 ;
  assign y15580 = n29888 ;
  assign y15581 = ~1'b0 ;
  assign y15582 = ~1'b0 ;
  assign y15583 = ~n29889 ;
  assign y15584 = n6671 ;
  assign y15585 = ~n29890 ;
  assign y15586 = ~n29893 ;
  assign y15587 = ~n29894 ;
  assign y15588 = ~1'b0 ;
  assign y15589 = ~n29897 ;
  assign y15590 = ~1'b0 ;
  assign y15591 = n29900 ;
  assign y15592 = ~n29905 ;
  assign y15593 = 1'b0 ;
  assign y15594 = ~n29908 ;
  assign y15595 = n29909 ;
  assign y15596 = ~n3671 ;
  assign y15597 = n29913 ;
  assign y15598 = ~n29914 ;
  assign y15599 = n29921 ;
  assign y15600 = ~n29923 ;
  assign y15601 = 1'b0 ;
  assign y15602 = n29925 ;
  assign y15603 = 1'b0 ;
  assign y15604 = ~n29927 ;
  assign y15605 = n11517 ;
  assign y15606 = ~n29929 ;
  assign y15607 = ~1'b0 ;
  assign y15608 = ~n29933 ;
  assign y15609 = n29936 ;
  assign y15610 = n29937 ;
  assign y15611 = ~n29941 ;
  assign y15612 = n29943 ;
  assign y15613 = ~1'b0 ;
  assign y15614 = n29947 ;
  assign y15615 = n29950 ;
  assign y15616 = ~n29952 ;
  assign y15617 = ~n29953 ;
  assign y15618 = n29955 ;
  assign y15619 = n29960 ;
  assign y15620 = ~n29962 ;
  assign y15621 = n29965 ;
  assign y15622 = ~1'b0 ;
  assign y15623 = ~n29970 ;
  assign y15624 = n29978 ;
  assign y15625 = ~n29981 ;
  assign y15626 = n29982 ;
  assign y15627 = ~1'b0 ;
  assign y15628 = n29984 ;
  assign y15629 = ~1'b0 ;
  assign y15630 = ~n29986 ;
  assign y15631 = n5396 ;
  assign y15632 = ~n29992 ;
  assign y15633 = n29994 ;
  assign y15634 = ~n15437 ;
  assign y15635 = ~n29997 ;
  assign y15636 = ~n29999 ;
  assign y15637 = ~1'b0 ;
  assign y15638 = n30000 ;
  assign y15639 = ~1'b0 ;
  assign y15640 = 1'b0 ;
  assign y15641 = n30005 ;
  assign y15642 = ~n30006 ;
  assign y15643 = ~1'b0 ;
  assign y15644 = n30007 ;
  assign y15645 = ~1'b0 ;
  assign y15646 = ~1'b0 ;
  assign y15647 = ~n30011 ;
  assign y15648 = ~1'b0 ;
  assign y15649 = ~1'b0 ;
  assign y15650 = ~n21276 ;
  assign y15651 = n30013 ;
  assign y15652 = ~1'b0 ;
  assign y15653 = ~n21027 ;
  assign y15654 = ~n30016 ;
  assign y15655 = ~n30019 ;
  assign y15656 = ~1'b0 ;
  assign y15657 = n30020 ;
  assign y15658 = ~n30022 ;
  assign y15659 = ~n30023 ;
  assign y15660 = ~1'b0 ;
  assign y15661 = n30024 ;
  assign y15662 = ~n30026 ;
  assign y15663 = ~n30030 ;
  assign y15664 = ~n30032 ;
  assign y15665 = ~n30034 ;
  assign y15666 = n30036 ;
  assign y15667 = ~n30037 ;
  assign y15668 = ~n30038 ;
  assign y15669 = n20291 ;
  assign y15670 = ~n30041 ;
  assign y15671 = n30045 ;
  assign y15672 = ~n30046 ;
  assign y15673 = n30047 ;
  assign y15674 = n30050 ;
  assign y15675 = n30054 ;
  assign y15676 = ~1'b0 ;
  assign y15677 = 1'b0 ;
  assign y15678 = ~n30058 ;
  assign y15679 = ~n30062 ;
  assign y15680 = ~n30063 ;
  assign y15681 = ~n30066 ;
  assign y15682 = ~1'b0 ;
  assign y15683 = ~1'b0 ;
  assign y15684 = ~n30067 ;
  assign y15685 = ~n30077 ;
  assign y15686 = n30079 ;
  assign y15687 = n30082 ;
  assign y15688 = ~n30083 ;
  assign y15689 = n30086 ;
  assign y15690 = ~1'b0 ;
  assign y15691 = ~n30088 ;
  assign y15692 = n30090 ;
  assign y15693 = ~n30092 ;
  assign y15694 = n30095 ;
  assign y15695 = n8978 ;
  assign y15696 = n27363 ;
  assign y15697 = ~n30096 ;
  assign y15698 = ~n30097 ;
  assign y15699 = ~n30100 ;
  assign y15700 = ~n30105 ;
  assign y15701 = ~1'b0 ;
  assign y15702 = ~1'b0 ;
  assign y15703 = ~n30106 ;
  assign y15704 = ~n30109 ;
  assign y15705 = ~n30110 ;
  assign y15706 = ~1'b0 ;
  assign y15707 = ~n8690 ;
  assign y15708 = ~1'b0 ;
  assign y15709 = ~n30113 ;
  assign y15710 = ~1'b0 ;
  assign y15711 = n30114 ;
  assign y15712 = ~n30117 ;
  assign y15713 = n30119 ;
  assign y15714 = ~n8404 ;
  assign y15715 = ~1'b0 ;
  assign y15716 = ~1'b0 ;
  assign y15717 = ~n30125 ;
  assign y15718 = n30127 ;
  assign y15719 = n30128 ;
  assign y15720 = n30129 ;
  assign y15721 = n30130 ;
  assign y15722 = ~n30132 ;
  assign y15723 = ~n30134 ;
  assign y15724 = n30138 ;
  assign y15725 = ~n30140 ;
  assign y15726 = n30142 ;
  assign y15727 = ~n30145 ;
  assign y15728 = ~n30148 ;
  assign y15729 = ~n30149 ;
  assign y15730 = ~1'b0 ;
  assign y15731 = 1'b0 ;
  assign y15732 = n30150 ;
  assign y15733 = ~1'b0 ;
  assign y15734 = ~n30153 ;
  assign y15735 = ~n30155 ;
  assign y15736 = n30158 ;
  assign y15737 = n30160 ;
  assign y15738 = ~n30161 ;
  assign y15739 = ~n30163 ;
  assign y15740 = ~1'b0 ;
  assign y15741 = ~1'b0 ;
  assign y15742 = n30165 ;
  assign y15743 = ~n30168 ;
  assign y15744 = ~n30169 ;
  assign y15745 = ~1'b0 ;
  assign y15746 = n30172 ;
  assign y15747 = ~n30176 ;
  assign y15748 = ~1'b0 ;
  assign y15749 = n30180 ;
  assign y15750 = ~1'b0 ;
  assign y15751 = ~n30181 ;
  assign y15752 = ~n30182 ;
  assign y15753 = n30185 ;
  assign y15754 = ~n30186 ;
  assign y15755 = n30189 ;
  assign y15756 = n30194 ;
  assign y15757 = ~n9048 ;
  assign y15758 = ~n30195 ;
  assign y15759 = ~1'b0 ;
  assign y15760 = n30196 ;
  assign y15761 = n501 ;
  assign y15762 = ~1'b0 ;
  assign y15763 = ~1'b0 ;
  assign y15764 = ~1'b0 ;
  assign y15765 = ~n30197 ;
  assign y15766 = ~1'b0 ;
  assign y15767 = ~n30198 ;
  assign y15768 = ~n30199 ;
  assign y15769 = n30204 ;
  assign y15770 = n30209 ;
  assign y15771 = ~1'b0 ;
  assign y15772 = n30210 ;
  assign y15773 = ~n30211 ;
  assign y15774 = ~n30213 ;
  assign y15775 = ~1'b0 ;
  assign y15776 = ~n30215 ;
  assign y15777 = n30218 ;
  assign y15778 = ~n30220 ;
  assign y15779 = n30224 ;
  assign y15780 = n30232 ;
  assign y15781 = ~n30235 ;
  assign y15782 = n21100 ;
  assign y15783 = ~1'b0 ;
  assign y15784 = n14192 ;
  assign y15785 = ~n30237 ;
  assign y15786 = ~1'b0 ;
  assign y15787 = n30239 ;
  assign y15788 = n30240 ;
  assign y15789 = ~n30241 ;
  assign y15790 = n12216 ;
  assign y15791 = n30242 ;
  assign y15792 = ~1'b0 ;
  assign y15793 = n30246 ;
  assign y15794 = ~n30250 ;
  assign y15795 = ~n30253 ;
  assign y15796 = ~1'b0 ;
  assign y15797 = ~n30254 ;
  assign y15798 = ~n30258 ;
  assign y15799 = n30260 ;
  assign y15800 = ~n30263 ;
  assign y15801 = n575 ;
  assign y15802 = ~n30270 ;
  assign y15803 = ~n30273 ;
  assign y15804 = n30276 ;
  assign y15805 = n30277 ;
  assign y15806 = ~n30279 ;
  assign y15807 = n24933 ;
  assign y15808 = n30280 ;
  assign y15809 = ~n30281 ;
  assign y15810 = ~n30283 ;
  assign y15811 = ~n30288 ;
  assign y15812 = n30289 ;
  assign y15813 = n30290 ;
  assign y15814 = n30291 ;
  assign y15815 = n27645 ;
  assign y15816 = ~n30292 ;
  assign y15817 = ~1'b0 ;
  assign y15818 = n30294 ;
  assign y15819 = n30298 ;
  assign y15820 = n30305 ;
  assign y15821 = n30309 ;
  assign y15822 = ~n30310 ;
  assign y15823 = ~n30311 ;
  assign y15824 = ~n30314 ;
  assign y15825 = n30327 ;
  assign y15826 = ~n30333 ;
  assign y15827 = ~n30334 ;
  assign y15828 = ~n30337 ;
  assign y15829 = n30338 ;
  assign y15830 = ~n30341 ;
  assign y15831 = ~1'b0 ;
  assign y15832 = n30342 ;
  assign y15833 = n30351 ;
  assign y15834 = ~n30352 ;
  assign y15835 = ~n30358 ;
  assign y15836 = n30366 ;
  assign y15837 = n30369 ;
  assign y15838 = n30374 ;
  assign y15839 = n30377 ;
  assign y15840 = n30381 ;
  assign y15841 = n30383 ;
  assign y15842 = n30386 ;
  assign y15843 = ~n30388 ;
  assign y15844 = ~n30390 ;
  assign y15845 = ~1'b0 ;
  assign y15846 = ~n30392 ;
  assign y15847 = ~n30393 ;
  assign y15848 = ~n30394 ;
  assign y15849 = n30395 ;
  assign y15850 = n30401 ;
  assign y15851 = ~n30406 ;
  assign y15852 = n30408 ;
  assign y15853 = ~1'b0 ;
  assign y15854 = ~1'b0 ;
  assign y15855 = n30416 ;
  assign y15856 = ~n30417 ;
  assign y15857 = n30419 ;
  assign y15858 = n30422 ;
  assign y15859 = ~1'b0 ;
  assign y15860 = ~1'b0 ;
  assign y15861 = ~1'b0 ;
  assign y15862 = ~n30427 ;
  assign y15863 = 1'b0 ;
  assign y15864 = ~1'b0 ;
  assign y15865 = ~n30430 ;
  assign y15866 = ~n30432 ;
  assign y15867 = n30437 ;
  assign y15868 = ~1'b0 ;
  assign y15869 = ~1'b0 ;
  assign y15870 = n30438 ;
  assign y15871 = n30439 ;
  assign y15872 = n15881 ;
  assign y15873 = n30442 ;
  assign y15874 = n30446 ;
  assign y15875 = ~n30449 ;
  assign y15876 = ~n30450 ;
  assign y15877 = n30452 ;
  assign y15878 = 1'b0 ;
  assign y15879 = n30453 ;
  assign y15880 = ~n30457 ;
  assign y15881 = ~n30462 ;
  assign y15882 = n30463 ;
  assign y15883 = n30466 ;
  assign y15884 = ~n30468 ;
  assign y15885 = n30470 ;
  assign y15886 = ~n30476 ;
  assign y15887 = ~n6272 ;
  assign y15888 = n30480 ;
  assign y15889 = n30491 ;
  assign y15890 = ~n30493 ;
  assign y15891 = n30498 ;
  assign y15892 = ~n1660 ;
  assign y15893 = ~n30499 ;
  assign y15894 = ~n30500 ;
  assign y15895 = ~1'b0 ;
  assign y15896 = ~1'b0 ;
  assign y15897 = n30508 ;
  assign y15898 = ~1'b0 ;
  assign y15899 = n30509 ;
  assign y15900 = ~n30511 ;
  assign y15901 = n30513 ;
  assign y15902 = n30514 ;
  assign y15903 = n30515 ;
  assign y15904 = n30516 ;
  assign y15905 = ~1'b0 ;
  assign y15906 = n30518 ;
  assign y15907 = ~n30521 ;
  assign y15908 = ~n30522 ;
  assign y15909 = 1'b0 ;
  assign y15910 = ~1'b0 ;
  assign y15911 = ~1'b0 ;
  assign y15912 = ~1'b0 ;
  assign y15913 = ~n30524 ;
  assign y15914 = ~n30526 ;
  assign y15915 = ~1'b0 ;
  assign y15916 = ~n30528 ;
  assign y15917 = ~1'b0 ;
  assign y15918 = ~n30529 ;
  assign y15919 = ~1'b0 ;
  assign y15920 = ~1'b0 ;
  assign y15921 = n30532 ;
  assign y15922 = ~n30534 ;
  assign y15923 = n30538 ;
  assign y15924 = n30539 ;
  assign y15925 = ~1'b0 ;
  assign y15926 = ~n30542 ;
  assign y15927 = n30543 ;
  assign y15928 = n30545 ;
  assign y15929 = ~1'b0 ;
  assign y15930 = ~1'b0 ;
  assign y15931 = n30547 ;
  assign y15932 = n30548 ;
  assign y15933 = n30551 ;
  assign y15934 = ~n30552 ;
  assign y15935 = ~n30554 ;
  assign y15936 = n15485 ;
  assign y15937 = n23633 ;
  assign y15938 = n30555 ;
  assign y15939 = ~n10582 ;
  assign y15940 = ~n30557 ;
  assign y15941 = ~1'b0 ;
  assign y15942 = n30559 ;
  assign y15943 = ~n28586 ;
  assign y15944 = n30560 ;
  assign y15945 = ~1'b0 ;
  assign y15946 = ~1'b0 ;
  assign y15947 = ~1'b0 ;
  assign y15948 = ~1'b0 ;
  assign y15949 = ~n30562 ;
  assign y15950 = ~1'b0 ;
  assign y15951 = n5039 ;
  assign y15952 = ~1'b0 ;
  assign y15953 = ~1'b0 ;
  assign y15954 = ~n18946 ;
  assign y15955 = ~n30564 ;
  assign y15956 = ~n30569 ;
  assign y15957 = ~n30573 ;
  assign y15958 = n27797 ;
  assign y15959 = n30575 ;
  assign y15960 = ~n6812 ;
  assign y15961 = ~n30578 ;
  assign y15962 = n30579 ;
  assign y15963 = n30580 ;
  assign y15964 = ~n30585 ;
  assign y15965 = ~n30590 ;
  assign y15966 = n862 ;
  assign y15967 = ~1'b0 ;
  assign y15968 = 1'b0 ;
  assign y15969 = n30595 ;
  assign y15970 = ~n30597 ;
  assign y15971 = ~n30601 ;
  assign y15972 = ~n30602 ;
  assign y15973 = n30603 ;
  assign y15974 = n30607 ;
  assign y15975 = n30608 ;
  assign y15976 = n30610 ;
  assign y15977 = ~n30612 ;
  assign y15978 = ~1'b0 ;
  assign y15979 = n5404 ;
  assign y15980 = ~n30614 ;
  assign y15981 = n30616 ;
  assign y15982 = 1'b0 ;
  assign y15983 = ~1'b0 ;
  assign y15984 = ~n30620 ;
  assign y15985 = n30622 ;
  assign y15986 = ~1'b0 ;
  assign y15987 = ~n30623 ;
  assign y15988 = ~1'b0 ;
  assign y15989 = ~1'b0 ;
  assign y15990 = ~n30625 ;
  assign y15991 = ~n30630 ;
  assign y15992 = 1'b0 ;
  assign y15993 = 1'b0 ;
  assign y15994 = ~1'b0 ;
  assign y15995 = ~n30633 ;
  assign y15996 = ~n30637 ;
  assign y15997 = ~1'b0 ;
  assign y15998 = ~1'b0 ;
  assign y15999 = ~1'b0 ;
  assign y16000 = n30641 ;
  assign y16001 = ~1'b0 ;
  assign y16002 = n9367 ;
  assign y16003 = ~1'b0 ;
  assign y16004 = n30645 ;
  assign y16005 = ~1'b0 ;
  assign y16006 = ~1'b0 ;
  assign y16007 = ~1'b0 ;
  assign y16008 = ~n30646 ;
  assign y16009 = n30650 ;
  assign y16010 = n30652 ;
  assign y16011 = ~n30655 ;
  assign y16012 = ~n30656 ;
  assign y16013 = ~1'b0 ;
  assign y16014 = ~n30658 ;
  assign y16015 = n30664 ;
  assign y16016 = n30666 ;
  assign y16017 = n30667 ;
  assign y16018 = ~n30670 ;
  assign y16019 = ~1'b0 ;
  assign y16020 = ~n30672 ;
  assign y16021 = ~1'b0 ;
  assign y16022 = n30673 ;
  assign y16023 = ~1'b0 ;
  assign y16024 = n30676 ;
  assign y16025 = n30680 ;
  assign y16026 = n30681 ;
  assign y16027 = ~n30694 ;
  assign y16028 = n30699 ;
  assign y16029 = n29745 ;
  assign y16030 = n30701 ;
  assign y16031 = n30704 ;
  assign y16032 = ~n8333 ;
  assign y16033 = ~n30705 ;
  assign y16034 = ~1'b0 ;
  assign y16035 = ~n29011 ;
  assign y16036 = n30706 ;
  assign y16037 = ~n30707 ;
  assign y16038 = ~n3837 ;
  assign y16039 = ~1'b0 ;
  assign y16040 = ~n30708 ;
  assign y16041 = ~1'b0 ;
  assign y16042 = ~1'b0 ;
  assign y16043 = ~1'b0 ;
  assign y16044 = ~n30710 ;
  assign y16045 = ~1'b0 ;
  assign y16046 = n30715 ;
  assign y16047 = ~n30719 ;
  assign y16048 = ~n30720 ;
  assign y16049 = n30727 ;
  assign y16050 = ~n30731 ;
  assign y16051 = ~1'b0 ;
  assign y16052 = ~1'b0 ;
  assign y16053 = ~n30732 ;
  assign y16054 = ~1'b0 ;
  assign y16055 = n30734 ;
  assign y16056 = ~1'b0 ;
  assign y16057 = 1'b0 ;
  assign y16058 = n30736 ;
  assign y16059 = ~1'b0 ;
  assign y16060 = n30737 ;
  assign y16061 = n30738 ;
  assign y16062 = ~n30740 ;
  assign y16063 = n30741 ;
  assign y16064 = ~1'b0 ;
  assign y16065 = ~n30743 ;
  assign y16066 = ~n30744 ;
  assign y16067 = n993 ;
  assign y16068 = ~1'b0 ;
  assign y16069 = ~n30745 ;
  assign y16070 = ~1'b0 ;
  assign y16071 = ~n30746 ;
  assign y16072 = ~n6049 ;
  assign y16073 = ~n30747 ;
  assign y16074 = n30748 ;
  assign y16075 = n30750 ;
  assign y16076 = ~1'b0 ;
  assign y16077 = ~n30753 ;
  assign y16078 = ~n30759 ;
  assign y16079 = ~n30762 ;
  assign y16080 = n30764 ;
  assign y16081 = 1'b0 ;
  assign y16082 = n30767 ;
  assign y16083 = n30770 ;
  assign y16084 = n30771 ;
  assign y16085 = ~n30774 ;
  assign y16086 = n30776 ;
  assign y16087 = ~n30782 ;
  assign y16088 = n30783 ;
  assign y16089 = 1'b0 ;
  assign y16090 = ~1'b0 ;
  assign y16091 = ~n30785 ;
  assign y16092 = ~n30788 ;
  assign y16093 = n30789 ;
  assign y16094 = ~n30793 ;
  assign y16095 = ~1'b0 ;
  assign y16096 = n30795 ;
  assign y16097 = ~n30796 ;
  assign y16098 = ~n16519 ;
  assign y16099 = n30801 ;
  assign y16100 = ~1'b0 ;
  assign y16101 = n30805 ;
  assign y16102 = ~1'b0 ;
  assign y16103 = ~1'b0 ;
  assign y16104 = 1'b0 ;
  assign y16105 = n30807 ;
  assign y16106 = n30809 ;
  assign y16107 = ~n30816 ;
  assign y16108 = ~1'b0 ;
  assign y16109 = ~1'b0 ;
  assign y16110 = ~1'b0 ;
  assign y16111 = ~n30819 ;
  assign y16112 = ~1'b0 ;
  assign y16113 = ~n30820 ;
  assign y16114 = ~n30823 ;
  assign y16115 = ~n9081 ;
  assign y16116 = n30824 ;
  assign y16117 = ~1'b0 ;
  assign y16118 = ~n29377 ;
  assign y16119 = n30825 ;
  assign y16120 = ~1'b0 ;
  assign y16121 = ~n30826 ;
  assign y16122 = n30827 ;
  assign y16123 = ~1'b0 ;
  assign y16124 = ~n30830 ;
  assign y16125 = ~n30835 ;
  assign y16126 = ~1'b0 ;
  assign y16127 = ~1'b0 ;
  assign y16128 = ~1'b0 ;
  assign y16129 = ~1'b0 ;
  assign y16130 = ~1'b0 ;
  assign y16131 = ~n30836 ;
  assign y16132 = ~1'b0 ;
  assign y16133 = n30838 ;
  assign y16134 = n30844 ;
  assign y16135 = ~1'b0 ;
  assign y16136 = ~1'b0 ;
  assign y16137 = n13051 ;
  assign y16138 = ~n30847 ;
  assign y16139 = ~n30848 ;
  assign y16140 = ~n30849 ;
  assign y16141 = ~n1073 ;
  assign y16142 = ~n30850 ;
  assign y16143 = n30857 ;
  assign y16144 = n30859 ;
  assign y16145 = n30861 ;
  assign y16146 = ~n30863 ;
  assign y16147 = ~n30867 ;
  assign y16148 = ~n30869 ;
  assign y16149 = ~1'b0 ;
  assign y16150 = ~1'b0 ;
  assign y16151 = n30875 ;
  assign y16152 = n22144 ;
  assign y16153 = n30876 ;
  assign y16154 = n1553 ;
  assign y16155 = ~n30911 ;
  assign y16156 = ~1'b0 ;
  assign y16157 = ~1'b0 ;
  assign y16158 = n30913 ;
  assign y16159 = n30916 ;
  assign y16160 = n30923 ;
  assign y16161 = n30925 ;
  assign y16162 = ~1'b0 ;
  assign y16163 = ~1'b0 ;
  assign y16164 = ~n7818 ;
  assign y16165 = ~1'b0 ;
  assign y16166 = n30927 ;
  assign y16167 = n15752 ;
  assign y16168 = n11344 ;
  assign y16169 = n30928 ;
  assign y16170 = ~1'b0 ;
  assign y16171 = ~n30931 ;
  assign y16172 = ~1'b0 ;
  assign y16173 = ~n30934 ;
  assign y16174 = ~n30936 ;
  assign y16175 = ~n30937 ;
  assign y16176 = ~n30939 ;
  assign y16177 = n30941 ;
  assign y16178 = ~n30942 ;
  assign y16179 = ~n30944 ;
  assign y16180 = ~n30945 ;
  assign y16181 = n30946 ;
  assign y16182 = n30950 ;
  assign y16183 = ~n30951 ;
  assign y16184 = ~n30952 ;
  assign y16185 = ~1'b0 ;
  assign y16186 = ~1'b0 ;
  assign y16187 = ~n30955 ;
  assign y16188 = ~1'b0 ;
  assign y16189 = ~n30956 ;
  assign y16190 = ~1'b0 ;
  assign y16191 = n30960 ;
  assign y16192 = n30962 ;
  assign y16193 = ~n30963 ;
  assign y16194 = n30966 ;
  assign y16195 = ~1'b0 ;
  assign y16196 = n30968 ;
  assign y16197 = ~1'b0 ;
  assign y16198 = n30969 ;
  assign y16199 = n30973 ;
  assign y16200 = ~n30982 ;
  assign y16201 = n30983 ;
  assign y16202 = n30986 ;
  assign y16203 = n30989 ;
  assign y16204 = ~n30990 ;
  assign y16205 = n30992 ;
  assign y16206 = ~n30995 ;
  assign y16207 = ~1'b0 ;
  assign y16208 = ~1'b0 ;
  assign y16209 = ~1'b0 ;
  assign y16210 = ~1'b0 ;
  assign y16211 = n25499 ;
  assign y16212 = ~n30997 ;
  assign y16213 = ~n31004 ;
  assign y16214 = ~n31005 ;
  assign y16215 = ~n31006 ;
  assign y16216 = n31011 ;
  assign y16217 = ~1'b0 ;
  assign y16218 = ~1'b0 ;
  assign y16219 = ~n31014 ;
  assign y16220 = ~1'b0 ;
  assign y16221 = ~n31017 ;
  assign y16222 = ~n31018 ;
  assign y16223 = ~n31020 ;
  assign y16224 = n31021 ;
  assign y16225 = ~n31022 ;
  assign y16226 = ~1'b0 ;
  assign y16227 = ~1'b0 ;
  assign y16228 = ~1'b0 ;
  assign y16229 = ~n31023 ;
  assign y16230 = n31024 ;
  assign y16231 = ~1'b0 ;
  assign y16232 = n31025 ;
  assign y16233 = ~n31028 ;
  assign y16234 = ~1'b0 ;
  assign y16235 = n31029 ;
  assign y16236 = ~n31030 ;
  assign y16237 = n31033 ;
  assign y16238 = n31035 ;
  assign y16239 = n31038 ;
  assign y16240 = ~1'b0 ;
  assign y16241 = 1'b0 ;
  assign y16242 = n31039 ;
  assign y16243 = ~n31040 ;
  assign y16244 = n31042 ;
  assign y16245 = n3016 ;
  assign y16246 = ~1'b0 ;
  assign y16247 = ~n31045 ;
  assign y16248 = ~n31047 ;
  assign y16249 = n31049 ;
  assign y16250 = ~1'b0 ;
  assign y16251 = ~n31050 ;
  assign y16252 = ~1'b0 ;
  assign y16253 = n31053 ;
  assign y16254 = n31055 ;
  assign y16255 = ~n31058 ;
  assign y16256 = ~n31062 ;
  assign y16257 = n31067 ;
  assign y16258 = n31068 ;
  assign y16259 = ~1'b0 ;
  assign y16260 = ~1'b0 ;
  assign y16261 = ~n31070 ;
  assign y16262 = ~n31072 ;
  assign y16263 = ~1'b0 ;
  assign y16264 = n31073 ;
  assign y16265 = ~1'b0 ;
  assign y16266 = ~1'b0 ;
  assign y16267 = ~n31076 ;
  assign y16268 = ~1'b0 ;
  assign y16269 = n31077 ;
  assign y16270 = ~n31078 ;
  assign y16271 = ~1'b0 ;
  assign y16272 = n31080 ;
  assign y16273 = ~n31081 ;
  assign y16274 = n27201 ;
  assign y16275 = ~n31086 ;
  assign y16276 = n31089 ;
  assign y16277 = n31095 ;
  assign y16278 = n31096 ;
  assign y16279 = ~n31097 ;
  assign y16280 = n31099 ;
  assign y16281 = ~n2002 ;
  assign y16282 = n31101 ;
  assign y16283 = ~n1630 ;
  assign y16284 = ~1'b0 ;
  assign y16285 = n31104 ;
  assign y16286 = ~1'b0 ;
  assign y16287 = n31105 ;
  assign y16288 = ~1'b0 ;
  assign y16289 = ~1'b0 ;
  assign y16290 = ~1'b0 ;
  assign y16291 = ~1'b0 ;
  assign y16292 = 1'b0 ;
  assign y16293 = ~n31113 ;
  assign y16294 = ~1'b0 ;
  assign y16295 = ~n31114 ;
  assign y16296 = ~1'b0 ;
  assign y16297 = ~n31118 ;
  assign y16298 = ~1'b0 ;
  assign y16299 = n1962 ;
  assign y16300 = n31119 ;
  assign y16301 = ~n31121 ;
  assign y16302 = ~1'b0 ;
  assign y16303 = n31122 ;
  assign y16304 = ~1'b0 ;
  assign y16305 = n31123 ;
  assign y16306 = ~1'b0 ;
  assign y16307 = n31126 ;
  assign y16308 = ~n31127 ;
  assign y16309 = n13164 ;
  assign y16310 = n31129 ;
  assign y16311 = ~n31132 ;
  assign y16312 = n31134 ;
  assign y16313 = ~n31140 ;
  assign y16314 = n31142 ;
  assign y16315 = n31144 ;
  assign y16316 = ~n31145 ;
  assign y16317 = n31146 ;
  assign y16318 = 1'b0 ;
  assign y16319 = ~n31148 ;
  assign y16320 = n22721 ;
  assign y16321 = ~1'b0 ;
  assign y16322 = ~1'b0 ;
  assign y16323 = ~n31150 ;
  assign y16324 = ~n30784 ;
  assign y16325 = ~n28544 ;
  assign y16326 = n31151 ;
  assign y16327 = ~n3023 ;
  assign y16328 = ~n31154 ;
  assign y16329 = ~1'b0 ;
  assign y16330 = ~n31158 ;
  assign y16331 = ~1'b0 ;
  assign y16332 = ~n31161 ;
  assign y16333 = ~1'b0 ;
  assign y16334 = n31163 ;
  assign y16335 = 1'b0 ;
  assign y16336 = ~n31165 ;
  assign y16337 = ~1'b0 ;
  assign y16338 = n31168 ;
  assign y16339 = ~n31171 ;
  assign y16340 = n31172 ;
  assign y16341 = n31173 ;
  assign y16342 = n31177 ;
  assign y16343 = n31178 ;
  assign y16344 = ~n31181 ;
  assign y16345 = ~1'b0 ;
  assign y16346 = ~n31184 ;
  assign y16347 = n31185 ;
  assign y16348 = ~n31187 ;
  assign y16349 = ~1'b0 ;
  assign y16350 = n5811 ;
  assign y16351 = n31195 ;
  assign y16352 = ~n31201 ;
  assign y16353 = n31206 ;
  assign y16354 = ~1'b0 ;
  assign y16355 = ~n31209 ;
  assign y16356 = ~n31210 ;
  assign y16357 = ~1'b0 ;
  assign y16358 = n31213 ;
  assign y16359 = ~n31214 ;
  assign y16360 = n31216 ;
  assign y16361 = ~1'b0 ;
  assign y16362 = ~n31220 ;
  assign y16363 = ~1'b0 ;
  assign y16364 = n24519 ;
  assign y16365 = ~1'b0 ;
  assign y16366 = ~n31224 ;
  assign y16367 = ~n31230 ;
  assign y16368 = ~n31232 ;
  assign y16369 = ~1'b0 ;
  assign y16370 = ~n31237 ;
  assign y16371 = ~n31238 ;
  assign y16372 = 1'b0 ;
  assign y16373 = ~1'b0 ;
  assign y16374 = n31239 ;
  assign y16375 = ~1'b0 ;
  assign y16376 = ~1'b0 ;
  assign y16377 = ~1'b0 ;
  assign y16378 = ~n31241 ;
  assign y16379 = ~1'b0 ;
  assign y16380 = ~1'b0 ;
  assign y16381 = ~1'b0 ;
  assign y16382 = ~n31243 ;
  assign y16383 = ~n31244 ;
  assign y16384 = ~1'b0 ;
  assign y16385 = ~1'b0 ;
  assign y16386 = ~1'b0 ;
  assign y16387 = ~n31246 ;
  assign y16388 = n31247 ;
  assign y16389 = ~n31248 ;
  assign y16390 = n31251 ;
  assign y16391 = ~n31256 ;
  assign y16392 = n31257 ;
  assign y16393 = ~n31259 ;
  assign y16394 = 1'b0 ;
  assign y16395 = ~1'b0 ;
  assign y16396 = n31262 ;
  assign y16397 = n31263 ;
  assign y16398 = ~1'b0 ;
  assign y16399 = ~1'b0 ;
  assign y16400 = n31268 ;
  assign y16401 = n31270 ;
  assign y16402 = ~1'b0 ;
  assign y16403 = ~1'b0 ;
  assign y16404 = n31274 ;
  assign y16405 = ~1'b0 ;
  assign y16406 = ~n31276 ;
  assign y16407 = ~n31279 ;
  assign y16408 = ~n31283 ;
  assign y16409 = ~n31287 ;
  assign y16410 = ~n31291 ;
  assign y16411 = ~1'b0 ;
  assign y16412 = ~n31292 ;
  assign y16413 = ~1'b0 ;
  assign y16414 = n31295 ;
  assign y16415 = 1'b0 ;
  assign y16416 = n31297 ;
  assign y16417 = ~1'b0 ;
  assign y16418 = ~1'b0 ;
  assign y16419 = ~1'b0 ;
  assign y16420 = n31299 ;
  assign y16421 = ~n31300 ;
  assign y16422 = ~n31301 ;
  assign y16423 = ~1'b0 ;
  assign y16424 = n31302 ;
  assign y16425 = ~1'b0 ;
  assign y16426 = ~1'b0 ;
  assign y16427 = n31306 ;
  assign y16428 = ~n31307 ;
  assign y16429 = ~n31310 ;
  assign y16430 = n31312 ;
  assign y16431 = ~1'b0 ;
  assign y16432 = ~1'b0 ;
  assign y16433 = n31316 ;
  assign y16434 = ~n31318 ;
  assign y16435 = n31323 ;
  assign y16436 = n31326 ;
  assign y16437 = ~1'b0 ;
  assign y16438 = n31329 ;
  assign y16439 = ~n31331 ;
  assign y16440 = n31333 ;
  assign y16441 = n31334 ;
  assign y16442 = ~1'b0 ;
  assign y16443 = n31338 ;
  assign y16444 = ~1'b0 ;
  assign y16445 = n31340 ;
  assign y16446 = ~n31341 ;
  assign y16447 = n31347 ;
  assign y16448 = n31349 ;
  assign y16449 = n31350 ;
  assign y16450 = ~1'b0 ;
  assign y16451 = n31351 ;
  assign y16452 = ~1'b0 ;
  assign y16453 = n31354 ;
  assign y16454 = n31356 ;
  assign y16455 = ~n31358 ;
  assign y16456 = ~n31359 ;
  assign y16457 = n31360 ;
  assign y16458 = ~n6943 ;
  assign y16459 = n31361 ;
  assign y16460 = ~n31363 ;
  assign y16461 = ~n31364 ;
  assign y16462 = n31365 ;
  assign y16463 = ~1'b0 ;
  assign y16464 = n31366 ;
  assign y16465 = n31367 ;
  assign y16466 = ~1'b0 ;
  assign y16467 = n31372 ;
  assign y16468 = n31374 ;
  assign y16469 = ~1'b0 ;
  assign y16470 = ~1'b0 ;
  assign y16471 = n31379 ;
  assign y16472 = ~1'b0 ;
  assign y16473 = n31380 ;
  assign y16474 = ~n31387 ;
  assign y16475 = n31388 ;
  assign y16476 = ~1'b0 ;
  assign y16477 = ~n31389 ;
  assign y16478 = n31391 ;
  assign y16479 = n23314 ;
  assign y16480 = ~1'b0 ;
  assign y16481 = ~1'b0 ;
  assign y16482 = ~1'b0 ;
  assign y16483 = ~1'b0 ;
  assign y16484 = ~n31392 ;
  assign y16485 = ~1'b0 ;
  assign y16486 = n31398 ;
  assign y16487 = ~n31399 ;
  assign y16488 = ~1'b0 ;
  assign y16489 = ~1'b0 ;
  assign y16490 = n14068 ;
  assign y16491 = ~n31400 ;
  assign y16492 = n31401 ;
  assign y16493 = n31403 ;
  assign y16494 = ~n31404 ;
  assign y16495 = ~1'b0 ;
  assign y16496 = ~n31406 ;
  assign y16497 = n31410 ;
  assign y16498 = ~1'b0 ;
  assign y16499 = ~n31411 ;
  assign y16500 = 1'b0 ;
  assign y16501 = ~1'b0 ;
  assign y16502 = n31412 ;
  assign y16503 = ~n31414 ;
  assign y16504 = ~1'b0 ;
  assign y16505 = n31415 ;
  assign y16506 = n31416 ;
  assign y16507 = ~n31417 ;
  assign y16508 = ~n31420 ;
  assign y16509 = n11040 ;
  assign y16510 = ~1'b0 ;
  assign y16511 = n31421 ;
  assign y16512 = n31019 ;
  assign y16513 = n31427 ;
  assign y16514 = ~n31428 ;
  assign y16515 = n31430 ;
  assign y16516 = n31433 ;
  assign y16517 = n31435 ;
  assign y16518 = n31436 ;
  assign y16519 = n31439 ;
  assign y16520 = ~n31442 ;
  assign y16521 = n31444 ;
  assign y16522 = ~1'b0 ;
  assign y16523 = ~1'b0 ;
  assign y16524 = n31449 ;
  assign y16525 = ~n31450 ;
  assign y16526 = n31452 ;
  assign y16527 = n19175 ;
  assign y16528 = ~n31453 ;
  assign y16529 = ~n31456 ;
  assign y16530 = ~1'b0 ;
  assign y16531 = ~n31460 ;
  assign y16532 = ~n31462 ;
  assign y16533 = n31464 ;
  assign y16534 = n31469 ;
  assign y16535 = n31474 ;
  assign y16536 = ~n31482 ;
  assign y16537 = n31483 ;
  assign y16538 = ~1'b0 ;
  assign y16539 = ~n31487 ;
  assign y16540 = ~1'b0 ;
  assign y16541 = ~n31488 ;
  assign y16542 = ~n5696 ;
  assign y16543 = n31489 ;
  assign y16544 = ~1'b0 ;
  assign y16545 = n31491 ;
  assign y16546 = n31493 ;
  assign y16547 = ~n31496 ;
  assign y16548 = n31497 ;
  assign y16549 = ~1'b0 ;
  assign y16550 = ~n30121 ;
  assign y16551 = ~x19 ;
  assign y16552 = ~1'b0 ;
  assign y16553 = n31500 ;
  assign y16554 = n31503 ;
  assign y16555 = n31505 ;
  assign y16556 = ~n31510 ;
  assign y16557 = n31511 ;
  assign y16558 = ~n9905 ;
  assign y16559 = ~1'b0 ;
  assign y16560 = ~n31512 ;
  assign y16561 = ~n25983 ;
  assign y16562 = ~1'b0 ;
  assign y16563 = n31513 ;
  assign y16564 = n31514 ;
  assign y16565 = ~1'b0 ;
  assign y16566 = n31515 ;
  assign y16567 = n31516 ;
  assign y16568 = n7027 ;
  assign y16569 = ~n31519 ;
  assign y16570 = ~n31522 ;
  assign y16571 = n31523 ;
  assign y16572 = n31528 ;
  assign y16573 = ~n31530 ;
  assign y16574 = ~1'b0 ;
  assign y16575 = ~1'b0 ;
  assign y16576 = ~n31531 ;
  assign y16577 = ~n31534 ;
  assign y16578 = ~1'b0 ;
  assign y16579 = ~1'b0 ;
  assign y16580 = ~1'b0 ;
  assign y16581 = ~n31535 ;
  assign y16582 = n5382 ;
  assign y16583 = n31536 ;
  assign y16584 = ~1'b0 ;
  assign y16585 = ~1'b0 ;
  assign y16586 = ~n31538 ;
  assign y16587 = ~1'b0 ;
  assign y16588 = n31539 ;
  assign y16589 = ~1'b0 ;
  assign y16590 = ~1'b0 ;
  assign y16591 = ~n31540 ;
  assign y16592 = n31541 ;
  assign y16593 = ~1'b0 ;
  assign y16594 = ~n31543 ;
  assign y16595 = n31547 ;
  assign y16596 = n31551 ;
  assign y16597 = ~1'b0 ;
  assign y16598 = n31552 ;
  assign y16599 = n31553 ;
  assign y16600 = ~1'b0 ;
  assign y16601 = ~n31556 ;
  assign y16602 = n31557 ;
  assign y16603 = ~1'b0 ;
  assign y16604 = n31563 ;
  assign y16605 = n31565 ;
  assign y16606 = n31567 ;
  assign y16607 = n31568 ;
  assign y16608 = n31570 ;
  assign y16609 = n31571 ;
  assign y16610 = ~n31574 ;
  assign y16611 = ~1'b0 ;
  assign y16612 = ~n31575 ;
  assign y16613 = n31580 ;
  assign y16614 = n31590 ;
  assign y16615 = ~1'b0 ;
  assign y16616 = ~n31595 ;
  assign y16617 = ~1'b0 ;
  assign y16618 = ~n31596 ;
  assign y16619 = n31603 ;
  assign y16620 = n31604 ;
  assign y16621 = ~n31605 ;
  assign y16622 = n31612 ;
  assign y16623 = ~n31614 ;
  assign y16624 = n31618 ;
  assign y16625 = n31621 ;
  assign y16626 = n31622 ;
  assign y16627 = ~n31624 ;
  assign y16628 = ~n31626 ;
  assign y16629 = ~n31629 ;
  assign y16630 = n31632 ;
  assign y16631 = ~n12079 ;
  assign y16632 = ~n31634 ;
  assign y16633 = ~n31635 ;
  assign y16634 = ~n31637 ;
  assign y16635 = n31639 ;
  assign y16636 = n31644 ;
  assign y16637 = n31648 ;
  assign y16638 = n31650 ;
  assign y16639 = ~1'b0 ;
  assign y16640 = n31651 ;
  assign y16641 = n31652 ;
  assign y16642 = ~n31653 ;
  assign y16643 = ~n31655 ;
  assign y16644 = ~1'b0 ;
  assign y16645 = n31657 ;
  assign y16646 = ~n31658 ;
  assign y16647 = n31659 ;
  assign y16648 = ~1'b0 ;
  assign y16649 = n31660 ;
  assign y16650 = ~n9814 ;
  assign y16651 = ~n31661 ;
  assign y16652 = ~1'b0 ;
  assign y16653 = 1'b0 ;
  assign y16654 = ~n31670 ;
  assign y16655 = 1'b0 ;
  assign y16656 = ~n31671 ;
  assign y16657 = ~1'b0 ;
  assign y16658 = n6155 ;
  assign y16659 = n31672 ;
  assign y16660 = ~1'b0 ;
  assign y16661 = ~n31680 ;
  assign y16662 = n31683 ;
  assign y16663 = ~1'b0 ;
  assign y16664 = n31685 ;
  assign y16665 = ~1'b0 ;
  assign y16666 = ~n31689 ;
  assign y16667 = ~1'b0 ;
  assign y16668 = n31693 ;
  assign y16669 = n31695 ;
  assign y16670 = 1'b0 ;
  assign y16671 = n31696 ;
  assign y16672 = ~1'b0 ;
  assign y16673 = n31702 ;
  assign y16674 = ~1'b0 ;
  assign y16675 = ~n31705 ;
  assign y16676 = ~n31706 ;
  assign y16677 = ~n31708 ;
  assign y16678 = n31710 ;
  assign y16679 = n31712 ;
  assign y16680 = n31713 ;
  assign y16681 = n31714 ;
  assign y16682 = ~1'b0 ;
  assign y16683 = ~1'b0 ;
  assign y16684 = n31715 ;
  assign y16685 = n31716 ;
  assign y16686 = ~n31719 ;
  assign y16687 = ~n31723 ;
  assign y16688 = ~n8254 ;
  assign y16689 = n11162 ;
  assign y16690 = n31726 ;
  assign y16691 = ~1'b0 ;
  assign y16692 = ~n31729 ;
  assign y16693 = 1'b0 ;
  assign y16694 = n31730 ;
  assign y16695 = n31732 ;
  assign y16696 = ~1'b0 ;
  assign y16697 = n31739 ;
  assign y16698 = n31744 ;
  assign y16699 = n31745 ;
  assign y16700 = 1'b0 ;
  assign y16701 = ~1'b0 ;
  assign y16702 = 1'b0 ;
  assign y16703 = ~n31748 ;
  assign y16704 = ~x212 ;
  assign y16705 = n31750 ;
  assign y16706 = ~n20633 ;
  assign y16707 = n21004 ;
  assign y16708 = n31751 ;
  assign y16709 = ~n31753 ;
  assign y16710 = n31756 ;
  assign y16711 = ~n7679 ;
  assign y16712 = ~n31758 ;
  assign y16713 = n31763 ;
  assign y16714 = n31765 ;
  assign y16715 = n31766 ;
  assign y16716 = n31769 ;
  assign y16717 = n31771 ;
  assign y16718 = n4934 ;
  assign y16719 = n31772 ;
  assign y16720 = ~n31774 ;
  assign y16721 = n31776 ;
  assign y16722 = n31779 ;
  assign y16723 = n31781 ;
  assign y16724 = ~1'b0 ;
  assign y16725 = n31791 ;
  assign y16726 = n31792 ;
  assign y16727 = ~n31793 ;
  assign y16728 = ~1'b0 ;
  assign y16729 = n31795 ;
  assign y16730 = ~1'b0 ;
  assign y16731 = ~n31799 ;
  assign y16732 = ~n31803 ;
  assign y16733 = ~1'b0 ;
  assign y16734 = ~n31808 ;
  assign y16735 = n31811 ;
  assign y16736 = ~1'b0 ;
  assign y16737 = n31815 ;
  assign y16738 = n31818 ;
  assign y16739 = ~1'b0 ;
  assign y16740 = ~1'b0 ;
  assign y16741 = ~n31820 ;
  assign y16742 = ~n31826 ;
  assign y16743 = n31830 ;
  assign y16744 = ~n31832 ;
  assign y16745 = ~1'b0 ;
  assign y16746 = n31835 ;
  assign y16747 = ~1'b0 ;
  assign y16748 = ~1'b0 ;
  assign y16749 = 1'b0 ;
  assign y16750 = ~1'b0 ;
  assign y16751 = ~n8270 ;
  assign y16752 = ~n31847 ;
  assign y16753 = ~1'b0 ;
  assign y16754 = ~n31848 ;
  assign y16755 = ~n31851 ;
  assign y16756 = ~n31854 ;
  assign y16757 = ~1'b0 ;
  assign y16758 = n31859 ;
  assign y16759 = n31862 ;
  assign y16760 = n31863 ;
  assign y16761 = ~1'b0 ;
  assign y16762 = ~n1088 ;
  assign y16763 = ~n31868 ;
  assign y16764 = n31872 ;
  assign y16765 = ~n31874 ;
  assign y16766 = ~n31877 ;
  assign y16767 = ~n4426 ;
  assign y16768 = ~1'b0 ;
  assign y16769 = n31878 ;
  assign y16770 = ~1'b0 ;
  assign y16771 = n31879 ;
  assign y16772 = ~n31881 ;
  assign y16773 = ~1'b0 ;
  assign y16774 = ~1'b0 ;
  assign y16775 = ~n31883 ;
  assign y16776 = ~1'b0 ;
  assign y16777 = ~n31887 ;
  assign y16778 = ~n31889 ;
  assign y16779 = ~1'b0 ;
  assign y16780 = ~n31893 ;
  assign y16781 = n31895 ;
  assign y16782 = n2414 ;
  assign y16783 = ~1'b0 ;
  assign y16784 = ~n31896 ;
  assign y16785 = ~1'b0 ;
  assign y16786 = ~1'b0 ;
  assign y16787 = ~n31897 ;
  assign y16788 = n31898 ;
  assign y16789 = n31899 ;
  assign y16790 = n31900 ;
  assign y16791 = n31904 ;
  assign y16792 = ~1'b0 ;
  assign y16793 = ~1'b0 ;
  assign y16794 = ~1'b0 ;
  assign y16795 = ~1'b0 ;
  assign y16796 = ~1'b0 ;
  assign y16797 = ~n31909 ;
  assign y16798 = n31912 ;
  assign y16799 = ~n18472 ;
  assign y16800 = n31915 ;
  assign y16801 = ~1'b0 ;
  assign y16802 = ~n31916 ;
  assign y16803 = ~1'b0 ;
  assign y16804 = n31926 ;
  assign y16805 = n31928 ;
  assign y16806 = ~n31929 ;
  assign y16807 = ~n31931 ;
  assign y16808 = ~1'b0 ;
  assign y16809 = ~1'b0 ;
  assign y16810 = ~1'b0 ;
  assign y16811 = ~1'b0 ;
  assign y16812 = n31934 ;
  assign y16813 = ~n31935 ;
  assign y16814 = ~1'b0 ;
  assign y16815 = ~n31948 ;
  assign y16816 = n31953 ;
  assign y16817 = ~n31954 ;
  assign y16818 = ~n31957 ;
  assign y16819 = n2194 ;
  assign y16820 = ~1'b0 ;
  assign y16821 = n31960 ;
  assign y16822 = ~1'b0 ;
  assign y16823 = n31961 ;
  assign y16824 = ~n31963 ;
  assign y16825 = ~n31968 ;
  assign y16826 = ~n31971 ;
  assign y16827 = n13414 ;
  assign y16828 = ~n31976 ;
  assign y16829 = ~1'b0 ;
  assign y16830 = ~1'b0 ;
  assign y16831 = n31977 ;
  assign y16832 = ~n31978 ;
  assign y16833 = 1'b0 ;
  assign y16834 = ~n31980 ;
  assign y16835 = n31981 ;
  assign y16836 = ~n31982 ;
  assign y16837 = n31985 ;
  assign y16838 = n31989 ;
  assign y16839 = ~1'b0 ;
  assign y16840 = ~1'b0 ;
  assign y16841 = ~n31992 ;
  assign y16842 = ~1'b0 ;
  assign y16843 = ~1'b0 ;
  assign y16844 = ~n31993 ;
  assign y16845 = ~n31994 ;
  assign y16846 = n31997 ;
  assign y16847 = n31999 ;
  assign y16848 = n32000 ;
  assign y16849 = ~n32001 ;
  assign y16850 = ~1'b0 ;
  assign y16851 = ~1'b0 ;
  assign y16852 = ~n32004 ;
  assign y16853 = n32005 ;
  assign y16854 = ~1'b0 ;
  assign y16855 = ~1'b0 ;
  assign y16856 = ~1'b0 ;
  assign y16857 = ~1'b0 ;
  assign y16858 = 1'b0 ;
  assign y16859 = n32006 ;
  assign y16860 = ~n32008 ;
  assign y16861 = n32009 ;
  assign y16862 = ~1'b0 ;
  assign y16863 = ~1'b0 ;
  assign y16864 = ~n32011 ;
  assign y16865 = ~1'b0 ;
  assign y16866 = ~1'b0 ;
  assign y16867 = n25926 ;
  assign y16868 = n28627 ;
  assign y16869 = ~n32014 ;
  assign y16870 = ~n32018 ;
  assign y16871 = ~n32022 ;
  assign y16872 = ~1'b0 ;
  assign y16873 = n32026 ;
  assign y16874 = ~1'b0 ;
  assign y16875 = n32027 ;
  assign y16876 = n32028 ;
  assign y16877 = ~n32030 ;
  assign y16878 = n32032 ;
  assign y16879 = ~1'b0 ;
  assign y16880 = ~n32038 ;
  assign y16881 = n32044 ;
  assign y16882 = 1'b0 ;
  assign y16883 = ~1'b0 ;
  assign y16884 = n32048 ;
  assign y16885 = ~1'b0 ;
  assign y16886 = n32052 ;
  assign y16887 = ~n32053 ;
  assign y16888 = n32056 ;
  assign y16889 = n18188 ;
  assign y16890 = n32057 ;
  assign y16891 = ~1'b0 ;
  assign y16892 = ~1'b0 ;
  assign y16893 = n32059 ;
  assign y16894 = ~n32061 ;
  assign y16895 = ~1'b0 ;
  assign y16896 = n32063 ;
  assign y16897 = ~1'b0 ;
  assign y16898 = ~n32065 ;
  assign y16899 = n32067 ;
  assign y16900 = n32069 ;
  assign y16901 = n32071 ;
  assign y16902 = n32073 ;
  assign y16903 = ~1'b0 ;
  assign y16904 = ~1'b0 ;
  assign y16905 = ~n32075 ;
  assign y16906 = ~1'b0 ;
  assign y16907 = n32076 ;
  assign y16908 = n32077 ;
  assign y16909 = ~1'b0 ;
  assign y16910 = ~1'b0 ;
  assign y16911 = ~n32078 ;
  assign y16912 = n32079 ;
  assign y16913 = n32080 ;
  assign y16914 = 1'b0 ;
  assign y16915 = n32083 ;
  assign y16916 = ~n32089 ;
  assign y16917 = ~n32091 ;
  assign y16918 = ~n535 ;
  assign y16919 = ~n32092 ;
  assign y16920 = ~n32095 ;
  assign y16921 = ~1'b0 ;
  assign y16922 = n32097 ;
  assign y16923 = n32102 ;
  assign y16924 = ~1'b0 ;
  assign y16925 = ~1'b0 ;
  assign y16926 = ~1'b0 ;
  assign y16927 = ~1'b0 ;
  assign y16928 = ~1'b0 ;
  assign y16929 = n32104 ;
  assign y16930 = ~1'b0 ;
  assign y16931 = ~1'b0 ;
  assign y16932 = ~n32109 ;
  assign y16933 = ~1'b0 ;
  assign y16934 = ~n32112 ;
  assign y16935 = ~1'b0 ;
  assign y16936 = n32120 ;
  assign y16937 = ~1'b0 ;
  assign y16938 = ~1'b0 ;
  assign y16939 = n32123 ;
  assign y16940 = ~n32126 ;
  assign y16941 = n32128 ;
  assign y16942 = n32129 ;
  assign y16943 = n32133 ;
  assign y16944 = ~1'b0 ;
  assign y16945 = ~n32135 ;
  assign y16946 = ~1'b0 ;
  assign y16947 = n32137 ;
  assign y16948 = ~1'b0 ;
  assign y16949 = ~n10174 ;
  assign y16950 = ~n32140 ;
  assign y16951 = ~n32143 ;
  assign y16952 = n32149 ;
  assign y16953 = n32153 ;
  assign y16954 = n32157 ;
  assign y16955 = ~n32160 ;
  assign y16956 = ~1'b0 ;
  assign y16957 = ~n32164 ;
  assign y16958 = ~n32165 ;
  assign y16959 = ~n32168 ;
  assign y16960 = ~n32173 ;
  assign y16961 = ~n32177 ;
  assign y16962 = ~1'b0 ;
  assign y16963 = n32178 ;
  assign y16964 = n32179 ;
  assign y16965 = n32181 ;
  assign y16966 = ~1'b0 ;
  assign y16967 = ~n32186 ;
  assign y16968 = ~1'b0 ;
  assign y16969 = n32187 ;
  assign y16970 = ~1'b0 ;
  assign y16971 = ~1'b0 ;
  assign y16972 = ~1'b0 ;
  assign y16973 = ~1'b0 ;
  assign y16974 = ~n32189 ;
  assign y16975 = ~n11818 ;
  assign y16976 = n32191 ;
  assign y16977 = ~1'b0 ;
  assign y16978 = n32192 ;
  assign y16979 = ~n32196 ;
  assign y16980 = ~1'b0 ;
  assign y16981 = n32197 ;
  assign y16982 = ~n32199 ;
  assign y16983 = n32201 ;
  assign y16984 = n32203 ;
  assign y16985 = ~1'b0 ;
  assign y16986 = ~1'b0 ;
  assign y16987 = n32204 ;
  assign y16988 = n32206 ;
  assign y16989 = ~n32212 ;
  assign y16990 = n32213 ;
  assign y16991 = ~n32215 ;
  assign y16992 = n32217 ;
  assign y16993 = ~1'b0 ;
  assign y16994 = ~n32220 ;
  assign y16995 = ~n32223 ;
  assign y16996 = ~n25708 ;
  assign y16997 = ~1'b0 ;
  assign y16998 = n31376 ;
  assign y16999 = ~n32224 ;
  assign y17000 = n32225 ;
  assign y17001 = ~1'b0 ;
  assign y17002 = ~n32229 ;
  assign y17003 = ~n28745 ;
  assign y17004 = ~n32230 ;
  assign y17005 = ~n32234 ;
  assign y17006 = n32236 ;
  assign y17007 = ~n32238 ;
  assign y17008 = n32240 ;
  assign y17009 = ~n6164 ;
  assign y17010 = n32242 ;
  assign y17011 = ~n32243 ;
  assign y17012 = ~n32245 ;
  assign y17013 = n32247 ;
  assign y17014 = 1'b0 ;
  assign y17015 = n32250 ;
  assign y17016 = ~n32253 ;
  assign y17017 = ~n10926 ;
  assign y17018 = n32254 ;
  assign y17019 = n32256 ;
  assign y17020 = ~n32258 ;
  assign y17021 = ~n32260 ;
  assign y17022 = ~n32261 ;
  assign y17023 = ~n32265 ;
  assign y17024 = ~1'b0 ;
  assign y17025 = n32268 ;
  assign y17026 = ~n32269 ;
  assign y17027 = ~n32271 ;
  assign y17028 = ~1'b0 ;
  assign y17029 = ~1'b0 ;
  assign y17030 = ~n32272 ;
  assign y17031 = n32274 ;
  assign y17032 = 1'b0 ;
  assign y17033 = n18229 ;
  assign y17034 = n32276 ;
  assign y17035 = ~1'b0 ;
  assign y17036 = ~n32277 ;
  assign y17037 = ~n32280 ;
  assign y17038 = n32283 ;
  assign y17039 = ~n32284 ;
  assign y17040 = ~n32287 ;
  assign y17041 = ~1'b0 ;
  assign y17042 = n32288 ;
  assign y17043 = ~1'b0 ;
  assign y17044 = n32291 ;
  assign y17045 = ~1'b0 ;
  assign y17046 = n32293 ;
  assign y17047 = ~n27615 ;
  assign y17048 = ~n32295 ;
  assign y17049 = n15180 ;
  assign y17050 = n32296 ;
  assign y17051 = ~n32301 ;
  assign y17052 = ~1'b0 ;
  assign y17053 = 1'b0 ;
  assign y17054 = n32303 ;
  assign y17055 = n32305 ;
  assign y17056 = ~n32307 ;
  assign y17057 = ~n32309 ;
  assign y17058 = ~n4305 ;
  assign y17059 = ~1'b0 ;
  assign y17060 = ~n32312 ;
  assign y17061 = ~n32314 ;
  assign y17062 = ~n32316 ;
  assign y17063 = ~n32318 ;
  assign y17064 = ~1'b0 ;
  assign y17065 = n32319 ;
  assign y17066 = n32320 ;
  assign y17067 = ~1'b0 ;
  assign y17068 = ~1'b0 ;
  assign y17069 = n32322 ;
  assign y17070 = ~1'b0 ;
  assign y17071 = ~n32324 ;
  assign y17072 = ~1'b0 ;
  assign y17073 = ~1'b0 ;
  assign y17074 = n32325 ;
  assign y17075 = ~1'b0 ;
  assign y17076 = ~n32326 ;
  assign y17077 = ~n32329 ;
  assign y17078 = ~n32332 ;
  assign y17079 = n32333 ;
  assign y17080 = n32334 ;
  assign y17081 = ~1'b0 ;
  assign y17082 = ~n32340 ;
  assign y17083 = ~1'b0 ;
  assign y17084 = ~n32350 ;
  assign y17085 = 1'b0 ;
  assign y17086 = ~n32352 ;
  assign y17087 = 1'b0 ;
  assign y17088 = ~n32354 ;
  assign y17089 = n32355 ;
  assign y17090 = ~n32356 ;
  assign y17091 = n32358 ;
  assign y17092 = n32359 ;
  assign y17093 = ~n32360 ;
  assign y17094 = n32361 ;
  assign y17095 = ~n32366 ;
  assign y17096 = n32367 ;
  assign y17097 = ~1'b0 ;
  assign y17098 = ~n32369 ;
  assign y17099 = ~n32373 ;
  assign y17100 = n5291 ;
  assign y17101 = n32374 ;
  assign y17102 = ~1'b0 ;
  assign y17103 = n32375 ;
  assign y17104 = ~n32377 ;
  assign y17105 = n6990 ;
  assign y17106 = n32379 ;
  assign y17107 = ~n32381 ;
  assign y17108 = ~1'b0 ;
  assign y17109 = ~n32382 ;
  assign y17110 = ~n32383 ;
  assign y17111 = ~1'b0 ;
  assign y17112 = ~n9416 ;
  assign y17113 = ~1'b0 ;
  assign y17114 = n32390 ;
  assign y17115 = ~1'b0 ;
  assign y17116 = n32393 ;
  assign y17117 = n32396 ;
  assign y17118 = ~1'b0 ;
  assign y17119 = n32398 ;
  assign y17120 = 1'b0 ;
  assign y17121 = ~n32404 ;
  assign y17122 = n32408 ;
  assign y17123 = ~1'b0 ;
  assign y17124 = ~n32411 ;
  assign y17125 = n32412 ;
  assign y17126 = ~n32414 ;
  assign y17127 = n32415 ;
  assign y17128 = ~1'b0 ;
  assign y17129 = ~1'b0 ;
  assign y17130 = n17338 ;
  assign y17131 = ~1'b0 ;
  assign y17132 = ~1'b0 ;
  assign y17133 = ~1'b0 ;
  assign y17134 = ~n32416 ;
  assign y17135 = n32417 ;
  assign y17136 = ~n32419 ;
  assign y17137 = n32421 ;
  assign y17138 = ~n32423 ;
  assign y17139 = n32424 ;
  assign y17140 = ~n32427 ;
  assign y17141 = ~1'b0 ;
  assign y17142 = ~1'b0 ;
  assign y17143 = ~n32428 ;
  assign y17144 = ~n32434 ;
  assign y17145 = ~1'b0 ;
  assign y17146 = ~n32438 ;
  assign y17147 = n8933 ;
  assign y17148 = ~n32439 ;
  assign y17149 = ~1'b0 ;
  assign y17150 = ~1'b0 ;
  assign y17151 = ~1'b0 ;
  assign y17152 = n32440 ;
  assign y17153 = n32441 ;
  assign y17154 = ~1'b0 ;
  assign y17155 = n32443 ;
  assign y17156 = ~1'b0 ;
  assign y17157 = ~n32444 ;
  assign y17158 = ~1'b0 ;
  assign y17159 = ~1'b0 ;
  assign y17160 = n32445 ;
  assign y17161 = n4852 ;
  assign y17162 = n25858 ;
  assign y17163 = ~n32446 ;
  assign y17164 = n32447 ;
  assign y17165 = n32448 ;
  assign y17166 = ~n32452 ;
  assign y17167 = ~n32453 ;
  assign y17168 = ~1'b0 ;
  assign y17169 = ~1'b0 ;
  assign y17170 = n32458 ;
  assign y17171 = ~n32459 ;
  assign y17172 = n32460 ;
  assign y17173 = ~1'b0 ;
  assign y17174 = ~1'b0 ;
  assign y17175 = ~1'b0 ;
  assign y17176 = ~n20298 ;
  assign y17177 = ~1'b0 ;
  assign y17178 = 1'b0 ;
  assign y17179 = ~1'b0 ;
  assign y17180 = ~1'b0 ;
  assign y17181 = ~n32467 ;
  assign y17182 = ~n32472 ;
  assign y17183 = n32473 ;
  assign y17184 = ~n32474 ;
  assign y17185 = ~1'b0 ;
  assign y17186 = n32476 ;
  assign y17187 = ~n32478 ;
  assign y17188 = ~n32482 ;
  assign y17189 = ~n32484 ;
  assign y17190 = ~1'b0 ;
  assign y17191 = ~n32487 ;
  assign y17192 = ~1'b0 ;
  assign y17193 = ~n32491 ;
  assign y17194 = n32492 ;
  assign y17195 = ~1'b0 ;
  assign y17196 = n32494 ;
  assign y17197 = ~1'b0 ;
  assign y17198 = n32495 ;
  assign y17199 = ~1'b0 ;
  assign y17200 = ~1'b0 ;
  assign y17201 = n32502 ;
  assign y17202 = ~1'b0 ;
  assign y17203 = ~n32508 ;
  assign y17204 = ~n32510 ;
  assign y17205 = n32513 ;
  assign y17206 = ~n32515 ;
  assign y17207 = n32517 ;
  assign y17208 = n32518 ;
  assign y17209 = ~n32521 ;
  assign y17210 = n32529 ;
  assign y17211 = n32531 ;
  assign y17212 = ~1'b0 ;
  assign y17213 = ~1'b0 ;
  assign y17214 = ~1'b0 ;
  assign y17215 = n32532 ;
  assign y17216 = ~1'b0 ;
  assign y17217 = n32534 ;
  assign y17218 = n32538 ;
  assign y17219 = ~n32539 ;
  assign y17220 = ~1'b0 ;
  assign y17221 = ~n32541 ;
  assign y17222 = ~1'b0 ;
  assign y17223 = ~n32542 ;
  assign y17224 = n32543 ;
  assign y17225 = n32546 ;
  assign y17226 = ~1'b0 ;
  assign y17227 = ~n32553 ;
  assign y17228 = ~1'b0 ;
  assign y17229 = ~n32557 ;
  assign y17230 = ~1'b0 ;
  assign y17231 = n32558 ;
  assign y17232 = ~n32559 ;
  assign y17233 = ~1'b0 ;
  assign y17234 = ~1'b0 ;
  assign y17235 = ~1'b0 ;
  assign y17236 = n32560 ;
  assign y17237 = ~n32562 ;
  assign y17238 = ~n32565 ;
  assign y17239 = ~1'b0 ;
  assign y17240 = n21191 ;
  assign y17241 = ~n10529 ;
  assign y17242 = ~n32566 ;
  assign y17243 = n32567 ;
  assign y17244 = ~1'b0 ;
  assign y17245 = ~n32572 ;
  assign y17246 = n32573 ;
  assign y17247 = ~n32576 ;
  assign y17248 = n32578 ;
  assign y17249 = ~n32581 ;
  assign y17250 = n32586 ;
  assign y17251 = ~n32593 ;
  assign y17252 = ~n32594 ;
  assign y17253 = ~n32596 ;
  assign y17254 = n25700 ;
  assign y17255 = ~n32600 ;
  assign y17256 = ~n32602 ;
  assign y17257 = n32604 ;
  assign y17258 = ~n32606 ;
  assign y17259 = ~1'b0 ;
  assign y17260 = ~1'b0 ;
  assign y17261 = 1'b0 ;
  assign y17262 = ~1'b0 ;
  assign y17263 = ~n32608 ;
  assign y17264 = ~n25147 ;
  assign y17265 = n32612 ;
  assign y17266 = n32615 ;
  assign y17267 = ~1'b0 ;
  assign y17268 = ~n32616 ;
  assign y17269 = ~1'b0 ;
  assign y17270 = ~n32619 ;
  assign y17271 = n32622 ;
  assign y17272 = ~1'b0 ;
  assign y17273 = ~n32627 ;
  assign y17274 = n32628 ;
  assign y17275 = ~1'b0 ;
  assign y17276 = n32630 ;
  assign y17277 = ~n32632 ;
  assign y17278 = ~n6397 ;
  assign y17279 = n32633 ;
  assign y17280 = ~1'b0 ;
  assign y17281 = ~n32634 ;
  assign y17282 = n32640 ;
  assign y17283 = ~n32642 ;
  assign y17284 = 1'b0 ;
  assign y17285 = ~n32644 ;
  assign y17286 = ~1'b0 ;
  assign y17287 = n32647 ;
  assign y17288 = ~n32650 ;
  assign y17289 = ~n32653 ;
  assign y17290 = n32656 ;
  assign y17291 = ~n32657 ;
  assign y17292 = ~1'b0 ;
  assign y17293 = ~n32658 ;
  assign y17294 = ~1'b0 ;
  assign y17295 = n32663 ;
  assign y17296 = ~n32664 ;
  assign y17297 = n32665 ;
  assign y17298 = ~n5118 ;
  assign y17299 = ~n32666 ;
  assign y17300 = ~n32674 ;
  assign y17301 = ~n32676 ;
  assign y17302 = ~1'b0 ;
  assign y17303 = n32679 ;
  assign y17304 = n32681 ;
  assign y17305 = ~1'b0 ;
  assign y17306 = n32684 ;
  assign y17307 = ~1'b0 ;
  assign y17308 = ~n32688 ;
  assign y17309 = n32690 ;
  assign y17310 = ~n32692 ;
  assign y17311 = ~1'b0 ;
  assign y17312 = n14543 ;
  assign y17313 = n32693 ;
  assign y17314 = ~n32695 ;
  assign y17315 = ~1'b0 ;
  assign y17316 = ~1'b0 ;
  assign y17317 = ~1'b0 ;
  assign y17318 = n32696 ;
  assign y17319 = ~1'b0 ;
  assign y17320 = n32698 ;
  assign y17321 = n32702 ;
  assign y17322 = ~n32706 ;
  assign y17323 = ~n32708 ;
  assign y17324 = ~n21829 ;
  assign y17325 = ~1'b0 ;
  assign y17326 = ~n32710 ;
  assign y17327 = ~n32712 ;
  assign y17328 = ~1'b0 ;
  assign y17329 = ~n32716 ;
  assign y17330 = ~n32720 ;
  assign y17331 = ~n32721 ;
  assign y17332 = ~n32722 ;
  assign y17333 = ~1'b0 ;
  assign y17334 = n32724 ;
  assign y17335 = 1'b0 ;
  assign y17336 = 1'b0 ;
  assign y17337 = ~1'b0 ;
  assign y17338 = 1'b0 ;
  assign y17339 = n32725 ;
  assign y17340 = ~n32731 ;
  assign y17341 = n32735 ;
  assign y17342 = ~1'b0 ;
  assign y17343 = ~n11127 ;
  assign y17344 = ~1'b0 ;
  assign y17345 = ~1'b0 ;
  assign y17346 = ~n10608 ;
  assign y17347 = n31605 ;
  assign y17348 = ~n32736 ;
  assign y17349 = ~n32737 ;
  assign y17350 = 1'b0 ;
  assign y17351 = n32740 ;
  assign y17352 = ~n32742 ;
  assign y17353 = n32743 ;
  assign y17354 = ~n32746 ;
  assign y17355 = ~n32748 ;
  assign y17356 = n32752 ;
  assign y17357 = n32754 ;
  assign y17358 = ~1'b0 ;
  assign y17359 = n32755 ;
  assign y17360 = ~n32756 ;
  assign y17361 = n32761 ;
  assign y17362 = ~1'b0 ;
  assign y17363 = ~n32763 ;
  assign y17364 = ~n32764 ;
  assign y17365 = n32766 ;
  assign y17366 = ~n32769 ;
  assign y17367 = ~1'b0 ;
  assign y17368 = ~n32771 ;
  assign y17369 = ~1'b0 ;
  assign y17370 = n32772 ;
  assign y17371 = ~n32777 ;
  assign y17372 = ~n17250 ;
  assign y17373 = n32783 ;
  assign y17374 = 1'b0 ;
  assign y17375 = n20001 ;
  assign y17376 = ~n20896 ;
  assign y17377 = ~n24917 ;
  assign y17378 = ~n32787 ;
  assign y17379 = ~n30762 ;
  assign y17380 = 1'b0 ;
  assign y17381 = ~1'b0 ;
  assign y17382 = ~n32792 ;
  assign y17383 = ~n32793 ;
  assign y17384 = n32794 ;
  assign y17385 = ~n32797 ;
  assign y17386 = n32799 ;
  assign y17387 = ~n32806 ;
  assign y17388 = ~1'b0 ;
  assign y17389 = ~1'b0 ;
  assign y17390 = 1'b0 ;
  assign y17391 = n12712 ;
  assign y17392 = ~1'b0 ;
  assign y17393 = ~n32809 ;
  assign y17394 = ~n32811 ;
  assign y17395 = n19381 ;
  assign y17396 = n32814 ;
  assign y17397 = n9758 ;
  assign y17398 = ~n32816 ;
  assign y17399 = n32817 ;
  assign y17400 = n32826 ;
  assign y17401 = ~1'b0 ;
  assign y17402 = ~n16348 ;
  assign y17403 = ~1'b0 ;
  assign y17404 = ~n32827 ;
  assign y17405 = n32830 ;
  assign y17406 = n32836 ;
  assign y17407 = n32837 ;
  assign y17408 = ~n32838 ;
  assign y17409 = ~n32840 ;
  assign y17410 = ~n32841 ;
  assign y17411 = ~1'b0 ;
  assign y17412 = 1'b0 ;
  assign y17413 = n32842 ;
  assign y17414 = ~n32843 ;
  assign y17415 = ~n32844 ;
  assign y17416 = ~1'b0 ;
  assign y17417 = n32847 ;
  assign y17418 = ~1'b0 ;
  assign y17419 = n32851 ;
  assign y17420 = ~n32855 ;
  assign y17421 = ~1'b0 ;
  assign y17422 = n32859 ;
  assign y17423 = n32860 ;
  assign y17424 = n32864 ;
  assign y17425 = ~n32865 ;
  assign y17426 = n32872 ;
  assign y17427 = ~1'b0 ;
  assign y17428 = ~n32876 ;
  assign y17429 = n32881 ;
  assign y17430 = ~1'b0 ;
  assign y17431 = ~n32882 ;
  assign y17432 = n32886 ;
  assign y17433 = ~n32888 ;
  assign y17434 = ~n32890 ;
  assign y17435 = n32891 ;
  assign y17436 = ~1'b0 ;
  assign y17437 = n32892 ;
  assign y17438 = n32894 ;
  assign y17439 = ~1'b0 ;
  assign y17440 = ~1'b0 ;
  assign y17441 = ~n32896 ;
  assign y17442 = n32900 ;
  assign y17443 = ~n32902 ;
  assign y17444 = ~1'b0 ;
  assign y17445 = ~n32905 ;
  assign y17446 = ~n32906 ;
  assign y17447 = n32910 ;
  assign y17448 = ~1'b0 ;
  assign y17449 = ~n32912 ;
  assign y17450 = ~1'b0 ;
  assign y17451 = ~1'b0 ;
  assign y17452 = ~n32917 ;
  assign y17453 = n32918 ;
  assign y17454 = 1'b0 ;
  assign y17455 = n32920 ;
  assign y17456 = ~n32922 ;
  assign y17457 = ~n32926 ;
  assign y17458 = ~n32929 ;
  assign y17459 = ~1'b0 ;
  assign y17460 = ~n32930 ;
  assign y17461 = n32932 ;
  assign y17462 = ~n32936 ;
  assign y17463 = n32937 ;
  assign y17464 = 1'b0 ;
  assign y17465 = 1'b0 ;
  assign y17466 = ~1'b0 ;
  assign y17467 = ~n4835 ;
  assign y17468 = ~n32938 ;
  assign y17469 = n18094 ;
  assign y17470 = n32942 ;
  assign y17471 = ~1'b0 ;
  assign y17472 = 1'b0 ;
  assign y17473 = ~n32944 ;
  assign y17474 = n32947 ;
  assign y17475 = n32948 ;
  assign y17476 = ~1'b0 ;
  assign y17477 = ~n32949 ;
  assign y17478 = ~1'b0 ;
  assign y17479 = x98 ;
  assign y17480 = ~1'b0 ;
  assign y17481 = ~1'b0 ;
  assign y17482 = n32950 ;
  assign y17483 = n32951 ;
  assign y17484 = n32957 ;
  assign y17485 = ~n32958 ;
  assign y17486 = ~1'b0 ;
  assign y17487 = ~n32959 ;
  assign y17488 = ~1'b0 ;
  assign y17489 = ~1'b0 ;
  assign y17490 = ~1'b0 ;
  assign y17491 = ~n32961 ;
  assign y17492 = ~n32963 ;
  assign y17493 = ~n32965 ;
  assign y17494 = ~n32968 ;
  assign y17495 = ~1'b0 ;
  assign y17496 = ~n32971 ;
  assign y17497 = n32976 ;
  assign y17498 = ~1'b0 ;
  assign y17499 = n32978 ;
  assign y17500 = ~1'b0 ;
  assign y17501 = ~n32979 ;
  assign y17502 = n2113 ;
  assign y17503 = ~n32984 ;
  assign y17504 = n32985 ;
  assign y17505 = ~1'b0 ;
  assign y17506 = n32986 ;
  assign y17507 = n32994 ;
  assign y17508 = ~n32995 ;
  assign y17509 = ~1'b0 ;
  assign y17510 = ~1'b0 ;
  assign y17511 = ~n32998 ;
  assign y17512 = ~n22665 ;
  assign y17513 = ~n33001 ;
  assign y17514 = ~n33004 ;
  assign y17515 = ~1'b0 ;
  assign y17516 = n24695 ;
  assign y17517 = ~1'b0 ;
  assign y17518 = ~1'b0 ;
  assign y17519 = n33016 ;
  assign y17520 = n33017 ;
  assign y17521 = ~1'b0 ;
  assign y17522 = n33022 ;
  assign y17523 = n33026 ;
  assign y17524 = n33028 ;
  assign y17525 = ~n33029 ;
  assign y17526 = ~1'b0 ;
  assign y17527 = ~n33030 ;
  assign y17528 = ~1'b0 ;
  assign y17529 = ~n33032 ;
  assign y17530 = ~1'b0 ;
  assign y17531 = n33036 ;
  assign y17532 = ~n33040 ;
  assign y17533 = ~n33044 ;
  assign y17534 = ~1'b0 ;
  assign y17535 = n33046 ;
  assign y17536 = n33047 ;
  assign y17537 = n33048 ;
  assign y17538 = n33050 ;
  assign y17539 = n33054 ;
  assign y17540 = ~n33056 ;
  assign y17541 = n33058 ;
  assign y17542 = ~n33060 ;
  assign y17543 = ~n33061 ;
  assign y17544 = ~1'b0 ;
  assign y17545 = n33063 ;
  assign y17546 = ~n26787 ;
  assign y17547 = n33066 ;
  assign y17548 = ~1'b0 ;
  assign y17549 = ~n12965 ;
  assign y17550 = ~1'b0 ;
  assign y17551 = ~n33070 ;
  assign y17552 = n33072 ;
  assign y17553 = n33076 ;
  assign y17554 = 1'b0 ;
  assign y17555 = ~1'b0 ;
  assign y17556 = n33077 ;
  assign y17557 = ~n33078 ;
  assign y17558 = ~n33083 ;
  assign y17559 = n33084 ;
  assign y17560 = ~n33086 ;
  assign y17561 = n33088 ;
  assign y17562 = n33093 ;
  assign y17563 = ~n33095 ;
  assign y17564 = ~n33097 ;
  assign y17565 = ~n33099 ;
  assign y17566 = n33100 ;
  assign y17567 = ~1'b0 ;
  assign y17568 = n33101 ;
  assign y17569 = n33103 ;
  assign y17570 = n13409 ;
  assign y17571 = n33105 ;
  assign y17572 = ~n33108 ;
  assign y17573 = n33112 ;
  assign y17574 = n16031 ;
  assign y17575 = ~n33115 ;
  assign y17576 = ~n33120 ;
  assign y17577 = ~1'b0 ;
  assign y17578 = ~1'b0 ;
  assign y17579 = ~n33124 ;
  assign y17580 = ~1'b0 ;
  assign y17581 = ~n33126 ;
  assign y17582 = n33127 ;
  assign y17583 = ~1'b0 ;
  assign y17584 = ~n33128 ;
  assign y17585 = ~n33132 ;
  assign y17586 = n33134 ;
  assign y17587 = ~1'b0 ;
  assign y17588 = ~1'b0 ;
  assign y17589 = n33136 ;
  assign y17590 = n33139 ;
  assign y17591 = ~n33140 ;
  assign y17592 = ~n33141 ;
  assign y17593 = ~n33143 ;
  assign y17594 = n33146 ;
  assign y17595 = ~n33148 ;
  assign y17596 = n33149 ;
  assign y17597 = ~1'b0 ;
  assign y17598 = ~1'b0 ;
  assign y17599 = ~1'b0 ;
  assign y17600 = n33151 ;
  assign y17601 = n33154 ;
  assign y17602 = n33155 ;
  assign y17603 = n33157 ;
  assign y17604 = ~n33158 ;
  assign y17605 = ~n33159 ;
  assign y17606 = ~1'b0 ;
  assign y17607 = n33161 ;
  assign y17608 = ~n33162 ;
  assign y17609 = ~1'b0 ;
  assign y17610 = n33164 ;
  assign y17611 = ~1'b0 ;
  assign y17612 = ~1'b0 ;
  assign y17613 = n18254 ;
  assign y17614 = n33167 ;
  assign y17615 = n33168 ;
  assign y17616 = ~n33171 ;
  assign y17617 = n33172 ;
  assign y17618 = n33175 ;
  assign y17619 = n33177 ;
  assign y17620 = ~1'b0 ;
  assign y17621 = n33178 ;
  assign y17622 = ~n33180 ;
  assign y17623 = ~1'b0 ;
  assign y17624 = n33181 ;
  assign y17625 = n33183 ;
  assign y17626 = ~n33184 ;
  assign y17627 = n33185 ;
  assign y17628 = ~1'b0 ;
  assign y17629 = 1'b0 ;
  assign y17630 = ~n33187 ;
  assign y17631 = ~n33189 ;
  assign y17632 = n33191 ;
  assign y17633 = ~n33193 ;
  assign y17634 = n33196 ;
  assign y17635 = ~1'b0 ;
  assign y17636 = n33197 ;
  assign y17637 = ~n33199 ;
  assign y17638 = ~1'b0 ;
  assign y17639 = n33200 ;
  assign y17640 = ~1'b0 ;
  assign y17641 = 1'b0 ;
  assign y17642 = n33202 ;
  assign y17643 = n33207 ;
  assign y17644 = ~1'b0 ;
  assign y17645 = 1'b0 ;
  assign y17646 = n33209 ;
  assign y17647 = n33212 ;
  assign y17648 = ~n33213 ;
  assign y17649 = n33217 ;
  assign y17650 = n33219 ;
  assign y17651 = n33220 ;
  assign y17652 = ~1'b0 ;
  assign y17653 = ~n33228 ;
  assign y17654 = ~n33229 ;
  assign y17655 = ~1'b0 ;
  assign y17656 = ~1'b0 ;
  assign y17657 = ~1'b0 ;
  assign y17658 = n33231 ;
  assign y17659 = ~1'b0 ;
  assign y17660 = ~1'b0 ;
  assign y17661 = ~n8746 ;
  assign y17662 = ~n33234 ;
  assign y17663 = n33235 ;
  assign y17664 = ~n33236 ;
  assign y17665 = 1'b0 ;
  assign y17666 = ~n33237 ;
  assign y17667 = n33238 ;
  assign y17668 = ~n33240 ;
  assign y17669 = n33242 ;
  assign y17670 = ~n30404 ;
  assign y17671 = ~1'b0 ;
  assign y17672 = ~n33243 ;
  assign y17673 = n33245 ;
  assign y17674 = ~n33247 ;
  assign y17675 = n33248 ;
  assign y17676 = ~n26136 ;
  assign y17677 = ~n33251 ;
  assign y17678 = ~1'b0 ;
  assign y17679 = n33252 ;
  assign y17680 = ~1'b0 ;
  assign y17681 = n33254 ;
  assign y17682 = ~n33256 ;
  assign y17683 = ~1'b0 ;
  assign y17684 = ~n33257 ;
  assign y17685 = n33261 ;
  assign y17686 = ~n33263 ;
  assign y17687 = n33265 ;
  assign y17688 = ~n33267 ;
  assign y17689 = ~n33269 ;
  assign y17690 = ~1'b0 ;
  assign y17691 = ~1'b0 ;
  assign y17692 = ~n33271 ;
  assign y17693 = ~n33272 ;
  assign y17694 = n33273 ;
  assign y17695 = ~n33275 ;
  assign y17696 = n33278 ;
  assign y17697 = ~1'b0 ;
  assign y17698 = n33279 ;
  assign y17699 = ~n33283 ;
  assign y17700 = n33285 ;
  assign y17701 = ~1'b0 ;
  assign y17702 = n33286 ;
  assign y17703 = n33288 ;
  assign y17704 = ~n33291 ;
  assign y17705 = n33292 ;
  assign y17706 = 1'b0 ;
  assign y17707 = ~n33293 ;
  assign y17708 = n33294 ;
  assign y17709 = ~1'b0 ;
  assign y17710 = ~n33297 ;
  assign y17711 = n33299 ;
  assign y17712 = ~1'b0 ;
  assign y17713 = n33300 ;
  assign y17714 = n33301 ;
  assign y17715 = ~n33303 ;
  assign y17716 = ~1'b0 ;
  assign y17717 = ~1'b0 ;
  assign y17718 = n33306 ;
  assign y17719 = ~n33307 ;
  assign y17720 = n33309 ;
  assign y17721 = ~1'b0 ;
  assign y17722 = ~1'b0 ;
  assign y17723 = n33310 ;
  assign y17724 = ~n12864 ;
  assign y17725 = ~n33313 ;
  assign y17726 = ~n33317 ;
  assign y17727 = n33323 ;
  assign y17728 = ~n33324 ;
  assign y17729 = 1'b0 ;
  assign y17730 = n33328 ;
  assign y17731 = ~1'b0 ;
  assign y17732 = ~n33334 ;
  assign y17733 = n33335 ;
  assign y17734 = ~n33337 ;
  assign y17735 = n18849 ;
  assign y17736 = ~n33339 ;
  assign y17737 = ~n33344 ;
  assign y17738 = ~1'b0 ;
  assign y17739 = ~n33348 ;
  assign y17740 = ~1'b0 ;
  assign y17741 = n33352 ;
  assign y17742 = ~n33353 ;
  assign y17743 = ~1'b0 ;
  assign y17744 = ~1'b0 ;
  assign y17745 = ~1'b0 ;
  assign y17746 = ~n33355 ;
  assign y17747 = ~1'b0 ;
  assign y17748 = ~n33356 ;
  assign y17749 = ~1'b0 ;
  assign y17750 = ~n33358 ;
  assign y17751 = n33360 ;
  assign y17752 = ~n11369 ;
  assign y17753 = ~n33362 ;
  assign y17754 = n33363 ;
  assign y17755 = n33365 ;
  assign y17756 = ~1'b0 ;
  assign y17757 = n33366 ;
  assign y17758 = n33368 ;
  assign y17759 = n33370 ;
  assign y17760 = ~1'b0 ;
  assign y17761 = ~n33372 ;
  assign y17762 = n33378 ;
  assign y17763 = ~n33381 ;
  assign y17764 = ~n33382 ;
  assign y17765 = ~n33383 ;
  assign y17766 = ~1'b0 ;
  assign y17767 = n33384 ;
  assign y17768 = ~1'b0 ;
  assign y17769 = n33386 ;
  assign y17770 = ~1'b0 ;
  assign y17771 = n33387 ;
  assign y17772 = n33388 ;
  assign y17773 = ~n33389 ;
  assign y17774 = ~1'b0 ;
  assign y17775 = n33391 ;
  assign y17776 = ~n33392 ;
  assign y17777 = ~1'b0 ;
  assign y17778 = ~1'b0 ;
  assign y17779 = ~n33394 ;
  assign y17780 = ~n33396 ;
  assign y17781 = n33401 ;
  assign y17782 = ~1'b0 ;
  assign y17783 = n33403 ;
  assign y17784 = ~n1482 ;
  assign y17785 = ~n33404 ;
  assign y17786 = n33406 ;
  assign y17787 = ~n33411 ;
  assign y17788 = ~1'b0 ;
  assign y17789 = ~1'b0 ;
  assign y17790 = ~n19628 ;
  assign y17791 = ~n33413 ;
  assign y17792 = ~n33415 ;
  assign y17793 = n33416 ;
  assign y17794 = n33417 ;
  assign y17795 = 1'b0 ;
  assign y17796 = n33418 ;
  assign y17797 = ~1'b0 ;
  assign y17798 = ~1'b0 ;
  assign y17799 = ~n33422 ;
  assign y17800 = ~n33424 ;
  assign y17801 = ~n33425 ;
  assign y17802 = n33429 ;
  assign y17803 = ~n33430 ;
  assign y17804 = n3805 ;
  assign y17805 = ~1'b0 ;
  assign y17806 = n33432 ;
  assign y17807 = ~1'b0 ;
  assign y17808 = 1'b0 ;
  assign y17809 = ~n33433 ;
  assign y17810 = ~1'b0 ;
  assign y17811 = ~n33435 ;
  assign y17812 = ~1'b0 ;
  assign y17813 = 1'b0 ;
  assign y17814 = ~n33437 ;
  assign y17815 = ~1'b0 ;
  assign y17816 = ~1'b0 ;
  assign y17817 = n33439 ;
  assign y17818 = n22913 ;
  assign y17819 = ~1'b0 ;
  assign y17820 = ~1'b0 ;
  assign y17821 = ~n33441 ;
  assign y17822 = ~1'b0 ;
  assign y17823 = ~1'b0 ;
  assign y17824 = n33442 ;
  assign y17825 = ~n33446 ;
  assign y17826 = ~n33447 ;
  assign y17827 = ~1'b0 ;
  assign y17828 = n33448 ;
  assign y17829 = ~1'b0 ;
  assign y17830 = n33449 ;
  assign y17831 = ~n33453 ;
  assign y17832 = ~n33455 ;
  assign y17833 = n16236 ;
  assign y17834 = ~n33457 ;
  assign y17835 = ~n33459 ;
  assign y17836 = n33460 ;
  assign y17837 = ~n33462 ;
  assign y17838 = n33463 ;
  assign y17839 = ~1'b0 ;
  assign y17840 = ~n33464 ;
  assign y17841 = n33465 ;
  assign y17842 = ~n33470 ;
  assign y17843 = ~n33472 ;
  assign y17844 = 1'b0 ;
  assign y17845 = n33474 ;
  assign y17846 = ~1'b0 ;
  assign y17847 = n28924 ;
  assign y17848 = ~1'b0 ;
  assign y17849 = n33475 ;
  assign y17850 = ~1'b0 ;
  assign y17851 = n33477 ;
  assign y17852 = ~n33480 ;
  assign y17853 = ~n33487 ;
  assign y17854 = n33491 ;
  assign y17855 = ~1'b0 ;
  assign y17856 = ~n33492 ;
  assign y17857 = ~n33493 ;
  assign y17858 = ~1'b0 ;
  assign y17859 = ~n33498 ;
  assign y17860 = n33502 ;
  assign y17861 = n33504 ;
  assign y17862 = ~1'b0 ;
  assign y17863 = n33510 ;
  assign y17864 = ~n33514 ;
  assign y17865 = ~n33517 ;
  assign y17866 = ~n33518 ;
  assign y17867 = ~1'b0 ;
  assign y17868 = ~n33520 ;
  assign y17869 = ~1'b0 ;
  assign y17870 = ~1'b0 ;
  assign y17871 = ~1'b0 ;
  assign y17872 = n33522 ;
  assign y17873 = n33525 ;
  assign y17874 = ~1'b0 ;
  assign y17875 = n33528 ;
  assign y17876 = ~n1255 ;
  assign y17877 = ~n33531 ;
  assign y17878 = ~n1935 ;
  assign y17879 = ~1'b0 ;
  assign y17880 = ~1'b0 ;
  assign y17881 = ~1'b0 ;
  assign y17882 = n33537 ;
  assign y17883 = ~1'b0 ;
  assign y17884 = n33539 ;
  assign y17885 = ~n33541 ;
  assign y17886 = n4778 ;
  assign y17887 = n33545 ;
  assign y17888 = n33546 ;
  assign y17889 = 1'b0 ;
  assign y17890 = 1'b0 ;
  assign y17891 = n33550 ;
  assign y17892 = n33552 ;
  assign y17893 = n33554 ;
  assign y17894 = ~n33556 ;
  assign y17895 = n33557 ;
  assign y17896 = n33558 ;
  assign y17897 = ~1'b0 ;
  assign y17898 = ~n33562 ;
  assign y17899 = n33565 ;
  assign y17900 = ~1'b0 ;
  assign y17901 = 1'b0 ;
  assign y17902 = ~n33567 ;
  assign y17903 = ~n33568 ;
  assign y17904 = n24626 ;
  assign y17905 = ~n6294 ;
  assign y17906 = n33577 ;
  assign y17907 = n17848 ;
  assign y17908 = n33582 ;
  assign y17909 = n2584 ;
  assign y17910 = ~1'b0 ;
  assign y17911 = ~1'b0 ;
  assign y17912 = ~1'b0 ;
  assign y17913 = ~n33583 ;
  assign y17914 = ~n33584 ;
  assign y17915 = ~1'b0 ;
  assign y17916 = 1'b0 ;
  assign y17917 = ~1'b0 ;
  assign y17918 = n33588 ;
  assign y17919 = ~n33589 ;
  assign y17920 = ~1'b0 ;
  assign y17921 = ~1'b0 ;
  assign y17922 = ~n33592 ;
  assign y17923 = ~1'b0 ;
  assign y17924 = n33593 ;
  assign y17925 = ~n33596 ;
  assign y17926 = ~1'b0 ;
  assign y17927 = n33597 ;
  assign y17928 = ~n33599 ;
  assign y17929 = ~n30519 ;
  assign y17930 = ~n33602 ;
  assign y17931 = ~1'b0 ;
  assign y17932 = ~n33603 ;
  assign y17933 = 1'b0 ;
  assign y17934 = ~n33604 ;
  assign y17935 = n33608 ;
  assign y17936 = ~1'b0 ;
  assign y17937 = ~1'b0 ;
  assign y17938 = ~n18169 ;
  assign y17939 = n13765 ;
  assign y17940 = n33610 ;
  assign y17941 = ~1'b0 ;
  assign y17942 = ~n33611 ;
  assign y17943 = n33615 ;
  assign y17944 = n33616 ;
  assign y17945 = n33618 ;
  assign y17946 = n33620 ;
  assign y17947 = ~1'b0 ;
  assign y17948 = ~n33623 ;
  assign y17949 = ~1'b0 ;
  assign y17950 = ~1'b0 ;
  assign y17951 = ~1'b0 ;
  assign y17952 = ~n33628 ;
  assign y17953 = ~1'b0 ;
  assign y17954 = ~1'b0 ;
  assign y17955 = n33629 ;
  assign y17956 = ~n33630 ;
  assign y17957 = ~n33631 ;
  assign y17958 = ~n33634 ;
  assign y17959 = ~n33640 ;
  assign y17960 = n33641 ;
  assign y17961 = ~1'b0 ;
  assign y17962 = ~n33642 ;
  assign y17963 = n33644 ;
  assign y17964 = n33646 ;
  assign y17965 = ~n9957 ;
  assign y17966 = n33650 ;
  assign y17967 = ~n33652 ;
  assign y17968 = ~n20282 ;
  assign y17969 = n8220 ;
  assign y17970 = n33671 ;
  assign y17971 = n33672 ;
  assign y17972 = n33673 ;
  assign y17973 = ~1'b0 ;
  assign y17974 = ~1'b0 ;
  assign y17975 = n33676 ;
  assign y17976 = ~n33678 ;
  assign y17977 = n33680 ;
  assign y17978 = ~n33681 ;
  assign y17979 = ~n33683 ;
  assign y17980 = n33684 ;
  assign y17981 = ~n33686 ;
  assign y17982 = ~n33690 ;
  assign y17983 = ~1'b0 ;
  assign y17984 = n33692 ;
  assign y17985 = ~1'b0 ;
  assign y17986 = 1'b0 ;
  assign y17987 = n33693 ;
  assign y17988 = ~n33694 ;
  assign y17989 = ~1'b0 ;
  assign y17990 = ~n33699 ;
  assign y17991 = n33700 ;
  assign y17992 = ~1'b0 ;
  assign y17993 = ~n1364 ;
  assign y17994 = ~n33701 ;
  assign y17995 = n3114 ;
  assign y17996 = n33703 ;
  assign y17997 = ~n33706 ;
  assign y17998 = n13657 ;
  assign y17999 = ~n18092 ;
  assign y18000 = n33707 ;
  assign y18001 = n33717 ;
  assign y18002 = ~1'b0 ;
  assign y18003 = ~1'b0 ;
  assign y18004 = n33719 ;
  assign y18005 = ~1'b0 ;
  assign y18006 = n33720 ;
  assign y18007 = n33721 ;
  assign y18008 = ~n33723 ;
  assign y18009 = n2550 ;
  assign y18010 = ~1'b0 ;
  assign y18011 = ~n33727 ;
  assign y18012 = ~n33729 ;
  assign y18013 = n33732 ;
  assign y18014 = n33734 ;
  assign y18015 = n33736 ;
  assign y18016 = ~1'b0 ;
  assign y18017 = ~n33737 ;
  assign y18018 = ~n33740 ;
  assign y18019 = ~n33741 ;
  assign y18020 = n33743 ;
  assign y18021 = ~1'b0 ;
  assign y18022 = n33744 ;
  assign y18023 = ~1'b0 ;
  assign y18024 = n33745 ;
  assign y18025 = ~n33751 ;
  assign y18026 = ~1'b0 ;
  assign y18027 = ~n33759 ;
  assign y18028 = ~n33762 ;
  assign y18029 = ~1'b0 ;
  assign y18030 = ~n33763 ;
  assign y18031 = ~n33766 ;
  assign y18032 = ~n33768 ;
  assign y18033 = ~n33773 ;
  assign y18034 = ~n33774 ;
  assign y18035 = ~1'b0 ;
  assign y18036 = ~n33778 ;
  assign y18037 = ~1'b0 ;
  assign y18038 = ~n33781 ;
  assign y18039 = ~n10608 ;
  assign y18040 = n33783 ;
  assign y18041 = 1'b0 ;
  assign y18042 = n33786 ;
  assign y18043 = n33787 ;
  assign y18044 = ~n33790 ;
  assign y18045 = n33791 ;
  assign y18046 = n33792 ;
  assign y18047 = ~n948 ;
  assign y18048 = ~n33794 ;
  assign y18049 = n33798 ;
  assign y18050 = ~1'b0 ;
  assign y18051 = n33799 ;
  assign y18052 = ~n33804 ;
  assign y18053 = ~n33807 ;
  assign y18054 = ~1'b0 ;
  assign y18055 = n33810 ;
  assign y18056 = ~1'b0 ;
  assign y18057 = ~1'b0 ;
  assign y18058 = n33811 ;
  assign y18059 = ~n33813 ;
  assign y18060 = n33814 ;
  assign y18061 = ~n33816 ;
  assign y18062 = ~n33819 ;
  assign y18063 = ~n33822 ;
  assign y18064 = ~1'b0 ;
  assign y18065 = ~n33825 ;
  assign y18066 = ~n33826 ;
  assign y18067 = ~1'b0 ;
  assign y18068 = ~n33829 ;
  assign y18069 = ~n33836 ;
  assign y18070 = ~1'b0 ;
  assign y18071 = ~1'b0 ;
  assign y18072 = ~n33837 ;
  assign y18073 = ~n33838 ;
  assign y18074 = ~n33844 ;
  assign y18075 = ~n33848 ;
  assign y18076 = n33851 ;
  assign y18077 = ~1'b0 ;
  assign y18078 = ~n33854 ;
  assign y18079 = ~1'b0 ;
  assign y18080 = ~1'b0 ;
  assign y18081 = ~1'b0 ;
  assign y18082 = ~n33857 ;
  assign y18083 = ~n33861 ;
  assign y18084 = ~n33862 ;
  assign y18085 = n33864 ;
  assign y18086 = ~n33865 ;
  assign y18087 = ~n33874 ;
  assign y18088 = 1'b0 ;
  assign y18089 = n33877 ;
  assign y18090 = n33880 ;
  assign y18091 = ~1'b0 ;
  assign y18092 = ~n33882 ;
  assign y18093 = ~n33883 ;
  assign y18094 = n6243 ;
  assign y18095 = ~1'b0 ;
  assign y18096 = ~n6986 ;
  assign y18097 = n33886 ;
  assign y18098 = n33888 ;
  assign y18099 = n33889 ;
  assign y18100 = n33890 ;
  assign y18101 = 1'b0 ;
  assign y18102 = n19916 ;
  assign y18103 = ~1'b0 ;
  assign y18104 = ~n33895 ;
  assign y18105 = ~n33899 ;
  assign y18106 = ~n33902 ;
  assign y18107 = ~n33911 ;
  assign y18108 = n33914 ;
  assign y18109 = ~1'b0 ;
  assign y18110 = ~n33915 ;
  assign y18111 = ~n33916 ;
  assign y18112 = 1'b0 ;
  assign y18113 = n33919 ;
  assign y18114 = ~1'b0 ;
  assign y18115 = ~n33920 ;
  assign y18116 = n33921 ;
  assign y18117 = n13121 ;
  assign y18118 = 1'b0 ;
  assign y18119 = n33925 ;
  assign y18120 = ~n464 ;
  assign y18121 = ~1'b0 ;
  assign y18122 = n33928 ;
  assign y18123 = ~n33191 ;
  assign y18124 = n33929 ;
  assign y18125 = n33932 ;
  assign y18126 = n2439 ;
  assign y18127 = n33933 ;
  assign y18128 = ~n33936 ;
  assign y18129 = ~n33939 ;
  assign y18130 = ~1'b0 ;
  assign y18131 = ~n16739 ;
  assign y18132 = ~n33942 ;
  assign y18133 = ~n2189 ;
  assign y18134 = n33945 ;
  assign y18135 = n18934 ;
  assign y18136 = ~1'b0 ;
  assign y18137 = ~n33948 ;
  assign y18138 = n33951 ;
  assign y18139 = ~1'b0 ;
  assign y18140 = ~1'b0 ;
  assign y18141 = ~1'b0 ;
  assign y18142 = n33953 ;
  assign y18143 = n33954 ;
  assign y18144 = ~n33959 ;
  assign y18145 = n33963 ;
  assign y18146 = ~n33969 ;
  assign y18147 = n33973 ;
  assign y18148 = ~n33977 ;
  assign y18149 = ~1'b0 ;
  assign y18150 = n33980 ;
  assign y18151 = n33982 ;
  assign y18152 = ~n33985 ;
  assign y18153 = n19757 ;
  assign y18154 = ~n33988 ;
  assign y18155 = 1'b0 ;
  assign y18156 = ~1'b0 ;
  assign y18157 = ~n16402 ;
  assign y18158 = n33991 ;
  assign y18159 = ~1'b0 ;
  assign y18160 = ~n33992 ;
  assign y18161 = n33994 ;
  assign y18162 = ~n33998 ;
  assign y18163 = n7584 ;
  assign y18164 = ~1'b0 ;
  assign y18165 = n34002 ;
  assign y18166 = ~1'b0 ;
  assign y18167 = ~n34006 ;
  assign y18168 = ~1'b0 ;
  assign y18169 = ~n34008 ;
  assign y18170 = ~1'b0 ;
  assign y18171 = ~n20619 ;
  assign y18172 = ~1'b0 ;
  assign y18173 = n34014 ;
  assign y18174 = ~n16037 ;
  assign y18175 = 1'b0 ;
  assign y18176 = ~n34015 ;
  assign y18177 = ~1'b0 ;
  assign y18178 = n34016 ;
  assign y18179 = n34017 ;
  assign y18180 = n26315 ;
  assign y18181 = n34019 ;
  assign y18182 = ~1'b0 ;
  assign y18183 = ~1'b0 ;
  assign y18184 = ~1'b0 ;
  assign y18185 = ~1'b0 ;
  assign y18186 = n34020 ;
  assign y18187 = ~n13490 ;
  assign y18188 = ~1'b0 ;
  assign y18189 = n34021 ;
  assign y18190 = n34029 ;
  assign y18191 = n34030 ;
  assign y18192 = ~1'b0 ;
  assign y18193 = n34032 ;
  assign y18194 = ~n34036 ;
  assign y18195 = ~1'b0 ;
  assign y18196 = ~n34037 ;
  assign y18197 = n34038 ;
  assign y18198 = ~1'b0 ;
  assign y18199 = ~n34040 ;
  assign y18200 = ~n27847 ;
  assign y18201 = n34042 ;
  assign y18202 = n25031 ;
  assign y18203 = ~n17877 ;
  assign y18204 = ~n34045 ;
  assign y18205 = ~1'b0 ;
  assign y18206 = ~n34046 ;
  assign y18207 = 1'b0 ;
  assign y18208 = 1'b0 ;
  assign y18209 = ~n34048 ;
  assign y18210 = ~1'b0 ;
  assign y18211 = n19888 ;
  assign y18212 = ~1'b0 ;
  assign y18213 = ~1'b0 ;
  assign y18214 = ~n34050 ;
  assign y18215 = ~n34053 ;
  assign y18216 = ~n7863 ;
  assign y18217 = ~1'b0 ;
  assign y18218 = ~1'b0 ;
  assign y18219 = ~n34059 ;
  assign y18220 = ~1'b0 ;
  assign y18221 = ~n34060 ;
  assign y18222 = ~n34062 ;
  assign y18223 = n34063 ;
  assign y18224 = n34065 ;
  assign y18225 = ~n33189 ;
  assign y18226 = n8513 ;
  assign y18227 = ~1'b0 ;
  assign y18228 = ~n34067 ;
  assign y18229 = ~1'b0 ;
  assign y18230 = ~n34074 ;
  assign y18231 = n28292 ;
  assign y18232 = ~n34077 ;
  assign y18233 = ~1'b0 ;
  assign y18234 = n34078 ;
  assign y18235 = ~n34080 ;
  assign y18236 = ~1'b0 ;
  assign y18237 = ~n34082 ;
  assign y18238 = n34084 ;
  assign y18239 = ~n34086 ;
  assign y18240 = ~1'b0 ;
  assign y18241 = ~n34087 ;
  assign y18242 = ~1'b0 ;
  assign y18243 = n34089 ;
  assign y18244 = ~1'b0 ;
  assign y18245 = ~n34091 ;
  assign y18246 = ~1'b0 ;
  assign y18247 = ~n5072 ;
  assign y18248 = ~1'b0 ;
  assign y18249 = n34095 ;
  assign y18250 = n34098 ;
  assign y18251 = n34101 ;
  assign y18252 = ~1'b0 ;
  assign y18253 = 1'b0 ;
  assign y18254 = n34103 ;
  assign y18255 = n34104 ;
  assign y18256 = ~1'b0 ;
  assign y18257 = ~n34108 ;
  assign y18258 = n34109 ;
  assign y18259 = ~n34110 ;
  assign y18260 = n34111 ;
  assign y18261 = ~1'b0 ;
  assign y18262 = ~1'b0 ;
  assign y18263 = n34113 ;
  assign y18264 = n34114 ;
  assign y18265 = ~n34119 ;
  assign y18266 = n32337 ;
  assign y18267 = n34121 ;
  assign y18268 = n34122 ;
  assign y18269 = n34124 ;
  assign y18270 = n34125 ;
  assign y18271 = ~1'b0 ;
  assign y18272 = ~n34133 ;
  assign y18273 = ~1'b0 ;
  assign y18274 = n34135 ;
  assign y18275 = ~n34141 ;
  assign y18276 = ~n34142 ;
  assign y18277 = n34150 ;
  assign y18278 = ~n1525 ;
  assign y18279 = ~n34152 ;
  assign y18280 = ~n34154 ;
  assign y18281 = ~n34156 ;
  assign y18282 = ~n34158 ;
  assign y18283 = ~n34159 ;
  assign y18284 = ~n34163 ;
  assign y18285 = ~1'b0 ;
  assign y18286 = n34165 ;
  assign y18287 = ~n34170 ;
  assign y18288 = n34173 ;
  assign y18289 = n34174 ;
  assign y18290 = ~n34177 ;
  assign y18291 = n34178 ;
  assign y18292 = ~1'b0 ;
  assign y18293 = ~n34179 ;
  assign y18294 = ~n34180 ;
  assign y18295 = n34183 ;
  assign y18296 = n34187 ;
  assign y18297 = ~n34189 ;
  assign y18298 = n34193 ;
  assign y18299 = n34198 ;
  assign y18300 = n34200 ;
  assign y18301 = n7203 ;
  assign y18302 = ~n34201 ;
  assign y18303 = ~n34202 ;
  assign y18304 = n34205 ;
  assign y18305 = ~1'b0 ;
  assign y18306 = ~n34206 ;
  assign y18307 = n34208 ;
  assign y18308 = ~n29031 ;
  assign y18309 = ~1'b0 ;
  assign y18310 = ~1'b0 ;
  assign y18311 = n34209 ;
  assign y18312 = n34210 ;
  assign y18313 = n34214 ;
  assign y18314 = n34217 ;
  assign y18315 = ~n34219 ;
  assign y18316 = n34224 ;
  assign y18317 = n34225 ;
  assign y18318 = n34234 ;
  assign y18319 = n34238 ;
  assign y18320 = n34242 ;
  assign y18321 = ~1'b0 ;
  assign y18322 = ~n34244 ;
  assign y18323 = ~n34247 ;
  assign y18324 = n34248 ;
  assign y18325 = 1'b0 ;
  assign y18326 = n34249 ;
  assign y18327 = ~n34251 ;
  assign y18328 = n34252 ;
  assign y18329 = ~1'b0 ;
  assign y18330 = n13838 ;
  assign y18331 = ~n34253 ;
  assign y18332 = ~1'b0 ;
  assign y18333 = n34254 ;
  assign y18334 = n34255 ;
  assign y18335 = ~1'b0 ;
  assign y18336 = ~1'b0 ;
  assign y18337 = ~n34259 ;
  assign y18338 = ~1'b0 ;
  assign y18339 = ~1'b0 ;
  assign y18340 = ~n34264 ;
  assign y18341 = ~n18948 ;
  assign y18342 = ~1'b0 ;
  assign y18343 = n34267 ;
  assign y18344 = ~n34271 ;
  assign y18345 = ~n34274 ;
  assign y18346 = n34276 ;
  assign y18347 = n34280 ;
  assign y18348 = n34283 ;
  assign y18349 = ~1'b0 ;
  assign y18350 = n34286 ;
  assign y18351 = ~n34288 ;
  assign y18352 = n34293 ;
  assign y18353 = n34294 ;
  assign y18354 = ~n34295 ;
  assign y18355 = ~n34300 ;
  assign y18356 = ~1'b0 ;
  assign y18357 = ~n34301 ;
  assign y18358 = ~n34304 ;
  assign y18359 = n34308 ;
  assign y18360 = n34309 ;
  assign y18361 = ~n1377 ;
  assign y18362 = ~n34310 ;
  assign y18363 = n19318 ;
  assign y18364 = ~n34312 ;
  assign y18365 = n34315 ;
  assign y18366 = n34320 ;
  assign y18367 = ~n34321 ;
  assign y18368 = 1'b0 ;
  assign y18369 = n34323 ;
  assign y18370 = n34326 ;
  assign y18371 = n34329 ;
  assign y18372 = ~1'b0 ;
  assign y18373 = ~1'b0 ;
  assign y18374 = n34331 ;
  assign y18375 = n34337 ;
  assign y18376 = n3628 ;
  assign y18377 = ~1'b0 ;
  assign y18378 = n34338 ;
  assign y18379 = ~1'b0 ;
  assign y18380 = ~1'b0 ;
  assign y18381 = ~n34342 ;
  assign y18382 = ~1'b0 ;
  assign y18383 = ~n34343 ;
  assign y18384 = n34345 ;
  assign y18385 = n34346 ;
  assign y18386 = ~n34348 ;
  assign y18387 = n34349 ;
  assign y18388 = n34350 ;
  assign y18389 = ~1'b0 ;
  assign y18390 = n34360 ;
  assign y18391 = n34362 ;
  assign y18392 = n34364 ;
  assign y18393 = n34366 ;
  assign y18394 = n34367 ;
  assign y18395 = ~1'b0 ;
  assign y18396 = ~n34369 ;
  assign y18397 = ~n34370 ;
  assign y18398 = ~1'b0 ;
  assign y18399 = ~n34371 ;
  assign y18400 = ~n34374 ;
  assign y18401 = ~n34377 ;
  assign y18402 = ~1'b0 ;
  assign y18403 = ~1'b0 ;
  assign y18404 = ~1'b0 ;
  assign y18405 = ~1'b0 ;
  assign y18406 = n34379 ;
  assign y18407 = n34381 ;
  assign y18408 = ~1'b0 ;
  assign y18409 = ~1'b0 ;
  assign y18410 = n5392 ;
  assign y18411 = n34384 ;
  assign y18412 = ~1'b0 ;
  assign y18413 = ~n34385 ;
  assign y18414 = ~n34386 ;
  assign y18415 = n34388 ;
  assign y18416 = ~n34390 ;
  assign y18417 = ~1'b0 ;
  assign y18418 = ~n34391 ;
  assign y18419 = n34392 ;
  assign y18420 = ~n34396 ;
  assign y18421 = 1'b0 ;
  assign y18422 = ~1'b0 ;
  assign y18423 = n34397 ;
  assign y18424 = ~1'b0 ;
  assign y18425 = ~1'b0 ;
  assign y18426 = ~n34399 ;
  assign y18427 = ~n31044 ;
  assign y18428 = n34400 ;
  assign y18429 = ~1'b0 ;
  assign y18430 = ~1'b0 ;
  assign y18431 = n34401 ;
  assign y18432 = ~n34402 ;
  assign y18433 = ~1'b0 ;
  assign y18434 = 1'b0 ;
  assign y18435 = ~1'b0 ;
  assign y18436 = ~n34404 ;
  assign y18437 = ~n34405 ;
  assign y18438 = n5726 ;
  assign y18439 = n34407 ;
  assign y18440 = ~1'b0 ;
  assign y18441 = ~n34410 ;
  assign y18442 = ~1'b0 ;
  assign y18443 = ~1'b0 ;
  assign y18444 = n34413 ;
  assign y18445 = ~n34414 ;
  assign y18446 = n34421 ;
  assign y18447 = n34422 ;
  assign y18448 = n34423 ;
  assign y18449 = ~n34425 ;
  assign y18450 = ~n34431 ;
  assign y18451 = ~n34435 ;
  assign y18452 = ~1'b0 ;
  assign y18453 = ~n34438 ;
  assign y18454 = n34440 ;
  assign y18455 = n28999 ;
  assign y18456 = ~n31743 ;
  assign y18457 = ~n34441 ;
  assign y18458 = ~1'b0 ;
  assign y18459 = n34443 ;
  assign y18460 = n34446 ;
  assign y18461 = ~1'b0 ;
  assign y18462 = ~n34447 ;
  assign y18463 = ~1'b0 ;
  assign y18464 = n34449 ;
  assign y18465 = ~n34453 ;
  assign y18466 = ~1'b0 ;
  assign y18467 = ~n10211 ;
  assign y18468 = ~1'b0 ;
  assign y18469 = ~n34454 ;
  assign y18470 = ~n34459 ;
  assign y18471 = ~1'b0 ;
  assign y18472 = n34462 ;
  assign y18473 = ~n34463 ;
  assign y18474 = ~1'b0 ;
  assign y18475 = ~1'b0 ;
  assign y18476 = n34472 ;
  assign y18477 = ~1'b0 ;
  assign y18478 = n34473 ;
  assign y18479 = ~n34476 ;
  assign y18480 = n34478 ;
  assign y18481 = n34480 ;
  assign y18482 = ~n34488 ;
  assign y18483 = ~1'b0 ;
  assign y18484 = ~n679 ;
  assign y18485 = ~n34489 ;
  assign y18486 = ~n34492 ;
  assign y18487 = ~n9110 ;
  assign y18488 = n34493 ;
  assign y18489 = ~1'b0 ;
  assign y18490 = ~n34498 ;
  assign y18491 = ~1'b0 ;
  assign y18492 = n34505 ;
  assign y18493 = 1'b0 ;
  assign y18494 = ~n34508 ;
  assign y18495 = ~1'b0 ;
  assign y18496 = ~1'b0 ;
  assign y18497 = ~n34512 ;
  assign y18498 = n34516 ;
  assign y18499 = ~1'b0 ;
  assign y18500 = ~n34519 ;
  assign y18501 = n34521 ;
  assign y18502 = n34524 ;
  assign y18503 = n34526 ;
  assign y18504 = ~1'b0 ;
  assign y18505 = ~n34528 ;
  assign y18506 = ~n13003 ;
  assign y18507 = ~n34529 ;
  assign y18508 = n34530 ;
  assign y18509 = n34533 ;
  assign y18510 = n34534 ;
  assign y18511 = ~n34536 ;
  assign y18512 = ~1'b0 ;
  assign y18513 = n34537 ;
  assign y18514 = ~n34538 ;
  assign y18515 = ~1'b0 ;
  assign y18516 = ~n34539 ;
  assign y18517 = n34540 ;
  assign y18518 = ~1'b0 ;
  assign y18519 = ~n34542 ;
  assign y18520 = n34544 ;
  assign y18521 = n34546 ;
  assign y18522 = n34551 ;
  assign y18523 = ~1'b0 ;
  assign y18524 = n34555 ;
  assign y18525 = n34558 ;
  assign y18526 = n34560 ;
  assign y18527 = ~1'b0 ;
  assign y18528 = ~n34563 ;
  assign y18529 = ~n34564 ;
  assign y18530 = 1'b0 ;
  assign y18531 = ~1'b0 ;
  assign y18532 = n34567 ;
  assign y18533 = n34569 ;
  assign y18534 = n34570 ;
  assign y18535 = ~n34572 ;
  assign y18536 = ~1'b0 ;
  assign y18537 = ~n34577 ;
  assign y18538 = n34578 ;
  assign y18539 = ~n34583 ;
  assign y18540 = ~n34587 ;
  assign y18541 = n34588 ;
  assign y18542 = n34589 ;
  assign y18543 = n34591 ;
  assign y18544 = n34594 ;
  assign y18545 = ~n31777 ;
  assign y18546 = ~n34595 ;
  assign y18547 = ~n34596 ;
  assign y18548 = n34600 ;
  assign y18549 = n34601 ;
  assign y18550 = n34602 ;
  assign y18551 = n32935 ;
  assign y18552 = ~n34603 ;
  assign y18553 = ~n34605 ;
  assign y18554 = n34607 ;
  assign y18555 = n18894 ;
  assign y18556 = ~n34608 ;
  assign y18557 = ~1'b0 ;
  assign y18558 = ~n34609 ;
  assign y18559 = n34610 ;
  assign y18560 = ~1'b0 ;
  assign y18561 = ~1'b0 ;
  assign y18562 = ~n34616 ;
  assign y18563 = n34617 ;
  assign y18564 = ~n34618 ;
  assign y18565 = ~n34619 ;
  assign y18566 = ~n34620 ;
  assign y18567 = n34623 ;
  assign y18568 = ~n34624 ;
  assign y18569 = n34625 ;
  assign y18570 = ~n34629 ;
  assign y18571 = ~1'b0 ;
  assign y18572 = ~n34630 ;
  assign y18573 = ~1'b0 ;
  assign y18574 = ~1'b0 ;
  assign y18575 = n34631 ;
  assign y18576 = n23852 ;
  assign y18577 = ~n34632 ;
  assign y18578 = ~n34635 ;
  assign y18579 = n34636 ;
  assign y18580 = n34639 ;
  assign y18581 = n34642 ;
  assign y18582 = n34644 ;
  assign y18583 = ~1'b0 ;
  assign y18584 = ~n34646 ;
  assign y18585 = ~1'b0 ;
  assign y18586 = n34647 ;
  assign y18587 = ~n34649 ;
  assign y18588 = ~1'b0 ;
  assign y18589 = n34651 ;
  assign y18590 = ~n34653 ;
  assign y18591 = ~n34655 ;
  assign y18592 = n17694 ;
  assign y18593 = n34656 ;
  assign y18594 = ~1'b0 ;
  assign y18595 = n34659 ;
  assign y18596 = ~1'b0 ;
  assign y18597 = ~n34661 ;
  assign y18598 = n34664 ;
  assign y18599 = ~n34666 ;
  assign y18600 = ~n34673 ;
  assign y18601 = ~n34675 ;
  assign y18602 = ~n34679 ;
  assign y18603 = n34680 ;
  assign y18604 = ~1'b0 ;
  assign y18605 = ~n34686 ;
  assign y18606 = n34688 ;
  assign y18607 = ~1'b0 ;
  assign y18608 = ~1'b0 ;
  assign y18609 = ~n34690 ;
  assign y18610 = 1'b0 ;
  assign y18611 = n34693 ;
  assign y18612 = ~n34694 ;
  assign y18613 = n34695 ;
  assign y18614 = ~1'b0 ;
  assign y18615 = n34698 ;
  assign y18616 = n34701 ;
  assign y18617 = n34703 ;
  assign y18618 = n34704 ;
  assign y18619 = ~1'b0 ;
  assign y18620 = ~1'b0 ;
  assign y18621 = n34705 ;
  assign y18622 = n34707 ;
  assign y18623 = n34709 ;
  assign y18624 = n34710 ;
  assign y18625 = ~n27787 ;
  assign y18626 = ~n34714 ;
  assign y18627 = ~1'b0 ;
  assign y18628 = n34715 ;
  assign y18629 = n34716 ;
  assign y18630 = ~n34720 ;
  assign y18631 = n34723 ;
  assign y18632 = n34724 ;
  assign y18633 = ~n34725 ;
  assign y18634 = n34730 ;
  assign y18635 = ~n34733 ;
  assign y18636 = ~1'b0 ;
  assign y18637 = ~n34736 ;
  assign y18638 = ~1'b0 ;
  assign y18639 = ~n34737 ;
  assign y18640 = n34742 ;
  assign y18641 = ~n29523 ;
  assign y18642 = ~n34744 ;
  assign y18643 = ~1'b0 ;
  assign y18644 = n34745 ;
  assign y18645 = ~n34750 ;
  assign y18646 = n34752 ;
  assign y18647 = n34753 ;
  assign y18648 = ~n16532 ;
  assign y18649 = n34754 ;
  assign y18650 = n34758 ;
  assign y18651 = ~n34762 ;
  assign y18652 = ~1'b0 ;
  assign y18653 = ~1'b0 ;
  assign y18654 = ~1'b0 ;
  assign y18655 = ~n34763 ;
  assign y18656 = ~n34765 ;
  assign y18657 = ~1'b0 ;
  assign y18658 = ~1'b0 ;
  assign y18659 = ~1'b0 ;
  assign y18660 = ~1'b0 ;
  assign y18661 = ~n34768 ;
  assign y18662 = ~1'b0 ;
  assign y18663 = n34769 ;
  assign y18664 = ~n34773 ;
  assign y18665 = n34774 ;
  assign y18666 = ~n34780 ;
  assign y18667 = ~n34786 ;
  assign y18668 = ~1'b0 ;
  assign y18669 = n34788 ;
  assign y18670 = ~1'b0 ;
  assign y18671 = ~n34790 ;
  assign y18672 = n34791 ;
  assign y18673 = ~1'b0 ;
  assign y18674 = ~n34792 ;
  assign y18675 = ~1'b0 ;
  assign y18676 = n34795 ;
  assign y18677 = n34797 ;
  assign y18678 = n34799 ;
  assign y18679 = ~1'b0 ;
  assign y18680 = n1674 ;
  assign y18681 = ~1'b0 ;
  assign y18682 = ~n34800 ;
  assign y18683 = ~n34802 ;
  assign y18684 = ~n34808 ;
  assign y18685 = n34813 ;
  assign y18686 = ~n7516 ;
  assign y18687 = ~1'b0 ;
  assign y18688 = ~n34816 ;
  assign y18689 = ~n34818 ;
  assign y18690 = n34822 ;
  assign y18691 = n34823 ;
  assign y18692 = 1'b0 ;
  assign y18693 = n3087 ;
  assign y18694 = ~1'b0 ;
  assign y18695 = n34825 ;
  assign y18696 = n34826 ;
  assign y18697 = ~1'b0 ;
  assign y18698 = ~1'b0 ;
  assign y18699 = n26212 ;
  assign y18700 = ~n34827 ;
  assign y18701 = n34831 ;
  assign y18702 = n34835 ;
  assign y18703 = ~n34836 ;
  assign y18704 = ~1'b0 ;
  assign y18705 = ~1'b0 ;
  assign y18706 = ~n34841 ;
  assign y18707 = ~n34844 ;
  assign y18708 = ~n34848 ;
  assign y18709 = ~n34851 ;
  assign y18710 = ~1'b0 ;
  assign y18711 = ~n34852 ;
  assign y18712 = ~n34853 ;
  assign y18713 = n34855 ;
  assign y18714 = n34858 ;
  assign y18715 = ~n34859 ;
  assign y18716 = n34863 ;
  assign y18717 = n34864 ;
  assign y18718 = ~1'b0 ;
  assign y18719 = ~1'b0 ;
  assign y18720 = ~n34865 ;
  assign y18721 = ~n34866 ;
  assign y18722 = ~n34868 ;
  assign y18723 = n34870 ;
  assign y18724 = n34873 ;
  assign y18725 = ~n34877 ;
  assign y18726 = ~1'b0 ;
  assign y18727 = n29639 ;
  assign y18728 = ~n34884 ;
  assign y18729 = n34888 ;
  assign y18730 = n5519 ;
  assign y18731 = ~n34890 ;
  assign y18732 = ~n34891 ;
  assign y18733 = ~n34893 ;
  assign y18734 = n34895 ;
  assign y18735 = ~1'b0 ;
  assign y18736 = ~n34900 ;
  assign y18737 = ~1'b0 ;
  assign y18738 = ~1'b0 ;
  assign y18739 = ~n34901 ;
  assign y18740 = n34907 ;
  assign y18741 = ~1'b0 ;
  assign y18742 = n34908 ;
  assign y18743 = 1'b0 ;
  assign y18744 = n34911 ;
  assign y18745 = ~n34913 ;
  assign y18746 = ~1'b0 ;
  assign y18747 = n34915 ;
  assign y18748 = n34917 ;
  assign y18749 = ~1'b0 ;
  assign y18750 = ~1'b0 ;
  assign y18751 = ~n34918 ;
  assign y18752 = n34920 ;
  assign y18753 = ~1'b0 ;
  assign y18754 = ~n17910 ;
  assign y18755 = n3312 ;
  assign y18756 = n34921 ;
  assign y18757 = n34922 ;
  assign y18758 = ~n34924 ;
  assign y18759 = ~1'b0 ;
  assign y18760 = ~1'b0 ;
  assign y18761 = n34928 ;
  assign y18762 = ~n34931 ;
  assign y18763 = ~n34934 ;
  assign y18764 = ~n34935 ;
  assign y18765 = ~n34947 ;
  assign y18766 = ~1'b0 ;
  assign y18767 = ~1'b0 ;
  assign y18768 = ~n34954 ;
  assign y18769 = ~n34955 ;
  assign y18770 = n34956 ;
  assign y18771 = ~1'b0 ;
  assign y18772 = n34958 ;
  assign y18773 = ~n34963 ;
  assign y18774 = ~n34967 ;
  assign y18775 = n2265 ;
  assign y18776 = ~n34968 ;
  assign y18777 = ~n34971 ;
  assign y18778 = ~1'b0 ;
  assign y18779 = ~n34973 ;
  assign y18780 = ~n34974 ;
  assign y18781 = ~n34976 ;
  assign y18782 = x91 ;
  assign y18783 = ~1'b0 ;
  assign y18784 = ~n11772 ;
  assign y18785 = ~n34977 ;
  assign y18786 = n34978 ;
  assign y18787 = n16085 ;
  assign y18788 = n34979 ;
  assign y18789 = n34981 ;
  assign y18790 = ~1'b0 ;
  assign y18791 = ~1'b0 ;
  assign y18792 = ~n34983 ;
  assign y18793 = ~1'b0 ;
  assign y18794 = ~n34987 ;
  assign y18795 = ~n34988 ;
  assign y18796 = ~1'b0 ;
  assign y18797 = n34990 ;
  assign y18798 = ~1'b0 ;
  assign y18799 = ~n3372 ;
  assign y18800 = ~1'b0 ;
  assign y18801 = ~1'b0 ;
  assign y18802 = ~n34994 ;
  assign y18803 = n35000 ;
  assign y18804 = ~n35002 ;
  assign y18805 = n9673 ;
  assign y18806 = n35003 ;
  assign y18807 = ~n35005 ;
  assign y18808 = ~1'b0 ;
  assign y18809 = n35008 ;
  assign y18810 = n35010 ;
  assign y18811 = ~n7863 ;
  assign y18812 = ~n35011 ;
  assign y18813 = n35013 ;
  assign y18814 = n35018 ;
  assign y18815 = ~1'b0 ;
  assign y18816 = ~1'b0 ;
  assign y18817 = n35021 ;
  assign y18818 = ~1'b0 ;
  assign y18819 = n35024 ;
  assign y18820 = ~n35026 ;
  assign y18821 = 1'b0 ;
  assign y18822 = ~n35028 ;
  assign y18823 = ~n35032 ;
  assign y18824 = ~1'b0 ;
  assign y18825 = n35034 ;
  assign y18826 = ~1'b0 ;
  assign y18827 = ~1'b0 ;
  assign y18828 = ~n35036 ;
  assign y18829 = ~1'b0 ;
  assign y18830 = n35038 ;
  assign y18831 = n35043 ;
  assign y18832 = 1'b0 ;
  assign y18833 = ~n9702 ;
  assign y18834 = n35045 ;
  assign y18835 = ~1'b0 ;
  assign y18836 = ~1'b0 ;
  assign y18837 = ~1'b0 ;
  assign y18838 = n35047 ;
  assign y18839 = ~1'b0 ;
  assign y18840 = ~n35051 ;
  assign y18841 = ~n35053 ;
  assign y18842 = n35055 ;
  assign y18843 = ~n35056 ;
  assign y18844 = ~n35057 ;
  assign y18845 = ~1'b0 ;
  assign y18846 = ~1'b0 ;
  assign y18847 = n35060 ;
  assign y18848 = ~1'b0 ;
  assign y18849 = ~n35065 ;
  assign y18850 = n35067 ;
  assign y18851 = ~1'b0 ;
  assign y18852 = ~1'b0 ;
  assign y18853 = ~n35069 ;
  assign y18854 = ~1'b0 ;
  assign y18855 = ~1'b0 ;
  assign y18856 = n35071 ;
  assign y18857 = ~n35073 ;
  assign y18858 = ~n35076 ;
  assign y18859 = ~1'b0 ;
  assign y18860 = ~n35077 ;
  assign y18861 = n35078 ;
  assign y18862 = ~1'b0 ;
  assign y18863 = ~1'b0 ;
  assign y18864 = ~1'b0 ;
  assign y18865 = ~n35079 ;
  assign y18866 = ~1'b0 ;
  assign y18867 = n35080 ;
  assign y18868 = n35081 ;
  assign y18869 = n35084 ;
  assign y18870 = ~n35088 ;
  assign y18871 = ~1'b0 ;
  assign y18872 = n35094 ;
  assign y18873 = n35095 ;
  assign y18874 = ~n35100 ;
  assign y18875 = ~1'b0 ;
  assign y18876 = n35102 ;
  assign y18877 = n35103 ;
  assign y18878 = ~1'b0 ;
  assign y18879 = ~n28489 ;
  assign y18880 = ~n35106 ;
  assign y18881 = ~1'b0 ;
  assign y18882 = ~1'b0 ;
  assign y18883 = 1'b0 ;
  assign y18884 = n35110 ;
  assign y18885 = n35111 ;
  assign y18886 = ~n35113 ;
  assign y18887 = n35117 ;
  assign y18888 = 1'b0 ;
  assign y18889 = ~1'b0 ;
  assign y18890 = n35119 ;
  assign y18891 = ~n35120 ;
  assign y18892 = ~1'b0 ;
  assign y18893 = n35123 ;
  assign y18894 = ~n35124 ;
  assign y18895 = ~1'b0 ;
  assign y18896 = ~1'b0 ;
  assign y18897 = ~n35125 ;
  assign y18898 = ~1'b0 ;
  assign y18899 = ~n35126 ;
  assign y18900 = ~n35128 ;
  assign y18901 = ~n7086 ;
  assign y18902 = n35135 ;
  assign y18903 = ~1'b0 ;
  assign y18904 = ~1'b0 ;
  assign y18905 = ~1'b0 ;
  assign y18906 = ~1'b0 ;
  assign y18907 = ~n35139 ;
  assign y18908 = n35142 ;
  assign y18909 = ~n35148 ;
  assign y18910 = n35150 ;
  assign y18911 = n35155 ;
  assign y18912 = ~n32829 ;
  assign y18913 = ~1'b0 ;
  assign y18914 = ~n35158 ;
  assign y18915 = ~x143 ;
  assign y18916 = ~n35159 ;
  assign y18917 = ~1'b0 ;
  assign y18918 = ~1'b0 ;
  assign y18919 = ~n35161 ;
  assign y18920 = ~1'b0 ;
  assign y18921 = ~1'b0 ;
  assign y18922 = n35163 ;
  assign y18923 = n35168 ;
  assign y18924 = ~1'b0 ;
  assign y18925 = ~n35173 ;
  assign y18926 = n35175 ;
  assign y18927 = n35176 ;
  assign y18928 = ~1'b0 ;
  assign y18929 = ~1'b0 ;
  assign y18930 = ~n35178 ;
  assign y18931 = ~n35184 ;
  assign y18932 = ~n35187 ;
  assign y18933 = n35190 ;
  assign y18934 = n34068 ;
  assign y18935 = ~1'b0 ;
  assign y18936 = ~1'b0 ;
  assign y18937 = n35192 ;
  assign y18938 = ~n35193 ;
  assign y18939 = ~n35197 ;
  assign y18940 = ~1'b0 ;
  assign y18941 = ~1'b0 ;
  assign y18942 = ~n35198 ;
  assign y18943 = ~n35199 ;
  assign y18944 = n35201 ;
  assign y18945 = ~1'b0 ;
  assign y18946 = n35202 ;
  assign y18947 = ~n6655 ;
  assign y18948 = ~1'b0 ;
  assign y18949 = ~n35203 ;
  assign y18950 = ~1'b0 ;
  assign y18951 = ~n35204 ;
  assign y18952 = ~1'b0 ;
  assign y18953 = n35206 ;
  assign y18954 = ~n35212 ;
  assign y18955 = ~1'b0 ;
  assign y18956 = n15176 ;
  assign y18957 = ~1'b0 ;
  assign y18958 = ~n35216 ;
  assign y18959 = ~n35223 ;
  assign y18960 = ~n35225 ;
  assign y18961 = ~n35227 ;
  assign y18962 = ~1'b0 ;
  assign y18963 = n26403 ;
  assign y18964 = n35230 ;
  assign y18965 = n30813 ;
  assign y18966 = ~n11852 ;
  assign y18967 = ~n35233 ;
  assign y18968 = n35234 ;
  assign y18969 = ~n6243 ;
  assign y18970 = ~n35237 ;
  assign y18971 = ~1'b0 ;
  assign y18972 = ~1'b0 ;
  assign y18973 = n35239 ;
  assign y18974 = n35240 ;
  assign y18975 = ~1'b0 ;
  assign y18976 = ~1'b0 ;
  assign y18977 = n35241 ;
  assign y18978 = ~1'b0 ;
  assign y18979 = ~n35243 ;
  assign y18980 = ~n23963 ;
  assign y18981 = ~n35245 ;
  assign y18982 = n35249 ;
  assign y18983 = ~1'b0 ;
  assign y18984 = n35253 ;
  assign y18985 = ~1'b0 ;
  assign y18986 = n35255 ;
  assign y18987 = n3155 ;
  assign y18988 = n35258 ;
  assign y18989 = ~n35261 ;
  assign y18990 = ~1'b0 ;
  assign y18991 = ~n35263 ;
  assign y18992 = ~n35266 ;
  assign y18993 = ~1'b0 ;
  assign y18994 = n35268 ;
  assign y18995 = ~n35272 ;
  assign y18996 = ~1'b0 ;
  assign y18997 = n35273 ;
  assign y18998 = ~n13037 ;
  assign y18999 = n35275 ;
  assign y19000 = ~n35282 ;
  assign y19001 = ~n26640 ;
  assign y19002 = ~1'b0 ;
  assign y19003 = ~1'b0 ;
  assign y19004 = n35287 ;
  assign y19005 = ~n35288 ;
  assign y19006 = ~n35289 ;
  assign y19007 = ~1'b0 ;
  assign y19008 = n35293 ;
  assign y19009 = n14635 ;
  assign y19010 = n35294 ;
  assign y19011 = ~1'b0 ;
  assign y19012 = ~n35296 ;
  assign y19013 = n18255 ;
  assign y19014 = n35297 ;
  assign y19015 = ~n35298 ;
  assign y19016 = ~1'b0 ;
  assign y19017 = ~n35300 ;
  assign y19018 = n35304 ;
  assign y19019 = n35312 ;
  assign y19020 = ~1'b0 ;
  assign y19021 = ~1'b0 ;
  assign y19022 = ~n35313 ;
  assign y19023 = ~n35314 ;
  assign y19024 = n35318 ;
  assign y19025 = ~1'b0 ;
  assign y19026 = n35319 ;
  assign y19027 = ~1'b0 ;
  assign y19028 = ~n35320 ;
  assign y19029 = ~1'b0 ;
  assign y19030 = ~1'b0 ;
  assign y19031 = ~n35324 ;
  assign y19032 = n35325 ;
  assign y19033 = ~n35330 ;
  assign y19034 = ~n35331 ;
  assign y19035 = n21741 ;
  assign y19036 = n35336 ;
  assign y19037 = n35337 ;
  assign y19038 = ~1'b0 ;
  assign y19039 = ~1'b0 ;
  assign y19040 = ~1'b0 ;
  assign y19041 = n35340 ;
  assign y19042 = n308 ;
  assign y19043 = ~1'b0 ;
  assign y19044 = ~1'b0 ;
  assign y19045 = 1'b0 ;
  assign y19046 = n35341 ;
  assign y19047 = ~n35345 ;
  assign y19048 = ~n35348 ;
  assign y19049 = n35349 ;
  assign y19050 = ~n35350 ;
  assign y19051 = n8488 ;
  assign y19052 = ~n35351 ;
  assign y19053 = ~1'b0 ;
  assign y19054 = ~1'b0 ;
  assign y19055 = ~n35354 ;
  assign y19056 = ~1'b0 ;
  assign y19057 = ~1'b0 ;
  assign y19058 = ~1'b0 ;
  assign y19059 = ~1'b0 ;
  assign y19060 = ~n2125 ;
  assign y19061 = ~n32025 ;
  assign y19062 = ~n35356 ;
  assign y19063 = n35359 ;
  assign y19064 = ~n35361 ;
  assign y19065 = ~1'b0 ;
  assign y19066 = ~1'b0 ;
  assign y19067 = n35363 ;
  assign y19068 = ~n906 ;
  assign y19069 = ~1'b0 ;
  assign y19070 = n35366 ;
  assign y19071 = n35367 ;
  assign y19072 = ~n35371 ;
  assign y19073 = ~1'b0 ;
  assign y19074 = ~1'b0 ;
  assign y19075 = ~n35373 ;
  assign y19076 = ~n35374 ;
  assign y19077 = n35377 ;
  assign y19078 = n2106 ;
  assign y19079 = ~n35378 ;
  assign y19080 = 1'b0 ;
  assign y19081 = ~n35379 ;
  assign y19082 = n35381 ;
  assign y19083 = ~1'b0 ;
  assign y19084 = ~1'b0 ;
  assign y19085 = n35382 ;
  assign y19086 = ~1'b0 ;
  assign y19087 = n35383 ;
  assign y19088 = n35384 ;
  assign y19089 = n35385 ;
  assign y19090 = n12879 ;
  assign y19091 = ~n35387 ;
  assign y19092 = ~n35389 ;
  assign y19093 = n35391 ;
  assign y19094 = n35393 ;
  assign y19095 = n35395 ;
  assign y19096 = ~n35398 ;
  assign y19097 = ~n35402 ;
  assign y19098 = ~n35408 ;
  assign y19099 = ~n35413 ;
  assign y19100 = ~n35416 ;
  assign y19101 = n35417 ;
  assign y19102 = ~n35421 ;
  assign y19103 = n35423 ;
  assign y19104 = 1'b0 ;
  assign y19105 = ~1'b0 ;
  assign y19106 = ~1'b0 ;
  assign y19107 = ~n35424 ;
  assign y19108 = n35425 ;
  assign y19109 = ~n7067 ;
  assign y19110 = ~n35429 ;
  assign y19111 = n35431 ;
  assign y19112 = n35432 ;
  assign y19113 = n35436 ;
  assign y19114 = ~n35438 ;
  assign y19115 = ~1'b0 ;
  assign y19116 = ~n35442 ;
  assign y19117 = n35447 ;
  assign y19118 = ~1'b0 ;
  assign y19119 = ~n35450 ;
  assign y19120 = ~n35452 ;
  assign y19121 = n35456 ;
  assign y19122 = ~n35459 ;
  assign y19123 = n35460 ;
  assign y19124 = n35461 ;
  assign y19125 = n35462 ;
  assign y19126 = n2406 ;
  assign y19127 = n35463 ;
  assign y19128 = ~n35466 ;
  assign y19129 = ~1'b0 ;
  assign y19130 = ~1'b0 ;
  assign y19131 = n11177 ;
  assign y19132 = ~1'b0 ;
  assign y19133 = ~1'b0 ;
  assign y19134 = ~n35467 ;
  assign y19135 = ~1'b0 ;
  assign y19136 = ~1'b0 ;
  assign y19137 = ~1'b0 ;
  assign y19138 = ~n35470 ;
  assign y19139 = n35471 ;
  assign y19140 = n35472 ;
  assign y19141 = n35473 ;
  assign y19142 = ~n35479 ;
  assign y19143 = ~n35483 ;
  assign y19144 = n35497 ;
  assign y19145 = ~1'b0 ;
  assign y19146 = n6851 ;
  assign y19147 = n35498 ;
  assign y19148 = ~n35500 ;
  assign y19149 = ~n29055 ;
  assign y19150 = ~n35502 ;
  assign y19151 = n35504 ;
  assign y19152 = ~1'b0 ;
  assign y19153 = ~1'b0 ;
  assign y19154 = ~n35505 ;
  assign y19155 = ~n35507 ;
  assign y19156 = ~n35511 ;
  assign y19157 = ~1'b0 ;
  assign y19158 = ~n35515 ;
  assign y19159 = ~1'b0 ;
  assign y19160 = ~n35516 ;
  assign y19161 = ~n31101 ;
  assign y19162 = ~n35522 ;
  assign y19163 = 1'b0 ;
  assign y19164 = ~n35525 ;
  assign y19165 = n35527 ;
  assign y19166 = n35528 ;
  assign y19167 = ~n35530 ;
  assign y19168 = ~1'b0 ;
  assign y19169 = ~n35533 ;
  assign y19170 = ~1'b0 ;
  assign y19171 = ~n35535 ;
  assign y19172 = ~n27355 ;
  assign y19173 = n35539 ;
  assign y19174 = ~n35540 ;
  assign y19175 = n35542 ;
  assign y19176 = ~n35543 ;
  assign y19177 = n35544 ;
  assign y19178 = ~1'b0 ;
  assign y19179 = ~1'b0 ;
  assign y19180 = ~1'b0 ;
  assign y19181 = ~n3670 ;
  assign y19182 = ~1'b0 ;
  assign y19183 = ~n35546 ;
  assign y19184 = ~n35550 ;
  assign y19185 = n35555 ;
  assign y19186 = ~n35556 ;
  assign y19187 = ~n35558 ;
  assign y19188 = ~1'b0 ;
  assign y19189 = ~1'b0 ;
  assign y19190 = n32918 ;
  assign y19191 = n35559 ;
  assign y19192 = ~n35564 ;
  assign y19193 = n35565 ;
  assign y19194 = n35566 ;
  assign y19195 = n35568 ;
  assign y19196 = ~1'b0 ;
  assign y19197 = ~1'b0 ;
  assign y19198 = n35569 ;
  assign y19199 = ~n35572 ;
  assign y19200 = n35575 ;
  assign y19201 = ~n35577 ;
  assign y19202 = n6655 ;
  assign y19203 = n35580 ;
  assign y19204 = n35581 ;
  assign y19205 = ~1'b0 ;
  assign y19206 = ~n35584 ;
  assign y19207 = n35586 ;
  assign y19208 = n35589 ;
  assign y19209 = ~1'b0 ;
  assign y19210 = ~1'b0 ;
  assign y19211 = n35593 ;
  assign y19212 = ~1'b0 ;
  assign y19213 = ~n35595 ;
  assign y19214 = ~n35597 ;
  assign y19215 = n35599 ;
  assign y19216 = ~1'b0 ;
  assign y19217 = ~1'b0 ;
  assign y19218 = ~n35602 ;
  assign y19219 = ~n35605 ;
  assign y19220 = ~n35607 ;
  assign y19221 = ~1'b0 ;
  assign y19222 = n35610 ;
  assign y19223 = ~n33496 ;
  assign y19224 = ~1'b0 ;
  assign y19225 = n35613 ;
  assign y19226 = ~1'b0 ;
  assign y19227 = n35615 ;
  assign y19228 = n35619 ;
  assign y19229 = ~1'b0 ;
  assign y19230 = ~n35622 ;
  assign y19231 = n35624 ;
  assign y19232 = ~1'b0 ;
  assign y19233 = n35627 ;
  assign y19234 = n35628 ;
  assign y19235 = n35629 ;
  assign y19236 = ~1'b0 ;
  assign y19237 = 1'b0 ;
  assign y19238 = ~1'b0 ;
  assign y19239 = ~1'b0 ;
  assign y19240 = ~1'b0 ;
  assign y19241 = n35631 ;
  assign y19242 = ~1'b0 ;
  assign y19243 = ~n35634 ;
  assign y19244 = ~1'b0 ;
  assign y19245 = n35635 ;
  assign y19246 = n35636 ;
  assign y19247 = n35638 ;
  assign y19248 = ~1'b0 ;
  assign y19249 = ~1'b0 ;
  assign y19250 = ~1'b0 ;
  assign y19251 = ~n35639 ;
  assign y19252 = ~n35643 ;
  assign y19253 = n35644 ;
  assign y19254 = n35646 ;
  assign y19255 = n35647 ;
  assign y19256 = ~1'b0 ;
  assign y19257 = n35649 ;
  assign y19258 = n35650 ;
  assign y19259 = n35652 ;
  assign y19260 = ~n35654 ;
  assign y19261 = ~n35656 ;
  assign y19262 = ~n35657 ;
  assign y19263 = n35659 ;
  assign y19264 = ~1'b0 ;
  assign y19265 = ~n35661 ;
  assign y19266 = ~1'b0 ;
  assign y19267 = ~n35667 ;
  assign y19268 = ~n35672 ;
  assign y19269 = n35673 ;
  assign y19270 = ~n35675 ;
  assign y19271 = n35677 ;
  assign y19272 = ~1'b0 ;
  assign y19273 = ~n35678 ;
  assign y19274 = ~n35680 ;
  assign y19275 = ~n35683 ;
  assign y19276 = ~1'b0 ;
  assign y19277 = n35686 ;
  assign y19278 = ~n35687 ;
  assign y19279 = n35689 ;
  assign y19280 = n35691 ;
  assign y19281 = n35698 ;
  assign y19282 = ~1'b0 ;
  assign y19283 = ~1'b0 ;
  assign y19284 = ~1'b0 ;
  assign y19285 = n35701 ;
  assign y19286 = ~1'b0 ;
  assign y19287 = ~n1801 ;
  assign y19288 = n35704 ;
  assign y19289 = ~1'b0 ;
  assign y19290 = ~n35707 ;
  assign y19291 = ~1'b0 ;
  assign y19292 = ~n35712 ;
  assign y19293 = n35713 ;
  assign y19294 = ~n35715 ;
  assign y19295 = ~1'b0 ;
  assign y19296 = 1'b0 ;
  assign y19297 = ~n35717 ;
  assign y19298 = ~n35718 ;
  assign y19299 = ~n35720 ;
  assign y19300 = ~n35722 ;
  assign y19301 = ~n35726 ;
  assign y19302 = n35727 ;
  assign y19303 = ~1'b0 ;
  assign y19304 = n35729 ;
  assign y19305 = ~n35731 ;
  assign y19306 = n35734 ;
  assign y19307 = ~1'b0 ;
  assign y19308 = ~n35735 ;
  assign y19309 = ~n35736 ;
  assign y19310 = ~1'b0 ;
  assign y19311 = ~1'b0 ;
  assign y19312 = n35741 ;
  assign y19313 = ~n35742 ;
  assign y19314 = n35743 ;
  assign y19315 = ~1'b0 ;
  assign y19316 = ~1'b0 ;
  assign y19317 = ~1'b0 ;
  assign y19318 = ~n35745 ;
  assign y19319 = n24640 ;
  assign y19320 = ~1'b0 ;
  assign y19321 = ~1'b0 ;
  assign y19322 = ~n35749 ;
  assign y19323 = ~n35751 ;
  assign y19324 = ~1'b0 ;
  assign y19325 = n35753 ;
  assign y19326 = ~n35754 ;
  assign y19327 = ~n35765 ;
  assign y19328 = ~x130 ;
  assign y19329 = ~n26190 ;
  assign y19330 = n35766 ;
  assign y19331 = ~1'b0 ;
  assign y19332 = ~n35768 ;
  assign y19333 = ~n35773 ;
  assign y19334 = ~n35777 ;
  assign y19335 = ~1'b0 ;
  assign y19336 = ~n35782 ;
  assign y19337 = n35783 ;
  assign y19338 = n35786 ;
  assign y19339 = n35787 ;
  assign y19340 = ~n35788 ;
  assign y19341 = n35796 ;
  assign y19342 = ~1'b0 ;
  assign y19343 = n35797 ;
  assign y19344 = ~1'b0 ;
  assign y19345 = ~n35799 ;
  assign y19346 = n35800 ;
  assign y19347 = ~n35804 ;
  assign y19348 = ~n35805 ;
  assign y19349 = ~n9181 ;
  assign y19350 = ~1'b0 ;
  assign y19351 = ~1'b0 ;
  assign y19352 = ~1'b0 ;
  assign y19353 = ~1'b0 ;
  assign y19354 = ~n35809 ;
  assign y19355 = n35810 ;
  assign y19356 = n5402 ;
  assign y19357 = ~n35813 ;
  assign y19358 = ~n35816 ;
  assign y19359 = ~1'b0 ;
  assign y19360 = n4023 ;
  assign y19361 = n35817 ;
  assign y19362 = ~1'b0 ;
  assign y19363 = ~1'b0 ;
  assign y19364 = n35818 ;
  assign y19365 = n35819 ;
  assign y19366 = ~1'b0 ;
  assign y19367 = n35823 ;
  assign y19368 = n35824 ;
  assign y19369 = ~n35825 ;
  assign y19370 = n35826 ;
  assign y19371 = n35833 ;
  assign y19372 = ~n35835 ;
  assign y19373 = ~1'b0 ;
  assign y19374 = n35837 ;
  assign y19375 = ~1'b0 ;
  assign y19376 = ~n35840 ;
  assign y19377 = ~n11653 ;
  assign y19378 = 1'b0 ;
  assign y19379 = n35842 ;
  assign y19380 = n2045 ;
  assign y19381 = ~n35843 ;
  assign y19382 = ~1'b0 ;
  assign y19383 = n35844 ;
  assign y19384 = 1'b0 ;
  assign y19385 = n35846 ;
  assign y19386 = n35848 ;
  assign y19387 = ~n35850 ;
  assign y19388 = ~n35853 ;
  assign y19389 = ~n35854 ;
  assign y19390 = ~1'b0 ;
  assign y19391 = ~n35858 ;
  assign y19392 = ~n35859 ;
  assign y19393 = ~n2785 ;
  assign y19394 = ~n35861 ;
  assign y19395 = ~1'b0 ;
  assign y19396 = n35864 ;
  assign y19397 = ~n35866 ;
  assign y19398 = n35871 ;
  assign y19399 = ~n35877 ;
  assign y19400 = ~n35878 ;
  assign y19401 = ~n35885 ;
  assign y19402 = 1'b0 ;
  assign y19403 = 1'b0 ;
  assign y19404 = ~1'b0 ;
  assign y19405 = ~1'b0 ;
  assign y19406 = ~n35171 ;
  assign y19407 = ~1'b0 ;
  assign y19408 = n35889 ;
  assign y19409 = ~n35890 ;
  assign y19410 = n35894 ;
  assign y19411 = ~n35792 ;
  assign y19412 = ~n35896 ;
  assign y19413 = ~1'b0 ;
  assign y19414 = n35897 ;
  assign y19415 = ~n35898 ;
  assign y19416 = ~1'b0 ;
  assign y19417 = n35899 ;
  assign y19418 = 1'b0 ;
  assign y19419 = ~n35903 ;
  assign y19420 = n35906 ;
  assign y19421 = ~1'b0 ;
  assign y19422 = ~n35907 ;
  assign y19423 = ~n35908 ;
  assign y19424 = ~1'b0 ;
  assign y19425 = ~1'b0 ;
  assign y19426 = ~1'b0 ;
  assign y19427 = ~1'b0 ;
  assign y19428 = ~n35912 ;
  assign y19429 = n35913 ;
  assign y19430 = ~n35914 ;
  assign y19431 = ~1'b0 ;
  assign y19432 = n35916 ;
  assign y19433 = ~n35923 ;
  assign y19434 = ~n35924 ;
  assign y19435 = ~1'b0 ;
  assign y19436 = ~n35925 ;
  assign y19437 = n35926 ;
  assign y19438 = ~n35928 ;
  assign y19439 = ~1'b0 ;
  assign y19440 = n35931 ;
  assign y19441 = ~1'b0 ;
  assign y19442 = ~1'b0 ;
  assign y19443 = ~1'b0 ;
  assign y19444 = ~n26841 ;
  assign y19445 = ~1'b0 ;
  assign y19446 = ~n35932 ;
  assign y19447 = n35934 ;
  assign y19448 = ~1'b0 ;
  assign y19449 = 1'b0 ;
  assign y19450 = n35936 ;
  assign y19451 = ~n35938 ;
  assign y19452 = ~1'b0 ;
  assign y19453 = n35949 ;
  assign y19454 = n35952 ;
  assign y19455 = ~n35955 ;
  assign y19456 = n35957 ;
  assign y19457 = ~1'b0 ;
  assign y19458 = ~n35959 ;
  assign y19459 = ~n35963 ;
  assign y19460 = ~n35965 ;
  assign y19461 = ~n35966 ;
  assign y19462 = ~1'b0 ;
  assign y19463 = ~n35969 ;
  assign y19464 = ~1'b0 ;
  assign y19465 = n35973 ;
  assign y19466 = ~n35974 ;
  assign y19467 = n25142 ;
  assign y19468 = ~1'b0 ;
  assign y19469 = n35976 ;
  assign y19470 = n35980 ;
  assign y19471 = ~1'b0 ;
  assign y19472 = n35985 ;
  assign y19473 = n35986 ;
  assign y19474 = ~n35988 ;
  assign y19475 = n14470 ;
  assign y19476 = n35989 ;
  assign y19477 = n35991 ;
  assign y19478 = ~1'b0 ;
  assign y19479 = n35992 ;
  assign y19480 = ~n35995 ;
  assign y19481 = n35996 ;
  assign y19482 = ~n35998 ;
  assign y19483 = n36001 ;
  assign y19484 = ~n36002 ;
  assign y19485 = ~n36003 ;
  assign y19486 = ~1'b0 ;
  assign y19487 = ~1'b0 ;
  assign y19488 = n858 ;
  assign y19489 = ~1'b0 ;
  assign y19490 = ~n23389 ;
  assign y19491 = ~n36008 ;
  assign y19492 = ~n36010 ;
  assign y19493 = ~1'b0 ;
  assign y19494 = ~1'b0 ;
  assign y19495 = n36014 ;
  assign y19496 = n13613 ;
  assign y19497 = ~n36019 ;
  assign y19498 = ~1'b0 ;
  assign y19499 = n36022 ;
  assign y19500 = n36023 ;
  assign y19501 = n36024 ;
  assign y19502 = n36033 ;
  assign y19503 = ~1'b0 ;
  assign y19504 = ~n36035 ;
  assign y19505 = ~1'b0 ;
  assign y19506 = ~n36038 ;
  assign y19507 = ~n36042 ;
  assign y19508 = ~1'b0 ;
  assign y19509 = 1'b0 ;
  assign y19510 = n36046 ;
  assign y19511 = ~n36050 ;
  assign y19512 = n36051 ;
  assign y19513 = ~1'b0 ;
  assign y19514 = ~n26515 ;
  assign y19515 = ~1'b0 ;
  assign y19516 = n36053 ;
  assign y19517 = ~1'b0 ;
  assign y19518 = ~n36054 ;
  assign y19519 = ~n36058 ;
  assign y19520 = n36060 ;
  assign y19521 = n36061 ;
  assign y19522 = ~1'b0 ;
  assign y19523 = n36063 ;
  assign y19524 = ~1'b0 ;
  assign y19525 = n32866 ;
  assign y19526 = n36064 ;
  assign y19527 = ~1'b0 ;
  assign y19528 = ~n36066 ;
  assign y19529 = n20204 ;
  assign y19530 = n36067 ;
  assign y19531 = ~1'b0 ;
  assign y19532 = n36069 ;
  assign y19533 = ~1'b0 ;
  assign y19534 = n36073 ;
  assign y19535 = n36076 ;
  assign y19536 = ~1'b0 ;
  assign y19537 = ~1'b0 ;
  assign y19538 = ~1'b0 ;
  assign y19539 = ~1'b0 ;
  assign y19540 = ~n36077 ;
  assign y19541 = n16023 ;
  assign y19542 = ~n36080 ;
  assign y19543 = ~1'b0 ;
  assign y19544 = ~n29289 ;
  assign y19545 = n36084 ;
  assign y19546 = n36085 ;
  assign y19547 = ~n36088 ;
  assign y19548 = ~n36089 ;
  assign y19549 = n36090 ;
  assign y19550 = ~n36091 ;
  assign y19551 = ~n36093 ;
  assign y19552 = ~1'b0 ;
  assign y19553 = ~1'b0 ;
  assign y19554 = n36098 ;
  assign y19555 = n36099 ;
  assign y19556 = ~n36103 ;
  assign y19557 = n36105 ;
  assign y19558 = ~n36106 ;
  assign y19559 = n36109 ;
  assign y19560 = n36112 ;
  assign y19561 = ~n36113 ;
  assign y19562 = 1'b0 ;
  assign y19563 = n36114 ;
  assign y19564 = n36116 ;
  assign y19565 = 1'b0 ;
  assign y19566 = n36117 ;
  assign y19567 = n36120 ;
  assign y19568 = ~1'b0 ;
  assign y19569 = ~1'b0 ;
  assign y19570 = ~1'b0 ;
  assign y19571 = n36122 ;
  assign y19572 = ~1'b0 ;
  assign y19573 = n36123 ;
  assign y19574 = n36124 ;
  assign y19575 = n36125 ;
  assign y19576 = ~1'b0 ;
  assign y19577 = ~n36130 ;
  assign y19578 = n36131 ;
  assign y19579 = ~n36133 ;
  assign y19580 = ~n36137 ;
  assign y19581 = ~n8763 ;
  assign y19582 = n36138 ;
  assign y19583 = n36139 ;
  assign y19584 = ~n36140 ;
  assign y19585 = ~n36143 ;
  assign y19586 = n36145 ;
  assign y19587 = n36151 ;
  assign y19588 = ~n36152 ;
  assign y19589 = ~1'b0 ;
  assign y19590 = ~1'b0 ;
  assign y19591 = ~n36154 ;
  assign y19592 = n36158 ;
  assign y19593 = ~n36159 ;
  assign y19594 = n36163 ;
  assign y19595 = 1'b0 ;
  assign y19596 = n36165 ;
  assign y19597 = ~1'b0 ;
  assign y19598 = ~n36168 ;
  assign y19599 = ~1'b0 ;
  assign y19600 = ~1'b0 ;
  assign y19601 = ~n21373 ;
  assign y19602 = n36170 ;
  assign y19603 = n36173 ;
  assign y19604 = n36175 ;
  assign y19605 = ~1'b0 ;
  assign y19606 = ~x86 ;
  assign y19607 = ~1'b0 ;
  assign y19608 = ~n36178 ;
  assign y19609 = ~1'b0 ;
  assign y19610 = n36183 ;
  assign y19611 = ~1'b0 ;
  assign y19612 = ~n36187 ;
  assign y19613 = n36188 ;
  assign y19614 = ~n36192 ;
  assign y19615 = n36195 ;
  assign y19616 = ~1'b0 ;
  assign y19617 = n36200 ;
  assign y19618 = n36204 ;
  assign y19619 = n36206 ;
  assign y19620 = n36207 ;
  assign y19621 = ~1'b0 ;
  assign y19622 = ~n36209 ;
  assign y19623 = ~n36211 ;
  assign y19624 = ~n36215 ;
  assign y19625 = n36218 ;
  assign y19626 = ~n36219 ;
  assign y19627 = ~1'b0 ;
  assign y19628 = ~n36222 ;
  assign y19629 = ~1'b0 ;
  assign y19630 = n36223 ;
  assign y19631 = n36226 ;
  assign y19632 = n36227 ;
  assign y19633 = ~n36228 ;
  assign y19634 = n36230 ;
  assign y19635 = ~n36231 ;
  assign y19636 = ~n36232 ;
  assign y19637 = ~1'b0 ;
  assign y19638 = ~1'b0 ;
  assign y19639 = n1404 ;
  assign y19640 = n36234 ;
  assign y19641 = ~n36235 ;
  assign y19642 = n36240 ;
  assign y19643 = ~1'b0 ;
  assign y19644 = ~n3828 ;
  assign y19645 = ~n36246 ;
  assign y19646 = ~1'b0 ;
  assign y19647 = ~1'b0 ;
  assign y19648 = ~1'b0 ;
  assign y19649 = ~1'b0 ;
  assign y19650 = ~n36247 ;
  assign y19651 = ~n35835 ;
  assign y19652 = ~n22461 ;
  assign y19653 = ~1'b0 ;
  assign y19654 = ~1'b0 ;
  assign y19655 = n36249 ;
  assign y19656 = ~1'b0 ;
  assign y19657 = n36252 ;
  assign y19658 = 1'b0 ;
  assign y19659 = ~1'b0 ;
  assign y19660 = ~n36256 ;
  assign y19661 = ~n36257 ;
  assign y19662 = ~1'b0 ;
  assign y19663 = ~n36259 ;
  assign y19664 = ~n36261 ;
  assign y19665 = ~1'b0 ;
  assign y19666 = ~n36263 ;
  assign y19667 = n36264 ;
  assign y19668 = ~n36266 ;
  assign y19669 = ~1'b0 ;
  assign y19670 = ~n36269 ;
  assign y19671 = ~n36270 ;
  assign y19672 = ~n36272 ;
  assign y19673 = ~1'b0 ;
  assign y19674 = n36277 ;
  assign y19675 = ~1'b0 ;
  assign y19676 = ~1'b0 ;
  assign y19677 = n36281 ;
  assign y19678 = ~1'b0 ;
  assign y19679 = n36283 ;
  assign y19680 = n36286 ;
  assign y19681 = n36291 ;
  assign y19682 = n36294 ;
  assign y19683 = ~1'b0 ;
  assign y19684 = ~1'b0 ;
  assign y19685 = n36298 ;
  assign y19686 = ~1'b0 ;
  assign y19687 = ~n36303 ;
  assign y19688 = n36306 ;
  assign y19689 = n36307 ;
  assign y19690 = ~n36312 ;
  assign y19691 = n36313 ;
  assign y19692 = ~n36317 ;
  assign y19693 = n36318 ;
  assign y19694 = ~1'b0 ;
  assign y19695 = ~1'b0 ;
  assign y19696 = ~n36322 ;
  assign y19697 = ~1'b0 ;
  assign y19698 = ~n36323 ;
  assign y19699 = 1'b0 ;
  assign y19700 = ~n36329 ;
  assign y19701 = ~n36334 ;
  assign y19702 = n36337 ;
  assign y19703 = ~n36339 ;
  assign y19704 = ~n36341 ;
  assign y19705 = ~n36344 ;
  assign y19706 = ~1'b0 ;
  assign y19707 = n36345 ;
  assign y19708 = n36353 ;
  assign y19709 = n36356 ;
  assign y19710 = ~1'b0 ;
  assign y19711 = n6446 ;
  assign y19712 = n36358 ;
  assign y19713 = ~1'b0 ;
  assign y19714 = ~1'b0 ;
  assign y19715 = ~n36360 ;
  assign y19716 = 1'b0 ;
  assign y19717 = ~n36361 ;
  assign y19718 = ~n36362 ;
  assign y19719 = ~n36365 ;
  assign y19720 = ~1'b0 ;
  assign y19721 = n9322 ;
  assign y19722 = ~1'b0 ;
  assign y19723 = n36366 ;
  assign y19724 = n36370 ;
  assign y19725 = ~1'b0 ;
  assign y19726 = ~n36373 ;
  assign y19727 = ~n36374 ;
  assign y19728 = ~1'b0 ;
  assign y19729 = ~1'b0 ;
  assign y19730 = ~1'b0 ;
  assign y19731 = ~n36376 ;
  assign y19732 = ~1'b0 ;
  assign y19733 = ~1'b0 ;
  assign y19734 = n36379 ;
  assign y19735 = ~n36380 ;
  assign y19736 = ~1'b0 ;
  assign y19737 = ~1'b0 ;
  assign y19738 = n36382 ;
  assign y19739 = n36383 ;
  assign y19740 = ~n36384 ;
  assign y19741 = n36386 ;
  assign y19742 = n36392 ;
  assign y19743 = n36393 ;
  assign y19744 = ~n29295 ;
  assign y19745 = ~n36395 ;
  assign y19746 = ~1'b0 ;
  assign y19747 = n36396 ;
  assign y19748 = n36398 ;
  assign y19749 = ~n36400 ;
  assign y19750 = n36403 ;
  assign y19751 = ~n36406 ;
  assign y19752 = ~1'b0 ;
  assign y19753 = ~n36411 ;
  assign y19754 = n36414 ;
  assign y19755 = ~1'b0 ;
  assign y19756 = ~n36416 ;
  assign y19757 = ~n36418 ;
  assign y19758 = ~1'b0 ;
  assign y19759 = n36421 ;
  assign y19760 = n36427 ;
  assign y19761 = n31776 ;
  assign y19762 = ~n36428 ;
  assign y19763 = n36430 ;
  assign y19764 = n36432 ;
  assign y19765 = 1'b0 ;
  assign y19766 = ~n36435 ;
  assign y19767 = ~1'b0 ;
  assign y19768 = ~1'b0 ;
  assign y19769 = n18847 ;
  assign y19770 = ~1'b0 ;
  assign y19771 = ~n36437 ;
  assign y19772 = n36439 ;
  assign y19773 = n36443 ;
  assign y19774 = ~n36447 ;
  assign y19775 = ~n36449 ;
  assign y19776 = n36453 ;
  assign y19777 = ~n36455 ;
  assign y19778 = ~1'b0 ;
  assign y19779 = ~n36458 ;
  assign y19780 = n36459 ;
  assign y19781 = ~1'b0 ;
  assign y19782 = n36461 ;
  assign y19783 = n786 ;
  assign y19784 = ~1'b0 ;
  assign y19785 = n36465 ;
  assign y19786 = n36467 ;
  assign y19787 = n36474 ;
  assign y19788 = n36475 ;
  assign y19789 = ~1'b0 ;
  assign y19790 = ~n36476 ;
  assign y19791 = 1'b0 ;
  assign y19792 = ~1'b0 ;
  assign y19793 = ~1'b0 ;
  assign y19794 = n36477 ;
  assign y19795 = ~1'b0 ;
  assign y19796 = 1'b0 ;
  assign y19797 = ~n36478 ;
  assign y19798 = ~1'b0 ;
  assign y19799 = ~n36479 ;
  assign y19800 = 1'b0 ;
  assign y19801 = ~n16866 ;
  assign y19802 = ~n36481 ;
  assign y19803 = n36485 ;
  assign y19804 = n36487 ;
  assign y19805 = ~n36493 ;
  assign y19806 = ~n36497 ;
  assign y19807 = ~n36501 ;
  assign y19808 = ~1'b0 ;
  assign y19809 = n36503 ;
  assign y19810 = ~1'b0 ;
  assign y19811 = ~1'b0 ;
  assign y19812 = ~1'b0 ;
  assign y19813 = ~1'b0 ;
  assign y19814 = ~1'b0 ;
  assign y19815 = ~n36509 ;
  assign y19816 = ~n36511 ;
  assign y19817 = ~1'b0 ;
  assign y19818 = ~1'b0 ;
  assign y19819 = ~1'b0 ;
  assign y19820 = ~1'b0 ;
  assign y19821 = n36519 ;
  assign y19822 = ~1'b0 ;
  assign y19823 = ~n36520 ;
  assign y19824 = ~n36521 ;
  assign y19825 = n36522 ;
  assign y19826 = ~n36525 ;
  assign y19827 = ~1'b0 ;
  assign y19828 = ~n36527 ;
  assign y19829 = ~1'b0 ;
  assign y19830 = ~n36531 ;
  assign y19831 = ~1'b0 ;
  assign y19832 = n36533 ;
  assign y19833 = ~n36534 ;
  assign y19834 = ~n7594 ;
  assign y19835 = ~1'b0 ;
  assign y19836 = n36535 ;
  assign y19837 = n36538 ;
  assign y19838 = ~1'b0 ;
  assign y19839 = ~1'b0 ;
  assign y19840 = n36540 ;
  assign y19841 = ~n36543 ;
  assign y19842 = ~1'b0 ;
  assign y19843 = n36544 ;
  assign y19844 = ~1'b0 ;
  assign y19845 = ~n36546 ;
  assign y19846 = ~n36549 ;
  assign y19847 = ~1'b0 ;
  assign y19848 = ~n36550 ;
  assign y19849 = ~n36554 ;
  assign y19850 = n36555 ;
  assign y19851 = n36556 ;
  assign y19852 = n9507 ;
  assign y19853 = n14805 ;
  assign y19854 = n29611 ;
  assign y19855 = n36557 ;
  assign y19856 = ~n36560 ;
  assign y19857 = ~1'b0 ;
  assign y19858 = ~1'b0 ;
  assign y19859 = ~n36563 ;
  assign y19860 = ~n36565 ;
  assign y19861 = ~n13025 ;
  assign y19862 = n36566 ;
  assign y19863 = ~1'b0 ;
  assign y19864 = n36567 ;
  assign y19865 = ~n36568 ;
  assign y19866 = ~n36571 ;
  assign y19867 = ~n36573 ;
  assign y19868 = ~n36574 ;
  assign y19869 = ~n36575 ;
  assign y19870 = ~1'b0 ;
  assign y19871 = ~n36576 ;
  assign y19872 = ~1'b0 ;
  assign y19873 = n36577 ;
  assign y19874 = n36581 ;
  assign y19875 = ~n36582 ;
  assign y19876 = ~1'b0 ;
  assign y19877 = ~1'b0 ;
  assign y19878 = ~1'b0 ;
  assign y19879 = n29541 ;
  assign y19880 = ~n36585 ;
  assign y19881 = n36586 ;
  assign y19882 = ~1'b0 ;
  assign y19883 = ~1'b0 ;
  assign y19884 = ~1'b0 ;
  assign y19885 = ~n14790 ;
  assign y19886 = 1'b0 ;
  assign y19887 = ~1'b0 ;
  assign y19888 = ~n36590 ;
  assign y19889 = n6090 ;
  assign y19890 = ~n36595 ;
  assign y19891 = ~1'b0 ;
  assign y19892 = n36599 ;
  assign y19893 = n36603 ;
  assign y19894 = n36604 ;
  assign y19895 = ~1'b0 ;
  assign y19896 = n36605 ;
  assign y19897 = ~n33721 ;
  assign y19898 = ~n36606 ;
  assign y19899 = ~n36607 ;
  assign y19900 = n36608 ;
  assign y19901 = n36610 ;
  assign y19902 = ~n36612 ;
  assign y19903 = n36614 ;
  assign y19904 = n36617 ;
  assign y19905 = n36621 ;
  assign y19906 = ~n36624 ;
  assign y19907 = ~n36625 ;
  assign y19908 = ~1'b0 ;
  assign y19909 = ~n36627 ;
  assign y19910 = n36628 ;
  assign y19911 = n36629 ;
  assign y19912 = ~n36630 ;
  assign y19913 = n36632 ;
  assign y19914 = ~1'b0 ;
  assign y19915 = n36633 ;
  assign y19916 = ~1'b0 ;
  assign y19917 = ~n36634 ;
  assign y19918 = ~n36635 ;
  assign y19919 = ~1'b0 ;
  assign y19920 = n36636 ;
  assign y19921 = ~n36641 ;
  assign y19922 = ~1'b0 ;
  assign y19923 = ~1'b0 ;
  assign y19924 = ~n36642 ;
  assign y19925 = n36647 ;
  assign y19926 = ~n36649 ;
  assign y19927 = ~1'b0 ;
  assign y19928 = ~n36652 ;
  assign y19929 = ~1'b0 ;
  assign y19930 = ~n36653 ;
  assign y19931 = n36654 ;
  assign y19932 = ~n36657 ;
  assign y19933 = ~n16214 ;
  assign y19934 = ~n36660 ;
  assign y19935 = ~1'b0 ;
  assign y19936 = n36661 ;
  assign y19937 = ~n36662 ;
  assign y19938 = n36666 ;
  assign y19939 = ~1'b0 ;
  assign y19940 = ~n1392 ;
  assign y19941 = n36667 ;
  assign y19942 = ~n36668 ;
  assign y19943 = n36670 ;
  assign y19944 = ~1'b0 ;
  assign y19945 = n24369 ;
  assign y19946 = n36671 ;
  assign y19947 = n36673 ;
  assign y19948 = n36675 ;
  assign y19949 = n20174 ;
  assign y19950 = ~n36678 ;
  assign y19951 = ~n36683 ;
  assign y19952 = ~1'b0 ;
  assign y19953 = n36689 ;
  assign y19954 = n36694 ;
  assign y19955 = ~1'b0 ;
  assign y19956 = ~n36695 ;
  assign y19957 = 1'b0 ;
  assign y19958 = ~n36697 ;
  assign y19959 = ~n36698 ;
  assign y19960 = n36700 ;
  assign y19961 = ~n4500 ;
  assign y19962 = n36705 ;
  assign y19963 = ~n36707 ;
  assign y19964 = n36711 ;
  assign y19965 = ~n36712 ;
  assign y19966 = ~1'b0 ;
  assign y19967 = ~1'b0 ;
  assign y19968 = ~n36713 ;
  assign y19969 = ~n18741 ;
  assign y19970 = ~n36718 ;
  assign y19971 = ~1'b0 ;
  assign y19972 = 1'b0 ;
  assign y19973 = ~1'b0 ;
  assign y19974 = n36719 ;
  assign y19975 = ~n36723 ;
  assign y19976 = ~1'b0 ;
  assign y19977 = ~1'b0 ;
  assign y19978 = n18150 ;
  assign y19979 = n36724 ;
  assign y19980 = ~n36725 ;
  assign y19981 = ~n36726 ;
  assign y19982 = ~n36727 ;
  assign y19983 = ~n20708 ;
  assign y19984 = ~n36728 ;
  assign y19985 = n23554 ;
  assign y19986 = ~n36731 ;
  assign y19987 = ~1'b0 ;
  assign y19988 = ~n36732 ;
  assign y19989 = n36739 ;
  assign y19990 = ~1'b0 ;
  assign y19991 = ~1'b0 ;
  assign y19992 = ~1'b0 ;
  assign y19993 = ~1'b0 ;
  assign y19994 = ~1'b0 ;
  assign y19995 = 1'b0 ;
  assign y19996 = ~n36743 ;
  assign y19997 = ~1'b0 ;
  assign y19998 = ~n36745 ;
  assign y19999 = ~1'b0 ;
  assign y20000 = n36749 ;
  assign y20001 = ~n36751 ;
  assign y20002 = ~n36754 ;
  assign y20003 = ~n12239 ;
  assign y20004 = ~n36756 ;
  assign y20005 = n36758 ;
  assign y20006 = n36760 ;
  assign y20007 = ~1'b0 ;
  assign y20008 = n36770 ;
  assign y20009 = ~n36772 ;
  assign y20010 = n8550 ;
  assign y20011 = ~n36774 ;
  assign y20012 = ~1'b0 ;
  assign y20013 = ~n36777 ;
  assign y20014 = ~1'b0 ;
  assign y20015 = n36778 ;
  assign y20016 = ~x207 ;
  assign y20017 = ~n36781 ;
  assign y20018 = n36782 ;
  assign y20019 = n36783 ;
  assign y20020 = ~1'b0 ;
  assign y20021 = ~1'b0 ;
  assign y20022 = n36787 ;
  assign y20023 = x112 ;
  assign y20024 = ~n36788 ;
  assign y20025 = ~n36791 ;
  assign y20026 = ~n36793 ;
  assign y20027 = ~1'b0 ;
  assign y20028 = ~1'b0 ;
  assign y20029 = ~1'b0 ;
  assign y20030 = ~n36795 ;
  assign y20031 = ~n36796 ;
  assign y20032 = ~n36804 ;
  assign y20033 = n36805 ;
  assign y20034 = ~1'b0 ;
  assign y20035 = ~1'b0 ;
  assign y20036 = ~n36808 ;
  assign y20037 = 1'b0 ;
  assign y20038 = ~n36809 ;
  assign y20039 = ~1'b0 ;
  assign y20040 = n36810 ;
  assign y20041 = n27740 ;
  assign y20042 = n36815 ;
  assign y20043 = n36819 ;
  assign y20044 = ~1'b0 ;
  assign y20045 = n36821 ;
  assign y20046 = ~1'b0 ;
  assign y20047 = n36823 ;
  assign y20048 = ~n36825 ;
  assign y20049 = ~1'b0 ;
  assign y20050 = ~n36827 ;
  assign y20051 = ~n36829 ;
  assign y20052 = ~n36830 ;
  assign y20053 = ~1'b0 ;
  assign y20054 = ~n36832 ;
  assign y20055 = n36833 ;
  assign y20056 = ~1'b0 ;
  assign y20057 = ~1'b0 ;
  assign y20058 = ~1'b0 ;
  assign y20059 = ~1'b0 ;
  assign y20060 = ~1'b0 ;
  assign y20061 = 1'b0 ;
  assign y20062 = ~n36834 ;
  assign y20063 = n36837 ;
  assign y20064 = n36839 ;
  assign y20065 = ~n36840 ;
  assign y20066 = ~1'b0 ;
  assign y20067 = ~n36841 ;
  assign y20068 = ~n36842 ;
  assign y20069 = ~1'b0 ;
  assign y20070 = n36844 ;
  assign y20071 = ~n36845 ;
  assign y20072 = ~n36847 ;
  assign y20073 = ~n3912 ;
  assign y20074 = ~1'b0 ;
  assign y20075 = ~1'b0 ;
  assign y20076 = n36849 ;
  assign y20077 = ~n36850 ;
  assign y20078 = ~1'b0 ;
  assign y20079 = n36851 ;
  assign y20080 = ~x249 ;
  assign y20081 = n36852 ;
  assign y20082 = ~n36855 ;
  assign y20083 = n25511 ;
  assign y20084 = ~1'b0 ;
  assign y20085 = ~n36857 ;
  assign y20086 = n36866 ;
  assign y20087 = ~n36867 ;
  assign y20088 = ~1'b0 ;
  assign y20089 = ~1'b0 ;
  assign y20090 = n36868 ;
  assign y20091 = ~n36870 ;
  assign y20092 = n36875 ;
  assign y20093 = ~1'b0 ;
  assign y20094 = ~1'b0 ;
  assign y20095 = ~1'b0 ;
  assign y20096 = ~n36876 ;
  assign y20097 = ~n21152 ;
  assign y20098 = n36877 ;
  assign y20099 = ~1'b0 ;
  assign y20100 = ~1'b0 ;
  assign y20101 = ~n36878 ;
  assign y20102 = ~n36882 ;
  assign y20103 = n36884 ;
  assign y20104 = ~1'b0 ;
  assign y20105 = n36885 ;
  assign y20106 = n36887 ;
  assign y20107 = ~n36888 ;
  assign y20108 = n36889 ;
  assign y20109 = n36892 ;
  assign y20110 = n36897 ;
  assign y20111 = n36898 ;
  assign y20112 = ~1'b0 ;
  assign y20113 = ~n36900 ;
  assign y20114 = ~n36903 ;
  assign y20115 = n36904 ;
  assign y20116 = n36909 ;
  assign y20117 = ~1'b0 ;
  assign y20118 = ~1'b0 ;
  assign y20119 = ~n36911 ;
  assign y20120 = ~n36912 ;
  assign y20121 = ~1'b0 ;
  assign y20122 = ~1'b0 ;
  assign y20123 = n36914 ;
  assign y20124 = n36917 ;
  assign y20125 = ~1'b0 ;
  assign y20126 = ~n36919 ;
  assign y20127 = ~n36921 ;
  assign y20128 = n36926 ;
  assign y20129 = n36927 ;
  assign y20130 = n36928 ;
  assign y20131 = n36929 ;
  assign y20132 = ~n36933 ;
  assign y20133 = ~n36935 ;
  assign y20134 = ~1'b0 ;
  assign y20135 = ~1'b0 ;
  assign y20136 = n19138 ;
  assign y20137 = ~1'b0 ;
  assign y20138 = n36944 ;
  assign y20139 = ~n36945 ;
  assign y20140 = ~1'b0 ;
  assign y20141 = ~n36949 ;
  assign y20142 = ~n36950 ;
  assign y20143 = ~1'b0 ;
  assign y20144 = ~1'b0 ;
  assign y20145 = ~n2010 ;
  assign y20146 = ~n36952 ;
  assign y20147 = ~n36953 ;
  assign y20148 = ~n36955 ;
  assign y20149 = n16673 ;
  assign y20150 = n36956 ;
  assign y20151 = n36963 ;
  assign y20152 = ~n36964 ;
  assign y20153 = n36966 ;
  assign y20154 = ~1'b0 ;
  assign y20155 = n8523 ;
  assign y20156 = ~1'b0 ;
  assign y20157 = ~n36967 ;
  assign y20158 = ~1'b0 ;
  assign y20159 = n36971 ;
  assign y20160 = ~n36972 ;
  assign y20161 = ~1'b0 ;
  assign y20162 = ~n7398 ;
  assign y20163 = ~n36975 ;
  assign y20164 = n11532 ;
  assign y20165 = 1'b0 ;
  assign y20166 = n36977 ;
  assign y20167 = ~1'b0 ;
  assign y20168 = ~n36981 ;
  assign y20169 = ~n36983 ;
  assign y20170 = ~1'b0 ;
  assign y20171 = n36987 ;
  assign y20172 = ~n36988 ;
  assign y20173 = n36989 ;
  assign y20174 = n36992 ;
  assign y20175 = ~1'b0 ;
  assign y20176 = n36993 ;
  assign y20177 = n36994 ;
  assign y20178 = n36995 ;
  assign y20179 = ~1'b0 ;
  assign y20180 = ~1'b0 ;
  assign y20181 = ~n37000 ;
  assign y20182 = ~1'b0 ;
  assign y20183 = n37002 ;
  assign y20184 = n37004 ;
  assign y20185 = n37007 ;
  assign y20186 = ~1'b0 ;
  assign y20187 = ~1'b0 ;
  assign y20188 = ~1'b0 ;
  assign y20189 = ~1'b0 ;
  assign y20190 = ~1'b0 ;
  assign y20191 = n37010 ;
  assign y20192 = ~1'b0 ;
  assign y20193 = ~n37011 ;
  assign y20194 = ~1'b0 ;
  assign y20195 = ~n37012 ;
  assign y20196 = ~n37015 ;
  assign y20197 = ~1'b0 ;
  assign y20198 = ~1'b0 ;
  assign y20199 = ~1'b0 ;
  assign y20200 = ~n37016 ;
  assign y20201 = ~1'b0 ;
  assign y20202 = ~n37018 ;
  assign y20203 = n37020 ;
  assign y20204 = ~1'b0 ;
  assign y20205 = ~n37022 ;
  assign y20206 = ~n37027 ;
  assign y20207 = ~n37030 ;
  assign y20208 = ~1'b0 ;
  assign y20209 = n37031 ;
  assign y20210 = n37033 ;
  assign y20211 = ~n37035 ;
  assign y20212 = ~1'b0 ;
  assign y20213 = n37036 ;
  assign y20214 = n37041 ;
  assign y20215 = n37047 ;
  assign y20216 = ~n37049 ;
  assign y20217 = n37052 ;
  assign y20218 = ~n37059 ;
  assign y20219 = ~n37060 ;
  assign y20220 = ~1'b0 ;
  assign y20221 = n37063 ;
  assign y20222 = n37064 ;
  assign y20223 = n37065 ;
  assign y20224 = ~n37066 ;
  assign y20225 = n37072 ;
  assign y20226 = ~1'b0 ;
  assign y20227 = ~n37073 ;
  assign y20228 = ~1'b0 ;
  assign y20229 = ~n37074 ;
  assign y20230 = n32106 ;
  assign y20231 = ~1'b0 ;
  assign y20232 = n37078 ;
  assign y20233 = ~1'b0 ;
  assign y20234 = ~n37079 ;
  assign y20235 = n37084 ;
  assign y20236 = ~n37085 ;
  assign y20237 = n37086 ;
  assign y20238 = n37095 ;
  assign y20239 = x9 ;
  assign y20240 = ~1'b0 ;
  assign y20241 = n37099 ;
  assign y20242 = n37103 ;
  assign y20243 = ~n37105 ;
  assign y20244 = ~1'b0 ;
  assign y20245 = ~1'b0 ;
  assign y20246 = n37108 ;
  assign y20247 = ~1'b0 ;
  assign y20248 = n37109 ;
  assign y20249 = n37111 ;
  assign y20250 = ~1'b0 ;
  assign y20251 = ~1'b0 ;
  assign y20252 = n37114 ;
  assign y20253 = ~1'b0 ;
  assign y20254 = ~1'b0 ;
  assign y20255 = ~1'b0 ;
  assign y20256 = ~1'b0 ;
  assign y20257 = ~1'b0 ;
  assign y20258 = ~n37117 ;
  assign y20259 = n37118 ;
  assign y20260 = n37119 ;
  assign y20261 = n37126 ;
  assign y20262 = ~n37129 ;
  assign y20263 = ~n11963 ;
  assign y20264 = ~n37130 ;
  assign y20265 = n37131 ;
  assign y20266 = ~n37132 ;
  assign y20267 = ~1'b0 ;
  assign y20268 = n37133 ;
  assign y20269 = ~n37134 ;
  assign y20270 = ~n37135 ;
  assign y20271 = n37136 ;
  assign y20272 = ~n37140 ;
  assign y20273 = n16144 ;
  assign y20274 = ~1'b0 ;
  assign y20275 = n37144 ;
  assign y20276 = ~1'b0 ;
  assign y20277 = ~n8382 ;
  assign y20278 = ~1'b0 ;
  assign y20279 = n37147 ;
  assign y20280 = n37149 ;
  assign y20281 = ~1'b0 ;
  assign y20282 = n37154 ;
  assign y20283 = ~n37157 ;
  assign y20284 = ~n37161 ;
  assign y20285 = n37166 ;
  assign y20286 = ~1'b0 ;
  assign y20287 = n32380 ;
  assign y20288 = n37167 ;
  assign y20289 = ~n37169 ;
  assign y20290 = ~n10966 ;
  assign y20291 = n37171 ;
  assign y20292 = ~n37175 ;
  assign y20293 = ~n37177 ;
  assign y20294 = ~1'b0 ;
  assign y20295 = ~1'b0 ;
  assign y20296 = ~1'b0 ;
  assign y20297 = ~n37178 ;
  assign y20298 = n13479 ;
  assign y20299 = n30025 ;
  assign y20300 = ~n37180 ;
  assign y20301 = n37182 ;
  assign y20302 = n37184 ;
  assign y20303 = n37185 ;
  assign y20304 = ~n37188 ;
  assign y20305 = ~1'b0 ;
  assign y20306 = ~1'b0 ;
  assign y20307 = n37189 ;
  assign y20308 = n15042 ;
  assign y20309 = ~1'b0 ;
  assign y20310 = ~1'b0 ;
  assign y20311 = ~n37191 ;
  assign y20312 = ~1'b0 ;
  assign y20313 = ~n9706 ;
  assign y20314 = ~n37192 ;
  assign y20315 = n37196 ;
  assign y20316 = n37197 ;
  assign y20317 = ~1'b0 ;
  assign y20318 = n37199 ;
  assign y20319 = 1'b0 ;
  assign y20320 = ~n37201 ;
  assign y20321 = ~1'b0 ;
  assign y20322 = ~n37202 ;
  assign y20323 = ~n37203 ;
  assign y20324 = ~n37205 ;
  assign y20325 = ~n37206 ;
  assign y20326 = n36895 ;
  assign y20327 = ~1'b0 ;
  assign y20328 = 1'b0 ;
  assign y20329 = ~n37207 ;
  assign y20330 = ~n37209 ;
  assign y20331 = n37210 ;
  assign y20332 = ~1'b0 ;
  assign y20333 = ~1'b0 ;
  assign y20334 = ~1'b0 ;
  assign y20335 = ~n37214 ;
  assign y20336 = ~1'b0 ;
  assign y20337 = n37216 ;
  assign y20338 = ~n37217 ;
  assign y20339 = ~n37218 ;
  assign y20340 = ~n37219 ;
  assign y20341 = ~n37223 ;
  assign y20342 = ~1'b0 ;
  assign y20343 = n31425 ;
  assign y20344 = ~n37229 ;
  assign y20345 = ~1'b0 ;
  assign y20346 = ~n37231 ;
  assign y20347 = ~1'b0 ;
  assign y20348 = n37234 ;
  assign y20349 = ~n37235 ;
  assign y20350 = n31337 ;
  assign y20351 = ~1'b0 ;
  assign y20352 = ~1'b0 ;
  assign y20353 = ~n37239 ;
  assign y20354 = n37240 ;
  assign y20355 = ~n37241 ;
  assign y20356 = n6479 ;
  assign y20357 = ~n37248 ;
  assign y20358 = n11287 ;
  assign y20359 = ~n37249 ;
  assign y20360 = ~n37252 ;
  assign y20361 = ~1'b0 ;
  assign y20362 = 1'b0 ;
  assign y20363 = ~n37257 ;
  assign y20364 = ~n37259 ;
  assign y20365 = ~1'b0 ;
  assign y20366 = ~1'b0 ;
  assign y20367 = ~n37260 ;
  assign y20368 = n37265 ;
  assign y20369 = ~1'b0 ;
  assign y20370 = n9538 ;
  assign y20371 = ~1'b0 ;
  assign y20372 = ~1'b0 ;
  assign y20373 = ~n37267 ;
  assign y20374 = ~n37270 ;
  assign y20375 = n37272 ;
  assign y20376 = n37273 ;
  assign y20377 = ~n37276 ;
  assign y20378 = n37277 ;
  assign y20379 = ~n37282 ;
  assign y20380 = n37286 ;
  assign y20381 = ~1'b0 ;
  assign y20382 = ~1'b0 ;
  assign y20383 = ~n37288 ;
  assign y20384 = n37289 ;
  assign y20385 = ~1'b0 ;
  assign y20386 = ~1'b0 ;
  assign y20387 = ~1'b0 ;
  assign y20388 = n37292 ;
  assign y20389 = ~n37294 ;
  assign y20390 = ~n37299 ;
  assign y20391 = ~n37301 ;
  assign y20392 = n37319 ;
  assign y20393 = ~n37321 ;
  assign y20394 = ~n37324 ;
  assign y20395 = ~n13768 ;
  assign y20396 = ~1'b0 ;
  assign y20397 = ~n37326 ;
  assign y20398 = ~1'b0 ;
  assign y20399 = n10443 ;
  assign y20400 = n37327 ;
  assign y20401 = n37331 ;
  assign y20402 = ~1'b0 ;
  assign y20403 = ~1'b0 ;
  assign y20404 = ~1'b0 ;
  assign y20405 = ~1'b0 ;
  assign y20406 = ~n37332 ;
  assign y20407 = n37334 ;
  assign y20408 = ~n37336 ;
  assign y20409 = n37337 ;
  assign y20410 = ~n37342 ;
  assign y20411 = ~1'b0 ;
  assign y20412 = ~1'b0 ;
  assign y20413 = n37345 ;
  assign y20414 = n37349 ;
  assign y20415 = ~n2296 ;
  assign y20416 = ~1'b0 ;
  assign y20417 = n37350 ;
  assign y20418 = ~1'b0 ;
  assign y20419 = n37354 ;
  assign y20420 = ~n34207 ;
  assign y20421 = ~1'b0 ;
  assign y20422 = n37357 ;
  assign y20423 = ~n37358 ;
  assign y20424 = ~1'b0 ;
  assign y20425 = n37363 ;
  assign y20426 = n4753 ;
  assign y20427 = n37370 ;
  assign y20428 = ~1'b0 ;
  assign y20429 = ~1'b0 ;
  assign y20430 = ~n37375 ;
  assign y20431 = ~n37380 ;
  assign y20432 = ~1'b0 ;
  assign y20433 = ~n37381 ;
  assign y20434 = 1'b0 ;
  assign y20435 = n37389 ;
  assign y20436 = ~n2848 ;
  assign y20437 = ~n37392 ;
  assign y20438 = n37395 ;
  assign y20439 = n37397 ;
  assign y20440 = ~n37401 ;
  assign y20441 = ~n37402 ;
  assign y20442 = ~n3379 ;
  assign y20443 = n37404 ;
  assign y20444 = ~n37407 ;
  assign y20445 = ~n8166 ;
  assign y20446 = ~1'b0 ;
  assign y20447 = ~1'b0 ;
  assign y20448 = ~1'b0 ;
  assign y20449 = ~n37408 ;
  assign y20450 = n16167 ;
  assign y20451 = n37409 ;
  assign y20452 = ~1'b0 ;
  assign y20453 = ~n37413 ;
  assign y20454 = n37414 ;
  assign y20455 = n37419 ;
  assign y20456 = ~n37420 ;
  assign y20457 = ~1'b0 ;
  assign y20458 = ~n37423 ;
  assign y20459 = ~n37424 ;
  assign y20460 = ~n37428 ;
  assign y20461 = ~1'b0 ;
  assign y20462 = n380 ;
  assign y20463 = ~1'b0 ;
  assign y20464 = n37437 ;
  assign y20465 = ~n37438 ;
  assign y20466 = ~n37439 ;
  assign y20467 = ~n37441 ;
  assign y20468 = ~1'b0 ;
  assign y20469 = ~n37442 ;
  assign y20470 = ~n21786 ;
  assign y20471 = n37443 ;
  assign y20472 = ~n37444 ;
  assign y20473 = ~n37445 ;
  assign y20474 = ~1'b0 ;
  assign y20475 = n37446 ;
  assign y20476 = n37451 ;
  assign y20477 = ~n37452 ;
  assign y20478 = n37453 ;
  assign y20479 = n37466 ;
  assign y20480 = ~1'b0 ;
  assign y20481 = n37467 ;
  assign y20482 = ~1'b0 ;
  assign y20483 = ~n37468 ;
  assign y20484 = 1'b0 ;
  assign y20485 = ~n37472 ;
  assign y20486 = ~n37474 ;
  assign y20487 = ~n37476 ;
  assign y20488 = n37477 ;
  assign y20489 = n20590 ;
  assign y20490 = ~n37483 ;
  assign y20491 = n37486 ;
  assign y20492 = ~n37488 ;
  assign y20493 = ~1'b0 ;
  assign y20494 = ~n37491 ;
  assign y20495 = ~1'b0 ;
  assign y20496 = ~1'b0 ;
  assign y20497 = ~n37494 ;
  assign y20498 = n6169 ;
  assign y20499 = ~n37495 ;
  assign y20500 = ~n37497 ;
  assign y20501 = ~1'b0 ;
  assign y20502 = n37502 ;
  assign y20503 = ~n37505 ;
  assign y20504 = ~1'b0 ;
  assign y20505 = ~1'b0 ;
  assign y20506 = ~n37506 ;
  assign y20507 = ~n37507 ;
  assign y20508 = 1'b0 ;
  assign y20509 = ~n37511 ;
  assign y20510 = ~n37513 ;
  assign y20511 = ~1'b0 ;
  assign y20512 = ~n37515 ;
  assign y20513 = n37519 ;
  assign y20514 = ~1'b0 ;
  assign y20515 = ~n37520 ;
  assign y20516 = ~n37521 ;
  assign y20517 = ~1'b0 ;
  assign y20518 = n37522 ;
  assign y20519 = ~n37524 ;
  assign y20520 = ~1'b0 ;
  assign y20521 = n37525 ;
  assign y20522 = ~n36881 ;
  assign y20523 = ~n37527 ;
  assign y20524 = ~n37528 ;
  assign y20525 = ~n37531 ;
  assign y20526 = n37532 ;
  assign y20527 = n37534 ;
  assign y20528 = ~1'b0 ;
  assign y20529 = ~n37535 ;
  assign y20530 = ~n37538 ;
  assign y20531 = ~1'b0 ;
  assign y20532 = ~1'b0 ;
  assign y20533 = ~n37539 ;
  assign y20534 = ~n37542 ;
  assign y20535 = ~1'b0 ;
  assign y20536 = n37548 ;
  assign y20537 = ~1'b0 ;
  assign y20538 = ~1'b0 ;
  assign y20539 = ~1'b0 ;
  assign y20540 = ~n37550 ;
  assign y20541 = ~1'b0 ;
  assign y20542 = ~n37551 ;
  assign y20543 = ~1'b0 ;
  assign y20544 = ~n37553 ;
  assign y20545 = ~1'b0 ;
  assign y20546 = n37554 ;
  assign y20547 = ~n37555 ;
  assign y20548 = n37556 ;
  assign y20549 = n37559 ;
  assign y20550 = ~1'b0 ;
  assign y20551 = ~1'b0 ;
  assign y20552 = ~n37562 ;
  assign y20553 = ~1'b0 ;
  assign y20554 = n37564 ;
  assign y20555 = ~n37565 ;
  assign y20556 = n37566 ;
  assign y20557 = ~1'b0 ;
  assign y20558 = n37567 ;
  assign y20559 = 1'b0 ;
  assign y20560 = ~n37572 ;
  assign y20561 = ~n5748 ;
  assign y20562 = ~1'b0 ;
  assign y20563 = n37579 ;
  assign y20564 = ~1'b0 ;
  assign y20565 = ~1'b0 ;
  assign y20566 = ~n6991 ;
  assign y20567 = ~n37582 ;
  assign y20568 = n37583 ;
  assign y20569 = n37584 ;
  assign y20570 = ~n37585 ;
  assign y20571 = ~1'b0 ;
  assign y20572 = ~n37587 ;
  assign y20573 = n37588 ;
  assign y20574 = n37593 ;
  assign y20575 = n24954 ;
  assign y20576 = ~1'b0 ;
  assign y20577 = ~1'b0 ;
  assign y20578 = n37596 ;
  assign y20579 = ~n37598 ;
  assign y20580 = n37599 ;
  assign y20581 = ~n37603 ;
  assign y20582 = ~1'b0 ;
  assign y20583 = ~1'b0 ;
  assign y20584 = n37605 ;
  assign y20585 = ~1'b0 ;
  assign y20586 = ~1'b0 ;
  assign y20587 = ~n37609 ;
  assign y20588 = ~n37610 ;
  assign y20589 = n37611 ;
  assign y20590 = ~n37613 ;
  assign y20591 = n37616 ;
  assign y20592 = ~n7420 ;
  assign y20593 = ~n37619 ;
  assign y20594 = ~1'b0 ;
  assign y20595 = ~1'b0 ;
  assign y20596 = ~1'b0 ;
  assign y20597 = n37620 ;
  assign y20598 = n31659 ;
  assign y20599 = ~1'b0 ;
  assign y20600 = n37622 ;
  assign y20601 = ~1'b0 ;
  assign y20602 = ~1'b0 ;
  assign y20603 = ~n37624 ;
  assign y20604 = ~1'b0 ;
  assign y20605 = ~1'b0 ;
  assign y20606 = ~1'b0 ;
  assign y20607 = ~n37629 ;
  assign y20608 = ~n37636 ;
  assign y20609 = 1'b0 ;
  assign y20610 = ~n31735 ;
  assign y20611 = n37638 ;
  assign y20612 = ~n37639 ;
  assign y20613 = ~1'b0 ;
  assign y20614 = ~1'b0 ;
  assign y20615 = n37645 ;
  assign y20616 = ~n37651 ;
  assign y20617 = ~n37653 ;
  assign y20618 = ~n37656 ;
  assign y20619 = n37657 ;
  assign y20620 = ~n37659 ;
  assign y20621 = n37662 ;
  assign y20622 = n18959 ;
  assign y20623 = ~n37663 ;
  assign y20624 = n37666 ;
  assign y20625 = ~n37669 ;
  assign y20626 = ~n37672 ;
  assign y20627 = ~1'b0 ;
  assign y20628 = n37673 ;
  assign y20629 = n37676 ;
  assign y20630 = ~n37678 ;
  assign y20631 = ~1'b0 ;
  assign y20632 = ~1'b0 ;
  assign y20633 = n37679 ;
  assign y20634 = ~1'b0 ;
  assign y20635 = n37682 ;
  assign y20636 = ~1'b0 ;
  assign y20637 = n37686 ;
  assign y20638 = ~n37689 ;
  assign y20639 = ~n26527 ;
  assign y20640 = n37690 ;
  assign y20641 = ~n37691 ;
  assign y20642 = n37693 ;
  assign y20643 = ~1'b0 ;
  assign y20644 = ~1'b0 ;
  assign y20645 = ~1'b0 ;
  assign y20646 = n37695 ;
  assign y20647 = ~n37698 ;
  assign y20648 = n37699 ;
  assign y20649 = ~n37700 ;
  assign y20650 = n37701 ;
  assign y20651 = ~1'b0 ;
  assign y20652 = n37703 ;
  assign y20653 = n37704 ;
  assign y20654 = n37706 ;
  assign y20655 = n37712 ;
  assign y20656 = n37713 ;
  assign y20657 = ~n37714 ;
  assign y20658 = n11476 ;
  assign y20659 = ~n37717 ;
  assign y20660 = ~n37719 ;
  assign y20661 = ~1'b0 ;
  assign y20662 = ~1'b0 ;
  assign y20663 = ~n37722 ;
  assign y20664 = n37724 ;
  assign y20665 = n37728 ;
  assign y20666 = ~n37732 ;
  assign y20667 = n37736 ;
  assign y20668 = ~n37738 ;
  assign y20669 = ~1'b0 ;
  assign y20670 = ~1'b0 ;
  assign y20671 = ~n37739 ;
  assign y20672 = ~1'b0 ;
  assign y20673 = ~1'b0 ;
  assign y20674 = n37740 ;
  assign y20675 = ~n37745 ;
  assign y20676 = ~n37747 ;
  assign y20677 = n37749 ;
  assign y20678 = ~1'b0 ;
  assign y20679 = n37750 ;
  assign y20680 = ~n37752 ;
  assign y20681 = ~1'b0 ;
  assign y20682 = ~n37756 ;
  assign y20683 = ~1'b0 ;
  assign y20684 = ~n37757 ;
  assign y20685 = ~1'b0 ;
  assign y20686 = ~n19081 ;
  assign y20687 = ~1'b0 ;
  assign y20688 = ~n37761 ;
  assign y20689 = ~n6654 ;
  assign y20690 = n37762 ;
  assign y20691 = n37763 ;
  assign y20692 = ~n37764 ;
  assign y20693 = ~1'b0 ;
  assign y20694 = n37766 ;
  assign y20695 = ~n18086 ;
  assign y20696 = n37767 ;
  assign y20697 = n37776 ;
  assign y20698 = n37777 ;
  assign y20699 = ~1'b0 ;
  assign y20700 = n37780 ;
  assign y20701 = ~n37781 ;
  assign y20702 = n37782 ;
  assign y20703 = ~1'b0 ;
  assign y20704 = n20501 ;
  assign y20705 = n37783 ;
  assign y20706 = ~1'b0 ;
  assign y20707 = ~1'b0 ;
  assign y20708 = n37784 ;
  assign y20709 = 1'b0 ;
  assign y20710 = ~n37788 ;
  assign y20711 = ~1'b0 ;
  assign y20712 = ~n37789 ;
  assign y20713 = n37790 ;
  assign y20714 = n37791 ;
  assign y20715 = ~1'b0 ;
  assign y20716 = n37801 ;
  assign y20717 = ~n37803 ;
  assign y20718 = n37806 ;
  assign y20719 = ~1'b0 ;
  assign y20720 = ~1'b0 ;
  assign y20721 = ~n37807 ;
  assign y20722 = ~n37808 ;
  assign y20723 = ~n37812 ;
  assign y20724 = n37813 ;
  assign y20725 = ~n37815 ;
  assign y20726 = ~n37816 ;
  assign y20727 = ~n37819 ;
  assign y20728 = ~1'b0 ;
  assign y20729 = ~n37820 ;
  assign y20730 = ~n37822 ;
  assign y20731 = ~1'b0 ;
  assign y20732 = n37826 ;
  assign y20733 = n18310 ;
  assign y20734 = ~1'b0 ;
  assign y20735 = ~n37829 ;
  assign y20736 = n37831 ;
  assign y20737 = ~1'b0 ;
  assign y20738 = ~n37833 ;
  assign y20739 = ~1'b0 ;
  assign y20740 = ~1'b0 ;
  assign y20741 = ~n37834 ;
  assign y20742 = ~n37835 ;
  assign y20743 = ~n37836 ;
  assign y20744 = ~1'b0 ;
  assign y20745 = n37837 ;
  assign y20746 = ~1'b0 ;
  assign y20747 = ~n14571 ;
  assign y20748 = ~1'b0 ;
  assign y20749 = ~1'b0 ;
  assign y20750 = ~1'b0 ;
  assign y20751 = ~n37838 ;
  assign y20752 = ~n37840 ;
  assign y20753 = ~1'b0 ;
  assign y20754 = 1'b0 ;
  assign y20755 = ~n37842 ;
  assign y20756 = n37845 ;
  assign y20757 = n37846 ;
  assign y20758 = n37849 ;
  assign y20759 = ~n16008 ;
  assign y20760 = ~1'b0 ;
  assign y20761 = n37851 ;
  assign y20762 = ~n37852 ;
  assign y20763 = n37854 ;
  assign y20764 = n37857 ;
  assign y20765 = ~1'b0 ;
  assign y20766 = ~n37858 ;
  assign y20767 = n37860 ;
  assign y20768 = ~1'b0 ;
  assign y20769 = ~1'b0 ;
  assign y20770 = ~n16037 ;
  assign y20771 = ~n37861 ;
  assign y20772 = ~n37871 ;
  assign y20773 = n37875 ;
  assign y20774 = n17369 ;
  assign y20775 = ~1'b0 ;
  assign y20776 = ~1'b0 ;
  assign y20777 = ~1'b0 ;
  assign y20778 = ~n37883 ;
  assign y20779 = n37884 ;
  assign y20780 = ~n37885 ;
  assign y20781 = n37887 ;
  assign y20782 = ~n37890 ;
  assign y20783 = ~n37892 ;
  assign y20784 = ~n37893 ;
  assign y20785 = n688 ;
  assign y20786 = n37897 ;
  assign y20787 = ~n37898 ;
  assign y20788 = 1'b0 ;
  assign y20789 = ~1'b0 ;
  assign y20790 = n37899 ;
  assign y20791 = ~n37906 ;
  assign y20792 = ~n37907 ;
  assign y20793 = ~1'b0 ;
  assign y20794 = n37909 ;
  assign y20795 = n37911 ;
  assign y20796 = ~1'b0 ;
  assign y20797 = n37914 ;
  assign y20798 = ~1'b0 ;
  assign y20799 = n37917 ;
  assign y20800 = ~1'b0 ;
  assign y20801 = n37918 ;
  assign y20802 = ~n37921 ;
  assign y20803 = ~n37923 ;
  assign y20804 = ~n37926 ;
  assign y20805 = n37930 ;
  assign y20806 = ~1'b0 ;
  assign y20807 = ~n37933 ;
  assign y20808 = ~1'b0 ;
  assign y20809 = ~n37938 ;
  assign y20810 = n37940 ;
  assign y20811 = n37941 ;
  assign y20812 = ~1'b0 ;
  assign y20813 = ~n37943 ;
  assign y20814 = ~1'b0 ;
  assign y20815 = ~n37946 ;
  assign y20816 = n37947 ;
  assign y20817 = ~n37950 ;
  assign y20818 = n37952 ;
  assign y20819 = ~1'b0 ;
  assign y20820 = ~n37956 ;
  assign y20821 = ~x203 ;
  assign y20822 = ~n37957 ;
  assign y20823 = ~n37958 ;
  assign y20824 = n37961 ;
  assign y20825 = n37962 ;
  assign y20826 = ~1'b0 ;
  assign y20827 = ~1'b0 ;
  assign y20828 = ~1'b0 ;
  assign y20829 = n4986 ;
  assign y20830 = ~n37965 ;
  assign y20831 = ~n37968 ;
  assign y20832 = n4255 ;
  assign y20833 = ~n37975 ;
  assign y20834 = ~n37977 ;
  assign y20835 = ~n37978 ;
  assign y20836 = n37982 ;
  assign y20837 = ~n37983 ;
  assign y20838 = ~n37985 ;
  assign y20839 = n37988 ;
  assign y20840 = 1'b0 ;
  assign y20841 = ~1'b0 ;
  assign y20842 = ~n37991 ;
  assign y20843 = ~n37992 ;
  assign y20844 = n37997 ;
  assign y20845 = ~n37999 ;
  assign y20846 = ~n38003 ;
  assign y20847 = ~n38004 ;
  assign y20848 = ~n38010 ;
  assign y20849 = ~n38012 ;
  assign y20850 = ~1'b0 ;
  assign y20851 = n38013 ;
  assign y20852 = n38014 ;
  assign y20853 = n38017 ;
  assign y20854 = n38019 ;
  assign y20855 = ~1'b0 ;
  assign y20856 = ~n38022 ;
  assign y20857 = n19645 ;
  assign y20858 = n38026 ;
  assign y20859 = ~n38027 ;
  assign y20860 = ~1'b0 ;
  assign y20861 = n38029 ;
  assign y20862 = ~n38031 ;
  assign y20863 = ~n38033 ;
  assign y20864 = n38034 ;
  assign y20865 = ~1'b0 ;
  assign y20866 = ~1'b0 ;
  assign y20867 = ~n38036 ;
  assign y20868 = n38038 ;
  assign y20869 = ~n11453 ;
  assign y20870 = ~n38040 ;
  assign y20871 = ~1'b0 ;
  assign y20872 = ~1'b0 ;
  assign y20873 = ~1'b0 ;
  assign y20874 = n38042 ;
  assign y20875 = 1'b0 ;
  assign y20876 = n38044 ;
  assign y20877 = 1'b0 ;
  assign y20878 = ~1'b0 ;
  assign y20879 = ~n38045 ;
  assign y20880 = n38046 ;
  assign y20881 = ~n38048 ;
  assign y20882 = n38049 ;
  assign y20883 = ~1'b0 ;
  assign y20884 = ~n38053 ;
  assign y20885 = 1'b0 ;
  assign y20886 = n38057 ;
  assign y20887 = ~n38059 ;
  assign y20888 = n38060 ;
  assign y20889 = ~1'b0 ;
  assign y20890 = n38061 ;
  assign y20891 = ~n38062 ;
  assign y20892 = n38063 ;
  assign y20893 = ~1'b0 ;
  assign y20894 = ~1'b0 ;
  assign y20895 = ~n38065 ;
  assign y20896 = n38067 ;
  assign y20897 = ~1'b0 ;
  assign y20898 = ~n38070 ;
  assign y20899 = ~n38075 ;
  assign y20900 = ~n38079 ;
  assign y20901 = ~n38081 ;
  assign y20902 = ~n9204 ;
  assign y20903 = n38083 ;
  assign y20904 = ~1'b0 ;
  assign y20905 = ~n38086 ;
  assign y20906 = ~n38088 ;
  assign y20907 = ~1'b0 ;
  assign y20908 = n38094 ;
  assign y20909 = ~n38095 ;
  assign y20910 = ~n38100 ;
  assign y20911 = ~1'b0 ;
  assign y20912 = ~1'b0 ;
  assign y20913 = ~n38104 ;
  assign y20914 = ~1'b0 ;
  assign y20915 = ~n38106 ;
  assign y20916 = ~1'b0 ;
  assign y20917 = n38107 ;
  assign y20918 = ~1'b0 ;
  assign y20919 = n38108 ;
  assign y20920 = ~n2182 ;
  assign y20921 = ~1'b0 ;
  assign y20922 = n18900 ;
  assign y20923 = ~1'b0 ;
  assign y20924 = ~1'b0 ;
  assign y20925 = ~n38110 ;
  assign y20926 = ~n38114 ;
  assign y20927 = n38118 ;
  assign y20928 = ~n38119 ;
  assign y20929 = n38122 ;
  assign y20930 = ~n38125 ;
  assign y20931 = ~n38127 ;
  assign y20932 = ~n38132 ;
  assign y20933 = ~n38135 ;
  assign y20934 = ~n38136 ;
  assign y20935 = ~1'b0 ;
  assign y20936 = ~n38138 ;
  assign y20937 = ~1'b0 ;
  assign y20938 = ~1'b0 ;
  assign y20939 = n3265 ;
  assign y20940 = n38139 ;
  assign y20941 = ~1'b0 ;
  assign y20942 = n38140 ;
  assign y20943 = ~1'b0 ;
  assign y20944 = ~n38141 ;
  assign y20945 = ~n38143 ;
  assign y20946 = ~1'b0 ;
  assign y20947 = ~n38144 ;
  assign y20948 = ~n38146 ;
  assign y20949 = n38148 ;
  assign y20950 = n38153 ;
  assign y20951 = ~n38154 ;
  assign y20952 = ~n38159 ;
  assign y20953 = ~n38161 ;
  assign y20954 = n38163 ;
  assign y20955 = ~n38165 ;
  assign y20956 = ~n38166 ;
  assign y20957 = ~n37719 ;
  assign y20958 = ~n38169 ;
  assign y20959 = ~1'b0 ;
  assign y20960 = n38174 ;
  assign y20961 = ~n38177 ;
  assign y20962 = ~n38178 ;
  assign y20963 = ~n38179 ;
  assign y20964 = ~n38181 ;
  assign y20965 = ~1'b0 ;
  assign y20966 = ~1'b0 ;
  assign y20967 = ~n38182 ;
  assign y20968 = 1'b0 ;
  assign y20969 = ~n38186 ;
  assign y20970 = ~1'b0 ;
  assign y20971 = ~n38188 ;
  assign y20972 = n38189 ;
  assign y20973 = n38190 ;
  assign y20974 = ~1'b0 ;
  assign y20975 = ~1'b0 ;
  assign y20976 = n38191 ;
  assign y20977 = ~1'b0 ;
  assign y20978 = ~1'b0 ;
  assign y20979 = ~1'b0 ;
  assign y20980 = ~1'b0 ;
  assign y20981 = n38193 ;
  assign y20982 = ~1'b0 ;
  assign y20983 = n38196 ;
  assign y20984 = ~n38197 ;
  assign y20985 = ~n38198 ;
  assign y20986 = n38202 ;
  assign y20987 = n38207 ;
  assign y20988 = ~n38212 ;
  assign y20989 = n38213 ;
  assign y20990 = ~1'b0 ;
  assign y20991 = ~n38225 ;
  assign y20992 = ~1'b0 ;
  assign y20993 = ~1'b0 ;
  assign y20994 = ~n38227 ;
  assign y20995 = ~n38229 ;
  assign y20996 = ~1'b0 ;
  assign y20997 = ~1'b0 ;
  assign y20998 = n38230 ;
  assign y20999 = n38231 ;
  assign y21000 = ~n38232 ;
  assign y21001 = ~1'b0 ;
  assign y21002 = n38233 ;
  assign y21003 = 1'b0 ;
  assign y21004 = n38236 ;
  assign y21005 = ~n38237 ;
  assign y21006 = n38242 ;
  assign y21007 = n38243 ;
  assign y21008 = n38244 ;
  assign y21009 = n38245 ;
  assign y21010 = n38247 ;
  assign y21011 = ~n38249 ;
  assign y21012 = ~n38250 ;
  assign y21013 = ~1'b0 ;
  assign y21014 = n38252 ;
  assign y21015 = ~1'b0 ;
  assign y21016 = ~n38253 ;
  assign y21017 = n38255 ;
  assign y21018 = ~1'b0 ;
  assign y21019 = ~1'b0 ;
  assign y21020 = ~1'b0 ;
  assign y21021 = ~n38257 ;
  assign y21022 = ~1'b0 ;
  assign y21023 = ~1'b0 ;
  assign y21024 = ~n38258 ;
  assign y21025 = n38266 ;
  assign y21026 = n38267 ;
  assign y21027 = n38268 ;
  assign y21028 = n38271 ;
  assign y21029 = n38273 ;
  assign y21030 = ~1'b0 ;
  assign y21031 = n38275 ;
  assign y21032 = ~1'b0 ;
  assign y21033 = ~n38279 ;
  assign y21034 = n38280 ;
  assign y21035 = ~1'b0 ;
  assign y21036 = ~n38283 ;
  assign y21037 = ~n38285 ;
  assign y21038 = ~n38289 ;
  assign y21039 = ~1'b0 ;
  assign y21040 = ~n38294 ;
  assign y21041 = n38296 ;
  assign y21042 = n38299 ;
  assign y21043 = ~n38300 ;
  assign y21044 = n38302 ;
  assign y21045 = ~1'b0 ;
  assign y21046 = ~n38303 ;
  assign y21047 = n38307 ;
  assign y21048 = n38308 ;
  assign y21049 = ~n38309 ;
  assign y21050 = ~1'b0 ;
  assign y21051 = ~1'b0 ;
  assign y21052 = n631 ;
  assign y21053 = ~n38310 ;
  assign y21054 = ~1'b0 ;
  assign y21055 = ~n38311 ;
  assign y21056 = n38315 ;
  assign y21057 = n38317 ;
  assign y21058 = ~n38319 ;
  assign y21059 = ~1'b0 ;
  assign y21060 = ~n38321 ;
  assign y21061 = n38322 ;
  assign y21062 = ~n38323 ;
  assign y21063 = ~n38324 ;
  assign y21064 = ~1'b0 ;
  assign y21065 = n38325 ;
  assign y21066 = ~1'b0 ;
  assign y21067 = ~n38327 ;
  assign y21068 = ~n38330 ;
  assign y21069 = ~1'b0 ;
  assign y21070 = ~n38332 ;
  assign y21071 = ~1'b0 ;
  assign y21072 = n21503 ;
  assign y21073 = n38338 ;
  assign y21074 = ~1'b0 ;
  assign y21075 = ~n38339 ;
  assign y21076 = ~1'b0 ;
  assign y21077 = ~1'b0 ;
  assign y21078 = ~1'b0 ;
  assign y21079 = ~n38340 ;
  assign y21080 = n38341 ;
  assign y21081 = ~1'b0 ;
  assign y21082 = ~n38345 ;
  assign y21083 = n38347 ;
  assign y21084 = ~1'b0 ;
  assign y21085 = ~1'b0 ;
  assign y21086 = n38114 ;
  assign y21087 = ~1'b0 ;
  assign y21088 = ~1'b0 ;
  assign y21089 = n38350 ;
  assign y21090 = ~1'b0 ;
  assign y21091 = ~n38353 ;
  assign y21092 = ~1'b0 ;
  assign y21093 = n38354 ;
  assign y21094 = n38355 ;
  assign y21095 = n38357 ;
  assign y21096 = 1'b0 ;
  assign y21097 = ~1'b0 ;
  assign y21098 = ~1'b0 ;
  assign y21099 = n8813 ;
  assign y21100 = 1'b0 ;
  assign y21101 = n38359 ;
  assign y21102 = ~1'b0 ;
  assign y21103 = n32028 ;
  assign y21104 = ~n38360 ;
  assign y21105 = ~n38361 ;
  assign y21106 = ~n38364 ;
  assign y21107 = n38365 ;
  assign y21108 = ~n38369 ;
  assign y21109 = ~n29050 ;
  assign y21110 = n38370 ;
  assign y21111 = ~1'b0 ;
  assign y21112 = ~1'b0 ;
  assign y21113 = n38372 ;
  assign y21114 = ~n38373 ;
  assign y21115 = ~n38374 ;
  assign y21116 = ~n38375 ;
  assign y21117 = ~1'b0 ;
  assign y21118 = ~n5565 ;
  assign y21119 = ~1'b0 ;
  assign y21120 = ~1'b0 ;
  assign y21121 = ~1'b0 ;
  assign y21122 = n38376 ;
  assign y21123 = n38377 ;
  assign y21124 = ~n38378 ;
  assign y21125 = n38379 ;
  assign y21126 = ~n38380 ;
  assign y21127 = ~n38382 ;
  assign y21128 = ~n38384 ;
  assign y21129 = ~n38386 ;
  assign y21130 = n38388 ;
  assign y21131 = n38389 ;
  assign y21132 = ~1'b0 ;
  assign y21133 = ~1'b0 ;
  assign y21134 = n38390 ;
  assign y21135 = ~1'b0 ;
  assign y21136 = ~1'b0 ;
  assign y21137 = ~1'b0 ;
  assign y21138 = ~n38393 ;
  assign y21139 = ~n38398 ;
  assign y21140 = n38400 ;
  assign y21141 = ~1'b0 ;
  assign y21142 = n38402 ;
  assign y21143 = ~n38405 ;
  assign y21144 = ~n38410 ;
  assign y21145 = ~n38413 ;
  assign y21146 = ~n38415 ;
  assign y21147 = ~1'b0 ;
  assign y21148 = ~1'b0 ;
  assign y21149 = n38416 ;
  assign y21150 = n38421 ;
  assign y21151 = ~n33936 ;
  assign y21152 = n38422 ;
  assign y21153 = ~n38423 ;
  assign y21154 = n38424 ;
  assign y21155 = ~1'b0 ;
  assign y21156 = ~n27619 ;
  assign y21157 = n38428 ;
  assign y21158 = ~1'b0 ;
  assign y21159 = ~1'b0 ;
  assign y21160 = ~n38431 ;
  assign y21161 = n38433 ;
  assign y21162 = n38435 ;
  assign y21163 = n38439 ;
  assign y21164 = ~n819 ;
  assign y21165 = ~1'b0 ;
  assign y21166 = n38440 ;
  assign y21167 = n38442 ;
  assign y21168 = ~n38443 ;
  assign y21169 = ~n38446 ;
  assign y21170 = ~1'b0 ;
  assign y21171 = n38448 ;
  assign y21172 = n38449 ;
  assign y21173 = ~n38450 ;
  assign y21174 = ~1'b0 ;
  assign y21175 = ~n38451 ;
  assign y21176 = ~n38453 ;
  assign y21177 = ~1'b0 ;
  assign y21178 = n38454 ;
  assign y21179 = n38455 ;
  assign y21180 = ~1'b0 ;
  assign y21181 = ~n38457 ;
  assign y21182 = ~1'b0 ;
  assign y21183 = ~n38458 ;
  assign y21184 = ~1'b0 ;
  assign y21185 = n38459 ;
  assign y21186 = n38463 ;
  assign y21187 = ~1'b0 ;
  assign y21188 = ~n38465 ;
  assign y21189 = ~1'b0 ;
  assign y21190 = ~1'b0 ;
  assign y21191 = n38469 ;
  assign y21192 = ~n32395 ;
  assign y21193 = n38472 ;
  assign y21194 = n38473 ;
  assign y21195 = ~1'b0 ;
  assign y21196 = ~1'b0 ;
  assign y21197 = ~1'b0 ;
  assign y21198 = ~1'b0 ;
  assign y21199 = n38474 ;
  assign y21200 = ~n34795 ;
  assign y21201 = n38475 ;
  assign y21202 = ~n38477 ;
  assign y21203 = n38478 ;
  assign y21204 = ~1'b0 ;
  assign y21205 = ~1'b0 ;
  assign y21206 = n38481 ;
  assign y21207 = n38484 ;
  assign y21208 = ~n38486 ;
  assign y21209 = n38489 ;
  assign y21210 = ~1'b0 ;
  assign y21211 = n38490 ;
  assign y21212 = n38493 ;
  assign y21213 = n22447 ;
  assign y21214 = n28925 ;
  assign y21215 = ~1'b0 ;
  assign y21216 = ~1'b0 ;
  assign y21217 = ~n38500 ;
  assign y21218 = 1'b0 ;
  assign y21219 = ~1'b0 ;
  assign y21220 = n38504 ;
  assign y21221 = n38505 ;
  assign y21222 = n38506 ;
  assign y21223 = ~n38509 ;
  assign y21224 = ~n38512 ;
  assign y21225 = n38514 ;
  assign y21226 = ~n38515 ;
  assign y21227 = n38516 ;
  assign y21228 = ~n38520 ;
  assign y21229 = ~1'b0 ;
  assign y21230 = n38522 ;
  assign y21231 = ~n38524 ;
  assign y21232 = n38526 ;
  assign y21233 = n38527 ;
  assign y21234 = n38534 ;
  assign y21235 = n38536 ;
  assign y21236 = n38538 ;
  assign y21237 = ~1'b0 ;
  assign y21238 = ~n38539 ;
  assign y21239 = ~n38543 ;
  assign y21240 = n38548 ;
  assign y21241 = ~1'b0 ;
  assign y21242 = ~n2593 ;
  assign y21243 = ~n38549 ;
  assign y21244 = ~n38551 ;
  assign y21245 = ~1'b0 ;
  assign y21246 = ~1'b0 ;
  assign y21247 = 1'b0 ;
  assign y21248 = ~n38552 ;
  assign y21249 = n38556 ;
  assign y21250 = ~n38558 ;
  assign y21251 = ~n38560 ;
  assign y21252 = ~n38561 ;
  assign y21253 = n838 ;
  assign y21254 = ~n38565 ;
  assign y21255 = n38568 ;
  assign y21256 = n38570 ;
  assign y21257 = ~n38575 ;
  assign y21258 = ~n38577 ;
  assign y21259 = ~1'b0 ;
  assign y21260 = ~n38578 ;
  assign y21261 = ~n38579 ;
  assign y21262 = n38581 ;
  assign y21263 = ~1'b0 ;
  assign y21264 = ~1'b0 ;
  assign y21265 = n38582 ;
  assign y21266 = n38583 ;
  assign y21267 = ~n38593 ;
  assign y21268 = ~1'b0 ;
  assign y21269 = ~n38596 ;
  assign y21270 = n38597 ;
  assign y21271 = n38601 ;
  assign y21272 = ~n38602 ;
  assign y21273 = ~1'b0 ;
  assign y21274 = ~1'b0 ;
  assign y21275 = ~1'b0 ;
  assign y21276 = n38603 ;
  assign y21277 = n38604 ;
  assign y21278 = n16794 ;
  assign y21279 = ~n38605 ;
  assign y21280 = n38608 ;
  assign y21281 = ~1'b0 ;
  assign y21282 = ~1'b0 ;
  assign y21283 = ~1'b0 ;
  assign y21284 = ~1'b0 ;
  assign y21285 = n38609 ;
  assign y21286 = n38610 ;
  assign y21287 = n38612 ;
  assign y21288 = ~n6352 ;
  assign y21289 = n38613 ;
  assign y21290 = ~n38614 ;
  assign y21291 = n38618 ;
  assign y21292 = ~n38619 ;
  assign y21293 = n38621 ;
  assign y21294 = ~1'b0 ;
  assign y21295 = n38622 ;
  assign y21296 = ~1'b0 ;
  assign y21297 = ~n38623 ;
  assign y21298 = ~1'b0 ;
  assign y21299 = n38626 ;
  assign y21300 = ~n38629 ;
  assign y21301 = n38631 ;
  assign y21302 = ~1'b0 ;
  assign y21303 = ~1'b0 ;
  assign y21304 = ~n38634 ;
  assign y21305 = ~1'b0 ;
  assign y21306 = ~n38636 ;
  assign y21307 = ~n38639 ;
  assign y21308 = ~1'b0 ;
  assign y21309 = n38641 ;
  assign y21310 = n38642 ;
  assign y21311 = n38650 ;
  assign y21312 = ~1'b0 ;
  assign y21313 = n38651 ;
  assign y21314 = ~n38654 ;
  assign y21315 = ~n38656 ;
  assign y21316 = ~1'b0 ;
  assign y21317 = n38657 ;
  assign y21318 = n38659 ;
  assign y21319 = ~1'b0 ;
  assign y21320 = ~n38662 ;
  assign y21321 = n6145 ;
  assign y21322 = ~n2286 ;
  assign y21323 = n38663 ;
  assign y21324 = ~1'b0 ;
  assign y21325 = n38664 ;
  assign y21326 = ~1'b0 ;
  assign y21327 = n38668 ;
  assign y21328 = ~1'b0 ;
  assign y21329 = ~1'b0 ;
  assign y21330 = n38669 ;
  assign y21331 = n38670 ;
  assign y21332 = ~1'b0 ;
  assign y21333 = ~n38672 ;
  assign y21334 = ~1'b0 ;
  assign y21335 = ~1'b0 ;
  assign y21336 = ~n38674 ;
  assign y21337 = ~1'b0 ;
  assign y21338 = ~1'b0 ;
  assign y21339 = n38677 ;
  assign y21340 = ~n38678 ;
  assign y21341 = ~n38683 ;
  assign y21342 = ~1'b0 ;
  assign y21343 = ~n38686 ;
  assign y21344 = ~n38687 ;
  assign y21345 = ~n38692 ;
  assign y21346 = ~n38694 ;
  assign y21347 = ~1'b0 ;
  assign y21348 = ~n38697 ;
  assign y21349 = ~n38698 ;
  assign y21350 = ~n38700 ;
  assign y21351 = ~n38701 ;
  assign y21352 = n38704 ;
  assign y21353 = n29568 ;
  assign y21354 = ~n38709 ;
  assign y21355 = n38710 ;
  assign y21356 = ~n38713 ;
  assign y21357 = ~n38715 ;
  assign y21358 = ~n38717 ;
  assign y21359 = n38719 ;
  assign y21360 = ~1'b0 ;
  assign y21361 = ~n38722 ;
  assign y21362 = ~1'b0 ;
  assign y21363 = ~n38725 ;
  assign y21364 = ~n38727 ;
  assign y21365 = ~1'b0 ;
  assign y21366 = ~n38729 ;
  assign y21367 = ~1'b0 ;
  assign y21368 = ~1'b0 ;
  assign y21369 = ~1'b0 ;
  assign y21370 = n38733 ;
  assign y21371 = n38734 ;
  assign y21372 = n38737 ;
  assign y21373 = ~1'b0 ;
  assign y21374 = ~1'b0 ;
  assign y21375 = ~n38739 ;
  assign y21376 = ~1'b0 ;
  assign y21377 = ~1'b0 ;
  assign y21378 = ~n38741 ;
  assign y21379 = n38743 ;
  assign y21380 = ~1'b0 ;
  assign y21381 = ~n38745 ;
  assign y21382 = ~1'b0 ;
  assign y21383 = ~n11689 ;
  assign y21384 = ~n38747 ;
  assign y21385 = ~1'b0 ;
  assign y21386 = ~n38748 ;
  assign y21387 = n38749 ;
  assign y21388 = n38755 ;
  assign y21389 = n38756 ;
  assign y21390 = n38758 ;
  assign y21391 = n38759 ;
  assign y21392 = n38760 ;
  assign y21393 = ~n38762 ;
  assign y21394 = n38763 ;
  assign y21395 = ~1'b0 ;
  assign y21396 = ~1'b0 ;
  assign y21397 = ~n38767 ;
  assign y21398 = ~1'b0 ;
  assign y21399 = 1'b0 ;
  assign y21400 = ~1'b0 ;
  assign y21401 = ~1'b0 ;
  assign y21402 = n38768 ;
  assign y21403 = ~n29150 ;
  assign y21404 = ~1'b0 ;
  assign y21405 = ~1'b0 ;
  assign y21406 = ~1'b0 ;
  assign y21407 = n38771 ;
  assign y21408 = 1'b0 ;
  assign y21409 = ~1'b0 ;
  assign y21410 = n38774 ;
  assign y21411 = n2939 ;
  assign y21412 = ~n38775 ;
  assign y21413 = ~n38777 ;
  assign y21414 = ~1'b0 ;
  assign y21415 = ~1'b0 ;
  assign y21416 = ~1'b0 ;
  assign y21417 = ~n38782 ;
  assign y21418 = ~n38198 ;
  assign y21419 = ~n38784 ;
  assign y21420 = ~1'b0 ;
  assign y21421 = ~n18700 ;
  assign y21422 = ~n38785 ;
  assign y21423 = n38786 ;
  assign y21424 = ~1'b0 ;
  assign y21425 = ~n38788 ;
  assign y21426 = ~n38790 ;
  assign y21427 = ~n38792 ;
  assign y21428 = n38793 ;
  assign y21429 = n38795 ;
  assign y21430 = n38797 ;
  assign y21431 = ~n38804 ;
  assign y21432 = ~n38805 ;
  assign y21433 = n38806 ;
  assign y21434 = ~n38808 ;
  assign y21435 = ~n38812 ;
  assign y21436 = ~n38818 ;
  assign y21437 = ~n38820 ;
  assign y21438 = ~1'b0 ;
  assign y21439 = n38825 ;
  assign y21440 = ~n38831 ;
  assign y21441 = ~1'b0 ;
  assign y21442 = ~n9070 ;
  assign y21443 = ~n38832 ;
  assign y21444 = ~1'b0 ;
  assign y21445 = n38833 ;
  assign y21446 = ~n38837 ;
  assign y21447 = ~n38841 ;
  assign y21448 = ~1'b0 ;
  assign y21449 = ~1'b0 ;
  assign y21450 = n38842 ;
  assign y21451 = n38847 ;
  assign y21452 = ~n38848 ;
  assign y21453 = ~n38849 ;
  assign y21454 = n38851 ;
  assign y21455 = ~1'b0 ;
  assign y21456 = n38853 ;
  assign y21457 = ~1'b0 ;
  assign y21458 = ~1'b0 ;
  assign y21459 = ~1'b0 ;
  assign y21460 = ~1'b0 ;
  assign y21461 = n11345 ;
  assign y21462 = n38854 ;
  assign y21463 = 1'b0 ;
  assign y21464 = n38855 ;
  assign y21465 = 1'b0 ;
  assign y21466 = n38856 ;
  assign y21467 = ~1'b0 ;
  assign y21468 = ~1'b0 ;
  assign y21469 = ~n38861 ;
  assign y21470 = n38863 ;
  assign y21471 = n38864 ;
  assign y21472 = n38865 ;
  assign y21473 = n38871 ;
  assign y21474 = n38873 ;
  assign y21475 = 1'b0 ;
  assign y21476 = ~1'b0 ;
  assign y21477 = ~1'b0 ;
  assign y21478 = ~1'b0 ;
  assign y21479 = ~1'b0 ;
  assign y21480 = ~1'b0 ;
  assign y21481 = ~1'b0 ;
  assign y21482 = ~1'b0 ;
  assign y21483 = n38874 ;
  assign y21484 = n38875 ;
  assign y21485 = n38876 ;
  assign y21486 = ~1'b0 ;
  assign y21487 = ~n38879 ;
  assign y21488 = n262 ;
  assign y21489 = ~n38881 ;
  assign y21490 = ~1'b0 ;
  assign y21491 = ~1'b0 ;
  assign y21492 = ~n38888 ;
  assign y21493 = ~n38889 ;
  assign y21494 = ~n38891 ;
  assign y21495 = ~1'b0 ;
  assign y21496 = ~n38893 ;
  assign y21497 = n12349 ;
  assign y21498 = ~1'b0 ;
  assign y21499 = ~1'b0 ;
  assign y21500 = ~1'b0 ;
  assign y21501 = n38894 ;
  assign y21502 = n38898 ;
  assign y21503 = n38899 ;
  assign y21504 = ~n38901 ;
  assign y21505 = ~1'b0 ;
  assign y21506 = ~n38903 ;
  assign y21507 = n38906 ;
  assign y21508 = ~1'b0 ;
  assign y21509 = ~n38907 ;
  assign y21510 = n38909 ;
  assign y21511 = n38911 ;
  assign y21512 = 1'b0 ;
  assign y21513 = ~1'b0 ;
  assign y21514 = ~1'b0 ;
  assign y21515 = ~n38912 ;
  assign y21516 = ~n38913 ;
  assign y21517 = ~n17302 ;
  assign y21518 = ~1'b0 ;
  assign y21519 = n38917 ;
  assign y21520 = ~n38919 ;
  assign y21521 = ~1'b0 ;
  assign y21522 = n1386 ;
  assign y21523 = n18399 ;
  assign y21524 = n38921 ;
  assign y21525 = ~n38923 ;
  assign y21526 = ~1'b0 ;
  assign y21527 = ~1'b0 ;
  assign y21528 = ~1'b0 ;
  assign y21529 = n38924 ;
  assign y21530 = n38927 ;
  assign y21531 = ~n38929 ;
  assign y21532 = ~n38934 ;
  assign y21533 = n38935 ;
  assign y21534 = ~1'b0 ;
  assign y21535 = ~n38941 ;
  assign y21536 = n38943 ;
  assign y21537 = ~1'b0 ;
  assign y21538 = n35369 ;
  assign y21539 = ~n38946 ;
  assign y21540 = ~1'b0 ;
  assign y21541 = ~n38951 ;
  assign y21542 = n38952 ;
  assign y21543 = ~1'b0 ;
  assign y21544 = ~n38956 ;
  assign y21545 = n38958 ;
  assign y21546 = ~1'b0 ;
  assign y21547 = ~n38959 ;
  assign y21548 = n38961 ;
  assign y21549 = n38962 ;
  assign y21550 = n38963 ;
  assign y21551 = ~1'b0 ;
  assign y21552 = ~n38968 ;
  assign y21553 = ~n38969 ;
  assign y21554 = n38972 ;
  assign y21555 = ~1'b0 ;
  assign y21556 = ~1'b0 ;
  assign y21557 = ~n38976 ;
  assign y21558 = ~1'b0 ;
  assign y21559 = n38979 ;
  assign y21560 = n38981 ;
  assign y21561 = n2296 ;
  assign y21562 = ~1'b0 ;
  assign y21563 = ~n38982 ;
  assign y21564 = 1'b0 ;
  assign y21565 = n20519 ;
  assign y21566 = n38983 ;
  assign y21567 = n38984 ;
  assign y21568 = ~n38985 ;
  assign y21569 = ~n38987 ;
  assign y21570 = ~1'b0 ;
  assign y21571 = ~1'b0 ;
  assign y21572 = ~1'b0 ;
  assign y21573 = n32170 ;
  assign y21574 = n38989 ;
  assign y21575 = x115 ;
  assign y21576 = n38994 ;
  assign y21577 = ~1'b0 ;
  assign y21578 = n38995 ;
  assign y21579 = ~n38996 ;
  assign y21580 = ~n38997 ;
  assign y21581 = n38998 ;
  assign y21582 = n38999 ;
  assign y21583 = ~n39001 ;
  assign y21584 = ~n39002 ;
  assign y21585 = ~1'b0 ;
  assign y21586 = ~1'b0 ;
  assign y21587 = 1'b0 ;
  assign y21588 = ~1'b0 ;
  assign y21589 = ~1'b0 ;
  assign y21590 = n39003 ;
  assign y21591 = n39005 ;
  assign y21592 = ~n39008 ;
  assign y21593 = 1'b0 ;
  assign y21594 = ~n39011 ;
  assign y21595 = n39014 ;
  assign y21596 = n39015 ;
  assign y21597 = ~1'b0 ;
  assign y21598 = n39019 ;
  assign y21599 = ~n39024 ;
  assign y21600 = ~1'b0 ;
  assign y21601 = ~n39026 ;
  assign y21602 = n39030 ;
  assign y21603 = n39031 ;
  assign y21604 = ~1'b0 ;
  assign y21605 = n39033 ;
  assign y21606 = n39035 ;
  assign y21607 = n39037 ;
  assign y21608 = n39038 ;
  assign y21609 = n39039 ;
  assign y21610 = n39042 ;
  assign y21611 = ~n39046 ;
  assign y21612 = ~n39050 ;
  assign y21613 = ~1'b0 ;
  assign y21614 = ~n39052 ;
  assign y21615 = ~1'b0 ;
  assign y21616 = ~n26263 ;
  assign y21617 = n39054 ;
  assign y21618 = ~1'b0 ;
  assign y21619 = ~n28511 ;
  assign y21620 = n39055 ;
  assign y21621 = ~n39058 ;
  assign y21622 = n39063 ;
  assign y21623 = ~1'b0 ;
  assign y21624 = ~n39064 ;
  assign y21625 = n39065 ;
  assign y21626 = ~n39067 ;
  assign y21627 = n39068 ;
  assign y21628 = ~n39075 ;
  assign y21629 = ~1'b0 ;
  assign y21630 = n39076 ;
  assign y21631 = n39077 ;
  assign y21632 = ~n39084 ;
  assign y21633 = ~1'b0 ;
  assign y21634 = n39085 ;
  assign y21635 = ~1'b0 ;
  assign y21636 = ~1'b0 ;
  assign y21637 = ~1'b0 ;
  assign y21638 = n39089 ;
  assign y21639 = n39093 ;
  assign y21640 = n39096 ;
  assign y21641 = ~n16603 ;
  assign y21642 = ~1'b0 ;
  assign y21643 = ~1'b0 ;
  assign y21644 = ~1'b0 ;
  assign y21645 = n17780 ;
  assign y21646 = n39098 ;
  assign y21647 = ~1'b0 ;
  assign y21648 = ~1'b0 ;
  assign y21649 = ~n39102 ;
  assign y21650 = n39104 ;
  assign y21651 = ~n39106 ;
  assign y21652 = ~n39108 ;
  assign y21653 = ~n39112 ;
  assign y21654 = ~1'b0 ;
  assign y21655 = ~n39116 ;
  assign y21656 = ~1'b0 ;
  assign y21657 = ~n39118 ;
  assign y21658 = ~n39120 ;
  assign y21659 = n39122 ;
  assign y21660 = ~1'b0 ;
  assign y21661 = n39124 ;
  assign y21662 = ~n39125 ;
  assign y21663 = 1'b0 ;
  assign y21664 = ~1'b0 ;
  assign y21665 = ~n12183 ;
  assign y21666 = 1'b0 ;
  assign y21667 = n39126 ;
  assign y21668 = ~1'b0 ;
  assign y21669 = ~n39127 ;
  assign y21670 = n16008 ;
  assign y21671 = ~1'b0 ;
  assign y21672 = n39131 ;
  assign y21673 = ~1'b0 ;
  assign y21674 = ~n39133 ;
  assign y21675 = ~1'b0 ;
  assign y21676 = ~1'b0 ;
  assign y21677 = ~1'b0 ;
  assign y21678 = n39135 ;
  assign y21679 = ~n39137 ;
  assign y21680 = ~1'b0 ;
  assign y21681 = ~n39138 ;
  assign y21682 = ~1'b0 ;
  assign y21683 = n39139 ;
  assign y21684 = n39142 ;
  assign y21685 = n39144 ;
  assign y21686 = ~1'b0 ;
  assign y21687 = n39147 ;
  assign y21688 = ~1'b0 ;
  assign y21689 = n7312 ;
  assign y21690 = ~n39149 ;
  assign y21691 = ~n39151 ;
  assign y21692 = 1'b0 ;
  assign y21693 = ~n39154 ;
  assign y21694 = 1'b0 ;
  assign y21695 = n39155 ;
  assign y21696 = n39156 ;
  assign y21697 = ~n3547 ;
  assign y21698 = ~1'b0 ;
  assign y21699 = ~n39159 ;
  assign y21700 = ~1'b0 ;
  assign y21701 = ~1'b0 ;
  assign y21702 = ~1'b0 ;
  assign y21703 = ~n39161 ;
  assign y21704 = n9744 ;
  assign y21705 = ~n39163 ;
  assign y21706 = n39164 ;
  assign y21707 = ~n39165 ;
  assign y21708 = ~n39166 ;
  assign y21709 = ~n39170 ;
  assign y21710 = ~1'b0 ;
  assign y21711 = ~n39171 ;
  assign y21712 = n39172 ;
  assign y21713 = 1'b0 ;
  assign y21714 = ~n39174 ;
  assign y21715 = ~1'b0 ;
  assign y21716 = ~n39178 ;
  assign y21717 = ~n39181 ;
  assign y21718 = ~1'b0 ;
  assign y21719 = n39182 ;
  assign y21720 = n39185 ;
  assign y21721 = ~n39187 ;
  assign y21722 = 1'b0 ;
  assign y21723 = n39188 ;
  assign y21724 = ~1'b0 ;
  assign y21725 = n18149 ;
  assign y21726 = n39194 ;
  assign y21727 = ~n39195 ;
  assign y21728 = n39197 ;
  assign y21729 = n39198 ;
  assign y21730 = ~n39201 ;
  assign y21731 = n39206 ;
  assign y21732 = ~1'b0 ;
  assign y21733 = n12133 ;
  assign y21734 = n39207 ;
  assign y21735 = ~1'b0 ;
  assign y21736 = n39210 ;
  assign y21737 = ~n39211 ;
  assign y21738 = n39212 ;
  assign y21739 = ~1'b0 ;
  assign y21740 = n39216 ;
  assign y21741 = n39218 ;
  assign y21742 = ~1'b0 ;
  assign y21743 = n39219 ;
  assign y21744 = ~1'b0 ;
  assign y21745 = ~n39225 ;
  assign y21746 = n39232 ;
  assign y21747 = n39233 ;
  assign y21748 = ~n8700 ;
  assign y21749 = ~1'b0 ;
  assign y21750 = ~n39235 ;
  assign y21751 = ~1'b0 ;
  assign y21752 = n39236 ;
  assign y21753 = n39240 ;
  assign y21754 = ~n39241 ;
  assign y21755 = ~n39242 ;
  assign y21756 = n39244 ;
  assign y21757 = n39249 ;
  assign y21758 = ~1'b0 ;
  assign y21759 = n14112 ;
  assign y21760 = n39252 ;
  assign y21761 = ~n39256 ;
  assign y21762 = n39258 ;
  assign y21763 = n39260 ;
  assign y21764 = ~1'b0 ;
  assign y21765 = ~1'b0 ;
  assign y21766 = n39261 ;
  assign y21767 = n39262 ;
  assign y21768 = ~n22416 ;
  assign y21769 = ~1'b0 ;
  assign y21770 = n39263 ;
  assign y21771 = ~n39266 ;
  assign y21772 = ~n39269 ;
  assign y21773 = n29524 ;
  assign y21774 = ~n39270 ;
  assign y21775 = n39271 ;
  assign y21776 = n39276 ;
  assign y21777 = n39279 ;
  assign y21778 = n39281 ;
  assign y21779 = ~1'b0 ;
  assign y21780 = ~1'b0 ;
  assign y21781 = ~1'b0 ;
  assign y21782 = ~n39284 ;
  assign y21783 = ~n39286 ;
  assign y21784 = n39292 ;
  assign y21785 = ~n39294 ;
  assign y21786 = n39295 ;
  assign y21787 = ~n39296 ;
  assign y21788 = n39299 ;
  assign y21789 = n39301 ;
  assign y21790 = ~1'b0 ;
  assign y21791 = ~1'b0 ;
  assign y21792 = n2916 ;
  assign y21793 = ~n39303 ;
  assign y21794 = ~1'b0 ;
  assign y21795 = ~n39305 ;
  assign y21796 = ~1'b0 ;
  assign y21797 = ~n39306 ;
  assign y21798 = ~n39313 ;
  assign y21799 = ~n39315 ;
  assign y21800 = ~1'b0 ;
  assign y21801 = ~n39317 ;
  assign y21802 = n39318 ;
  assign y21803 = ~1'b0 ;
  assign y21804 = ~1'b0 ;
  assign y21805 = ~1'b0 ;
  assign y21806 = n39320 ;
  assign y21807 = ~n39321 ;
  assign y21808 = ~1'b0 ;
  assign y21809 = ~1'b0 ;
  assign y21810 = n2356 ;
  assign y21811 = ~1'b0 ;
  assign y21812 = ~1'b0 ;
  assign y21813 = ~n39327 ;
  assign y21814 = n39328 ;
  assign y21815 = ~n39329 ;
  assign y21816 = n39332 ;
  assign y21817 = n39337 ;
  assign y21818 = ~1'b0 ;
  assign y21819 = n39340 ;
  assign y21820 = n3050 ;
  assign y21821 = ~n39342 ;
  assign y21822 = ~n39345 ;
  assign y21823 = ~n39347 ;
  assign y21824 = ~n39349 ;
  assign y21825 = ~n39350 ;
  assign y21826 = ~n39351 ;
  assign y21827 = ~n39352 ;
  assign y21828 = ~n39354 ;
  assign y21829 = ~n39359 ;
  assign y21830 = ~1'b0 ;
  assign y21831 = n39362 ;
  assign y21832 = ~1'b0 ;
  assign y21833 = ~n39363 ;
  assign y21834 = ~n39367 ;
  assign y21835 = 1'b0 ;
  assign y21836 = n39368 ;
  assign y21837 = ~n39369 ;
  assign y21838 = ~1'b0 ;
  assign y21839 = n39373 ;
  assign y21840 = n39378 ;
  assign y21841 = ~n39382 ;
  assign y21842 = n39389 ;
  assign y21843 = ~n39391 ;
  assign y21844 = n39393 ;
  assign y21845 = ~n39399 ;
  assign y21846 = n39402 ;
  assign y21847 = n39408 ;
  assign y21848 = ~n39411 ;
  assign y21849 = n39413 ;
  assign y21850 = n39414 ;
  assign y21851 = ~1'b0 ;
  assign y21852 = n39416 ;
  assign y21853 = n39421 ;
  assign y21854 = ~n15030 ;
  assign y21855 = n39422 ;
  assign y21856 = ~n39424 ;
  assign y21857 = ~1'b0 ;
  assign y21858 = n39425 ;
  assign y21859 = n39427 ;
  assign y21860 = ~1'b0 ;
  assign y21861 = ~1'b0 ;
  assign y21862 = n39429 ;
  assign y21863 = n39430 ;
  assign y21864 = ~n39433 ;
  assign y21865 = n4128 ;
  assign y21866 = ~n14421 ;
  assign y21867 = ~1'b0 ;
  assign y21868 = ~n39434 ;
  assign y21869 = ~1'b0 ;
  assign y21870 = n39441 ;
  assign y21871 = ~n39443 ;
  assign y21872 = ~1'b0 ;
  assign y21873 = ~n39447 ;
  assign y21874 = n21690 ;
  assign y21875 = n39448 ;
  assign y21876 = n39449 ;
  assign y21877 = ~n16269 ;
  assign y21878 = n9194 ;
  assign y21879 = n39450 ;
  assign y21880 = ~n36642 ;
  assign y21881 = ~1'b0 ;
  assign y21882 = n39452 ;
  assign y21883 = n39453 ;
  assign y21884 = ~1'b0 ;
  assign y21885 = ~1'b0 ;
  assign y21886 = ~n39458 ;
  assign y21887 = ~n39460 ;
  assign y21888 = ~n39461 ;
  assign y21889 = n39462 ;
  assign y21890 = ~1'b0 ;
  assign y21891 = ~n39466 ;
  assign y21892 = ~1'b0 ;
  assign y21893 = n39468 ;
  assign y21894 = ~1'b0 ;
  assign y21895 = n39469 ;
  assign y21896 = ~n39470 ;
  assign y21897 = ~n39471 ;
  assign y21898 = n1541 ;
  assign y21899 = ~n39480 ;
  assign y21900 = ~n39481 ;
  assign y21901 = n39483 ;
  assign y21902 = ~1'b0 ;
  assign y21903 = 1'b0 ;
  assign y21904 = ~1'b0 ;
  assign y21905 = ~n39485 ;
  assign y21906 = ~n39490 ;
  assign y21907 = ~n39493 ;
  assign y21908 = ~n19758 ;
  assign y21909 = ~n39498 ;
  assign y21910 = ~1'b0 ;
  assign y21911 = ~n39503 ;
  assign y21912 = n39505 ;
  assign y21913 = n39507 ;
  assign y21914 = ~1'b0 ;
  assign y21915 = ~n39508 ;
  assign y21916 = ~n11392 ;
  assign y21917 = ~1'b0 ;
  assign y21918 = ~n35005 ;
  assign y21919 = n39511 ;
  assign y21920 = n39512 ;
  assign y21921 = n39514 ;
  assign y21922 = ~1'b0 ;
  assign y21923 = ~n39516 ;
  assign y21924 = ~n20644 ;
  assign y21925 = ~n39518 ;
  assign y21926 = ~n39520 ;
  assign y21927 = ~n39522 ;
  assign y21928 = n39524 ;
  assign y21929 = ~n39525 ;
  assign y21930 = ~n39527 ;
  assign y21931 = ~n39529 ;
  assign y21932 = ~1'b0 ;
  assign y21933 = n39532 ;
  assign y21934 = ~n39533 ;
  assign y21935 = ~n39536 ;
  assign y21936 = ~1'b0 ;
  assign y21937 = ~1'b0 ;
  assign y21938 = 1'b0 ;
  assign y21939 = n39539 ;
  assign y21940 = ~1'b0 ;
  assign y21941 = n39541 ;
  assign y21942 = n25958 ;
  assign y21943 = ~1'b0 ;
  assign y21944 = ~1'b0 ;
  assign y21945 = ~1'b0 ;
  assign y21946 = ~n39544 ;
  assign y21947 = ~n39550 ;
  assign y21948 = n39556 ;
  assign y21949 = n39558 ;
  assign y21950 = ~1'b0 ;
  assign y21951 = n39561 ;
  assign y21952 = n39564 ;
  assign y21953 = ~n1185 ;
  assign y21954 = ~n39565 ;
  assign y21955 = ~n39570 ;
  assign y21956 = n39572 ;
  assign y21957 = ~1'b0 ;
  assign y21958 = n39576 ;
  assign y21959 = n39577 ;
  assign y21960 = ~n39581 ;
  assign y21961 = ~1'b0 ;
  assign y21962 = ~1'b0 ;
  assign y21963 = n39583 ;
  assign y21964 = n39585 ;
  assign y21965 = ~1'b0 ;
  assign y21966 = ~1'b0 ;
  assign y21967 = ~1'b0 ;
  assign y21968 = n39586 ;
  assign y21969 = ~n39587 ;
  assign y21970 = ~n39588 ;
  assign y21971 = ~1'b0 ;
  assign y21972 = n39590 ;
  assign y21973 = ~n39591 ;
  assign y21974 = ~n5382 ;
  assign y21975 = ~n39593 ;
  assign y21976 = ~1'b0 ;
  assign y21977 = n39596 ;
  assign y21978 = ~1'b0 ;
  assign y21979 = n39602 ;
  assign y21980 = n39606 ;
  assign y21981 = ~n39607 ;
  assign y21982 = n39608 ;
  assign y21983 = n39616 ;
  assign y21984 = ~1'b0 ;
  assign y21985 = 1'b0 ;
  assign y21986 = n39617 ;
  assign y21987 = ~1'b0 ;
  assign y21988 = ~n8382 ;
  assign y21989 = n39619 ;
  assign y21990 = n39620 ;
  assign y21991 = n2400 ;
  assign y21992 = n39622 ;
  assign y21993 = n39624 ;
  assign y21994 = ~1'b0 ;
  assign y21995 = n39629 ;
  assign y21996 = ~n39633 ;
  assign y21997 = n39637 ;
  assign y21998 = n39638 ;
  assign y21999 = n39639 ;
  assign y22000 = ~n39642 ;
  assign y22001 = ~n39645 ;
  assign y22002 = ~1'b0 ;
  assign y22003 = n39647 ;
  assign y22004 = ~1'b0 ;
  assign y22005 = ~1'b0 ;
  assign y22006 = ~1'b0 ;
  assign y22007 = ~1'b0 ;
  assign y22008 = n39648 ;
  assign y22009 = n39649 ;
  assign y22010 = ~1'b0 ;
  assign y22011 = ~n39652 ;
  assign y22012 = n39653 ;
  assign y22013 = ~1'b0 ;
  assign y22014 = ~1'b0 ;
  assign y22015 = ~1'b0 ;
  assign y22016 = ~n39654 ;
  assign y22017 = n6333 ;
  assign y22018 = ~1'b0 ;
  assign y22019 = ~1'b0 ;
  assign y22020 = ~n39655 ;
  assign y22021 = 1'b0 ;
  assign y22022 = ~n39657 ;
  assign y22023 = n1496 ;
  assign y22024 = ~1'b0 ;
  assign y22025 = n2528 ;
  assign y22026 = n39659 ;
  assign y22027 = n39660 ;
  assign y22028 = ~n39661 ;
  assign y22029 = ~n39662 ;
  assign y22030 = ~n39665 ;
  assign y22031 = ~n3549 ;
  assign y22032 = ~n39667 ;
  assign y22033 = ~1'b0 ;
  assign y22034 = ~1'b0 ;
  assign y22035 = n39673 ;
  assign y22036 = ~n39675 ;
  assign y22037 = n39677 ;
  assign y22038 = ~1'b0 ;
  assign y22039 = ~n39678 ;
  assign y22040 = ~n39682 ;
  assign y22041 = ~n39684 ;
  assign y22042 = ~1'b0 ;
  assign y22043 = n39686 ;
  assign y22044 = ~n39689 ;
  assign y22045 = ~1'b0 ;
  assign y22046 = ~1'b0 ;
  assign y22047 = ~1'b0 ;
  assign y22048 = n39694 ;
  assign y22049 = ~n39695 ;
  assign y22050 = n39698 ;
  assign y22051 = n39701 ;
  assign y22052 = ~n39703 ;
  assign y22053 = ~n39705 ;
  assign y22054 = n39706 ;
  assign y22055 = ~1'b0 ;
  assign y22056 = ~1'b0 ;
  assign y22057 = n39707 ;
  assign y22058 = n39709 ;
  assign y22059 = n8136 ;
  assign y22060 = ~1'b0 ;
  assign y22061 = ~n39713 ;
  assign y22062 = ~1'b0 ;
  assign y22063 = n39714 ;
  assign y22064 = ~n39716 ;
  assign y22065 = ~1'b0 ;
  assign y22066 = ~n31213 ;
  assign y22067 = n39718 ;
  assign y22068 = n39721 ;
  assign y22069 = n39724 ;
  assign y22070 = ~n39725 ;
  assign y22071 = n39729 ;
  assign y22072 = n39731 ;
  assign y22073 = ~1'b0 ;
  assign y22074 = ~1'b0 ;
  assign y22075 = ~n39733 ;
  assign y22076 = ~1'b0 ;
  assign y22077 = ~n39735 ;
  assign y22078 = n39737 ;
  assign y22079 = ~1'b0 ;
  assign y22080 = n39739 ;
  assign y22081 = ~n39741 ;
  assign y22082 = ~1'b0 ;
  assign y22083 = ~n39743 ;
  assign y22084 = ~n39749 ;
  assign y22085 = ~n39750 ;
  assign y22086 = n13734 ;
  assign y22087 = ~1'b0 ;
  assign y22088 = n39751 ;
  assign y22089 = ~n39752 ;
  assign y22090 = n39753 ;
  assign y22091 = n39755 ;
  assign y22092 = n39757 ;
  assign y22093 = 1'b0 ;
  assign y22094 = n39761 ;
  assign y22095 = ~n39763 ;
  assign y22096 = ~n28691 ;
  assign y22097 = ~n39765 ;
  assign y22098 = ~1'b0 ;
  assign y22099 = n39766 ;
  assign y22100 = n28269 ;
  assign y22101 = ~n39768 ;
  assign y22102 = n39772 ;
  assign y22103 = n39773 ;
  assign y22104 = ~1'b0 ;
  assign y22105 = ~1'b0 ;
  assign y22106 = ~n39775 ;
  assign y22107 = ~1'b0 ;
  assign y22108 = ~n39777 ;
  assign y22109 = n39778 ;
  assign y22110 = ~n39779 ;
  assign y22111 = ~n39784 ;
  assign y22112 = n39787 ;
  assign y22113 = n39790 ;
  assign y22114 = n4060 ;
  assign y22115 = ~n39792 ;
  assign y22116 = n39794 ;
  assign y22117 = ~1'b0 ;
  assign y22118 = n39796 ;
  assign y22119 = n39797 ;
  assign y22120 = n39798 ;
  assign y22121 = ~n39800 ;
  assign y22122 = ~n39803 ;
  assign y22123 = ~n39804 ;
  assign y22124 = ~n39811 ;
  assign y22125 = ~n39814 ;
  assign y22126 = ~1'b0 ;
  assign y22127 = ~n39817 ;
  assign y22128 = n39818 ;
  assign y22129 = n39821 ;
  assign y22130 = ~n39822 ;
  assign y22131 = n39826 ;
  assign y22132 = n39828 ;
  assign y22133 = n39830 ;
  assign y22134 = n39831 ;
  assign y22135 = ~n3115 ;
  assign y22136 = ~n39836 ;
  assign y22137 = ~1'b0 ;
  assign y22138 = ~n39838 ;
  assign y22139 = n39845 ;
  assign y22140 = ~n39848 ;
  assign y22141 = ~n39849 ;
  assign y22142 = ~1'b0 ;
  assign y22143 = ~n39850 ;
  assign y22144 = ~n39852 ;
  assign y22145 = ~1'b0 ;
  assign y22146 = ~1'b0 ;
  assign y22147 = n11777 ;
  assign y22148 = ~n39854 ;
  assign y22149 = ~1'b0 ;
  assign y22150 = ~1'b0 ;
  assign y22151 = ~n39856 ;
  assign y22152 = 1'b0 ;
  assign y22153 = ~1'b0 ;
  assign y22154 = ~1'b0 ;
  assign y22155 = n39860 ;
  assign y22156 = n39864 ;
  assign y22157 = n35011 ;
  assign y22158 = n39867 ;
  assign y22159 = ~n39875 ;
  assign y22160 = ~n39876 ;
  assign y22161 = ~n28840 ;
  assign y22162 = n39877 ;
  assign y22163 = ~n39879 ;
  assign y22164 = n39880 ;
  assign y22165 = n39883 ;
  assign y22166 = ~n39887 ;
  assign y22167 = n39889 ;
  assign y22168 = n39891 ;
  assign y22169 = n39896 ;
  assign y22170 = n39900 ;
  assign y22171 = ~1'b0 ;
  assign y22172 = n39902 ;
  assign y22173 = ~n39903 ;
  assign y22174 = n38818 ;
  assign y22175 = ~n39905 ;
  assign y22176 = ~1'b0 ;
  assign y22177 = n19071 ;
  assign y22178 = ~n39907 ;
  assign y22179 = ~1'b0 ;
  assign y22180 = n39908 ;
  assign y22181 = ~n39909 ;
  assign y22182 = ~n39911 ;
  assign y22183 = n39912 ;
  assign y22184 = ~1'b0 ;
  assign y22185 = ~1'b0 ;
  assign y22186 = 1'b0 ;
  assign y22187 = ~1'b0 ;
  assign y22188 = ~1'b0 ;
  assign y22189 = n39913 ;
  assign y22190 = n39914 ;
  assign y22191 = ~n39915 ;
  assign y22192 = ~1'b0 ;
  assign y22193 = ~1'b0 ;
  assign y22194 = ~1'b0 ;
  assign y22195 = ~1'b0 ;
  assign y22196 = ~n39921 ;
  assign y22197 = 1'b0 ;
  assign y22198 = ~n39922 ;
  assign y22199 = ~1'b0 ;
  assign y22200 = n39924 ;
  assign y22201 = ~n39930 ;
  assign y22202 = n39931 ;
  assign y22203 = ~1'b0 ;
  assign y22204 = ~n39932 ;
  assign y22205 = n39936 ;
  assign y22206 = ~1'b0 ;
  assign y22207 = ~1'b0 ;
  assign y22208 = n39940 ;
  assign y22209 = ~n25135 ;
  assign y22210 = ~n3305 ;
  assign y22211 = n39941 ;
  assign y22212 = n39942 ;
  assign y22213 = n39944 ;
  assign y22214 = ~1'b0 ;
  assign y22215 = n39947 ;
  assign y22216 = ~1'b0 ;
  assign y22217 = ~1'b0 ;
  assign y22218 = n39948 ;
  assign y22219 = ~n39953 ;
  assign y22220 = n39955 ;
  assign y22221 = n39956 ;
  assign y22222 = ~n39957 ;
  assign y22223 = n39958 ;
  assign y22224 = ~1'b0 ;
  assign y22225 = n39959 ;
  assign y22226 = ~n39960 ;
  assign y22227 = ~1'b0 ;
  assign y22228 = n39961 ;
  assign y22229 = n39964 ;
  assign y22230 = ~n39968 ;
  assign y22231 = ~n39969 ;
  assign y22232 = ~1'b0 ;
  assign y22233 = n39971 ;
  assign y22234 = n39972 ;
  assign y22235 = n39973 ;
  assign y22236 = n39977 ;
  assign y22237 = ~n22217 ;
  assign y22238 = ~n39978 ;
  assign y22239 = n39979 ;
  assign y22240 = ~n39983 ;
  assign y22241 = n39984 ;
  assign y22242 = ~n14619 ;
  assign y22243 = ~n39985 ;
  assign y22244 = ~n39986 ;
  assign y22245 = ~n39987 ;
  assign y22246 = ~n36078 ;
  assign y22247 = n39988 ;
  assign y22248 = n39989 ;
  assign y22249 = n39992 ;
  assign y22250 = ~n39995 ;
  assign y22251 = ~n39997 ;
  assign y22252 = ~1'b0 ;
  assign y22253 = ~1'b0 ;
  assign y22254 = ~n40001 ;
  assign y22255 = ~1'b0 ;
  assign y22256 = 1'b0 ;
  assign y22257 = ~n40003 ;
  assign y22258 = ~n40005 ;
  assign y22259 = n40010 ;
  assign y22260 = ~n40011 ;
  assign y22261 = n40012 ;
  assign y22262 = ~n40014 ;
  assign y22263 = n40015 ;
  assign y22264 = n40017 ;
  assign y22265 = n40021 ;
  assign y22266 = ~1'b0 ;
  assign y22267 = ~n40023 ;
  assign y22268 = n40024 ;
  assign y22269 = ~n40025 ;
  assign y22270 = ~n40026 ;
  assign y22271 = n40030 ;
  assign y22272 = n40032 ;
  assign y22273 = ~n1727 ;
  assign y22274 = n40033 ;
  assign y22275 = n40037 ;
  assign y22276 = ~1'b0 ;
  assign y22277 = n40038 ;
  assign y22278 = ~n40041 ;
  assign y22279 = n40045 ;
  assign y22280 = ~1'b0 ;
  assign y22281 = ~1'b0 ;
  assign y22282 = 1'b0 ;
  assign y22283 = ~1'b0 ;
  assign y22284 = ~n40049 ;
  assign y22285 = n40051 ;
  assign y22286 = n22787 ;
  assign y22287 = ~n40056 ;
  assign y22288 = n40059 ;
  assign y22289 = n40061 ;
  assign y22290 = ~n40063 ;
  assign y22291 = n40064 ;
  assign y22292 = ~n40066 ;
  assign y22293 = ~1'b0 ;
  assign y22294 = ~1'b0 ;
  assign y22295 = ~n40068 ;
  assign y22296 = ~n40070 ;
  assign y22297 = n40072 ;
  assign y22298 = ~n40073 ;
  assign y22299 = ~n5418 ;
  assign y22300 = n40078 ;
  assign y22301 = ~n40080 ;
  assign y22302 = n40081 ;
  assign y22303 = n40082 ;
  assign y22304 = n40083 ;
  assign y22305 = ~1'b0 ;
  assign y22306 = ~n11493 ;
  assign y22307 = n40087 ;
  assign y22308 = n40090 ;
  assign y22309 = ~n40093 ;
  assign y22310 = n40096 ;
  assign y22311 = n40100 ;
  assign y22312 = ~1'b0 ;
  assign y22313 = n40101 ;
  assign y22314 = ~n19444 ;
  assign y22315 = ~1'b0 ;
  assign y22316 = ~n40105 ;
  assign y22317 = ~1'b0 ;
  assign y22318 = ~1'b0 ;
  assign y22319 = n40108 ;
  assign y22320 = n40110 ;
  assign y22321 = ~n40111 ;
  assign y22322 = ~n4080 ;
  assign y22323 = ~1'b0 ;
  assign y22324 = ~n40116 ;
  assign y22325 = ~n20006 ;
  assign y22326 = ~1'b0 ;
  assign y22327 = ~1'b0 ;
  assign y22328 = ~1'b0 ;
  assign y22329 = n40117 ;
  assign y22330 = ~n40119 ;
  assign y22331 = n40121 ;
  assign y22332 = ~n40125 ;
  assign y22333 = n40128 ;
  assign y22334 = ~1'b0 ;
  assign y22335 = ~1'b0 ;
  assign y22336 = n40129 ;
  assign y22337 = ~1'b0 ;
  assign y22338 = ~1'b0 ;
  assign y22339 = ~1'b0 ;
  assign y22340 = n40132 ;
  assign y22341 = ~n40136 ;
  assign y22342 = n12832 ;
  assign y22343 = ~n32505 ;
  assign y22344 = n40140 ;
  assign y22345 = ~n40143 ;
  assign y22346 = ~n40145 ;
  assign y22347 = ~n40149 ;
  assign y22348 = ~1'b0 ;
  assign y22349 = n40151 ;
  assign y22350 = n40155 ;
  assign y22351 = n40157 ;
  assign y22352 = n40158 ;
  assign y22353 = ~n40160 ;
  assign y22354 = n40162 ;
  assign y22355 = n40163 ;
  assign y22356 = ~1'b0 ;
  assign y22357 = ~n40164 ;
  assign y22358 = ~1'b0 ;
  assign y22359 = ~1'b0 ;
  assign y22360 = ~n40167 ;
  assign y22361 = n40168 ;
  assign y22362 = ~1'b0 ;
  assign y22363 = ~n40172 ;
  assign y22364 = n40180 ;
  assign y22365 = n40182 ;
  assign y22366 = ~1'b0 ;
  assign y22367 = ~n40183 ;
  assign y22368 = ~n29894 ;
  assign y22369 = n40184 ;
  assign y22370 = ~n40189 ;
  assign y22371 = n40191 ;
  assign y22372 = ~n40194 ;
  assign y22373 = ~n40196 ;
  assign y22374 = ~n21122 ;
  assign y22375 = n40197 ;
  assign y22376 = ~1'b0 ;
  assign y22377 = n18279 ;
  assign y22378 = ~n40198 ;
  assign y22379 = n40199 ;
  assign y22380 = n8066 ;
  assign y22381 = ~n40200 ;
  assign y22382 = ~n40201 ;
  assign y22383 = ~n40203 ;
  assign y22384 = n40205 ;
  assign y22385 = n40206 ;
  assign y22386 = ~1'b0 ;
  assign y22387 = ~1'b0 ;
  assign y22388 = ~n40209 ;
  assign y22389 = ~n40213 ;
  assign y22390 = ~n40217 ;
  assign y22391 = ~n7906 ;
  assign y22392 = n40220 ;
  assign y22393 = ~1'b0 ;
  assign y22394 = n40221 ;
  assign y22395 = ~n40222 ;
  assign y22396 = 1'b0 ;
  assign y22397 = ~1'b0 ;
  assign y22398 = ~n40224 ;
  assign y22399 = ~1'b0 ;
  assign y22400 = ~n40225 ;
  assign y22401 = ~n40229 ;
  assign y22402 = ~n40230 ;
  assign y22403 = n40232 ;
  assign y22404 = ~1'b0 ;
  assign y22405 = n40234 ;
  assign y22406 = ~1'b0 ;
  assign y22407 = n40238 ;
  assign y22408 = n40241 ;
  assign y22409 = n40245 ;
  assign y22410 = n40246 ;
  assign y22411 = ~n40247 ;
  assign y22412 = 1'b0 ;
  assign y22413 = ~n40251 ;
  assign y22414 = ~n40259 ;
  assign y22415 = ~n40261 ;
  assign y22416 = ~1'b0 ;
  assign y22417 = ~n40263 ;
  assign y22418 = ~n1099 ;
  assign y22419 = ~n40264 ;
  assign y22420 = ~n40266 ;
  assign y22421 = n40267 ;
  assign y22422 = ~1'b0 ;
  assign y22423 = ~1'b0 ;
  assign y22424 = ~1'b0 ;
  assign y22425 = n40271 ;
  assign y22426 = ~n40277 ;
  assign y22427 = ~1'b0 ;
  assign y22428 = 1'b0 ;
  assign y22429 = ~1'b0 ;
  assign y22430 = n40283 ;
  assign y22431 = ~n40287 ;
  assign y22432 = ~n40290 ;
  assign y22433 = n17907 ;
  assign y22434 = ~1'b0 ;
  assign y22435 = n40294 ;
  assign y22436 = ~n40296 ;
  assign y22437 = ~1'b0 ;
  assign y22438 = ~1'b0 ;
  assign y22439 = ~n40297 ;
  assign y22440 = n40299 ;
  assign y22441 = n40303 ;
  assign y22442 = n40311 ;
  assign y22443 = ~1'b0 ;
  assign y22444 = ~1'b0 ;
  assign y22445 = ~n40312 ;
  assign y22446 = n40315 ;
  assign y22447 = ~1'b0 ;
  assign y22448 = ~n40316 ;
  assign y22449 = ~n40318 ;
  assign y22450 = ~n40320 ;
  assign y22451 = ~1'b0 ;
  assign y22452 = ~n40321 ;
  assign y22453 = ~n40322 ;
  assign y22454 = ~n40323 ;
  assign y22455 = n40325 ;
  assign y22456 = ~n26602 ;
  assign y22457 = ~1'b0 ;
  assign y22458 = ~1'b0 ;
  assign y22459 = n7798 ;
  assign y22460 = ~n40326 ;
  assign y22461 = ~1'b0 ;
  assign y22462 = n40327 ;
  assign y22463 = n40328 ;
  assign y22464 = ~n11416 ;
  assign y22465 = ~n40330 ;
  assign y22466 = n35174 ;
  assign y22467 = ~1'b0 ;
  assign y22468 = n40332 ;
  assign y22469 = ~n40334 ;
  assign y22470 = ~n40336 ;
  assign y22471 = ~n40340 ;
  assign y22472 = ~1'b0 ;
  assign y22473 = ~n40342 ;
  assign y22474 = n40343 ;
  assign y22475 = ~n40345 ;
  assign y22476 = 1'b0 ;
  assign y22477 = ~1'b0 ;
  assign y22478 = ~1'b0 ;
  assign y22479 = ~n40348 ;
  assign y22480 = ~1'b0 ;
  assign y22481 = n40349 ;
  assign y22482 = n40352 ;
  assign y22483 = ~1'b0 ;
  assign y22484 = ~n40359 ;
  assign y22485 = n40363 ;
  assign y22486 = 1'b0 ;
  assign y22487 = ~n40364 ;
  assign y22488 = n40365 ;
  assign y22489 = n40369 ;
  assign y22490 = ~n40370 ;
  assign y22491 = ~n40372 ;
  assign y22492 = ~n40375 ;
  assign y22493 = ~1'b0 ;
  assign y22494 = ~1'b0 ;
  assign y22495 = n40380 ;
  assign y22496 = n40381 ;
  assign y22497 = ~1'b0 ;
  assign y22498 = ~1'b0 ;
  assign y22499 = ~n40386 ;
  assign y22500 = ~n40387 ;
  assign y22501 = ~n40389 ;
  assign y22502 = ~n40391 ;
  assign y22503 = ~n40394 ;
  assign y22504 = ~n40396 ;
  assign y22505 = n40400 ;
  assign y22506 = ~1'b0 ;
  assign y22507 = ~n40406 ;
  assign y22508 = ~1'b0 ;
  assign y22509 = n40408 ;
  assign y22510 = n40410 ;
  assign y22511 = n40411 ;
  assign y22512 = ~n40413 ;
  assign y22513 = n40415 ;
  assign y22514 = ~1'b0 ;
  assign y22515 = ~n40418 ;
  assign y22516 = ~1'b0 ;
  assign y22517 = n40421 ;
  assign y22518 = n40422 ;
  assign y22519 = ~1'b0 ;
  assign y22520 = n40426 ;
  assign y22521 = ~n40430 ;
  assign y22522 = n10017 ;
  assign y22523 = ~1'b0 ;
  assign y22524 = ~1'b0 ;
  assign y22525 = 1'b0 ;
  assign y22526 = ~n40435 ;
  assign y22527 = ~n40440 ;
  assign y22528 = ~n40442 ;
  assign y22529 = ~n40444 ;
  assign y22530 = ~n37478 ;
  assign y22531 = n40447 ;
  assign y22532 = n40448 ;
  assign y22533 = ~n40451 ;
  assign y22534 = n40452 ;
  assign y22535 = ~1'b0 ;
  assign y22536 = n23794 ;
  assign y22537 = ~n40454 ;
  assign y22538 = ~1'b0 ;
  assign y22539 = n40456 ;
  assign y22540 = n40458 ;
  assign y22541 = n40461 ;
  assign y22542 = n40463 ;
  assign y22543 = ~n40464 ;
  assign y22544 = ~n40466 ;
  assign y22545 = n2925 ;
  assign y22546 = n40467 ;
  assign y22547 = ~1'b0 ;
  assign y22548 = n40468 ;
  assign y22549 = ~n40469 ;
  assign y22550 = ~1'b0 ;
  assign y22551 = ~n40471 ;
  assign y22552 = ~n40478 ;
  assign y22553 = n1109 ;
  assign y22554 = n40479 ;
  assign y22555 = ~n40480 ;
  assign y22556 = n40482 ;
  assign y22557 = ~1'b0 ;
  assign y22558 = n40484 ;
  assign y22559 = n40485 ;
  assign y22560 = n40488 ;
  assign y22561 = ~1'b0 ;
  assign y22562 = ~n40495 ;
  assign y22563 = n34782 ;
  assign y22564 = n40500 ;
  assign y22565 = ~n40505 ;
  assign y22566 = ~n14345 ;
  assign y22567 = n40508 ;
  assign y22568 = ~n40509 ;
  assign y22569 = ~n40511 ;
  assign y22570 = ~n4676 ;
  assign y22571 = n40516 ;
  assign y22572 = n40520 ;
  assign y22573 = ~n40522 ;
  assign y22574 = ~n40523 ;
  assign y22575 = n40524 ;
  assign y22576 = ~n40525 ;
  assign y22577 = ~n40526 ;
  assign y22578 = ~n40530 ;
  assign y22579 = ~n40532 ;
  assign y22580 = ~1'b0 ;
  assign y22581 = ~1'b0 ;
  assign y22582 = n40533 ;
  assign y22583 = 1'b0 ;
  assign y22584 = ~1'b0 ;
  assign y22585 = n40535 ;
  assign y22586 = ~1'b0 ;
  assign y22587 = ~1'b0 ;
  assign y22588 = ~n7016 ;
  assign y22589 = ~n40536 ;
  assign y22590 = ~1'b0 ;
  assign y22591 = n40538 ;
  assign y22592 = n40541 ;
  assign y22593 = n40545 ;
  assign y22594 = ~1'b0 ;
  assign y22595 = ~n2781 ;
  assign y22596 = ~1'b0 ;
  assign y22597 = ~1'b0 ;
  assign y22598 = ~n40548 ;
  assign y22599 = n40549 ;
  assign y22600 = ~1'b0 ;
  assign y22601 = ~1'b0 ;
  assign y22602 = ~1'b0 ;
  assign y22603 = ~1'b0 ;
  assign y22604 = ~n40552 ;
  assign y22605 = n19714 ;
  assign y22606 = ~n40554 ;
  assign y22607 = ~n40557 ;
  assign y22608 = ~1'b0 ;
  assign y22609 = n40561 ;
  assign y22610 = n40562 ;
  assign y22611 = ~n40563 ;
  assign y22612 = ~1'b0 ;
  assign y22613 = ~n40567 ;
  assign y22614 = n40571 ;
  assign y22615 = ~1'b0 ;
  assign y22616 = ~n40572 ;
  assign y22617 = ~n40575 ;
  assign y22618 = ~1'b0 ;
  assign y22619 = ~1'b0 ;
  assign y22620 = n40578 ;
  assign y22621 = n40581 ;
  assign y22622 = ~n40585 ;
  assign y22623 = ~n40586 ;
  assign y22624 = ~1'b0 ;
  assign y22625 = n40589 ;
  assign y22626 = n40591 ;
  assign y22627 = ~n40592 ;
  assign y22628 = n40595 ;
  assign y22629 = n27660 ;
  assign y22630 = n40596 ;
  assign y22631 = ~n40597 ;
  assign y22632 = n40598 ;
  assign y22633 = ~1'b0 ;
  assign y22634 = ~1'b0 ;
  assign y22635 = ~n40600 ;
  assign y22636 = ~1'b0 ;
  assign y22637 = ~n40602 ;
  assign y22638 = ~n40606 ;
  assign y22639 = ~1'b0 ;
  assign y22640 = n40609 ;
  assign y22641 = n40610 ;
  assign y22642 = ~n40612 ;
  assign y22643 = ~n40614 ;
  assign y22644 = n40616 ;
  assign y22645 = ~n40618 ;
  assign y22646 = ~1'b0 ;
  assign y22647 = ~n14878 ;
  assign y22648 = n40619 ;
  assign y22649 = n40620 ;
  assign y22650 = n40621 ;
  assign y22651 = n40624 ;
  assign y22652 = n40626 ;
  assign y22653 = ~1'b0 ;
  assign y22654 = ~n38236 ;
  assign y22655 = ~n40628 ;
  assign y22656 = n40630 ;
  assign y22657 = ~n40636 ;
  assign y22658 = n40640 ;
  assign y22659 = n13999 ;
  assign y22660 = ~1'b0 ;
  assign y22661 = n40641 ;
  assign y22662 = n40643 ;
  assign y22663 = n40644 ;
  assign y22664 = n40645 ;
  assign y22665 = n40646 ;
  assign y22666 = ~n40648 ;
  assign y22667 = n40654 ;
  assign y22668 = n40656 ;
  assign y22669 = n40660 ;
  assign y22670 = ~1'b0 ;
  assign y22671 = n40662 ;
  assign y22672 = ~1'b0 ;
  assign y22673 = n40663 ;
  assign y22674 = ~n40664 ;
  assign y22675 = ~1'b0 ;
  assign y22676 = ~1'b0 ;
  assign y22677 = n40665 ;
  assign y22678 = ~1'b0 ;
  assign y22679 = ~1'b0 ;
  assign y22680 = ~n40667 ;
  assign y22681 = ~n40673 ;
  assign y22682 = ~x135 ;
  assign y22683 = ~1'b0 ;
  assign y22684 = ~n40677 ;
  assign y22685 = ~n40678 ;
  assign y22686 = ~n8917 ;
  assign y22687 = ~n40679 ;
  assign y22688 = n40680 ;
  assign y22689 = ~1'b0 ;
  assign y22690 = n40682 ;
  assign y22691 = ~n18727 ;
  assign y22692 = ~1'b0 ;
  assign y22693 = ~n40683 ;
  assign y22694 = ~n40687 ;
  assign y22695 = n40688 ;
  assign y22696 = n38430 ;
  assign y22697 = ~n40690 ;
  assign y22698 = ~n40698 ;
  assign y22699 = n40700 ;
  assign y22700 = ~n40702 ;
  assign y22701 = n40703 ;
  assign y22702 = n40704 ;
  assign y22703 = n40707 ;
  assign y22704 = ~1'b0 ;
  assign y22705 = n40710 ;
  assign y22706 = ~n40714 ;
  assign y22707 = n40715 ;
  assign y22708 = n32505 ;
  assign y22709 = ~n9404 ;
  assign y22710 = ~1'b0 ;
  assign y22711 = ~n40716 ;
  assign y22712 = n40718 ;
  assign y22713 = ~n40720 ;
  assign y22714 = ~n40722 ;
  assign y22715 = n38023 ;
  assign y22716 = ~1'b0 ;
  assign y22717 = n40723 ;
  assign y22718 = ~n40724 ;
  assign y22719 = n40725 ;
  assign y22720 = n40726 ;
  assign y22721 = ~1'b0 ;
  assign y22722 = ~n40731 ;
  assign y22723 = ~1'b0 ;
  assign y22724 = n40732 ;
  assign y22725 = ~1'b0 ;
  assign y22726 = ~n40734 ;
  assign y22727 = ~n40738 ;
  assign y22728 = n40741 ;
  assign y22729 = n40744 ;
  assign y22730 = n40745 ;
  assign y22731 = n40746 ;
  assign y22732 = n40747 ;
  assign y22733 = ~n40749 ;
  assign y22734 = ~1'b0 ;
  assign y22735 = ~1'b0 ;
  assign y22736 = n40750 ;
  assign y22737 = ~n40753 ;
  assign y22738 = ~1'b0 ;
  assign y22739 = ~n13779 ;
  assign y22740 = n40754 ;
  assign y22741 = ~n40758 ;
  assign y22742 = n6235 ;
  assign y22743 = ~1'b0 ;
  assign y22744 = ~n40760 ;
  assign y22745 = ~n40762 ;
  assign y22746 = n40765 ;
  assign y22747 = n40767 ;
  assign y22748 = n40769 ;
  assign y22749 = ~n40771 ;
  assign y22750 = n40773 ;
  assign y22751 = n40774 ;
  assign y22752 = ~1'b0 ;
  assign y22753 = ~n40778 ;
  assign y22754 = ~n40779 ;
  assign y22755 = n6257 ;
  assign y22756 = ~1'b0 ;
  assign y22757 = n40784 ;
  assign y22758 = n40787 ;
  assign y22759 = ~1'b0 ;
  assign y22760 = n27016 ;
  assign y22761 = ~n40794 ;
  assign y22762 = ~1'b0 ;
  assign y22763 = ~n40795 ;
  assign y22764 = ~n40796 ;
  assign y22765 = n40798 ;
  assign y22766 = 1'b0 ;
  assign y22767 = n40800 ;
  assign y22768 = ~n40802 ;
  assign y22769 = n40803 ;
  assign y22770 = ~n40804 ;
  assign y22771 = ~n40806 ;
  assign y22772 = n40809 ;
  assign y22773 = ~n40811 ;
  assign y22774 = ~n40812 ;
  assign y22775 = 1'b0 ;
  assign y22776 = ~1'b0 ;
  assign y22777 = ~1'b0 ;
  assign y22778 = ~n40813 ;
  assign y22779 = ~n40818 ;
  assign y22780 = n40820 ;
  assign y22781 = ~1'b0 ;
  assign y22782 = ~n40823 ;
  assign y22783 = n2988 ;
  assign y22784 = n19169 ;
  assign y22785 = ~1'b0 ;
  assign y22786 = ~1'b0 ;
  assign y22787 = ~1'b0 ;
  assign y22788 = ~n40824 ;
  assign y22789 = ~1'b0 ;
  assign y22790 = n40825 ;
  assign y22791 = ~n12585 ;
  assign y22792 = ~1'b0 ;
  assign y22793 = n40826 ;
  assign y22794 = n40834 ;
  assign y22795 = n40838 ;
  assign y22796 = ~n40840 ;
  assign y22797 = ~n40841 ;
  assign y22798 = ~n40842 ;
  assign y22799 = ~1'b0 ;
  assign y22800 = n40846 ;
  assign y22801 = n40848 ;
  assign y22802 = n40849 ;
  assign y22803 = x145 ;
  assign y22804 = n40854 ;
  assign y22805 = ~n40857 ;
  assign y22806 = ~n40858 ;
  assign y22807 = ~1'b0 ;
  assign y22808 = ~1'b0 ;
  assign y22809 = 1'b0 ;
  assign y22810 = ~1'b0 ;
  assign y22811 = ~n40863 ;
  assign y22812 = ~1'b0 ;
  assign y22813 = n40864 ;
  assign y22814 = ~n40865 ;
  assign y22815 = ~n40869 ;
  assign y22816 = n40870 ;
  assign y22817 = ~n40871 ;
  assign y22818 = 1'b0 ;
  assign y22819 = ~1'b0 ;
  assign y22820 = n6405 ;
  assign y22821 = n15166 ;
  assign y22822 = ~n40872 ;
  assign y22823 = ~1'b0 ;
  assign y22824 = ~n40873 ;
  assign y22825 = ~n40877 ;
  assign y22826 = ~n40878 ;
  assign y22827 = ~1'b0 ;
  assign y22828 = ~1'b0 ;
  assign y22829 = n40881 ;
  assign y22830 = ~1'b0 ;
  assign y22831 = ~1'b0 ;
  assign y22832 = ~1'b0 ;
  assign y22833 = ~1'b0 ;
  assign y22834 = ~n40882 ;
  assign y22835 = ~n40883 ;
  assign y22836 = n40884 ;
  assign y22837 = ~n40887 ;
  assign y22838 = ~n40888 ;
  assign y22839 = ~n40889 ;
  assign y22840 = ~1'b0 ;
  assign y22841 = ~n40890 ;
  assign y22842 = n40892 ;
  assign y22843 = ~1'b0 ;
  assign y22844 = ~n40898 ;
  assign y22845 = ~1'b0 ;
  assign y22846 = ~1'b0 ;
  assign y22847 = ~n40899 ;
  assign y22848 = n40900 ;
  assign y22849 = n40901 ;
  assign y22850 = ~1'b0 ;
  assign y22851 = ~n34510 ;
  assign y22852 = n40904 ;
  assign y22853 = ~n40906 ;
  assign y22854 = n40912 ;
  assign y22855 = 1'b0 ;
  assign y22856 = ~1'b0 ;
  assign y22857 = ~1'b0 ;
  assign y22858 = ~n40914 ;
  assign y22859 = ~n40917 ;
  assign y22860 = ~n40918 ;
  assign y22861 = n40919 ;
  assign y22862 = n40921 ;
  assign y22863 = ~1'b0 ;
  assign y22864 = ~1'b0 ;
  assign y22865 = ~1'b0 ;
  assign y22866 = ~n40928 ;
  assign y22867 = ~1'b0 ;
  assign y22868 = ~n40931 ;
  assign y22869 = ~n40934 ;
  assign y22870 = n40935 ;
  assign y22871 = ~n40937 ;
  assign y22872 = n40939 ;
  assign y22873 = ~1'b0 ;
  assign y22874 = ~1'b0 ;
  assign y22875 = ~n40941 ;
  assign y22876 = n40942 ;
  assign y22877 = n19312 ;
  assign y22878 = ~1'b0 ;
  assign y22879 = n40944 ;
  assign y22880 = n40945 ;
  assign y22881 = ~n40946 ;
  assign y22882 = n11511 ;
  assign y22883 = n40947 ;
  assign y22884 = ~1'b0 ;
  assign y22885 = ~n22741 ;
  assign y22886 = ~n7783 ;
  assign y22887 = ~n40949 ;
  assign y22888 = ~1'b0 ;
  assign y22889 = ~n1405 ;
  assign y22890 = ~1'b0 ;
  assign y22891 = ~n40951 ;
  assign y22892 = ~n40953 ;
  assign y22893 = ~n9028 ;
  assign y22894 = n40954 ;
  assign y22895 = ~n40957 ;
  assign y22896 = n31171 ;
  assign y22897 = ~n40960 ;
  assign y22898 = ~n40961 ;
  assign y22899 = ~1'b0 ;
  assign y22900 = ~n40962 ;
  assign y22901 = ~1'b0 ;
  assign y22902 = n40963 ;
  assign y22903 = n40966 ;
  assign y22904 = ~1'b0 ;
  assign y22905 = ~n40969 ;
  assign y22906 = ~1'b0 ;
  assign y22907 = n40971 ;
  assign y22908 = ~1'b0 ;
  assign y22909 = ~1'b0 ;
  assign y22910 = n40972 ;
  assign y22911 = ~n40973 ;
  assign y22912 = ~n10777 ;
  assign y22913 = n40975 ;
  assign y22914 = n40976 ;
  assign y22915 = 1'b0 ;
  assign y22916 = ~1'b0 ;
  assign y22917 = n40977 ;
  assign y22918 = n40979 ;
  assign y22919 = ~n27165 ;
  assign y22920 = n40981 ;
  assign y22921 = n19496 ;
  assign y22922 = ~1'b0 ;
  assign y22923 = ~n40983 ;
  assign y22924 = n30042 ;
  assign y22925 = n19068 ;
  assign y22926 = ~n40987 ;
  assign y22927 = ~1'b0 ;
  assign y22928 = ~1'b0 ;
  assign y22929 = n40988 ;
  assign y22930 = ~n15968 ;
  assign y22931 = 1'b0 ;
  assign y22932 = ~n40992 ;
  assign y22933 = ~n40993 ;
  assign y22934 = ~n10042 ;
  assign y22935 = ~n40997 ;
  assign y22936 = n40998 ;
  assign y22937 = ~1'b0 ;
  assign y22938 = n41004 ;
  assign y22939 = ~1'b0 ;
  assign y22940 = n13612 ;
  assign y22941 = n41008 ;
  assign y22942 = ~n41009 ;
  assign y22943 = n41010 ;
  assign y22944 = n41013 ;
  assign y22945 = n41015 ;
  assign y22946 = n41019 ;
  assign y22947 = ~n41020 ;
  assign y22948 = n41022 ;
  assign y22949 = ~n41023 ;
  assign y22950 = ~1'b0 ;
  assign y22951 = n2016 ;
  assign y22952 = ~n41024 ;
  assign y22953 = n41025 ;
  assign y22954 = ~n41028 ;
  assign y22955 = n41029 ;
  assign y22956 = ~n41032 ;
  assign y22957 = ~n41033 ;
  assign y22958 = ~n41034 ;
  assign y22959 = ~n6805 ;
  assign y22960 = ~1'b0 ;
  assign y22961 = ~1'b0 ;
  assign y22962 = ~n41035 ;
  assign y22963 = ~n41036 ;
  assign y22964 = n41039 ;
  assign y22965 = ~1'b0 ;
  assign y22966 = ~1'b0 ;
  assign y22967 = ~1'b0 ;
  assign y22968 = n41040 ;
  assign y22969 = 1'b0 ;
  assign y22970 = ~1'b0 ;
  assign y22971 = ~n25809 ;
  assign y22972 = ~1'b0 ;
  assign y22973 = ~1'b0 ;
  assign y22974 = 1'b0 ;
  assign y22975 = n41041 ;
  assign y22976 = n41042 ;
  assign y22977 = ~n41043 ;
  assign y22978 = ~n41044 ;
  assign y22979 = ~n41046 ;
  assign y22980 = ~1'b0 ;
  assign y22981 = ~1'b0 ;
  assign y22982 = ~n41050 ;
  assign y22983 = n26689 ;
  assign y22984 = 1'b0 ;
  assign y22985 = ~n9872 ;
  assign y22986 = ~1'b0 ;
  assign y22987 = n41051 ;
  assign y22988 = ~n41054 ;
  assign y22989 = ~n41055 ;
  assign y22990 = ~1'b0 ;
  assign y22991 = ~n41060 ;
  assign y22992 = n41063 ;
  assign y22993 = ~n41064 ;
  assign y22994 = n41065 ;
  assign y22995 = n41067 ;
  assign y22996 = n41069 ;
  assign y22997 = ~1'b0 ;
  assign y22998 = ~1'b0 ;
  assign y22999 = ~n41074 ;
  assign y23000 = n41077 ;
  assign y23001 = n41079 ;
  assign y23002 = ~n41080 ;
  assign y23003 = ~n41081 ;
  assign y23004 = ~n41085 ;
  assign y23005 = ~1'b0 ;
  assign y23006 = ~n41086 ;
  assign y23007 = ~1'b0 ;
  assign y23008 = ~n41087 ;
  assign y23009 = n41089 ;
  assign y23010 = n41092 ;
  assign y23011 = ~n41093 ;
  assign y23012 = ~n41095 ;
  assign y23013 = ~1'b0 ;
  assign y23014 = ~n41098 ;
  assign y23015 = ~1'b0 ;
  assign y23016 = n41099 ;
  assign y23017 = n41101 ;
  assign y23018 = ~1'b0 ;
  assign y23019 = ~1'b0 ;
  assign y23020 = ~n41103 ;
  assign y23021 = n41104 ;
  assign y23022 = n41113 ;
  assign y23023 = ~n41114 ;
  assign y23024 = ~1'b0 ;
  assign y23025 = ~1'b0 ;
  assign y23026 = n41116 ;
  assign y23027 = n41118 ;
  assign y23028 = ~n41119 ;
  assign y23029 = ~1'b0 ;
  assign y23030 = n41124 ;
  assign y23031 = n41126 ;
  assign y23032 = ~1'b0 ;
  assign y23033 = n41129 ;
  assign y23034 = n41130 ;
  assign y23035 = ~1'b0 ;
  assign y23036 = ~1'b0 ;
  assign y23037 = n41131 ;
  assign y23038 = ~1'b0 ;
  assign y23039 = n41134 ;
  assign y23040 = ~n41137 ;
  assign y23041 = ~n41139 ;
  assign y23042 = ~n41145 ;
  assign y23043 = ~n41147 ;
  assign y23044 = n41150 ;
  assign y23045 = n41151 ;
  assign y23046 = ~1'b0 ;
  assign y23047 = ~1'b0 ;
  assign y23048 = ~n41155 ;
  assign y23049 = ~1'b0 ;
  assign y23050 = ~n41158 ;
  assign y23051 = ~n35198 ;
  assign y23052 = ~n41159 ;
  assign y23053 = n7679 ;
  assign y23054 = ~n41161 ;
  assign y23055 = ~1'b0 ;
  assign y23056 = n41163 ;
  assign y23057 = ~1'b0 ;
  assign y23058 = ~n41164 ;
  assign y23059 = ~n41166 ;
  assign y23060 = ~n41168 ;
  assign y23061 = ~1'b0 ;
  assign y23062 = n41173 ;
  assign y23063 = n41175 ;
  assign y23064 = ~n41178 ;
  assign y23065 = n41182 ;
  assign y23066 = ~1'b0 ;
  assign y23067 = ~n41184 ;
  assign y23068 = ~n41185 ;
  assign y23069 = ~n41188 ;
  assign y23070 = ~1'b0 ;
  assign y23071 = ~1'b0 ;
  assign y23072 = ~n41189 ;
  assign y23073 = ~n41190 ;
  assign y23074 = n41197 ;
  assign y23075 = ~n41198 ;
  assign y23076 = n41201 ;
  assign y23077 = ~1'b0 ;
  assign y23078 = n25051 ;
  assign y23079 = ~n41202 ;
  assign y23080 = ~1'b0 ;
  assign y23081 = 1'b0 ;
  assign y23082 = n41204 ;
  assign y23083 = n41205 ;
  assign y23084 = ~n11921 ;
  assign y23085 = n41210 ;
  assign y23086 = n41211 ;
  assign y23087 = ~1'b0 ;
  assign y23088 = ~n41217 ;
  assign y23089 = ~1'b0 ;
  assign y23090 = ~1'b0 ;
  assign y23091 = ~1'b0 ;
  assign y23092 = n41218 ;
  assign y23093 = ~1'b0 ;
  assign y23094 = n41220 ;
  assign y23095 = ~1'b0 ;
  assign y23096 = ~1'b0 ;
  assign y23097 = n41221 ;
  assign y23098 = ~1'b0 ;
  assign y23099 = ~1'b0 ;
  assign y23100 = ~1'b0 ;
  assign y23101 = n17412 ;
  assign y23102 = n41224 ;
  assign y23103 = ~1'b0 ;
  assign y23104 = ~n41229 ;
  assign y23105 = ~1'b0 ;
  assign y23106 = ~1'b0 ;
  assign y23107 = n41230 ;
  assign y23108 = ~n41238 ;
  assign y23109 = n22027 ;
  assign y23110 = ~n41241 ;
  assign y23111 = n41251 ;
  assign y23112 = ~1'b0 ;
  assign y23113 = ~1'b0 ;
  assign y23114 = ~1'b0 ;
  assign y23115 = n41255 ;
  assign y23116 = n41256 ;
  assign y23117 = ~1'b0 ;
  assign y23118 = ~n41259 ;
  assign y23119 = ~1'b0 ;
  assign y23120 = n41261 ;
  assign y23121 = n41265 ;
  assign y23122 = ~n41267 ;
  assign y23123 = ~1'b0 ;
  assign y23124 = ~1'b0 ;
  assign y23125 = ~n41270 ;
  assign y23126 = n26366 ;
  assign y23127 = ~1'b0 ;
  assign y23128 = ~1'b0 ;
  assign y23129 = ~n41276 ;
  assign y23130 = ~n41278 ;
  assign y23131 = 1'b0 ;
  assign y23132 = ~n41280 ;
  assign y23133 = ~1'b0 ;
  assign y23134 = n10487 ;
  assign y23135 = ~n41283 ;
  assign y23136 = ~n41284 ;
  assign y23137 = n2852 ;
  assign y23138 = ~n41286 ;
  assign y23139 = ~n41287 ;
  assign y23140 = 1'b0 ;
  assign y23141 = ~n41288 ;
  assign y23142 = ~1'b0 ;
  assign y23143 = ~1'b0 ;
  assign y23144 = ~n41291 ;
  assign y23145 = ~1'b0 ;
  assign y23146 = n22978 ;
  assign y23147 = ~1'b0 ;
  assign y23148 = ~n41294 ;
  assign y23149 = ~1'b0 ;
  assign y23150 = n7966 ;
  assign y23151 = n41296 ;
  assign y23152 = ~1'b0 ;
  assign y23153 = ~1'b0 ;
  assign y23154 = ~1'b0 ;
  assign y23155 = ~1'b0 ;
  assign y23156 = n41298 ;
  assign y23157 = n41300 ;
  assign y23158 = n41301 ;
  assign y23159 = n41302 ;
  assign y23160 = ~1'b0 ;
  assign y23161 = ~n41306 ;
  assign y23162 = n41311 ;
  assign y23163 = ~n41312 ;
  assign y23164 = n41313 ;
  assign y23165 = ~n41317 ;
  assign y23166 = ~1'b0 ;
  assign y23167 = n41320 ;
  assign y23168 = n41324 ;
  assign y23169 = n41325 ;
  assign y23170 = ~n34486 ;
  assign y23171 = ~n41332 ;
  assign y23172 = ~n41333 ;
  assign y23173 = n41335 ;
  assign y23174 = ~1'b0 ;
  assign y23175 = n41336 ;
  assign y23176 = ~n41337 ;
  assign y23177 = ~1'b0 ;
  assign y23178 = n41340 ;
  assign y23179 = ~n41342 ;
  assign y23180 = n41346 ;
  assign y23181 = ~n41351 ;
  assign y23182 = n41352 ;
  assign y23183 = n41354 ;
  assign y23184 = ~1'b0 ;
  assign y23185 = ~n41357 ;
  assign y23186 = n41359 ;
  assign y23187 = ~1'b0 ;
  assign y23188 = ~n41361 ;
  assign y23189 = ~n41363 ;
  assign y23190 = ~n41367 ;
  assign y23191 = ~1'b0 ;
  assign y23192 = n41370 ;
  assign y23193 = n41373 ;
  assign y23194 = ~1'b0 ;
  assign y23195 = n32964 ;
  assign y23196 = ~1'b0 ;
  assign y23197 = ~n41377 ;
  assign y23198 = ~n6793 ;
  assign y23199 = ~n23608 ;
  assign y23200 = ~1'b0 ;
  assign y23201 = n41379 ;
  assign y23202 = ~1'b0 ;
  assign y23203 = ~1'b0 ;
  assign y23204 = ~n41380 ;
  assign y23205 = n41381 ;
  assign y23206 = ~n41387 ;
  assign y23207 = ~n41389 ;
  assign y23208 = ~1'b0 ;
  assign y23209 = ~1'b0 ;
  assign y23210 = n40724 ;
  assign y23211 = ~n17639 ;
  assign y23212 = 1'b0 ;
  assign y23213 = ~n41390 ;
  assign y23214 = n41392 ;
  assign y23215 = ~n41396 ;
  assign y23216 = ~n41398 ;
  assign y23217 = ~n41399 ;
  assign y23218 = 1'b0 ;
  assign y23219 = ~n41403 ;
  assign y23220 = ~n41404 ;
  assign y23221 = n41405 ;
  assign y23222 = ~n41406 ;
  assign y23223 = ~1'b0 ;
  assign y23224 = n41411 ;
  assign y23225 = ~n41415 ;
  assign y23226 = n5308 ;
  assign y23227 = n41419 ;
  assign y23228 = ~n41420 ;
  assign y23229 = ~1'b0 ;
  assign y23230 = ~1'b0 ;
  assign y23231 = ~1'b0 ;
  assign y23232 = ~n41421 ;
  assign y23233 = ~1'b0 ;
  assign y23234 = ~1'b0 ;
  assign y23235 = n5954 ;
  assign y23236 = n41422 ;
  assign y23237 = ~n41424 ;
  assign y23238 = n41428 ;
  assign y23239 = n41431 ;
  assign y23240 = ~1'b0 ;
  assign y23241 = ~1'b0 ;
  assign y23242 = n41435 ;
  assign y23243 = n41439 ;
  assign y23244 = ~n41441 ;
  assign y23245 = n41442 ;
  assign y23246 = n41443 ;
  assign y23247 = n41446 ;
  assign y23248 = n41449 ;
  assign y23249 = ~n41451 ;
  assign y23250 = ~1'b0 ;
  assign y23251 = ~n41454 ;
  assign y23252 = ~n41455 ;
  assign y23253 = ~n41458 ;
  assign y23254 = ~n41461 ;
  assign y23255 = ~1'b0 ;
  assign y23256 = n41466 ;
  assign y23257 = ~n41467 ;
  assign y23258 = n41469 ;
  assign y23259 = n41474 ;
  assign y23260 = n41475 ;
  assign y23261 = n41485 ;
  assign y23262 = ~n7414 ;
  assign y23263 = ~1'b0 ;
  assign y23264 = ~n41486 ;
  assign y23265 = ~1'b0 ;
  assign y23266 = ~n41487 ;
  assign y23267 = ~n41491 ;
  assign y23268 = n41495 ;
  assign y23269 = n41496 ;
  assign y23270 = ~1'b0 ;
  assign y23271 = ~n41497 ;
  assign y23272 = ~n41501 ;
  assign y23273 = ~1'b0 ;
  assign y23274 = ~1'b0 ;
  assign y23275 = ~1'b0 ;
  assign y23276 = n41505 ;
  assign y23277 = n41508 ;
  assign y23278 = n41511 ;
  assign y23279 = n41512 ;
  assign y23280 = ~n41516 ;
  assign y23281 = ~n19199 ;
  assign y23282 = n3300 ;
  assign y23283 = ~n41520 ;
  assign y23284 = ~1'b0 ;
  assign y23285 = n41523 ;
  assign y23286 = ~1'b0 ;
  assign y23287 = ~1'b0 ;
  assign y23288 = ~1'b0 ;
  assign y23289 = ~n41524 ;
  assign y23290 = n41525 ;
  assign y23291 = ~1'b0 ;
  assign y23292 = n2348 ;
  assign y23293 = ~n37733 ;
  assign y23294 = ~n41529 ;
  assign y23295 = ~n41530 ;
  assign y23296 = n41531 ;
  assign y23297 = n25566 ;
  assign y23298 = ~1'b0 ;
  assign y23299 = n41532 ;
  assign y23300 = ~n41534 ;
  assign y23301 = ~n41541 ;
  assign y23302 = ~1'b0 ;
  assign y23303 = ~n41542 ;
  assign y23304 = ~1'b0 ;
  assign y23305 = ~1'b0 ;
  assign y23306 = ~n41543 ;
  assign y23307 = ~n41550 ;
  assign y23308 = ~n41551 ;
  assign y23309 = n41553 ;
  assign y23310 = ~n41554 ;
  assign y23311 = ~1'b0 ;
  assign y23312 = n41555 ;
  assign y23313 = ~1'b0 ;
  assign y23314 = ~n41556 ;
  assign y23315 = n41558 ;
  assign y23316 = ~n41567 ;
  assign y23317 = ~n2360 ;
  assign y23318 = ~n41568 ;
  assign y23319 = ~1'b0 ;
  assign y23320 = ~n41572 ;
  assign y23321 = n41579 ;
  assign y23322 = ~n41580 ;
  assign y23323 = ~1'b0 ;
  assign y23324 = n41581 ;
  assign y23325 = ~n41583 ;
  assign y23326 = n41586 ;
  assign y23327 = ~1'b0 ;
  assign y23328 = ~1'b0 ;
  assign y23329 = ~n41587 ;
  assign y23330 = n41588 ;
  assign y23331 = n41589 ;
  assign y23332 = 1'b0 ;
  assign y23333 = ~1'b0 ;
  assign y23334 = ~1'b0 ;
  assign y23335 = n41591 ;
  assign y23336 = n41595 ;
  assign y23337 = n36517 ;
  assign y23338 = ~n4933 ;
  assign y23339 = ~1'b0 ;
  assign y23340 = ~1'b0 ;
  assign y23341 = ~n41596 ;
  assign y23342 = n30751 ;
  assign y23343 = ~n41597 ;
  assign y23344 = n41598 ;
  assign y23345 = n41599 ;
  assign y23346 = n41604 ;
  assign y23347 = ~1'b0 ;
  assign y23348 = n41605 ;
  assign y23349 = ~n41606 ;
  assign y23350 = ~1'b0 ;
  assign y23351 = n41609 ;
  assign y23352 = n18180 ;
  assign y23353 = n37254 ;
  assign y23354 = n41610 ;
  assign y23355 = ~1'b0 ;
  assign y23356 = ~1'b0 ;
  assign y23357 = ~1'b0 ;
  assign y23358 = n25973 ;
  assign y23359 = ~n41612 ;
  assign y23360 = ~1'b0 ;
  assign y23361 = ~1'b0 ;
  assign y23362 = n41616 ;
  assign y23363 = ~n41620 ;
  assign y23364 = ~1'b0 ;
  assign y23365 = ~1'b0 ;
  assign y23366 = ~n41623 ;
  assign y23367 = ~1'b0 ;
  assign y23368 = ~n30583 ;
  assign y23369 = ~n41626 ;
  assign y23370 = ~1'b0 ;
  assign y23371 = n41629 ;
  assign y23372 = ~1'b0 ;
  assign y23373 = n41631 ;
  assign y23374 = n28952 ;
  assign y23375 = ~1'b0 ;
  assign y23376 = ~1'b0 ;
  assign y23377 = ~n41632 ;
  assign y23378 = ~n41636 ;
  assign y23379 = ~1'b0 ;
  assign y23380 = n41638 ;
  assign y23381 = n41640 ;
  assign y23382 = ~n41645 ;
  assign y23383 = n41647 ;
  assign y23384 = n41650 ;
  assign y23385 = n41651 ;
  assign y23386 = n41672 ;
  assign y23387 = n41676 ;
  assign y23388 = ~n41677 ;
  assign y23389 = ~1'b0 ;
  assign y23390 = ~1'b0 ;
  assign y23391 = ~1'b0 ;
  assign y23392 = 1'b0 ;
  assign y23393 = ~1'b0 ;
  assign y23394 = n41678 ;
  assign y23395 = n41681 ;
  assign y23396 = ~n41687 ;
  assign y23397 = n41693 ;
  assign y23398 = ~n41695 ;
  assign y23399 = ~n41699 ;
  assign y23400 = ~n41701 ;
  assign y23401 = ~n19222 ;
  assign y23402 = n41703 ;
  assign y23403 = ~1'b0 ;
  assign y23404 = n41704 ;
  assign y23405 = ~n41705 ;
  assign y23406 = n41707 ;
  assign y23407 = ~1'b0 ;
  assign y23408 = n41709 ;
  assign y23409 = 1'b0 ;
  assign y23410 = ~1'b0 ;
  assign y23411 = ~1'b0 ;
  assign y23412 = ~n41713 ;
  assign y23413 = n41714 ;
  assign y23414 = n41715 ;
  assign y23415 = n26744 ;
  assign y23416 = ~n41716 ;
  assign y23417 = ~n41717 ;
  assign y23418 = n41718 ;
  assign y23419 = n41723 ;
  assign y23420 = ~n41724 ;
  assign y23421 = ~1'b0 ;
  assign y23422 = ~n41726 ;
  assign y23423 = ~1'b0 ;
  assign y23424 = n41729 ;
  assign y23425 = n41733 ;
  assign y23426 = n41734 ;
  assign y23427 = ~n41735 ;
  assign y23428 = n9788 ;
  assign y23429 = ~1'b0 ;
  assign y23430 = n41736 ;
  assign y23431 = ~n41739 ;
  assign y23432 = ~1'b0 ;
  assign y23433 = ~1'b0 ;
  assign y23434 = ~1'b0 ;
  assign y23435 = n41741 ;
  assign y23436 = ~1'b0 ;
  assign y23437 = ~n41743 ;
  assign y23438 = n41746 ;
  assign y23439 = n41750 ;
  assign y23440 = n41752 ;
  assign y23441 = ~n29586 ;
  assign y23442 = ~n41754 ;
  assign y23443 = n41757 ;
  assign y23444 = ~n41758 ;
  assign y23445 = ~1'b0 ;
  assign y23446 = n41762 ;
  assign y23447 = ~1'b0 ;
  assign y23448 = n41763 ;
  assign y23449 = n37635 ;
  assign y23450 = 1'b0 ;
  assign y23451 = ~1'b0 ;
  assign y23452 = n41764 ;
  assign y23453 = n41765 ;
  assign y23454 = ~n41767 ;
  assign y23455 = ~1'b0 ;
  assign y23456 = n41774 ;
  assign y23457 = n41775 ;
  assign y23458 = ~n41779 ;
  assign y23459 = ~n41785 ;
  assign y23460 = ~n41786 ;
  assign y23461 = n1208 ;
  assign y23462 = ~n41788 ;
  assign y23463 = ~1'b0 ;
  assign y23464 = ~1'b0 ;
  assign y23465 = ~n41791 ;
  assign y23466 = ~1'b0 ;
  assign y23467 = ~1'b0 ;
  assign y23468 = ~n41792 ;
  assign y23469 = ~n41796 ;
  assign y23470 = ~1'b0 ;
  assign y23471 = n41800 ;
  assign y23472 = ~n5779 ;
  assign y23473 = n41801 ;
  assign y23474 = ~n41805 ;
  assign y23475 = ~1'b0 ;
  assign y23476 = ~1'b0 ;
  assign y23477 = ~n41807 ;
  assign y23478 = n41808 ;
  assign y23479 = ~n41812 ;
  assign y23480 = ~n41814 ;
  assign y23481 = ~n35620 ;
  assign y23482 = n41815 ;
  assign y23483 = ~n41816 ;
  assign y23484 = ~n41819 ;
  assign y23485 = ~n19654 ;
  assign y23486 = ~1'b0 ;
  assign y23487 = ~n41823 ;
  assign y23488 = ~n41827 ;
  assign y23489 = ~n41828 ;
  assign y23490 = ~n41830 ;
  assign y23491 = ~n41834 ;
  assign y23492 = n41835 ;
  assign y23493 = ~n41836 ;
  assign y23494 = n41837 ;
  assign y23495 = ~1'b0 ;
  assign y23496 = ~1'b0 ;
  assign y23497 = ~1'b0 ;
  assign y23498 = ~n41838 ;
  assign y23499 = ~n41840 ;
  assign y23500 = ~n41844 ;
  assign y23501 = ~n41846 ;
  assign y23502 = ~1'b0 ;
  assign y23503 = n41847 ;
  assign y23504 = n41850 ;
  assign y23505 = ~n36705 ;
  assign y23506 = ~1'b0 ;
  assign y23507 = ~n41852 ;
  assign y23508 = ~1'b0 ;
  assign y23509 = n41856 ;
  assign y23510 = ~n41859 ;
  assign y23511 = 1'b0 ;
  assign y23512 = n41860 ;
  assign y23513 = ~n41864 ;
  assign y23514 = ~n41868 ;
  assign y23515 = ~n41870 ;
  assign y23516 = n41873 ;
  assign y23517 = ~n41874 ;
  assign y23518 = n41875 ;
  assign y23519 = ~1'b0 ;
  assign y23520 = ~1'b0 ;
  assign y23521 = ~n41877 ;
  assign y23522 = ~1'b0 ;
  assign y23523 = ~n41878 ;
  assign y23524 = n41883 ;
  assign y23525 = ~n41885 ;
  assign y23526 = n41886 ;
  assign y23527 = n24648 ;
  assign y23528 = ~n41887 ;
  assign y23529 = n41888 ;
  assign y23530 = ~n41889 ;
  assign y23531 = n41893 ;
  assign y23532 = ~1'b0 ;
  assign y23533 = 1'b0 ;
  assign y23534 = n41895 ;
  assign y23535 = n41896 ;
  assign y23536 = ~n41897 ;
  assign y23537 = ~1'b0 ;
  assign y23538 = ~n41899 ;
  assign y23539 = ~n41901 ;
  assign y23540 = ~n41902 ;
  assign y23541 = ~n6662 ;
  assign y23542 = ~n29423 ;
  assign y23543 = ~1'b0 ;
  assign y23544 = ~n41904 ;
  assign y23545 = ~1'b0 ;
  assign y23546 = n41909 ;
  assign y23547 = ~n41912 ;
  assign y23548 = ~n41913 ;
  assign y23549 = 1'b0 ;
  assign y23550 = ~1'b0 ;
  assign y23551 = ~1'b0 ;
  assign y23552 = ~1'b0 ;
  assign y23553 = ~1'b0 ;
  assign y23554 = ~1'b0 ;
  assign y23555 = ~n41914 ;
  assign y23556 = ~n10189 ;
  assign y23557 = n41916 ;
  assign y23558 = n41919 ;
  assign y23559 = ~n41920 ;
  assign y23560 = n41921 ;
  assign y23561 = ~1'b0 ;
  assign y23562 = ~n41922 ;
  assign y23563 = ~n30330 ;
  assign y23564 = ~n41923 ;
  assign y23565 = ~1'b0 ;
  assign y23566 = ~1'b0 ;
  assign y23567 = ~n30256 ;
  assign y23568 = ~n41926 ;
  assign y23569 = ~n41927 ;
  assign y23570 = ~1'b0 ;
  assign y23571 = ~1'b0 ;
  assign y23572 = n41932 ;
  assign y23573 = ~n32202 ;
  assign y23574 = n41933 ;
  assign y23575 = n41936 ;
  assign y23576 = ~1'b0 ;
  assign y23577 = ~n10140 ;
  assign y23578 = n41938 ;
  assign y23579 = ~n41939 ;
  assign y23580 = n41940 ;
  assign y23581 = ~n41942 ;
  assign y23582 = ~1'b0 ;
  assign y23583 = ~n41943 ;
  assign y23584 = n41946 ;
  assign y23585 = n41952 ;
  assign y23586 = ~n41957 ;
  assign y23587 = ~n41962 ;
  assign y23588 = ~n41964 ;
  assign y23589 = ~n41965 ;
  assign y23590 = n41966 ;
  assign y23591 = ~1'b0 ;
  assign y23592 = n41967 ;
  assign y23593 = ~n41970 ;
  assign y23594 = 1'b0 ;
  assign y23595 = ~1'b0 ;
  assign y23596 = ~n41971 ;
  assign y23597 = ~n41972 ;
  assign y23598 = n41975 ;
  assign y23599 = ~n41978 ;
  assign y23600 = n41980 ;
  assign y23601 = n41981 ;
  assign y23602 = ~n41985 ;
  assign y23603 = ~n41986 ;
  assign y23604 = n41987 ;
  assign y23605 = ~1'b0 ;
  assign y23606 = n41989 ;
  assign y23607 = n529 ;
  assign y23608 = n36497 ;
  assign y23609 = ~1'b0 ;
  assign y23610 = n41991 ;
  assign y23611 = ~n41993 ;
  assign y23612 = ~n41995 ;
  assign y23613 = 1'b0 ;
  assign y23614 = ~n41998 ;
  assign y23615 = ~1'b0 ;
  assign y23616 = ~n42004 ;
  assign y23617 = ~1'b0 ;
  assign y23618 = ~n42008 ;
  assign y23619 = ~1'b0 ;
  assign y23620 = ~1'b0 ;
  assign y23621 = ~1'b0 ;
  assign y23622 = n42015 ;
  assign y23623 = n42017 ;
  assign y23624 = n42020 ;
  assign y23625 = ~1'b0 ;
  assign y23626 = ~1'b0 ;
  assign y23627 = n42021 ;
  assign y23628 = 1'b0 ;
  assign y23629 = ~n42022 ;
  assign y23630 = n42023 ;
  assign y23631 = n42026 ;
  assign y23632 = ~1'b0 ;
  assign y23633 = ~1'b0 ;
  assign y23634 = n3845 ;
  assign y23635 = ~1'b0 ;
  assign y23636 = n42027 ;
  assign y23637 = ~n42035 ;
  assign y23638 = ~1'b0 ;
  assign y23639 = n42036 ;
  assign y23640 = n42041 ;
  assign y23641 = ~1'b0 ;
  assign y23642 = n42045 ;
  assign y23643 = 1'b0 ;
  assign y23644 = n42048 ;
  assign y23645 = n42050 ;
  assign y23646 = ~1'b0 ;
  assign y23647 = ~1'b0 ;
  assign y23648 = ~1'b0 ;
  assign y23649 = n42053 ;
  assign y23650 = n1766 ;
  assign y23651 = ~1'b0 ;
  assign y23652 = ~n42055 ;
  assign y23653 = ~n42062 ;
  assign y23654 = ~n42064 ;
  assign y23655 = n42065 ;
  assign y23656 = n42075 ;
  assign y23657 = n27971 ;
  assign y23658 = n42077 ;
  assign y23659 = ~1'b0 ;
  assign y23660 = ~1'b0 ;
  assign y23661 = n42078 ;
  assign y23662 = ~1'b0 ;
  assign y23663 = n42079 ;
  assign y23664 = ~n42081 ;
  assign y23665 = ~n42085 ;
  assign y23666 = ~n42086 ;
  assign y23667 = n42090 ;
  assign y23668 = ~n42093 ;
  assign y23669 = ~1'b0 ;
  assign y23670 = n42094 ;
  assign y23671 = ~n42095 ;
  assign y23672 = ~1'b0 ;
  assign y23673 = ~1'b0 ;
  assign y23674 = ~1'b0 ;
  assign y23675 = ~n42100 ;
  assign y23676 = ~1'b0 ;
  assign y23677 = ~n42102 ;
  assign y23678 = n42104 ;
  assign y23679 = ~n42105 ;
  assign y23680 = ~n42106 ;
  assign y23681 = ~n42108 ;
  assign y23682 = n25122 ;
  assign y23683 = ~1'b0 ;
  assign y23684 = n42109 ;
  assign y23685 = ~1'b0 ;
  assign y23686 = ~n42111 ;
  assign y23687 = ~n42112 ;
  assign y23688 = n42116 ;
  assign y23689 = ~n42117 ;
  assign y23690 = n42118 ;
  assign y23691 = ~n42120 ;
  assign y23692 = n21351 ;
  assign y23693 = ~1'b0 ;
  assign y23694 = n42121 ;
  assign y23695 = ~1'b0 ;
  assign y23696 = ~1'b0 ;
  assign y23697 = ~1'b0 ;
  assign y23698 = n11196 ;
  assign y23699 = ~n42124 ;
  assign y23700 = ~n42126 ;
  assign y23701 = ~1'b0 ;
  assign y23702 = n42128 ;
  assign y23703 = n42129 ;
  assign y23704 = ~n42131 ;
  assign y23705 = ~n42133 ;
  assign y23706 = n42136 ;
  assign y23707 = n42137 ;
  assign y23708 = ~n42138 ;
  assign y23709 = ~1'b0 ;
  assign y23710 = n42141 ;
  assign y23711 = n42145 ;
  assign y23712 = 1'b0 ;
  assign y23713 = n42146 ;
  assign y23714 = ~1'b0 ;
  assign y23715 = n42148 ;
  assign y23716 = n36680 ;
  assign y23717 = n42149 ;
  assign y23718 = 1'b0 ;
  assign y23719 = ~1'b0 ;
  assign y23720 = ~1'b0 ;
  assign y23721 = n42150 ;
  assign y23722 = n42151 ;
  assign y23723 = ~n42153 ;
  assign y23724 = ~n42157 ;
  assign y23725 = n42159 ;
  assign y23726 = ~1'b0 ;
  assign y23727 = ~1'b0 ;
  assign y23728 = ~n42163 ;
  assign y23729 = ~n42168 ;
  assign y23730 = ~n42169 ;
  assign y23731 = ~1'b0 ;
  assign y23732 = ~1'b0 ;
  assign y23733 = ~n42171 ;
  assign y23734 = ~1'b0 ;
  assign y23735 = n2065 ;
  assign y23736 = ~1'b0 ;
  assign y23737 = ~1'b0 ;
  assign y23738 = ~1'b0 ;
  assign y23739 = ~1'b0 ;
  assign y23740 = ~1'b0 ;
  assign y23741 = ~n42172 ;
  assign y23742 = n42173 ;
  assign y23743 = ~n42174 ;
  assign y23744 = ~n42178 ;
  assign y23745 = ~1'b0 ;
  assign y23746 = ~1'b0 ;
  assign y23747 = ~n42179 ;
  assign y23748 = ~1'b0 ;
  assign y23749 = ~n42180 ;
  assign y23750 = ~1'b0 ;
  assign y23751 = ~n42181 ;
  assign y23752 = n42183 ;
  assign y23753 = n42184 ;
  assign y23754 = n42187 ;
  assign y23755 = ~n42188 ;
  assign y23756 = ~1'b0 ;
  assign y23757 = n42189 ;
  assign y23758 = ~n32585 ;
  assign y23759 = ~1'b0 ;
  assign y23760 = 1'b0 ;
  assign y23761 = ~n42191 ;
  assign y23762 = n42193 ;
  assign y23763 = ~1'b0 ;
  assign y23764 = ~n42195 ;
  assign y23765 = ~n42196 ;
  assign y23766 = ~n42197 ;
  assign y23767 = ~n42201 ;
  assign y23768 = ~1'b0 ;
  assign y23769 = 1'b0 ;
  assign y23770 = n42202 ;
  assign y23771 = ~1'b0 ;
  assign y23772 = ~n42207 ;
  assign y23773 = ~n42210 ;
  assign y23774 = n42211 ;
  assign y23775 = ~1'b0 ;
  assign y23776 = ~n42212 ;
  assign y23777 = n42213 ;
  assign y23778 = ~n42216 ;
  assign y23779 = n4230 ;
  assign y23780 = ~n42220 ;
  assign y23781 = ~n42224 ;
  assign y23782 = n42226 ;
  assign y23783 = n1213 ;
  assign y23784 = ~1'b0 ;
  assign y23785 = n42228 ;
  assign y23786 = ~n42232 ;
  assign y23787 = ~n42234 ;
  assign y23788 = n42236 ;
  assign y23789 = n42238 ;
  assign y23790 = n14376 ;
  assign y23791 = ~n42239 ;
  assign y23792 = ~1'b0 ;
  assign y23793 = ~n42242 ;
  assign y23794 = 1'b0 ;
  assign y23795 = ~1'b0 ;
  assign y23796 = ~n42243 ;
  assign y23797 = ~1'b0 ;
  assign y23798 = ~1'b0 ;
  assign y23799 = n42249 ;
  assign y23800 = ~1'b0 ;
  assign y23801 = ~1'b0 ;
  assign y23802 = ~n42251 ;
  assign y23803 = n42252 ;
  assign y23804 = n42255 ;
  assign y23805 = ~n1635 ;
endmodule
