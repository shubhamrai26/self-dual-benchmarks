module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 ;
  assign n129 = ( ~x43 & x77 ) | ( ~x43 & x106 ) | ( x77 & x106 ) ;
  assign n130 = ( ~x66 & x77 ) | ( ~x66 & x91 ) | ( x77 & x91 ) ;
  assign n131 = x81 ^ x40 ^ 1'b0 ;
  assign n132 = x122 & n131 ;
  assign n133 = x90 ^ x66 ^ 1'b0 ;
  assign n134 = x103 & n133 ;
  assign n135 = ( x101 & ~x107 ) | ( x101 & x124 ) | ( ~x107 & x124 ) ;
  assign n136 = ( x45 & x47 ) | ( x45 & ~n135 ) | ( x47 & ~n135 ) ;
  assign n137 = n136 ^ x97 ^ 1'b0 ;
  assign n138 = n130 & n137 ;
  assign n140 = x104 ^ x36 ^ 1'b0 ;
  assign n141 = x87 & n140 ;
  assign n139 = x70 & n134 ;
  assign n142 = n141 ^ n139 ^ 1'b0 ;
  assign n143 = ~x69 & n141 ;
  assign n144 = x61 ^ x40 ^ 1'b0 ;
  assign n145 = x28 & n144 ;
  assign n146 = x101 ^ x65 ^ 1'b0 ;
  assign n147 = x52 & n143 ;
  assign n148 = ~x47 & n147 ;
  assign n149 = x101 ^ x38 ^ x8 ;
  assign n150 = ( ~x7 & x9 ) | ( ~x7 & n141 ) | ( x9 & n141 ) ;
  assign n151 = x92 ^ x77 ^ x5 ;
  assign n152 = x121 ^ x111 ^ 1'b0 ;
  assign n153 = ~n151 & n152 ;
  assign n154 = x47 & n153 ;
  assign n155 = ~n150 & n154 ;
  assign n156 = ( x63 & x91 ) | ( x63 & ~x93 ) | ( x91 & ~x93 ) ;
  assign n157 = x61 & x81 ;
  assign n158 = n157 ^ x37 ^ 1'b0 ;
  assign n159 = x118 ^ x70 ^ x55 ;
  assign n160 = n159 ^ x64 ^ 1'b0 ;
  assign n161 = x87 & ~n160 ;
  assign n162 = x64 & n161 ;
  assign n163 = n149 & n162 ;
  assign n164 = x13 & ~n163 ;
  assign n165 = n164 ^ x14 ^ 1'b0 ;
  assign n166 = x104 ^ x84 ^ x46 ;
  assign n167 = ( x114 & ~x116 ) | ( x114 & n166 ) | ( ~x116 & n166 ) ;
  assign n168 = x94 & ~n167 ;
  assign n169 = ~x31 & n168 ;
  assign n170 = x30 ^ x4 ^ 1'b0 ;
  assign n171 = x33 & n170 ;
  assign n172 = x121 ^ x93 ^ 1'b0 ;
  assign n173 = n171 & n172 ;
  assign n174 = x90 ^ x74 ^ x46 ;
  assign n175 = x19 | n155 ;
  assign n176 = x54 & x68 ;
  assign n177 = x54 & ~n176 ;
  assign n178 = x96 & ~n177 ;
  assign n179 = n178 ^ n145 ^ 1'b0 ;
  assign n181 = x103 & n132 ;
  assign n182 = n158 & n181 ;
  assign n180 = x35 & x69 ;
  assign n183 = n182 ^ n180 ^ 1'b0 ;
  assign n184 = n169 ^ x56 ^ 1'b0 ;
  assign n185 = x37 & ~n184 ;
  assign n186 = ( ~n153 & n159 ) | ( ~n153 & n185 ) | ( n159 & n185 ) ;
  assign n187 = x52 ^ x1 ^ 1'b0 ;
  assign n188 = x56 & n187 ;
  assign n189 = n188 ^ x103 ^ 1'b0 ;
  assign n190 = x107 ^ x27 ^ x12 ;
  assign n191 = ( x35 & x47 ) | ( x35 & ~n130 ) | ( x47 & ~n130 ) ;
  assign n192 = n130 & n191 ;
  assign n193 = n190 & n192 ;
  assign n194 = n145 & n193 ;
  assign n196 = x125 ^ x123 ^ x35 ;
  assign n195 = x2 & x80 ;
  assign n197 = n196 ^ n195 ^ 1'b0 ;
  assign n198 = x2 & x36 ;
  assign n199 = n198 ^ x79 ^ 1'b0 ;
  assign n200 = x119 ^ x103 ^ x66 ;
  assign n201 = n142 ^ x3 ^ 1'b0 ;
  assign n202 = n200 | n201 ;
  assign n203 = x56 & x106 ;
  assign n204 = ~x5 & n203 ;
  assign n205 = x9 & ~n204 ;
  assign n206 = ~x59 & n205 ;
  assign n207 = n136 ^ x112 ^ 1'b0 ;
  assign n208 = n143 & n207 ;
  assign n209 = n208 ^ x124 ^ 1'b0 ;
  assign n210 = ~n206 & n209 ;
  assign n211 = x13 & n132 ;
  assign n212 = ~x46 & n211 ;
  assign n213 = x120 & ~n142 ;
  assign n214 = n213 ^ n135 ^ 1'b0 ;
  assign n215 = x32 & ~n214 ;
  assign n216 = n200 ^ n161 ^ x119 ;
  assign n217 = x124 ^ x28 ^ x7 ;
  assign n218 = ( ~x3 & x13 ) | ( ~x3 & x26 ) | ( x13 & x26 ) ;
  assign n219 = x56 & n194 ;
  assign n220 = ~x87 & n219 ;
  assign n221 = ~x44 & n220 ;
  assign n222 = n217 | n221 ;
  assign n223 = x108 | n222 ;
  assign n224 = x21 & x67 ;
  assign n225 = n224 ^ x20 ^ 1'b0 ;
  assign n226 = x20 & x90 ;
  assign n227 = n226 ^ x102 ^ 1'b0 ;
  assign n228 = x18 & x113 ;
  assign n229 = ~x96 & n228 ;
  assign n230 = x118 & ~n229 ;
  assign n231 = n227 & n230 ;
  assign n233 = x78 & x101 ;
  assign n234 = n233 ^ x38 ^ 1'b0 ;
  assign n235 = n234 ^ x20 ^ 1'b0 ;
  assign n232 = x7 & n153 ;
  assign n236 = n235 ^ n232 ^ 1'b0 ;
  assign n237 = x104 ^ x59 ^ x50 ;
  assign n238 = x123 & ~n237 ;
  assign n239 = n236 & n238 ;
  assign n240 = n218 & n239 ;
  assign n241 = x118 ^ x46 ^ 1'b0 ;
  assign n242 = ( x64 & n145 ) | ( x64 & n159 ) | ( n145 & n159 ) ;
  assign n243 = n242 ^ n173 ^ 1'b0 ;
  assign n244 = n193 ^ x122 ^ 1'b0 ;
  assign n245 = x39 & ~n244 ;
  assign n246 = x28 & ~n166 ;
  assign n247 = n246 ^ x63 ^ 1'b0 ;
  assign n248 = n247 ^ x92 ^ x75 ;
  assign n249 = n248 ^ x16 ^ 1'b0 ;
  assign n250 = n156 & n249 ;
  assign n251 = n250 ^ x11 ^ 1'b0 ;
  assign n252 = ~n234 & n251 ;
  assign n253 = x39 & x51 ;
  assign n254 = ~x102 & n253 ;
  assign n255 = x109 & ~n215 ;
  assign n256 = ~x9 & n255 ;
  assign n257 = x52 | n256 ;
  assign n258 = x116 & ~n166 ;
  assign n259 = x60 & ~n258 ;
  assign n260 = n132 & n215 ;
  assign n261 = x20 & n173 ;
  assign n262 = x88 | n155 ;
  assign n263 = x99 ^ x22 ^ 1'b0 ;
  assign n264 = n156 & n263 ;
  assign n265 = n264 ^ n138 ^ x33 ;
  assign n266 = n189 | n265 ;
  assign n267 = n182 & ~n266 ;
  assign n268 = x59 & n235 ;
  assign n269 = ~n153 & n268 ;
  assign n270 = n247 ^ n227 ^ 1'b0 ;
  assign n271 = ~n247 & n270 ;
  assign n272 = n173 & n271 ;
  assign n273 = n272 ^ x36 ^ 1'b0 ;
  assign n274 = n269 | n273 ;
  assign n275 = n274 ^ n221 ^ 1'b0 ;
  assign n276 = n229 ^ x62 ^ x9 ;
  assign n277 = n161 ^ x113 ^ 1'b0 ;
  assign n278 = n277 ^ x95 ^ 1'b0 ;
  assign n279 = n276 & ~n278 ;
  assign n280 = ( ~x121 & x122 ) | ( ~x121 & n191 ) | ( x122 & n191 ) ;
  assign n281 = n275 ^ x56 ^ 1'b0 ;
  assign n282 = n141 & ~n281 ;
  assign n283 = ( ~x117 & n191 ) | ( ~x117 & n242 ) | ( n191 & n242 ) ;
  assign n284 = x99 ^ x47 ^ 1'b0 ;
  assign n285 = n283 & n284 ;
  assign n286 = x29 & x115 ;
  assign n287 = n286 ^ n200 ^ 1'b0 ;
  assign n288 = n142 | n287 ;
  assign n289 = x119 & ~n288 ;
  assign n290 = ~n285 & n289 ;
  assign n292 = x56 & x99 ;
  assign n293 = ~x88 & n292 ;
  assign n294 = x77 & ~n293 ;
  assign n295 = n294 ^ x13 ^ 1'b0 ;
  assign n291 = x7 & ~n177 ;
  assign n296 = n295 ^ n291 ^ 1'b0 ;
  assign n297 = x68 ^ x38 ^ 1'b0 ;
  assign n298 = n297 ^ n197 ^ 1'b0 ;
  assign n299 = ~n158 & n298 ;
  assign n300 = n296 & n299 ;
  assign n301 = ~n194 & n300 ;
  assign n307 = x107 & x119 ;
  assign n305 = ( ~x31 & x53 ) | ( ~x31 & x106 ) | ( x53 & x106 ) ;
  assign n302 = x66 & x105 ;
  assign n303 = n302 ^ x10 ^ 1'b0 ;
  assign n304 = x61 & ~n303 ;
  assign n306 = n305 ^ n304 ^ 1'b0 ;
  assign n308 = n307 ^ n306 ^ n261 ;
  assign n309 = n308 ^ n212 ^ 1'b0 ;
  assign n310 = ~x4 & x115 ;
  assign n311 = x99 & n269 ;
  assign n312 = n311 ^ n151 ^ x0 ;
  assign n313 = n308 ^ x19 ^ 1'b0 ;
  assign n314 = x22 & n313 ;
  assign n315 = x44 & n314 ;
  assign n316 = n315 ^ x99 ^ 1'b0 ;
  assign n321 = x56 ^ x6 ^ 1'b0 ;
  assign n322 = x74 & n321 ;
  assign n323 = ( x76 & n142 ) | ( x76 & n322 ) | ( n142 & n322 ) ;
  assign n317 = x103 ^ x75 ^ x4 ;
  assign n324 = n323 ^ n317 ^ 1'b0 ;
  assign n318 = x84 & n145 ;
  assign n319 = ~x126 & n318 ;
  assign n320 = ( x13 & n317 ) | ( x13 & n319 ) | ( n317 & n319 ) ;
  assign n325 = n324 ^ n320 ^ 1'b0 ;
  assign n326 = n242 ^ x67 ^ x52 ;
  assign n327 = x30 | n326 ;
  assign n328 = ( x19 & x100 ) | ( x19 & ~n264 ) | ( x100 & ~n264 ) ;
  assign n329 = x10 & x112 ;
  assign n330 = ~n156 & n329 ;
  assign n331 = ( ~n132 & n328 ) | ( ~n132 & n330 ) | ( n328 & n330 ) ;
  assign n332 = ( x14 & x116 ) | ( x14 & n331 ) | ( x116 & n331 ) ;
  assign n333 = n332 ^ x39 ^ 1'b0 ;
  assign n334 = n333 ^ x45 ^ 1'b0 ;
  assign n335 = n327 & ~n334 ;
  assign n336 = n193 ^ x122 ^ x50 ;
  assign n337 = x102 & ~n229 ;
  assign n338 = ( n182 & n336 ) | ( n182 & ~n337 ) | ( n336 & ~n337 ) ;
  assign n339 = x28 & ~n338 ;
  assign n340 = n339 ^ n141 ^ 1'b0 ;
  assign n341 = ~x13 & x67 ;
  assign n342 = x77 ^ x51 ^ x1 ;
  assign n343 = n225 ^ n216 ^ x28 ;
  assign n344 = n343 ^ n130 ^ 1'b0 ;
  assign n345 = ~n342 & n344 ;
  assign n346 = ~x94 & n345 ;
  assign n347 = n341 & ~n346 ;
  assign n348 = ~x71 & n347 ;
  assign n349 = ~x34 & x44 ;
  assign n350 = ~x29 & x124 ;
  assign n351 = x71 ^ x67 ^ 1'b0 ;
  assign n352 = x77 & n351 ;
  assign n353 = ~x38 & n352 ;
  assign n354 = x90 & ~n293 ;
  assign n355 = n354 ^ n283 ^ 1'b0 ;
  assign n356 = n355 ^ x118 ^ 1'b0 ;
  assign n357 = n353 | n356 ;
  assign n358 = x75 & ~n166 ;
  assign n359 = n206 & n358 ;
  assign n360 = x89 & n134 ;
  assign n361 = n359 & n360 ;
  assign n362 = ( n156 & n296 ) | ( n156 & n317 ) | ( n296 & n317 ) ;
  assign n363 = ~x36 & x38 ;
  assign n365 = x32 & x113 ;
  assign n366 = ~n150 & n365 ;
  assign n364 = x114 & ~n166 ;
  assign n367 = n366 ^ n364 ^ 1'b0 ;
  assign n370 = x5 & x35 ;
  assign n368 = n161 ^ x126 ^ x77 ;
  assign n369 = ( x36 & ~x114 ) | ( x36 & n368 ) | ( ~x114 & n368 ) ;
  assign n371 = n370 ^ n369 ^ 1'b0 ;
  assign n372 = ~n220 & n237 ;
  assign n373 = ( x37 & ~x86 ) | ( x37 & x92 ) | ( ~x86 & x92 ) ;
  assign n374 = n373 ^ x18 ^ 1'b0 ;
  assign n375 = n374 ^ x31 ^ 1'b0 ;
  assign n376 = x5 & ~n375 ;
  assign n379 = n163 ^ x124 ^ x122 ;
  assign n377 = n335 ^ x116 ^ x113 ;
  assign n378 = n363 | n377 ;
  assign n380 = n379 ^ n378 ^ 1'b0 ;
  assign n381 = ~x23 & n156 ;
  assign n382 = x23 & ~n237 ;
  assign n383 = ~x14 & n382 ;
  assign n384 = x21 & ~n383 ;
  assign n385 = n384 ^ n169 ^ 1'b0 ;
  assign n386 = ( x79 & ~x118 ) | ( x79 & n385 ) | ( ~x118 & n385 ) ;
  assign n387 = x84 & x89 ;
  assign n388 = ( x34 & n146 ) | ( x34 & ~n185 ) | ( n146 & ~n185 ) ;
  assign n389 = ~n202 & n388 ;
  assign n390 = n389 ^ x17 ^ 1'b0 ;
  assign n391 = n293 ^ x43 ^ x35 ;
  assign n392 = x35 & x118 ;
  assign n393 = ~x34 & n392 ;
  assign n394 = x119 & ~n393 ;
  assign n395 = n394 ^ n242 ^ 1'b0 ;
  assign n396 = n130 & n395 ;
  assign n397 = n227 | n260 ;
  assign n398 = x58 | n397 ;
  assign n399 = ( n149 & n252 ) | ( n149 & ~n398 ) | ( n252 & ~n398 ) ;
  assign n400 = n370 ^ x94 ^ 1'b0 ;
  assign n401 = ~n167 & n400 ;
  assign n402 = n305 ^ n191 ^ 1'b0 ;
  assign n403 = ~n204 & n402 ;
  assign n404 = x9 | n330 ;
  assign n405 = n403 & n404 ;
  assign n406 = ~n275 & n405 ;
  assign n407 = n183 ^ x103 ^ x32 ;
  assign n408 = ( x29 & ~n306 ) | ( x29 & n407 ) | ( ~n306 & n407 ) ;
  assign n409 = ~x1 & n408 ;
  assign n410 = n145 & ~n227 ;
  assign n411 = n383 ^ n370 ^ n199 ;
  assign n417 = n175 ^ n143 ^ 1'b0 ;
  assign n418 = ~n297 & n417 ;
  assign n412 = x91 & x103 ;
  assign n413 = ~x26 & n412 ;
  assign n414 = n352 ^ x38 ^ 1'b0 ;
  assign n415 = ~n413 & n414 ;
  assign n416 = ( x20 & n225 ) | ( x20 & n415 ) | ( n225 & n415 ) ;
  assign n419 = n418 ^ n416 ^ x110 ;
  assign n421 = x36 & n194 ;
  assign n420 = x69 & n285 ;
  assign n422 = n421 ^ n420 ^ n404 ;
  assign n423 = n204 ^ x50 ^ 1'b0 ;
  assign n424 = x71 & ~n423 ;
  assign n425 = x94 & n161 ;
  assign n426 = n142 | n425 ;
  assign n427 = x9 | n426 ;
  assign n428 = n401 ^ x39 ^ 1'b0 ;
  assign n429 = n427 & n428 ;
  assign n432 = x48 ^ x16 ^ 1'b0 ;
  assign n433 = ~n200 & n432 ;
  assign n430 = n143 ^ x11 ^ 1'b0 ;
  assign n431 = n322 & n430 ;
  assign n434 = n433 ^ n431 ^ 1'b0 ;
  assign n435 = n176 & n434 ;
  assign n436 = n435 ^ x75 ^ 1'b0 ;
  assign n437 = x93 & n436 ;
  assign n438 = ~n408 & n437 ;
  assign n441 = n158 ^ x23 ^ 1'b0 ;
  assign n442 = n166 | n441 ;
  assign n439 = ~x74 & n435 ;
  assign n440 = n310 | n439 ;
  assign n443 = n442 ^ n440 ^ 1'b0 ;
  assign n444 = x109 & n129 ;
  assign n445 = n444 ^ x26 ^ 1'b0 ;
  assign n446 = n369 | n445 ;
  assign n447 = n446 ^ x50 ^ 1'b0 ;
  assign n448 = ~n442 & n447 ;
  assign n449 = n448 ^ x12 ^ 1'b0 ;
  assign n450 = ( x25 & ~n223 ) | ( x25 & n403 ) | ( ~n223 & n403 ) ;
  assign n451 = ( x62 & x76 ) | ( x62 & ~n450 ) | ( x76 & ~n450 ) ;
  assign n452 = n346 ^ x117 ^ x114 ;
  assign n453 = n416 ^ x33 ^ 1'b0 ;
  assign n454 = n452 & n453 ;
  assign n455 = x32 & ~n259 ;
  assign n456 = ~n454 & n455 ;
  assign n461 = ~x5 & n257 ;
  assign n457 = x58 ^ x28 ^ 1'b0 ;
  assign n458 = n297 & ~n405 ;
  assign n459 = ~n457 & n458 ;
  assign n460 = n259 | n459 ;
  assign n462 = n461 ^ n460 ^ 1'b0 ;
  assign n463 = x62 & n161 ;
  assign n465 = x88 & ~n167 ;
  assign n466 = n393 & n465 ;
  assign n464 = n182 | n234 ;
  assign n467 = n466 ^ n464 ^ 1'b0 ;
  assign n468 = x15 & n311 ;
  assign n469 = n468 ^ x86 ^ 1'b0 ;
  assign n470 = ( x14 & n275 ) | ( x14 & ~n469 ) | ( n275 & ~n469 ) ;
  assign n471 = ~n167 & n227 ;
  assign n472 = x48 & x73 ;
  assign n473 = ~x35 & n472 ;
  assign n474 = n473 ^ x120 ^ 1'b0 ;
  assign n475 = ~x4 & n474 ;
  assign n476 = n442 ^ n199 ^ 1'b0 ;
  assign n477 = n433 & n476 ;
  assign n478 = x105 & n477 ;
  assign n479 = ( x61 & ~n129 ) | ( x61 & n158 ) | ( ~n129 & n158 ) ;
  assign n480 = x47 & ~x69 ;
  assign n481 = n480 ^ x127 ^ 1'b0 ;
  assign n482 = n136 & ~n481 ;
  assign n483 = x101 & n482 ;
  assign n484 = n483 ^ n132 ^ 1'b0 ;
  assign n485 = ~x37 & n401 ;
  assign n486 = n261 ^ n218 ^ 1'b0 ;
  assign n488 = ( x24 & n336 ) | ( x24 & n425 ) | ( n336 & n425 ) ;
  assign n487 = n379 ^ x71 ^ 1'b0 ;
  assign n489 = n488 ^ n487 ^ 1'b0 ;
  assign n490 = ~n240 & n489 ;
  assign n491 = n202 ^ n158 ^ 1'b0 ;
  assign n492 = n245 & n491 ;
  assign n493 = n492 ^ x61 ^ 1'b0 ;
  assign n494 = n265 ^ n138 ^ 1'b0 ;
  assign n495 = x60 & ~n494 ;
  assign n496 = n319 & n495 ;
  assign n497 = x45 & n496 ;
  assign n498 = n254 ^ x115 ^ 1'b0 ;
  assign n502 = x77 ^ x9 ^ 1'b0 ;
  assign n499 = ~x56 & n403 ;
  assign n500 = n189 & n499 ;
  assign n501 = x57 & ~n500 ;
  assign n503 = n502 ^ n501 ^ 1'b0 ;
  assign n504 = x2 & n421 ;
  assign n505 = n504 ^ n269 ^ 1'b0 ;
  assign n506 = x1 & n505 ;
  assign n507 = n506 ^ n449 ^ 1'b0 ;
  assign n508 = n353 ^ x107 ^ 1'b0 ;
  assign n509 = ( x10 & n436 ) | ( x10 & n508 ) | ( n436 & n508 ) ;
  assign n512 = ~x4 & x36 ;
  assign n510 = n326 ^ n220 ^ 1'b0 ;
  assign n511 = x20 & n510 ;
  assign n513 = n512 ^ n511 ^ 1'b0 ;
  assign n514 = n325 & n513 ;
  assign n515 = ~n461 & n514 ;
  assign n517 = n469 ^ n223 ^ 1'b0 ;
  assign n516 = x105 & n457 ;
  assign n518 = n517 ^ n516 ^ 1'b0 ;
  assign n519 = ~n231 & n518 ;
  assign n520 = n312 ^ x65 ^ 1'b0 ;
  assign n521 = n519 & n520 ;
  assign n522 = n188 & n398 ;
  assign n523 = ~n314 & n522 ;
  assign n524 = n254 ^ x26 ^ x20 ;
  assign n525 = ~n518 & n524 ;
  assign n526 = n523 & n525 ;
  assign n528 = n155 | n225 ;
  assign n529 = n264 | n528 ;
  assign n527 = n312 ^ n241 ^ x52 ;
  assign n530 = n529 ^ n527 ^ x54 ;
  assign n531 = x26 & ~n190 ;
  assign n532 = n459 & n531 ;
  assign n533 = n532 ^ n408 ^ 1'b0 ;
  assign n534 = x36 & ~x77 ;
  assign n535 = n534 ^ x63 ^ 1'b0 ;
  assign n536 = n535 ^ n333 ^ x34 ;
  assign n537 = n177 | n536 ;
  assign n538 = n537 ^ n505 ^ 1'b0 ;
  assign n539 = ( x16 & x47 ) | ( x16 & ~n466 ) | ( x47 & ~n466 ) ;
  assign n540 = x29 & x86 ;
  assign n541 = n540 ^ n398 ^ 1'b0 ;
  assign n546 = x36 & x44 ;
  assign n547 = ~n130 & n546 ;
  assign n548 = ( n314 & n396 ) | ( n314 & n547 ) | ( n396 & n547 ) ;
  assign n542 = x103 ^ x49 ^ 1'b0 ;
  assign n543 = ~n393 & n542 ;
  assign n544 = n149 | n543 ;
  assign n545 = n362 & n544 ;
  assign n549 = n548 ^ n545 ^ 1'b0 ;
  assign n550 = n261 ^ x79 ^ 1'b0 ;
  assign n551 = x25 & n550 ;
  assign n552 = n376 & n454 ;
  assign n553 = ~x14 & n552 ;
  assign n554 = n474 & ~n553 ;
  assign n555 = ~n551 & n554 ;
  assign n564 = x72 ^ x33 ^ 1'b0 ;
  assign n565 = n564 ^ n330 ^ x22 ;
  assign n556 = n204 | n317 ;
  assign n557 = x91 | n556 ;
  assign n558 = n254 | n557 ;
  assign n559 = x17 ^ x5 ^ 1'b0 ;
  assign n560 = x127 & n559 ;
  assign n561 = ~n267 & n560 ;
  assign n562 = ~n173 & n561 ;
  assign n563 = n558 | n562 ;
  assign n566 = n565 ^ n563 ^ n297 ;
  assign n573 = x26 & x59 ;
  assign n574 = n237 & n573 ;
  assign n569 = n237 ^ x22 ^ 1'b0 ;
  assign n568 = ~n303 & n482 ;
  assign n570 = n569 ^ n568 ^ 1'b0 ;
  assign n567 = ( x13 & ~x86 ) | ( x13 & x107 ) | ( ~x86 & x107 ) ;
  assign n571 = n570 ^ n567 ^ x116 ;
  assign n572 = x88 & ~n571 ;
  assign n575 = n574 ^ n572 ^ 1'b0 ;
  assign n576 = n575 ^ x45 ^ x23 ;
  assign n577 = n576 ^ n357 ^ 1'b0 ;
  assign n578 = ( n196 & ~n283 ) | ( n196 & n474 ) | ( ~n283 & n474 ) ;
  assign n579 = n346 & n497 ;
  assign n580 = x71 & ~n306 ;
  assign n581 = ~x78 & n580 ;
  assign n582 = n581 ^ n239 ^ 1'b0 ;
  assign n583 = x28 & n141 ;
  assign n584 = n583 ^ n285 ^ 1'b0 ;
  assign n585 = n584 ^ x5 ^ 1'b0 ;
  assign n586 = n560 & ~n585 ;
  assign n587 = n547 ^ n381 ^ 1'b0 ;
  assign n588 = n336 & n587 ;
  assign n589 = n586 & n588 ;
  assign n590 = n132 & n589 ;
  assign n591 = n227 ^ n186 ^ 1'b0 ;
  assign n592 = ~n333 & n591 ;
  assign n593 = ( ~x90 & n415 ) | ( ~x90 & n592 ) | ( n415 & n592 ) ;
  assign n594 = ( ~x71 & x88 ) | ( ~x71 & n264 ) | ( x88 & n264 ) ;
  assign n595 = ~n359 & n451 ;
  assign n596 = n595 ^ n374 ^ 1'b0 ;
  assign n597 = n594 & n596 ;
  assign n598 = x116 & n597 ;
  assign n599 = n142 & n598 ;
  assign n600 = ~n363 & n433 ;
  assign n601 = n600 ^ x55 ^ 1'b0 ;
  assign n602 = n173 | n260 ;
  assign n603 = n602 ^ x88 ^ 1'b0 ;
  assign n604 = n443 ^ x25 ^ 1'b0 ;
  assign n605 = n215 | n604 ;
  assign n606 = n605 ^ n553 ^ x68 ;
  assign n607 = n413 ^ n353 ^ x42 ;
  assign n608 = ~x1 & n305 ;
  assign n609 = ~n320 & n608 ;
  assign n610 = n607 & n609 ;
  assign n611 = n586 ^ n376 ^ 1'b0 ;
  assign n612 = ~n610 & n611 ;
  assign n615 = n194 | n234 ;
  assign n613 = x100 ^ x86 ^ 1'b0 ;
  assign n614 = n575 & ~n613 ;
  assign n616 = n615 ^ n614 ^ 1'b0 ;
  assign n617 = n293 ^ n280 ^ 1'b0 ;
  assign n618 = x81 | n617 ;
  assign n619 = n618 ^ x75 ^ 1'b0 ;
  assign n620 = n216 & ~n416 ;
  assign n621 = n620 ^ n418 ^ x85 ;
  assign n630 = ( ~x91 & n188 ) | ( ~x91 & n275 ) | ( n188 & n275 ) ;
  assign n624 = n336 & ~n473 ;
  assign n625 = ~n286 & n624 ;
  assign n626 = n519 ^ n301 ^ 1'b0 ;
  assign n627 = n625 | n626 ;
  assign n623 = n303 ^ x89 ^ 1'b0 ;
  assign n628 = n627 ^ n623 ^ n271 ;
  assign n629 = x21 & ~n628 ;
  assign n631 = n630 ^ n629 ^ 1'b0 ;
  assign n622 = x117 & n433 ;
  assign n632 = n631 ^ n622 ^ 1'b0 ;
  assign n633 = n387 ^ x43 ^ 1'b0 ;
  assign n634 = x100 & x112 ;
  assign n635 = n229 & n634 ;
  assign n636 = n635 ^ n225 ^ 1'b0 ;
  assign n642 = n293 & n454 ;
  assign n637 = x94 & n296 ;
  assign n638 = n637 ^ x59 ^ 1'b0 ;
  assign n639 = x10 | n638 ;
  assign n640 = n639 ^ x18 ^ 1'b0 ;
  assign n641 = x11 & ~n640 ;
  assign n643 = n642 ^ n641 ^ 1'b0 ;
  assign n644 = n625 ^ n521 ^ n519 ;
  assign n645 = ( x88 & ~n264 ) | ( x88 & n405 ) | ( ~n264 & n405 ) ;
  assign n646 = n343 ^ n254 ^ 1'b0 ;
  assign n647 = x82 & x109 ;
  assign n648 = n148 & n647 ;
  assign n649 = n439 | n648 ;
  assign n650 = n649 ^ n486 ^ 1'b0 ;
  assign n651 = n142 | n404 ;
  assign n652 = n383 & ~n651 ;
  assign n653 = ( n323 & ~n651 ) | ( n323 & n652 ) | ( ~n651 & n652 ) ;
  assign n654 = n653 ^ x5 ^ 1'b0 ;
  assign n655 = x127 & n575 ;
  assign n662 = x74 & ~n277 ;
  assign n663 = n662 ^ n534 ^ 1'b0 ;
  assign n656 = n413 ^ n235 ^ 1'b0 ;
  assign n657 = n247 | n656 ;
  assign n658 = n136 ^ x119 ^ 1'b0 ;
  assign n659 = x109 & n658 ;
  assign n660 = ~n657 & n659 ;
  assign n661 = ~n146 & n660 ;
  assign n664 = n663 ^ n661 ^ x97 ;
  assign n665 = x110 & ~x123 ;
  assign n666 = x33 & x126 ;
  assign n667 = n666 ^ n345 ^ 1'b0 ;
  assign n668 = x62 & x102 ;
  assign n669 = x78 & n258 ;
  assign n670 = ~n173 & n669 ;
  assign n671 = n668 & ~n670 ;
  assign n672 = x59 & n202 ;
  assign n673 = n518 ^ x6 ^ 1'b0 ;
  assign n674 = ( x90 & n199 ) | ( x90 & ~n673 ) | ( n199 & ~n673 ) ;
  assign n675 = n551 & n674 ;
  assign n676 = n675 ^ n273 ^ 1'b0 ;
  assign n677 = n398 & ~n676 ;
  assign n678 = n146 & ~n189 ;
  assign n679 = ~n383 & n408 ;
  assign n680 = n508 & n679 ;
  assign n681 = n680 ^ n482 ^ 1'b0 ;
  assign n685 = n167 | n383 ;
  assign n686 = n685 ^ n177 ^ 1'b0 ;
  assign n687 = n355 & ~n686 ;
  assign n682 = n352 ^ n326 ^ 1'b0 ;
  assign n683 = x38 & ~n682 ;
  assign n684 = n672 & n683 ;
  assign n688 = n687 ^ n684 ^ 1'b0 ;
  assign n689 = n508 ^ x72 ^ 1'b0 ;
  assign n690 = n416 & ~n689 ;
  assign n691 = ( n193 & n433 ) | ( n193 & n488 ) | ( n433 & n488 ) ;
  assign n692 = n488 ^ x29 ^ 1'b0 ;
  assign n693 = n691 & n692 ;
  assign n694 = n693 ^ x70 ^ 1'b0 ;
  assign n695 = x41 & x45 ;
  assign n696 = n165 & n695 ;
  assign n697 = n696 ^ n664 ^ n461 ;
  assign n699 = x78 & x115 ;
  assign n700 = ~x29 & n699 ;
  assign n698 = ~x27 & n483 ;
  assign n701 = n700 ^ n698 ^ n558 ;
  assign n702 = n326 & ~n701 ;
  assign n710 = n385 & ~n558 ;
  assign n711 = n710 ^ n547 ^ 1'b0 ;
  assign n705 = x33 & n311 ;
  assign n706 = n306 & n705 ;
  assign n707 = ( x31 & ~n216 ) | ( x31 & n706 ) | ( ~n216 & n706 ) ;
  assign n708 = n620 & ~n707 ;
  assign n709 = x94 & n708 ;
  assign n712 = n711 ^ n709 ^ 1'b0 ;
  assign n703 = ~n242 & n529 ;
  assign n704 = n653 & n703 ;
  assign n713 = n712 ^ n704 ^ 1'b0 ;
  assign n715 = n385 ^ n286 ^ 1'b0 ;
  assign n716 = x98 & n715 ;
  assign n714 = x19 & ~n306 ;
  assign n717 = n716 ^ n714 ^ 1'b0 ;
  assign n718 = ( x49 & ~x100 ) | ( x49 & n215 ) | ( ~x100 & n215 ) ;
  assign n719 = ( x64 & n717 ) | ( x64 & ~n718 ) | ( n717 & ~n718 ) ;
  assign n720 = ( n361 & ~n372 ) | ( n361 & n477 ) | ( ~n372 & n477 ) ;
  assign n721 = n720 ^ x63 ^ 1'b0 ;
  assign n722 = ~n553 & n721 ;
  assign n723 = n722 ^ n673 ^ 1'b0 ;
  assign n724 = x87 & ~n723 ;
  assign n725 = ~x113 & n724 ;
  assign n726 = x28 & ~n403 ;
  assign n728 = n368 ^ x110 ^ x13 ;
  assign n727 = n457 & ~n696 ;
  assign n729 = n728 ^ n727 ^ 1'b0 ;
  assign n730 = n668 ^ x65 ^ 1'b0 ;
  assign n731 = n730 ^ n190 ^ x26 ;
  assign n732 = x117 & n136 ;
  assign n733 = n732 ^ x12 ^ 1'b0 ;
  assign n734 = ~x19 & n544 ;
  assign n735 = n734 ^ n332 ^ 1'b0 ;
  assign n736 = n733 | n735 ;
  assign n737 = n408 & n482 ;
  assign n738 = n736 & n737 ;
  assign n739 = ~n399 & n671 ;
  assign n743 = x95 & ~n407 ;
  assign n744 = ~n129 & n743 ;
  assign n740 = n214 ^ x70 ^ 1'b0 ;
  assign n741 = n740 ^ n462 ^ 1'b0 ;
  assign n742 = n220 | n741 ;
  assign n745 = n744 ^ n742 ^ x30 ;
  assign n746 = n673 & ~n691 ;
  assign n747 = x122 ^ x2 ^ 1'b0 ;
  assign n748 = x67 & n747 ;
  assign n749 = n748 ^ x101 ^ 1'b0 ;
  assign n750 = n487 & n749 ;
  assign n751 = x108 & ~n409 ;
  assign n752 = n751 ^ n387 ^ 1'b0 ;
  assign n753 = ( ~x19 & n750 ) | ( ~x19 & n752 ) | ( n750 & n752 ) ;
  assign n754 = n153 ^ x109 ^ 1'b0 ;
  assign n755 = n754 ^ n492 ^ n327 ;
  assign n756 = x112 | n755 ;
  assign n757 = ( n341 & ~n753 ) | ( n341 & n756 ) | ( ~n753 & n756 ) ;
  assign n758 = n746 & ~n757 ;
  assign n759 = n327 & n389 ;
  assign n760 = n759 ^ x66 ^ 1'b0 ;
  assign n761 = n186 | n648 ;
  assign n762 = n142 & ~n761 ;
  assign n763 = n762 ^ n744 ^ n651 ;
  assign n764 = ~x36 & x123 ;
  assign n765 = n562 ^ n290 ^ x100 ;
  assign n766 = n765 ^ x94 ^ 1'b0 ;
  assign n767 = n764 & n766 ;
  assign n768 = x62 & ~n635 ;
  assign n769 = n768 ^ n141 ^ 1'b0 ;
  assign n770 = n769 ^ n173 ^ 1'b0 ;
  assign n771 = ( x100 & ~n183 ) | ( x100 & n530 ) | ( ~n183 & n530 ) ;
  assign n772 = n771 ^ n508 ^ 1'b0 ;
  assign n773 = n197 & n772 ;
  assign n774 = n612 & n773 ;
  assign n775 = ~n770 & n774 ;
  assign n776 = n707 | n775 ;
  assign n777 = x91 | n776 ;
  assign n779 = ( x1 & ~x21 ) | ( x1 & x45 ) | ( ~x21 & x45 ) ;
  assign n778 = n553 ^ n418 ^ 1'b0 ;
  assign n780 = n779 ^ n778 ^ 1'b0 ;
  assign n781 = x47 & n780 ;
  assign n782 = n188 ^ x57 ^ 1'b0 ;
  assign n783 = ~n265 & n782 ;
  assign n784 = n484 & n783 ;
  assign n785 = n784 ^ x60 ^ 1'b0 ;
  assign n786 = ( n410 & ~n781 ) | ( n410 & n785 ) | ( ~n781 & n785 ) ;
  assign n787 = n618 ^ n416 ^ 1'b0 ;
  assign n788 = x40 & n787 ;
  assign n789 = n584 ^ n463 ^ 1'b0 ;
  assign n790 = n290 | n789 ;
  assign n793 = ( ~n146 & n311 ) | ( ~n146 & n413 ) | ( n311 & n413 ) ;
  assign n791 = x112 ^ x10 ^ 1'b0 ;
  assign n792 = n733 | n791 ;
  assign n794 = n793 ^ n792 ^ 1'b0 ;
  assign n795 = n794 ^ n231 ^ 1'b0 ;
  assign n796 = x1 & n795 ;
  assign n797 = ~n148 & n796 ;
  assign n798 = n797 ^ n286 ^ 1'b0 ;
  assign n799 = n467 & ~n584 ;
  assign n800 = n471 ^ x30 ^ 1'b0 ;
  assign n801 = x29 & ~n800 ;
  assign n802 = n264 & n801 ;
  assign n803 = n183 & n241 ;
  assign n804 = n803 ^ n286 ^ 1'b0 ;
  assign n805 = n535 ^ n250 ^ 1'b0 ;
  assign n806 = n427 ^ x106 ^ x25 ;
  assign n807 = n805 & ~n806 ;
  assign n808 = ~n379 & n807 ;
  assign n809 = n299 ^ x91 ^ 1'b0 ;
  assign n810 = n616 | n809 ;
  assign n811 = n810 ^ n574 ^ 1'b0 ;
  assign n812 = x5 & ~n214 ;
  assign n813 = n812 ^ n541 ^ n409 ;
  assign n814 = x37 ^ x26 ^ 1'b0 ;
  assign n815 = n452 & n814 ;
  assign n816 = n815 ^ n424 ^ 1'b0 ;
  assign n817 = n813 & n816 ;
  assign n818 = n308 ^ n190 ^ x16 ;
  assign n819 = n297 & n818 ;
  assign n820 = ~n306 & n819 ;
  assign n821 = n558 & n820 ;
  assign n822 = x109 & n250 ;
  assign n823 = n822 ^ n385 ^ 1'b0 ;
  assign n824 = n823 ^ n176 ^ 1'b0 ;
  assign n825 = n752 ^ n250 ^ 1'b0 ;
  assign n826 = n145 & ~n825 ;
  assign n827 = ~x94 & n248 ;
  assign n828 = ( n264 & n333 ) | ( n264 & n827 ) | ( n333 & n827 ) ;
  assign n829 = n828 ^ n678 ^ n130 ;
  assign n830 = n264 ^ n254 ^ n236 ;
  assign n831 = n691 ^ n190 ^ n141 ;
  assign n832 = n651 ^ n619 ^ n262 ;
  assign n834 = n635 ^ x93 ^ 1'b0 ;
  assign n835 = n197 & ~n834 ;
  assign n833 = x79 ^ x10 ^ 1'b0 ;
  assign n836 = n835 ^ n833 ^ 1'b0 ;
  assign n837 = n760 ^ x101 ^ 1'b0 ;
  assign n838 = ( ~x53 & x119 ) | ( ~x53 & n372 ) | ( x119 & n372 ) ;
  assign n839 = n838 ^ n527 ^ 1'b0 ;
  assign n840 = ~n331 & n839 ;
  assign n841 = ~n331 & n655 ;
  assign n842 = ~x66 & n841 ;
  assign n843 = x36 & n773 ;
  assign n844 = n843 ^ n661 ^ 1'b0 ;
  assign n853 = x31 & ~n229 ;
  assign n854 = ~x52 & n853 ;
  assign n855 = n854 ^ x94 ^ 1'b0 ;
  assign n856 = n254 | n855 ;
  assign n850 = x17 & n190 ;
  assign n851 = n369 | n850 ;
  assign n852 = n851 ^ n640 ^ 1'b0 ;
  assign n845 = n171 | n330 ;
  assign n846 = ~x81 & n779 ;
  assign n847 = n846 ^ n569 ^ 1'b0 ;
  assign n848 = n845 & ~n847 ;
  assign n849 = n387 & ~n848 ;
  assign n857 = n856 ^ n852 ^ n849 ;
  assign n858 = n411 ^ n150 ^ x3 ;
  assign n859 = ~n857 & n858 ;
  assign n860 = n518 ^ n303 ^ 1'b0 ;
  assign n861 = ~n217 & n860 ;
  assign n862 = n497 ^ n236 ^ 1'b0 ;
  assign n863 = n861 & ~n862 ;
  assign n864 = n863 ^ n527 ^ 1'b0 ;
  assign n865 = n856 | n864 ;
  assign n866 = n409 | n865 ;
  assign n867 = x42 | n866 ;
  assign n868 = n327 & ~n509 ;
  assign n869 = n868 ^ n500 ^ n202 ;
  assign n870 = x15 & ~n155 ;
  assign n871 = n870 ^ x49 ^ 1'b0 ;
  assign n872 = n871 ^ n499 ^ 1'b0 ;
  assign n873 = ( x78 & n391 ) | ( x78 & n872 ) | ( n391 & n872 ) ;
  assign n874 = n873 ^ n260 ^ 1'b0 ;
  assign n875 = n692 & ~n874 ;
  assign n876 = n875 ^ n736 ^ 1'b0 ;
  assign n877 = x40 ^ x7 ^ 1'b0 ;
  assign n878 = x86 & ~n830 ;
  assign n879 = ~x37 & n878 ;
  assign n880 = n879 ^ x84 ^ 1'b0 ;
  assign n881 = n742 | n880 ;
  assign n882 = n410 ^ n163 ^ 1'b0 ;
  assign n885 = x69 & n262 ;
  assign n886 = n885 ^ n319 ^ 1'b0 ;
  assign n883 = ~x3 & n835 ;
  assign n884 = n883 ^ x58 ^ x51 ;
  assign n887 = n886 ^ n884 ^ 1'b0 ;
  assign n888 = n663 & ~n887 ;
  assign n889 = x65 | n616 ;
  assign n890 = ( n200 & ~n771 ) | ( n200 & n889 ) | ( ~n771 & n889 ) ;
  assign n891 = ( ~x80 & x94 ) | ( ~x80 & n190 ) | ( x94 & n190 ) ;
  assign n892 = ( n129 & n190 ) | ( n129 & ~n891 ) | ( n190 & ~n891 ) ;
  assign n893 = n892 ^ n819 ^ 1'b0 ;
  assign n894 = x120 & ~n217 ;
  assign n895 = ~n893 & n894 ;
  assign n896 = ( n149 & n371 ) | ( n149 & ~n493 ) | ( n371 & ~n493 ) ;
  assign n897 = n896 ^ n256 ^ 1'b0 ;
  assign n898 = n176 & ~n576 ;
  assign n899 = n214 & n898 ;
  assign n900 = n899 ^ n310 ^ 1'b0 ;
  assign n901 = n433 & n900 ;
  assign n904 = n341 | n418 ;
  assign n905 = n904 ^ n848 ^ 1'b0 ;
  assign n902 = n530 ^ x54 ^ 1'b0 ;
  assign n903 = ~n842 & n902 ;
  assign n906 = n905 ^ n903 ^ 1'b0 ;
  assign n907 = n809 ^ n738 ^ 1'b0 ;
  assign n908 = ~x20 & n161 ;
  assign n909 = n355 ^ n242 ^ n132 ;
  assign n910 = n908 & n909 ;
  assign n911 = n478 ^ x63 ^ 1'b0 ;
  assign n912 = ~n696 & n911 ;
  assign n913 = n912 ^ n739 ^ 1'b0 ;
  assign n914 = ~n877 & n913 ;
  assign n916 = n293 ^ n235 ^ 1'b0 ;
  assign n917 = n409 | n916 ;
  assign n918 = n917 ^ x77 ^ 1'b0 ;
  assign n919 = x68 ^ x3 ^ 1'b0 ;
  assign n920 = n918 & ~n919 ;
  assign n921 = x24 & n920 ;
  assign n922 = ~n643 & n921 ;
  assign n915 = n697 | n769 ;
  assign n923 = n922 ^ n915 ^ 1'b0 ;
  assign n924 = n923 ^ n457 ^ 1'b0 ;
  assign n925 = x103 & ~n924 ;
  assign n926 = n590 ^ n533 ^ 1'b0 ;
  assign n927 = ~n896 & n926 ;
  assign n928 = n804 ^ n676 ^ n406 ;
  assign n929 = ~n149 & n341 ;
  assign n931 = x23 & x79 ;
  assign n932 = ~x49 & n931 ;
  assign n930 = n279 ^ n258 ^ 1'b0 ;
  assign n933 = n932 ^ n930 ^ 1'b0 ;
  assign n934 = n240 & ~n932 ;
  assign n935 = n889 | n934 ;
  assign n936 = ~n933 & n935 ;
  assign n937 = ~n929 & n936 ;
  assign n938 = x42 | n277 ;
  assign n939 = n938 ^ n746 ^ n636 ;
  assign n940 = x127 & n555 ;
  assign n941 = x29 & ~n706 ;
  assign n942 = n940 & n941 ;
  assign n943 = ( n456 & n485 ) | ( n456 & n919 ) | ( n485 & n919 ) ;
  assign n944 = n383 ^ n296 ^ x123 ;
  assign n945 = ~n362 & n944 ;
  assign n946 = n330 ^ x16 ^ 1'b0 ;
  assign n947 = ( x22 & x87 ) | ( x22 & n733 ) | ( x87 & n733 ) ;
  assign n948 = n947 ^ n179 ^ 1'b0 ;
  assign n949 = n374 & ~n948 ;
  assign n950 = n946 & n949 ;
  assign n951 = n349 | n377 ;
  assign n952 = n951 ^ n282 ^ 1'b0 ;
  assign n953 = ~n655 & n952 ;
  assign n954 = ( n311 & n405 ) | ( n311 & n648 ) | ( n405 & n648 ) ;
  assign n955 = ( x60 & n186 ) | ( x60 & n954 ) | ( n186 & n954 ) ;
  assign n956 = n891 ^ n706 ^ n297 ;
  assign n957 = n221 | n484 ;
  assign n958 = n645 ^ n451 ^ 1'b0 ;
  assign n959 = n584 | n958 ;
  assign n960 = x18 & ~n499 ;
  assign n961 = x36 & n960 ;
  assign n962 = n961 ^ n930 ^ n241 ;
  assign n963 = n944 ^ n261 ^ 1'b0 ;
  assign n964 = x120 & n963 ;
  assign n965 = n858 ^ n293 ^ 1'b0 ;
  assign n966 = n965 ^ n557 ^ 1'b0 ;
  assign n967 = n771 | n966 ;
  assign n968 = x49 & n322 ;
  assign n969 = n968 ^ x108 ^ 1'b0 ;
  assign n970 = n171 & n969 ;
  assign n971 = n970 ^ x15 ^ 1'b0 ;
  assign n972 = n413 | n971 ;
  assign n973 = ~n327 & n371 ;
  assign n974 = n973 ^ n348 ^ n145 ;
  assign n975 = n974 ^ n690 ^ 1'b0 ;
  assign n976 = n497 & ~n953 ;
  assign n977 = ~x113 & n976 ;
  assign n978 = n265 & n672 ;
  assign n979 = x29 & ~n188 ;
  assign n980 = n979 ^ n909 ^ 1'b0 ;
  assign n981 = n980 ^ n500 ^ 1'b0 ;
  assign n982 = n978 | n981 ;
  assign n983 = x21 & ~n191 ;
  assign n984 = n683 ^ n561 ^ 1'b0 ;
  assign n985 = x57 & ~n670 ;
  assign n986 = n725 & n985 ;
  assign n987 = ~n984 & n986 ;
  assign n988 = ( n459 & n605 ) | ( n459 & n987 ) | ( n605 & n987 ) ;
  assign n989 = n564 & n582 ;
  assign n990 = ~x124 & n989 ;
  assign n992 = x50 & n297 ;
  assign n993 = n488 & n992 ;
  assign n994 = n993 ^ n535 ^ 1'b0 ;
  assign n995 = n994 ^ n593 ^ 1'b0 ;
  assign n996 = x7 & n995 ;
  assign n991 = n370 & n683 ;
  assign n997 = n996 ^ n991 ^ 1'b0 ;
  assign n998 = ( ~n541 & n654 ) | ( ~n541 & n899 ) | ( n654 & n899 ) ;
  assign n999 = x57 & ~n186 ;
  assign n1000 = ~n889 & n999 ;
  assign n1001 = n1000 ^ n435 ^ n337 ;
  assign n1002 = n349 ^ n330 ^ 1'b0 ;
  assign n1003 = x58 | n494 ;
  assign n1004 = ( n821 & n1002 ) | ( n821 & ~n1003 ) | ( n1002 & ~n1003 ) ;
  assign n1005 = x75 ^ x38 ^ 1'b0 ;
  assign n1006 = n311 & n1005 ;
  assign n1007 = x118 & n312 ;
  assign n1008 = ~n370 & n1007 ;
  assign n1009 = n1006 & n1008 ;
  assign n1010 = x39 & n854 ;
  assign n1011 = x6 & ~n969 ;
  assign n1012 = n1011 ^ x1 ^ 1'b0 ;
  assign n1013 = ~n166 & n1012 ;
  assign n1014 = n439 & ~n707 ;
  assign n1015 = n143 & ~n1014 ;
  assign n1016 = n1015 ^ n497 ^ 1'b0 ;
  assign n1017 = ( n411 & n783 ) | ( n411 & ~n1016 ) | ( n783 & ~n1016 ) ;
  assign n1018 = n507 ^ x0 ^ 1'b0 ;
  assign n1019 = n668 & n1018 ;
  assign n1020 = n815 ^ n316 ^ 1'b0 ;
  assign n1021 = n1019 & ~n1020 ;
  assign n1022 = n319 ^ n275 ^ x86 ;
  assign n1023 = ( x4 & ~n690 ) | ( x4 & n1022 ) | ( ~n690 & n1022 ) ;
  assign n1024 = n601 | n1023 ;
  assign n1025 = n1021 | n1024 ;
  assign n1026 = n614 & ~n933 ;
  assign n1027 = n777 ^ n319 ^ 1'b0 ;
  assign n1028 = n493 ^ n159 ^ 1'b0 ;
  assign n1029 = x83 & ~n1028 ;
  assign n1030 = n653 & n1029 ;
  assign n1031 = ( n328 & ~n543 ) | ( n328 & n638 ) | ( ~n543 & n638 ) ;
  assign n1032 = x20 & x41 ;
  assign n1033 = n1032 ^ x21 ^ 1'b0 ;
  assign n1034 = n1033 ^ n138 ^ 1'b0 ;
  assign n1035 = n508 | n1034 ;
  assign n1036 = n129 | n1035 ;
  assign n1037 = n848 ^ n355 ^ 1'b0 ;
  assign n1038 = n383 | n1037 ;
  assign n1039 = x84 & n1038 ;
  assign n1040 = n248 | n1039 ;
  assign n1041 = n156 & n341 ;
  assign n1042 = n742 ^ n690 ^ n208 ;
  assign n1043 = n1041 & n1042 ;
  assign n1044 = ~n1040 & n1043 ;
  assign n1045 = n612 ^ n303 ^ 1'b0 ;
  assign n1046 = x67 & n541 ;
  assign n1047 = n132 & n1046 ;
  assign n1048 = ~n517 & n1047 ;
  assign n1049 = n1048 ^ n212 ^ 1'b0 ;
  assign n1050 = n1045 & n1049 ;
  assign n1051 = ~n703 & n1042 ;
  assign n1052 = n946 ^ n148 ^ 1'b0 ;
  assign n1053 = n661 & ~n1052 ;
  assign n1054 = ( n731 & n806 ) | ( n731 & ~n974 ) | ( n806 & ~n974 ) ;
  assign n1055 = n813 ^ n562 ^ 1'b0 ;
  assign n1056 = n1055 ^ n156 ^ 1'b0 ;
  assign n1057 = n1056 ^ n694 ^ 1'b0 ;
  assign n1060 = n342 ^ n130 ^ 1'b0 ;
  assign n1061 = x76 & ~n1060 ;
  assign n1058 = n309 & n668 ;
  assign n1059 = ~n417 & n1058 ;
  assign n1062 = n1061 ^ n1059 ^ 1'b0 ;
  assign n1063 = n817 & n1062 ;
  assign n1064 = ~x61 & n1063 ;
  assign n1065 = x66 | n1064 ;
  assign n1066 = x92 & x103 ;
  assign n1067 = ~x93 & n1066 ;
  assign n1068 = x53 & ~n1067 ;
  assign n1069 = n1039 & n1068 ;
  assign n1070 = n595 & ~n1069 ;
  assign n1071 = x69 & ~x110 ;
  assign n1072 = n1071 ^ n1061 ^ 1'b0 ;
  assign n1073 = n1072 ^ n234 ^ 1'b0 ;
  assign n1074 = ~n330 & n1073 ;
  assign n1075 = n396 & ~n933 ;
  assign n1076 = x72 & x119 ;
  assign n1077 = n1076 ^ x120 ^ 1'b0 ;
  assign n1078 = n469 | n1077 ;
  assign n1079 = n461 | n1078 ;
  assign n1080 = n161 & n561 ;
  assign n1081 = n241 ^ x84 ^ x33 ;
  assign n1082 = n1081 ^ n175 ^ x40 ;
  assign n1083 = x97 & ~n1082 ;
  assign n1084 = ( n1079 & n1080 ) | ( n1079 & ~n1083 ) | ( n1080 & ~n1083 ) ;
  assign n1085 = ( n239 & ~n756 ) | ( n239 & n1084 ) | ( ~n756 & n1084 ) ;
  assign n1088 = n595 & ~n620 ;
  assign n1086 = n533 ^ n158 ^ x43 ;
  assign n1087 = n812 | n1086 ;
  assign n1089 = n1088 ^ n1087 ^ 1'b0 ;
  assign n1090 = ( n409 & n447 ) | ( n409 & n479 ) | ( n447 & n479 ) ;
  assign n1091 = n597 & ~n1090 ;
  assign n1092 = n648 & n1091 ;
  assign n1093 = n186 | n353 ;
  assign n1094 = n269 & ~n1093 ;
  assign n1095 = x93 & ~n801 ;
  assign n1096 = n218 ^ x105 ^ 1'b0 ;
  assign n1097 = n328 & n1096 ;
  assign n1098 = x107 & n134 ;
  assign n1099 = ~n1097 & n1098 ;
  assign n1100 = n1095 & n1099 ;
  assign n1101 = n1055 ^ x102 ^ 1'b0 ;
  assign n1102 = n655 ^ n183 ^ 1'b0 ;
  assign n1103 = ~n363 & n1102 ;
  assign n1104 = n297 & ~n433 ;
  assign n1105 = n200 | n639 ;
  assign n1106 = n707 & ~n1105 ;
  assign n1107 = n306 | n353 ;
  assign n1108 = n1106 & ~n1107 ;
  assign n1110 = n499 ^ x40 ^ 1'b0 ;
  assign n1111 = n337 & n1110 ;
  assign n1109 = n590 ^ n461 ^ 1'b0 ;
  assign n1112 = n1111 ^ n1109 ^ 1'b0 ;
  assign n1113 = n1108 | n1112 ;
  assign n1114 = n691 & ~n850 ;
  assign n1115 = ~n1062 & n1114 ;
  assign n1116 = n1115 ^ x68 ^ 1'b0 ;
  assign n1117 = n1116 ^ n1053 ^ n306 ;
  assign n1118 = n635 ^ n229 ^ x40 ;
  assign n1119 = n1118 ^ x114 ^ 1'b0 ;
  assign n1120 = x78 & ~n1119 ;
  assign n1121 = n796 & ~n833 ;
  assign n1122 = ~n1120 & n1121 ;
  assign n1123 = n826 | n1122 ;
  assign n1124 = n651 & ~n1123 ;
  assign n1129 = n1059 ^ n368 ^ 1'b0 ;
  assign n1130 = n497 & n1129 ;
  assign n1125 = ~x74 & n429 ;
  assign n1126 = n1081 ^ n507 ^ 1'b0 ;
  assign n1127 = n969 | n1126 ;
  assign n1128 = n1125 & ~n1127 ;
  assign n1131 = n1130 ^ n1128 ^ 1'b0 ;
  assign n1132 = n1131 ^ n1030 ^ 1'b0 ;
  assign n1133 = n895 | n1132 ;
  assign n1134 = ( n250 & n262 ) | ( n250 & n1133 ) | ( n262 & n1133 ) ;
  assign n1135 = ~n239 & n984 ;
  assign n1136 = n380 ^ x42 ^ 1'b0 ;
  assign n1137 = n1136 ^ n937 ^ 1'b0 ;
  assign n1138 = n1135 | n1137 ;
  assign n1139 = n688 ^ n471 ^ 1'b0 ;
  assign n1140 = ~n793 & n801 ;
  assign n1141 = n243 | n509 ;
  assign n1142 = x104 & n322 ;
  assign n1143 = n1142 ^ n812 ^ 1'b0 ;
  assign n1144 = ~n132 & n1085 ;
  assign n1145 = n1143 & n1144 ;
  assign n1146 = x80 & n1082 ;
  assign n1147 = n1146 ^ n923 ^ 1'b0 ;
  assign n1148 = n417 & ~n610 ;
  assign n1149 = n269 & n1148 ;
  assign n1150 = x127 ^ x108 ^ 1'b0 ;
  assign n1151 = n1150 ^ n912 ^ n877 ;
  assign n1152 = n1151 ^ n994 ^ 1'b0 ;
  assign n1153 = ~n1149 & n1152 ;
  assign n1154 = n141 & n942 ;
  assign n1157 = ~n196 & n606 ;
  assign n1155 = ( n500 & n645 ) | ( n500 & n750 ) | ( n645 & n750 ) ;
  assign n1156 = ( ~n690 & n914 ) | ( ~n690 & n1155 ) | ( n914 & n1155 ) ;
  assign n1158 = n1157 ^ n1156 ^ 1'b0 ;
  assign n1159 = ~n148 & n1158 ;
  assign n1160 = n174 & n803 ;
  assign n1161 = n515 & n996 ;
  assign n1162 = n145 & ~n1161 ;
  assign n1163 = n844 ^ n651 ^ x49 ;
  assign n1164 = n286 & ~n1163 ;
  assign n1165 = n1164 ^ n1072 ^ 1'b0 ;
  assign n1166 = n896 ^ n742 ^ 1'b0 ;
  assign n1167 = n906 ^ n305 ^ 1'b0 ;
  assign n1168 = n1166 & n1167 ;
  assign n1169 = n1042 ^ x25 ^ 1'b0 ;
  assign n1170 = n1169 ^ n1030 ^ 1'b0 ;
  assign n1171 = n823 | n1170 ;
  assign n1172 = n377 & ~n584 ;
  assign n1174 = n1118 ^ n569 ^ 1'b0 ;
  assign n1175 = ~n277 & n1174 ;
  assign n1176 = x101 & n588 ;
  assign n1177 = ~n1175 & n1176 ;
  assign n1173 = n1094 ^ n879 ^ 1'b0 ;
  assign n1178 = n1177 ^ n1173 ^ 1'b0 ;
  assign n1179 = n914 & ~n1178 ;
  assign n1180 = n903 & n1179 ;
  assign n1181 = n1172 & n1180 ;
  assign n1182 = n762 | n859 ;
  assign n1183 = n379 ^ n202 ^ x107 ;
  assign n1184 = n1183 ^ n194 ^ n142 ;
  assign n1185 = n282 & ~n1184 ;
  assign n1186 = ( n183 & ~n607 ) | ( n183 & n1051 ) | ( ~n607 & n1051 ) ;
  assign n1187 = n362 & ~n763 ;
  assign n1188 = n383 & n1187 ;
  assign n1195 = n166 & ~n632 ;
  assign n1190 = n267 | n330 ;
  assign n1191 = n1190 ^ n852 ^ 1'b0 ;
  assign n1189 = n518 ^ n445 ^ x26 ;
  assign n1192 = n1191 ^ n1189 ^ n616 ;
  assign n1193 = ~n702 & n1192 ;
  assign n1194 = n264 & ~n1193 ;
  assign n1196 = n1195 ^ n1194 ^ 1'b0 ;
  assign n1197 = n1009 ^ n335 ^ 1'b0 ;
  assign n1198 = ~n355 & n563 ;
  assign n1199 = n418 | n744 ;
  assign n1200 = n1199 ^ n158 ^ 1'b0 ;
  assign n1201 = n1200 ^ n1046 ^ 1'b0 ;
  assign n1202 = n1198 | n1201 ;
  assign n1203 = n644 ^ n454 ^ 1'b0 ;
  assign n1205 = n391 ^ x70 ^ 1'b0 ;
  assign n1204 = ~n239 & n311 ;
  assign n1206 = n1205 ^ n1204 ^ 1'b0 ;
  assign n1207 = ~n802 & n1206 ;
  assign n1208 = ~n1203 & n1207 ;
  assign n1215 = x9 & ~n683 ;
  assign n1216 = n733 | n1215 ;
  assign n1217 = n1062 | n1216 ;
  assign n1218 = n1115 & n1217 ;
  assign n1209 = n640 ^ n380 ^ n368 ;
  assign n1211 = n730 ^ x36 ^ 1'b0 ;
  assign n1212 = x19 & ~n1211 ;
  assign n1210 = n254 | n932 ;
  assign n1213 = n1212 ^ n1210 ^ 1'b0 ;
  assign n1214 = ~n1209 & n1213 ;
  assign n1219 = n1218 ^ n1214 ^ 1'b0 ;
  assign n1220 = n1012 ^ x83 ^ 1'b0 ;
  assign n1221 = n1220 ^ n892 ^ 1'b0 ;
  assign n1222 = n719 & n1221 ;
  assign n1223 = n153 & ~n876 ;
  assign n1224 = ~n1222 & n1223 ;
  assign n1225 = ~n142 & n602 ;
  assign n1226 = n1225 ^ n241 ^ 1'b0 ;
  assign n1228 = n438 ^ n407 ^ 1'b0 ;
  assign n1227 = n702 & ~n756 ;
  assign n1229 = n1228 ^ n1227 ^ 1'b0 ;
  assign n1230 = ( ~n646 & n758 ) | ( ~n646 & n1229 ) | ( n758 & n1229 ) ;
  assign n1231 = ( n314 & ~n578 ) | ( n314 & n1230 ) | ( ~n578 & n1230 ) ;
  assign n1232 = n273 | n775 ;
  assign n1233 = x46 & n332 ;
  assign n1234 = n1232 & n1233 ;
  assign n1235 = n456 & ~n969 ;
  assign n1236 = n908 & n935 ;
  assign n1237 = ~n293 & n1184 ;
  assign n1238 = n720 ^ n496 ^ 1'b0 ;
  assign n1239 = ( n466 & n1237 ) | ( n466 & n1238 ) | ( n1237 & n1238 ) ;
  assign n1240 = ~n376 & n1239 ;
  assign n1242 = ~n380 & n1125 ;
  assign n1241 = n279 & ~n953 ;
  assign n1243 = n1242 ^ n1241 ^ 1'b0 ;
  assign n1244 = ~n236 & n488 ;
  assign n1245 = ( n275 & n1243 ) | ( n275 & ~n1244 ) | ( n1243 & ~n1244 ) ;
  assign n1246 = n519 ^ n463 ^ n290 ;
  assign n1247 = x67 & ~n179 ;
  assign n1248 = n1247 ^ n760 ^ 1'b0 ;
  assign n1249 = n1248 ^ n586 ^ 1'b0 ;
  assign n1250 = x98 & n1249 ;
  assign n1251 = n1250 ^ n340 ^ 1'b0 ;
  assign n1252 = n1067 ^ n990 ^ 1'b0 ;
  assign n1253 = ~n696 & n1252 ;
  assign n1254 = n672 ^ x44 ^ 1'b0 ;
  assign n1255 = n643 & ~n665 ;
  assign n1256 = ~n1254 & n1255 ;
  assign n1257 = ~n548 & n549 ;
  assign n1258 = ~n962 & n1257 ;
  assign n1259 = n345 & n955 ;
  assign n1260 = ~n1231 & n1259 ;
  assign n1261 = n883 ^ x86 ^ 1'b0 ;
  assign n1262 = n1261 ^ n937 ^ 1'b0 ;
  assign n1263 = ~n1232 & n1262 ;
  assign n1264 = n420 & n895 ;
  assign n1265 = ( n510 & n1179 ) | ( n510 & ~n1264 ) | ( n1179 & ~n1264 ) ;
  assign n1268 = x100 ^ x70 ^ 1'b0 ;
  assign n1266 = n563 ^ x32 ^ 1'b0 ;
  assign n1267 = n713 & n1266 ;
  assign n1269 = n1268 ^ n1267 ^ x64 ;
  assign n1270 = n1269 ^ n678 ^ 1'b0 ;
  assign n1271 = n1228 & ~n1270 ;
  assign n1272 = n422 ^ x123 ^ 1'b0 ;
  assign n1273 = n1272 ^ n510 ^ 1'b0 ;
  assign n1274 = n616 ^ n401 ^ 1'b0 ;
  assign n1275 = n371 & ~n1274 ;
  assign n1276 = n857 & ~n1275 ;
  assign n1277 = x99 & ~n379 ;
  assign n1278 = ( x55 & ~n950 ) | ( x55 & n1277 ) | ( ~n950 & n1277 ) ;
  assign n1279 = n422 ^ n341 ^ 1'b0 ;
  assign n1280 = n599 ^ n243 ^ 1'b0 ;
  assign n1281 = ~n533 & n1280 ;
  assign n1282 = n486 | n1013 ;
  assign n1283 = n1282 ^ n561 ^ 1'b0 ;
  assign n1289 = n812 & n1062 ;
  assign n1290 = n1289 ^ n823 ^ 1'b0 ;
  assign n1291 = n1290 ^ n593 ^ 1'b0 ;
  assign n1292 = x81 & ~n1291 ;
  assign n1284 = n610 | n796 ;
  assign n1285 = n452 & n1284 ;
  assign n1286 = n1285 ^ n252 ^ 1'b0 ;
  assign n1287 = n1286 ^ x71 ^ 1'b0 ;
  assign n1288 = n769 | n1287 ;
  assign n1293 = n1292 ^ n1288 ^ n1034 ;
  assign n1296 = x12 & n143 ;
  assign n1297 = ~n764 & n1296 ;
  assign n1294 = n764 ^ n592 ^ 1'b0 ;
  assign n1295 = n543 & n1294 ;
  assign n1298 = n1297 ^ n1295 ^ 1'b0 ;
  assign n1299 = n927 & ~n1298 ;
  assign n1300 = n1299 ^ n1254 ^ n564 ;
  assign n1301 = n953 ^ n524 ^ 1'b0 ;
  assign n1302 = n174 | n1301 ;
  assign n1303 = n418 & ~n872 ;
  assign n1304 = n1303 ^ n578 ^ 1'b0 ;
  assign n1305 = n757 & n1304 ;
  assign n1306 = n290 | n1305 ;
  assign n1307 = n488 ^ x58 ^ x28 ;
  assign n1308 = ( x67 & n265 ) | ( x67 & n1307 ) | ( n265 & n1307 ) ;
  assign n1309 = n1303 | n1308 ;
  assign n1310 = n1309 ^ n688 ^ 1'b0 ;
  assign n1311 = ~n1306 & n1310 ;
  assign n1312 = n954 ^ n467 ^ n257 ;
  assign n1313 = n1312 ^ n832 ^ 1'b0 ;
  assign n1317 = n510 & n857 ;
  assign n1318 = n167 & n1317 ;
  assign n1314 = x29 & n326 ;
  assign n1315 = n254 | n1133 ;
  assign n1316 = n1314 | n1315 ;
  assign n1319 = n1318 ^ n1316 ^ n478 ;
  assign n1320 = n838 ^ n132 ^ 1'b0 ;
  assign n1321 = x41 & ~n1065 ;
  assign n1322 = ~n1156 & n1195 ;
  assign n1323 = n1322 ^ n248 ^ 1'b0 ;
  assign n1324 = x14 & ~n307 ;
  assign n1325 = n1324 ^ n683 ^ 1'b0 ;
  assign n1326 = ~n578 & n1325 ;
  assign n1327 = n1326 ^ n532 ^ 1'b0 ;
  assign n1328 = ~n413 & n1168 ;
  assign n1329 = ~n1327 & n1328 ;
  assign n1330 = n1097 ^ n454 ^ n231 ;
  assign n1331 = n229 | n576 ;
  assign n1332 = n1033 & ~n1331 ;
  assign n1333 = ( n235 & ~n317 ) | ( n235 & n1332 ) | ( ~n317 & n1332 ) ;
  assign n1334 = n922 | n1055 ;
  assign n1335 = n1334 ^ n1082 ^ 1'b0 ;
  assign n1336 = ~n978 & n1335 ;
  assign n1337 = ~n1333 & n1336 ;
  assign n1338 = n576 | n1326 ;
  assign n1339 = n1209 ^ n129 ^ 1'b0 ;
  assign n1341 = n680 ^ n411 ^ 1'b0 ;
  assign n1340 = x19 & ~n1027 ;
  assign n1342 = n1341 ^ n1340 ^ 1'b0 ;
  assign n1343 = ~n310 & n652 ;
  assign n1344 = n733 ^ n717 ^ 1'b0 ;
  assign n1345 = ~n1343 & n1344 ;
  assign n1346 = ~n661 & n1345 ;
  assign n1347 = ~n544 & n1346 ;
  assign n1348 = n1347 ^ n1320 ^ 1'b0 ;
  assign n1349 = n1234 ^ n691 ^ 1'b0 ;
  assign n1350 = n960 | n1349 ;
  assign n1351 = n220 | n917 ;
  assign n1352 = n1351 ^ n134 ^ 1'b0 ;
  assign n1353 = ~n331 & n588 ;
  assign n1354 = n1353 ^ n369 ^ 1'b0 ;
  assign n1355 = n161 & ~n265 ;
  assign n1356 = n1355 ^ x45 ^ 1'b0 ;
  assign n1357 = n1140 ^ n438 ^ 1'b0 ;
  assign n1358 = n314 & ~n1357 ;
  assign n1359 = ~n808 & n1358 ;
  assign n1360 = n1356 & n1359 ;
  assign n1362 = n1122 ^ n668 ^ 1'b0 ;
  assign n1363 = n1362 ^ n399 ^ 1'b0 ;
  assign n1364 = ~n326 & n1363 ;
  assign n1361 = ~n338 & n888 ;
  assign n1365 = n1364 ^ n1361 ^ 1'b0 ;
  assign n1366 = n872 ^ x82 ^ 1'b0 ;
  assign n1367 = x110 & ~n1366 ;
  assign n1368 = ~n947 & n1367 ;
  assign n1369 = n1205 ^ n191 ^ 1'b0 ;
  assign n1370 = n707 | n1369 ;
  assign n1372 = n1041 ^ n557 ^ 1'b0 ;
  assign n1373 = n470 & ~n505 ;
  assign n1374 = ( ~n509 & n1372 ) | ( ~n509 & n1373 ) | ( n1372 & n1373 ) ;
  assign n1371 = x107 ^ x35 ^ 1'b0 ;
  assign n1375 = n1374 ^ n1371 ^ 1'b0 ;
  assign n1376 = n1293 ^ n588 ^ n325 ;
  assign n1377 = x8 & n454 ;
  assign n1378 = ~x17 & n1377 ;
  assign n1379 = n753 | n1378 ;
  assign n1380 = n565 ^ n353 ^ x64 ;
  assign n1381 = ~n361 & n1380 ;
  assign n1382 = n1379 & n1381 ;
  assign n1383 = n564 ^ n158 ^ 1'b0 ;
  assign n1384 = n331 | n1383 ;
  assign n1385 = n1117 ^ n606 ^ 1'b0 ;
  assign n1386 = n1385 ^ n738 ^ 1'b0 ;
  assign n1387 = ~n1384 & n1386 ;
  assign n1388 = ~n927 & n1192 ;
  assign n1389 = n773 ^ n482 ^ 1'b0 ;
  assign n1390 = ~n1362 & n1389 ;
  assign n1391 = n897 & n1390 ;
  assign n1392 = n1391 ^ n1085 ^ 1'b0 ;
  assign n1393 = n467 | n935 ;
  assign n1394 = n1000 & n1393 ;
  assign n1395 = ~n393 & n897 ;
  assign n1396 = n891 & n1395 ;
  assign n1397 = n1396 ^ n380 ^ 1'b0 ;
  assign n1398 = n492 & n1248 ;
  assign n1399 = ~x41 & n1398 ;
  assign n1400 = n1399 ^ n447 ^ 1'b0 ;
  assign n1401 = n876 | n1400 ;
  assign n1402 = x20 & n586 ;
  assign n1403 = ~x119 & n1402 ;
  assign n1404 = n1039 ^ n262 ^ 1'b0 ;
  assign n1405 = n1300 | n1404 ;
  assign n1406 = n1286 ^ n1220 ^ 1'b0 ;
  assign n1410 = ~n461 & n1009 ;
  assign n1407 = ( x46 & n594 ) | ( x46 & ~n818 ) | ( n594 & ~n818 ) ;
  assign n1408 = n628 | n1407 ;
  assign n1409 = n1343 & ~n1408 ;
  assign n1411 = n1410 ^ n1409 ^ 1'b0 ;
  assign n1412 = n770 ^ n637 ^ 1'b0 ;
  assign n1413 = ~x10 & x30 ;
  assign n1414 = ( n969 & ~n1412 ) | ( n969 & n1413 ) | ( ~n1412 & n1413 ) ;
  assign n1415 = n1155 | n1414 ;
  assign n1416 = ( x16 & ~x101 ) | ( x16 & n474 ) | ( ~x101 & n474 ) ;
  assign n1417 = n389 & n1416 ;
  assign n1418 = ~n875 & n1417 ;
  assign n1419 = ~n267 & n470 ;
  assign n1420 = ~n659 & n1419 ;
  assign n1421 = ~n206 & n1420 ;
  assign n1422 = n1421 ^ n1045 ^ 1'b0 ;
  assign n1423 = n1033 ^ n223 ^ 1'b0 ;
  assign n1424 = n914 ^ n764 ^ 1'b0 ;
  assign n1425 = n352 ^ n310 ^ 1'b0 ;
  assign n1426 = n707 ^ n355 ^ 1'b0 ;
  assign n1427 = n1079 & n1426 ;
  assign n1428 = x53 & n1427 ;
  assign n1429 = ~n169 & n1279 ;
  assign n1430 = ~n1330 & n1429 ;
  assign n1431 = n848 & n1147 ;
  assign n1432 = n1431 ^ n355 ^ 1'b0 ;
  assign n1433 = n1432 ^ n1111 ^ n543 ;
  assign n1434 = n605 ^ x76 ^ 1'b0 ;
  assign n1435 = ( n359 & n421 ) | ( n359 & ~n616 ) | ( n421 & ~n616 ) ;
  assign n1436 = n1435 ^ n1308 ^ 1'b0 ;
  assign n1437 = ~n1172 & n1436 ;
  assign n1438 = ~n713 & n1437 ;
  assign n1439 = n1149 ^ n466 ^ 1'b0 ;
  assign n1440 = n215 ^ n179 ^ 1'b0 ;
  assign n1441 = n135 & n322 ;
  assign n1442 = n1441 ^ n348 ^ 1'b0 ;
  assign n1443 = x92 & n1442 ;
  assign n1444 = n1443 ^ n1324 ^ 1'b0 ;
  assign n1445 = ~n1440 & n1444 ;
  assign n1446 = n1445 ^ n185 ^ 1'b0 ;
  assign n1447 = x73 & ~n342 ;
  assign n1448 = ~n557 & n1447 ;
  assign n1449 = n1448 ^ x25 ^ x14 ;
  assign n1450 = n1449 ^ n627 ^ 1'b0 ;
  assign n1451 = n1450 ^ n1299 ^ 1'b0 ;
  assign n1452 = n265 & ~n319 ;
  assign n1453 = n1120 ^ n538 ^ 1'b0 ;
  assign n1454 = ~n338 & n1453 ;
  assign n1455 = n917 ^ n295 ^ 1'b0 ;
  assign n1456 = n1454 & n1455 ;
  assign n1457 = n1452 & n1456 ;
  assign n1458 = x43 ^ x22 ^ 1'b0 ;
  assign n1459 = n949 & n1203 ;
  assign n1460 = n1458 & ~n1459 ;
  assign n1461 = n1457 & n1460 ;
  assign n1462 = n798 & ~n975 ;
  assign n1463 = n1462 ^ n199 ^ 1'b0 ;
  assign n1469 = x126 & ~n167 ;
  assign n1470 = ~n493 & n1469 ;
  assign n1464 = x113 & n469 ;
  assign n1465 = n1464 ^ n445 ^ 1'b0 ;
  assign n1466 = ~n231 & n643 ;
  assign n1467 = n1466 ^ n254 ^ 1'b0 ;
  assign n1468 = n1465 & n1467 ;
  assign n1471 = n1470 ^ n1468 ^ 1'b0 ;
  assign n1472 = x68 | n301 ;
  assign n1473 = n652 | n1013 ;
  assign n1474 = x101 & ~n1473 ;
  assign n1475 = n1474 ^ n150 ^ 1'b0 ;
  assign n1476 = n659 | n922 ;
  assign n1477 = n667 & n910 ;
  assign n1478 = n283 & ~n547 ;
  assign n1479 = n1478 ^ x109 ^ 1'b0 ;
  assign n1480 = n1479 ^ n961 ^ x74 ;
  assign n1481 = n1480 ^ n301 ^ 1'b0 ;
  assign n1482 = n225 ^ x68 ^ 1'b0 ;
  assign n1483 = n891 ^ x13 ^ 1'b0 ;
  assign n1484 = ~n1482 & n1483 ;
  assign n1485 = x6 & n884 ;
  assign n1486 = ( n535 & n922 ) | ( n535 & n1485 ) | ( n922 & n1485 ) ;
  assign n1489 = n1236 & n1480 ;
  assign n1487 = n933 ^ n728 ^ n177 ;
  assign n1488 = n1038 | n1487 ;
  assign n1490 = n1489 ^ n1488 ^ 1'b0 ;
  assign n1496 = n1479 ^ n1175 ^ 1'b0 ;
  assign n1497 = ~n212 & n1496 ;
  assign n1498 = n1497 ^ x9 ^ 1'b0 ;
  assign n1499 = n1498 ^ n569 ^ 1'b0 ;
  assign n1491 = n1002 ^ x95 ^ 1'b0 ;
  assign n1492 = n204 | n1491 ;
  assign n1493 = x64 & n214 ;
  assign n1494 = n1061 | n1493 ;
  assign n1495 = n1492 | n1494 ;
  assign n1500 = n1499 ^ n1495 ^ 1'b0 ;
  assign n1501 = ~n197 & n299 ;
  assign n1502 = n1033 | n1376 ;
  assign n1503 = n1025 | n1502 ;
  assign n1504 = n258 ^ x41 ^ 1'b0 ;
  assign n1505 = n1465 ^ n840 ^ 1'b0 ;
  assign n1506 = ( n252 & n562 ) | ( n252 & ~n1371 ) | ( n562 & ~n1371 ) ;
  assign n1507 = n1505 | n1506 ;
  assign n1511 = ~x33 & n141 ;
  assign n1512 = n1511 ^ x12 ^ 1'b0 ;
  assign n1508 = n461 & ~n606 ;
  assign n1509 = n1508 ^ n1222 ^ 1'b0 ;
  assign n1510 = n311 & ~n1509 ;
  assign n1513 = n1512 ^ n1510 ^ 1'b0 ;
  assign n1514 = n871 ^ n673 ^ 1'b0 ;
  assign n1515 = n480 | n1514 ;
  assign n1516 = n1515 ^ n1307 ^ 1'b0 ;
  assign n1517 = ~n254 & n753 ;
  assign n1518 = n1276 & ~n1517 ;
  assign n1519 = ~n690 & n1518 ;
  assign n1521 = n338 ^ x96 ^ 1'b0 ;
  assign n1520 = ( ~n161 & n681 ) | ( ~n161 & n1021 ) | ( n681 & n1021 ) ;
  assign n1522 = n1521 ^ n1520 ^ n728 ;
  assign n1524 = n929 ^ n577 ^ 1'b0 ;
  assign n1525 = x23 & n1524 ;
  assign n1523 = n603 & ~n1230 ;
  assign n1526 = n1525 ^ n1523 ^ 1'b0 ;
  assign n1527 = x57 | n301 ;
  assign n1528 = n1217 ^ n877 ^ n799 ;
  assign n1529 = ~n812 & n939 ;
  assign n1530 = n1407 | n1529 ;
  assign n1531 = x50 & n1530 ;
  assign n1532 = n1531 ^ x23 ^ 1'b0 ;
  assign n1533 = x92 & ~n996 ;
  assign n1534 = ~n1162 & n1533 ;
  assign n1535 = n1165 ^ n1012 ^ 1'b0 ;
  assign n1536 = n1083 ^ n422 ^ 1'b0 ;
  assign n1537 = ~n277 & n1536 ;
  assign n1538 = x78 & ~n1065 ;
  assign n1539 = ~n746 & n1538 ;
  assign n1540 = n1539 ^ n252 ^ 1'b0 ;
  assign n1541 = x3 & ~n1384 ;
  assign n1542 = n1541 ^ n130 ^ 1'b0 ;
  assign n1543 = n1542 ^ n690 ^ n535 ;
  assign n1544 = n202 | n1543 ;
  assign n1545 = n920 | n1544 ;
  assign n1546 = n1353 & n1545 ;
  assign n1547 = n229 & n1546 ;
  assign n1548 = n690 ^ n645 ^ 1'b0 ;
  assign n1549 = x117 & ~n1548 ;
  assign n1550 = n494 & ~n1272 ;
  assign n1551 = n1549 & n1550 ;
  assign n1552 = n1551 ^ n1506 ^ 1'b0 ;
  assign n1554 = ~n479 & n652 ;
  assign n1553 = n1086 ^ n560 ^ n243 ;
  assign n1555 = n1554 ^ n1553 ^ 1'b0 ;
  assign n1556 = x111 ^ x29 ^ 1'b0 ;
  assign n1557 = x14 & n1556 ;
  assign n1558 = n1557 ^ n954 ^ 1'b0 ;
  assign n1559 = ~n979 & n1558 ;
  assign n1560 = n748 & n767 ;
  assign n1561 = ( ~x41 & n1559 ) | ( ~x41 & n1560 ) | ( n1559 & n1560 ) ;
  assign n1562 = n644 | n670 ;
  assign n1563 = n343 & ~n812 ;
  assign n1564 = n1563 ^ n330 ^ 1'b0 ;
  assign n1565 = n1564 ^ n794 ^ 1'b0 ;
  assign n1566 = n891 ^ n225 ^ n200 ;
  assign n1567 = n718 | n1566 ;
  assign n1568 = n1567 ^ n388 ^ x56 ;
  assign n1569 = ~n640 & n1568 ;
  assign n1570 = ~n417 & n1569 ;
  assign n1571 = ( ~n290 & n616 ) | ( ~n290 & n690 ) | ( n616 & n690 ) ;
  assign n1572 = ( n899 & n901 ) | ( n899 & ~n1571 ) | ( n901 & ~n1571 ) ;
  assign n1573 = n1572 ^ n1288 ^ 1'b0 ;
  assign n1574 = n496 ^ n273 ^ 1'b0 ;
  assign n1575 = ~n1573 & n1574 ;
  assign n1576 = n938 ^ n627 ^ n571 ;
  assign n1577 = n466 ^ n254 ^ 1'b0 ;
  assign n1578 = n659 & n1577 ;
  assign n1579 = n459 ^ n449 ^ 1'b0 ;
  assign n1580 = ~n969 & n1579 ;
  assign n1581 = ( n1576 & n1578 ) | ( n1576 & n1580 ) | ( n1578 & n1580 ) ;
  assign n1582 = n1581 ^ n928 ^ 1'b0 ;
  assign n1583 = n793 ^ x34 ^ 1'b0 ;
  assign n1584 = ( x51 & ~n535 ) | ( x51 & n1583 ) | ( ~n535 & n1583 ) ;
  assign n1585 = ~n563 & n1584 ;
  assign n1586 = n1462 & n1585 ;
  assign n1587 = n845 ^ n477 ^ n159 ;
  assign n1588 = n788 & ~n1587 ;
  assign n1589 = ( n618 & n652 ) | ( n618 & ~n928 ) | ( n652 & ~n928 ) ;
  assign n1590 = n1154 & n1589 ;
  assign n1591 = x109 ^ x7 ^ 1'b0 ;
  assign n1592 = ~n320 & n333 ;
  assign n1593 = n1592 ^ n269 ^ 1'b0 ;
  assign n1594 = n332 & n1593 ;
  assign n1595 = n1594 ^ n664 ^ 1'b0 ;
  assign n1596 = n141 & ~n1595 ;
  assign n1597 = ( ~n1041 & n1591 ) | ( ~n1041 & n1596 ) | ( n1591 & n1596 ) ;
  assign n1598 = ~n275 & n461 ;
  assign n1599 = n456 & n1598 ;
  assign n1600 = n1599 ^ n754 ^ n200 ;
  assign n1601 = n1600 ^ n980 ^ 1'b0 ;
  assign n1605 = n239 & n417 ;
  assign n1606 = n1553 | n1605 ;
  assign n1607 = n1606 ^ n433 ^ 1'b0 ;
  assign n1608 = x116 & ~n1607 ;
  assign n1602 = n231 & ~n895 ;
  assign n1603 = n563 & n1602 ;
  assign n1604 = n707 | n1603 ;
  assign n1609 = n1608 ^ n1604 ^ 1'b0 ;
  assign n1610 = n1594 ^ n461 ^ 1'b0 ;
  assign n1611 = ( n191 & ~n619 ) | ( n191 & n959 ) | ( ~n619 & n959 ) ;
  assign n1612 = ~n670 & n952 ;
  assign n1613 = n1611 & n1612 ;
  assign n1614 = n480 | n907 ;
  assign n1615 = x25 | n584 ;
  assign n1616 = x52 & n1615 ;
  assign n1617 = n293 & n1616 ;
  assign n1618 = x61 & ~n849 ;
  assign n1619 = ~n507 & n1618 ;
  assign n1620 = n1356 | n1619 ;
  assign n1621 = n1620 ^ n1463 ^ 1'b0 ;
  assign n1622 = n1621 ^ n1059 ^ 1'b0 ;
  assign n1623 = n955 & ~n1622 ;
  assign n1624 = n338 ^ n328 ^ n134 ;
  assign n1625 = n1624 ^ x51 ^ 1'b0 ;
  assign n1626 = x121 & n1625 ;
  assign n1627 = ( n405 & n518 ) | ( n405 & n1571 ) | ( n518 & n1571 ) ;
  assign n1628 = ( ~n620 & n1626 ) | ( ~n620 & n1627 ) | ( n1626 & n1627 ) ;
  assign n1629 = n1507 ^ n1041 ^ 1'b0 ;
  assign n1630 = n1127 & ~n1629 ;
  assign n1631 = n1030 ^ x86 ^ 1'b0 ;
  assign n1632 = n1090 ^ x13 ^ 1'b0 ;
  assign n1633 = n324 & ~n1600 ;
  assign n1634 = n310 | n1633 ;
  assign n1635 = ~n548 & n930 ;
  assign n1636 = n923 & n1635 ;
  assign n1637 = n1636 ^ n1321 ^ 1'b0 ;
  assign n1638 = n1193 ^ n788 ^ x55 ;
  assign n1639 = n1637 & n1638 ;
  assign n1640 = ~n355 & n1019 ;
  assign n1641 = n1640 ^ n707 ^ 1'b0 ;
  assign n1642 = n516 & n1641 ;
  assign n1643 = n1642 ^ n254 ^ 1'b0 ;
  assign n1644 = n1151 & n1643 ;
  assign n1645 = n389 & ~n1571 ;
  assign n1646 = n1645 ^ n277 ^ 1'b0 ;
  assign n1647 = n176 & ~n1022 ;
  assign n1648 = n1647 ^ x90 ^ 1'b0 ;
  assign n1649 = ~x100 & n827 ;
  assign n1650 = ( n286 & n1648 ) | ( n286 & ~n1649 ) | ( n1648 & ~n1649 ) ;
  assign n1651 = n945 | n1124 ;
  assign n1652 = n1021 | n1651 ;
  assign n1653 = n914 & n1237 ;
  assign n1654 = n581 & n1653 ;
  assign n1655 = n216 & n1059 ;
  assign n1656 = ( n293 & ~n1149 ) | ( n293 & n1554 ) | ( ~n1149 & n1554 ) ;
  assign n1657 = n794 ^ x91 ^ 1'b0 ;
  assign n1658 = n1480 | n1657 ;
  assign n1659 = x43 & ~n487 ;
  assign n1660 = n1658 & n1659 ;
  assign n1661 = ( x117 & ~n683 ) | ( x117 & n786 ) | ( ~n683 & n786 ) ;
  assign n1662 = n593 & ~n701 ;
  assign n1663 = ~n703 & n1662 ;
  assign n1664 = n513 & ~n952 ;
  assign n1665 = n1664 ^ n1200 ^ 1'b0 ;
  assign n1666 = ~n1663 & n1665 ;
  assign n1667 = n570 & ~n1564 ;
  assign n1668 = n1217 ^ n1215 ^ n706 ;
  assign n1669 = n788 & n1668 ;
  assign n1670 = n1669 ^ n1562 ^ 1'b0 ;
  assign n1671 = ( n350 & n1371 ) | ( n350 & ~n1379 ) | ( n1371 & ~n1379 ) ;
  assign n1672 = n777 & n1671 ;
  assign n1673 = n1672 ^ x70 ^ 1'b0 ;
  assign n1674 = n686 ^ x64 ^ 1'b0 ;
  assign n1675 = ( n350 & ~n756 ) | ( n350 & n1674 ) | ( ~n756 & n1674 ) ;
  assign n1676 = ~n498 & n1675 ;
  assign n1677 = n1676 ^ n312 ^ 1'b0 ;
  assign n1678 = n425 | n1677 ;
  assign n1679 = n424 | n1678 ;
  assign n1680 = n445 & ~n494 ;
  assign n1681 = n379 ^ n179 ^ 1'b0 ;
  assign n1682 = ( n1034 & ~n1680 ) | ( n1034 & n1681 ) | ( ~n1680 & n1681 ) ;
  assign n1683 = ~x97 & n1435 ;
  assign n1684 = ( n906 & n1649 ) | ( n906 & n1683 ) | ( n1649 & n1683 ) ;
  assign n1686 = n526 ^ x77 ^ 1'b0 ;
  assign n1685 = n190 & n802 ;
  assign n1687 = n1686 ^ n1685 ^ 1'b0 ;
  assign n1688 = n1414 ^ n734 ^ 1'b0 ;
  assign n1689 = n1688 ^ x100 ^ 1'b0 ;
  assign n1690 = n886 & ~n1248 ;
  assign n1691 = n1689 & ~n1690 ;
  assign n1692 = ~n1284 & n1691 ;
  assign n1693 = n1220 & n1576 ;
  assign n1694 = ( n319 & ~n790 ) | ( n319 & n1693 ) | ( ~n790 & n1693 ) ;
  assign n1695 = n1694 ^ n541 ^ n499 ;
  assign n1696 = n322 ^ x85 ^ 1'b0 ;
  assign n1697 = ~n872 & n1696 ;
  assign n1698 = n1697 ^ n243 ^ 1'b0 ;
  assign n1699 = ~n473 & n819 ;
  assign n1700 = n355 & n1699 ;
  assign n1701 = n1698 & ~n1700 ;
  assign n1702 = n1701 ^ x62 ^ 1'b0 ;
  assign n1703 = ~n320 & n1525 ;
  assign n1704 = ~n1702 & n1703 ;
  assign n1705 = ~n750 & n1704 ;
  assign n1706 = n1184 ^ n646 ^ n632 ;
  assign n1707 = n1423 ^ x13 ^ 1'b0 ;
  assign n1708 = n1706 & n1707 ;
  assign n1709 = n1629 ^ n130 ^ 1'b0 ;
  assign n1710 = n416 & ~n1709 ;
  assign n1711 = ( ~n671 & n720 ) | ( ~n671 & n1251 ) | ( n720 & n1251 ) ;
  assign n1712 = x82 & n1711 ;
  assign n1713 = n1712 ^ n770 ^ 1'b0 ;
  assign n1714 = ( n959 & n1371 ) | ( n959 & n1422 ) | ( n1371 & n1422 ) ;
  assign n1715 = x47 & ~n696 ;
  assign n1716 = n1715 ^ n1572 ^ 1'b0 ;
  assign n1717 = n398 & n746 ;
  assign n1718 = ~n726 & n1717 ;
  assign n1719 = n753 ^ n371 ^ 1'b0 ;
  assign n1720 = n362 & ~n1719 ;
  assign n1721 = n220 & n1720 ;
  assign n1722 = n1297 ^ n145 ^ x66 ;
  assign n1723 = n664 ^ n576 ^ 1'b0 ;
  assign n1724 = n381 & ~n1723 ;
  assign n1725 = n1724 ^ n603 ^ 1'b0 ;
  assign n1726 = n1250 & n1725 ;
  assign n1727 = x94 & ~n1169 ;
  assign n1728 = ~n386 & n1727 ;
  assign n1729 = n1451 ^ n1160 ^ 1'b0 ;
  assign n1730 = ~n1728 & n1729 ;
  assign n1731 = n1730 ^ n1554 ^ 1'b0 ;
  assign n1732 = n614 & ~n1731 ;
  assign n1733 = n1263 ^ n248 ^ 1'b0 ;
  assign n1734 = ~n1108 & n1733 ;
  assign n1735 = n1686 ^ n1684 ^ 1'b0 ;
  assign n1736 = n332 & ~n1735 ;
  assign n1737 = x35 & n796 ;
  assign n1738 = n1737 ^ n346 ^ 1'b0 ;
  assign n1739 = n852 | n1738 ;
  assign n1740 = ~x12 & n655 ;
  assign n1741 = ~n1182 & n1740 ;
  assign n1742 = n497 ^ x11 ^ 1'b0 ;
  assign n1743 = ~n388 & n1134 ;
  assign n1744 = n1743 ^ n171 ^ 1'b0 ;
  assign n1745 = n1742 & ~n1744 ;
  assign n1746 = ( n401 & ~n482 ) | ( n401 & n592 ) | ( ~n482 & n592 ) ;
  assign n1747 = ( x40 & ~n678 ) | ( x40 & n1746 ) | ( ~n678 & n1746 ) ;
  assign n1748 = n1516 ^ n661 ^ 1'b0 ;
  assign n1749 = ~n896 & n1748 ;
  assign n1750 = n1458 & n1686 ;
  assign n1751 = ~n1217 & n1750 ;
  assign n1752 = n1751 ^ n654 ^ 1'b0 ;
  assign n1753 = ~n1242 & n1384 ;
  assign n1756 = n408 & n463 ;
  assign n1757 = ~n421 & n1756 ;
  assign n1754 = ( n742 & ~n1600 ) | ( n742 & n1740 ) | ( ~n1600 & n1740 ) ;
  assign n1755 = n819 & n1754 ;
  assign n1758 = n1757 ^ n1755 ^ 1'b0 ;
  assign n1759 = n1758 ^ n612 ^ 1'b0 ;
  assign n1760 = n210 & n1759 ;
  assign n1761 = n1290 ^ n467 ^ 1'b0 ;
  assign n1762 = n1761 ^ n1711 ^ 1'b0 ;
  assign n1765 = n499 ^ n425 ^ x29 ;
  assign n1763 = n796 & ~n837 ;
  assign n1764 = n707 & n1763 ;
  assign n1766 = n1765 ^ n1764 ^ n1083 ;
  assign n1767 = n1766 ^ n781 ^ n612 ;
  assign n1768 = n1767 ^ n1470 ^ n427 ;
  assign n1769 = n1768 ^ n708 ^ n456 ;
  assign n1770 = x3 & n1422 ;
  assign n1771 = n1770 ^ n330 ^ 1'b0 ;
  assign n1772 = n606 & n1771 ;
  assign n1773 = n1040 & ~n1479 ;
  assign n1774 = n1773 ^ n722 ^ 1'b0 ;
  assign n1775 = x103 ^ x86 ^ 1'b0 ;
  assign n1776 = n1775 ^ n1300 ^ x122 ;
  assign n1777 = n930 & ~n1019 ;
  assign n1778 = x7 & n992 ;
  assign n1779 = n1778 ^ n290 ^ 1'b0 ;
  assign n1780 = n1324 & ~n1779 ;
  assign n1781 = ( ~x15 & n477 ) | ( ~x15 & n1780 ) | ( n477 & n1780 ) ;
  assign n1782 = n581 ^ n532 ^ n150 ;
  assign n1783 = ~n405 & n615 ;
  assign n1784 = ~n362 & n1783 ;
  assign n1785 = n1782 | n1784 ;
  assign n1786 = n393 ^ n129 ^ 1'b0 ;
  assign n1787 = x123 & ~n1645 ;
  assign n1788 = n1787 ^ n1687 ^ 1'b0 ;
  assign n1789 = n720 ^ n717 ^ n241 ;
  assign n1790 = n770 & n1789 ;
  assign n1791 = n1790 ^ n1482 ^ 1'b0 ;
  assign n1792 = n717 ^ n279 ^ x70 ;
  assign n1793 = n1792 ^ n1455 ^ 1'b0 ;
  assign n1794 = n844 & n1793 ;
  assign n1795 = n1794 ^ n194 ^ x19 ;
  assign n1796 = ~n466 & n1795 ;
  assign n1797 = n616 | n1796 ;
  assign n1798 = n1797 ^ n730 ^ 1'b0 ;
  assign n1799 = n886 ^ n627 ^ 1'b0 ;
  assign n1800 = n206 | n801 ;
  assign n1805 = n961 ^ x13 ^ 1'b0 ;
  assign n1801 = n487 ^ n380 ^ 1'b0 ;
  assign n1802 = ~n896 & n1801 ;
  assign n1803 = x76 & ~n1802 ;
  assign n1804 = n1326 & n1803 ;
  assign n1806 = n1805 ^ n1804 ^ 1'b0 ;
  assign n1807 = n1800 & n1806 ;
  assign n1808 = ~n1388 & n1807 ;
  assign n1809 = x118 | n872 ;
  assign n1810 = ( n974 & n1674 ) | ( n974 & n1809 ) | ( n1674 & n1809 ) ;
  assign n1811 = n1810 ^ x27 ^ 1'b0 ;
  assign n1812 = ~n381 & n1706 ;
  assign n1813 = n1812 ^ n1371 ^ 1'b0 ;
  assign n1814 = n1379 ^ n1273 ^ 1'b0 ;
  assign n1815 = n757 & n1814 ;
  assign n1816 = x51 & n1815 ;
  assign n1817 = ~n1670 & n1816 ;
  assign n1818 = n696 | n1172 ;
  assign n1819 = n1362 ^ n707 ^ 1'b0 ;
  assign n1820 = ( n1054 & ~n1532 ) | ( n1054 & n1819 ) | ( ~n1532 & n1819 ) ;
  assign n1821 = n1820 ^ n439 ^ 1'b0 ;
  assign n1822 = n197 & n886 ;
  assign n1823 = n1457 & n1822 ;
  assign n1824 = n943 ^ n837 ^ 1'b0 ;
  assign n1825 = n1824 ^ n854 ^ 1'b0 ;
  assign n1826 = n1442 & ~n1825 ;
  assign n1827 = ~n175 & n335 ;
  assign n1828 = n1827 ^ n1010 ^ 1'b0 ;
  assign n1829 = n785 ^ n740 ^ 1'b0 ;
  assign n1831 = n206 | n733 ;
  assign n1832 = n1831 ^ n1686 ^ 1'b0 ;
  assign n1830 = ~n982 & n1432 ;
  assign n1833 = n1832 ^ n1830 ^ 1'b0 ;
  assign n1834 = n1833 ^ n595 ^ 1'b0 ;
  assign n1835 = n1829 | n1834 ;
  assign n1836 = n1525 ^ n610 ^ x119 ;
  assign n1837 = n1449 & n1539 ;
  assign n1838 = n983 | n1837 ;
  assign n1839 = n1836 | n1838 ;
  assign n1840 = n1064 ^ n336 ^ 1'b0 ;
  assign n1841 = n1840 ^ n1420 ^ 1'b0 ;
  assign n1842 = n132 | n1841 ;
  assign n1843 = n225 & n314 ;
  assign n1844 = n1008 ^ n375 ^ 1'b0 ;
  assign n1845 = n1844 ^ n1530 ^ 1'b0 ;
  assign n1846 = ~n1843 & n1845 ;
  assign n1847 = n1842 | n1846 ;
  assign n1850 = n698 | n1619 ;
  assign n1848 = n1085 ^ n663 ^ x100 ;
  assign n1849 = ( ~n407 & n946 ) | ( ~n407 & n1848 ) | ( n946 & n1848 ) ;
  assign n1851 = n1850 ^ n1849 ^ n1589 ;
  assign n1852 = n370 & ~n1307 ;
  assign n1853 = n1852 ^ n1600 ^ 1'b0 ;
  assign n1854 = ( n254 & n551 ) | ( n254 & ~n663 ) | ( n551 & ~n663 ) ;
  assign n1855 = n395 & ~n1854 ;
  assign n1856 = n138 | n254 ;
  assign n1857 = n1266 ^ x119 ^ 1'b0 ;
  assign n1858 = ~n1856 & n1857 ;
  assign n1859 = n802 & ~n1636 ;
  assign n1860 = n1859 ^ n1345 ^ 1'b0 ;
  assign n1861 = ( ~n1379 & n1858 ) | ( ~n1379 & n1860 ) | ( n1858 & n1860 ) ;
  assign n1862 = n517 ^ n240 ^ 1'b0 ;
  assign n1863 = n362 & ~n1862 ;
  assign n1864 = n1568 & n1863 ;
  assign n1865 = n277 | n1480 ;
  assign n1866 = n1865 ^ n1594 ^ 1'b0 ;
  assign n1868 = n659 ^ n204 ^ n163 ;
  assign n1869 = n1868 ^ x49 ^ 1'b0 ;
  assign n1867 = x10 & n1829 ;
  assign n1870 = n1869 ^ n1867 ^ 1'b0 ;
  assign n1871 = n581 & n1424 ;
  assign n1872 = n262 & ~n892 ;
  assign n1873 = n359 | n1197 ;
  assign n1874 = n1854 & ~n1873 ;
  assign n1875 = n319 ^ n265 ^ x95 ;
  assign n1876 = n1583 & ~n1875 ;
  assign n1877 = n829 & ~n1876 ;
  assign n1878 = n1877 ^ n1246 ^ 1'b0 ;
  assign n1879 = n1874 | n1878 ;
  assign n1880 = ~n1687 & n1842 ;
  assign n1881 = n688 | n790 ;
  assign n1882 = n259 & ~n1881 ;
  assign n1883 = n1882 ^ n603 ^ 1'b0 ;
  assign n1884 = x20 & ~n1883 ;
  assign n1885 = n1614 ^ n1499 ^ n730 ;
  assign n1886 = n1641 ^ n1168 ^ n1046 ;
  assign n1887 = n1800 ^ n1034 ^ 1'b0 ;
  assign n1888 = x101 | n1409 ;
  assign n1889 = n739 & ~n1888 ;
  assign n1890 = n639 & n1889 ;
  assign n1891 = n1890 ^ n1554 ^ 1'b0 ;
  assign n1892 = ~n206 & n1891 ;
  assign n1893 = n361 | n1850 ;
  assign n1894 = n1893 ^ n273 ^ 1'b0 ;
  assign n1895 = n1894 ^ n1062 ^ 1'b0 ;
  assign n1896 = n1521 ^ n1046 ^ 1'b0 ;
  assign n1897 = n1895 & ~n1896 ;
  assign n1898 = n949 & n1897 ;
  assign n1899 = ~n1892 & n1898 ;
  assign n1900 = x74 & ~n1885 ;
  assign n1901 = ~n1496 & n1900 ;
  assign n1902 = ~n260 & n671 ;
  assign n1903 = n1902 ^ x16 ^ 1'b0 ;
  assign n1904 = n1903 ^ n499 ^ 1'b0 ;
  assign n1905 = ~n922 & n1904 ;
  assign n1906 = ( ~x27 & x30 ) | ( ~x27 & n449 ) | ( x30 & n449 ) ;
  assign n1907 = ( ~n1231 & n1905 ) | ( ~n1231 & n1906 ) | ( n1905 & n1906 ) ;
  assign n1908 = ~n837 & n952 ;
  assign n1909 = n1908 ^ n1149 ^ 1'b0 ;
  assign n1910 = n1291 ^ n891 ^ 1'b0 ;
  assign n1911 = n463 & ~n1910 ;
  assign n1912 = n1911 ^ n1690 ^ n130 ;
  assign n1913 = x61 ^ x50 ^ 1'b0 ;
  assign n1914 = ~n895 & n1053 ;
  assign n1915 = ~n1372 & n1914 ;
  assign n1916 = n1915 ^ n1821 ^ 1'b0 ;
  assign n1917 = n1913 | n1916 ;
  assign n1918 = n668 ^ n308 ^ x79 ;
  assign n1919 = n1918 ^ n817 ^ n264 ;
  assign n1920 = n712 ^ n323 ^ 1'b0 ;
  assign n1921 = n1680 ^ n953 ^ 1'b0 ;
  assign n1922 = ~n1920 & n1921 ;
  assign n1923 = ( n1332 & ~n1919 ) | ( n1332 & n1922 ) | ( ~n1919 & n1922 ) ;
  assign n1924 = x125 & n1923 ;
  assign n1925 = n1061 ^ n1030 ^ 1'b0 ;
  assign n1926 = x61 & ~n680 ;
  assign n1927 = n1926 ^ n1191 ^ 1'b0 ;
  assign n1928 = n1927 ^ n736 ^ n237 ;
  assign n1929 = n1928 ^ n466 ^ 1'b0 ;
  assign n1930 = ( n888 & ~n1251 ) | ( n888 & n1929 ) | ( ~n1251 & n1929 ) ;
  assign n1931 = n383 & ~n1930 ;
  assign n1932 = n939 ^ n831 ^ 1'b0 ;
  assign n1933 = n469 & n1932 ;
  assign n1934 = n805 & ~n1654 ;
  assign n1935 = ~n1933 & n1934 ;
  assign n1936 = n740 ^ n703 ^ x11 ;
  assign n1937 = n1936 ^ n1242 ^ 1'b0 ;
  assign n1938 = n990 & ~n1937 ;
  assign n1939 = n1789 ^ n564 ^ 1'b0 ;
  assign n1940 = n526 | n602 ;
  assign n1941 = x103 & n1940 ;
  assign n1942 = n413 | n1827 ;
  assign n1943 = n1942 ^ x68 ^ 1'b0 ;
  assign n1944 = n1424 ^ n1323 ^ n773 ;
  assign n1945 = ( x70 & n1019 ) | ( x70 & n1633 ) | ( n1019 & n1633 ) ;
  assign n1946 = n1945 ^ n380 ^ 1'b0 ;
  assign n1947 = ( ~n277 & n713 ) | ( ~n277 & n1124 ) | ( n713 & n1124 ) ;
  assign n1948 = ~n1879 & n1947 ;
  assign n1955 = ( n610 & n871 ) | ( n610 & ~n922 ) | ( n871 & ~n922 ) ;
  assign n1956 = n1416 & ~n1955 ;
  assign n1957 = n1956 ^ n1408 ^ 1'b0 ;
  assign n1953 = ( x5 & n757 ) | ( x5 & ~n1034 ) | ( n757 & ~n1034 ) ;
  assign n1949 = n1088 | n1149 ;
  assign n1950 = n1012 & ~n1949 ;
  assign n1951 = x21 & ~n1065 ;
  assign n1952 = ~n1950 & n1951 ;
  assign n1954 = n1953 ^ n1952 ^ n1394 ;
  assign n1958 = n1957 ^ n1954 ^ 1'b0 ;
  assign n1961 = n861 ^ n189 ^ 1'b0 ;
  assign n1960 = n677 | n775 ;
  assign n1962 = n1961 ^ n1960 ^ 1'b0 ;
  assign n1959 = n1143 ^ n508 ^ 1'b0 ;
  assign n1963 = n1962 ^ n1959 ^ 1'b0 ;
  assign n1964 = n831 & n1476 ;
  assign n1965 = n1848 & n1964 ;
  assign n1966 = ( n519 & ~n1693 ) | ( n519 & n1965 ) | ( ~n1693 & n1965 ) ;
  assign n1967 = n1072 ^ n543 ^ n415 ;
  assign n1968 = n922 | n1967 ;
  assign n1969 = n1162 & ~n1968 ;
  assign n1970 = ~n1966 & n1969 ;
  assign n1971 = ( n854 & n929 ) | ( n854 & n1099 ) | ( n929 & n1099 ) ;
  assign n1972 = ( ~n725 & n1463 ) | ( ~n725 & n1765 ) | ( n1463 & n1765 ) ;
  assign n1973 = n1399 ^ n1111 ^ 1'b0 ;
  assign n1974 = ( x57 & n631 ) | ( x57 & ~n1324 ) | ( n631 & ~n1324 ) ;
  assign n1975 = ~n359 & n1974 ;
  assign n1976 = n1973 & n1975 ;
  assign n1977 = n1976 ^ n1288 ^ n273 ;
  assign n1978 = n804 & n930 ;
  assign n1979 = n1978 ^ n890 ^ 1'b0 ;
  assign n1980 = n1979 ^ n1022 ^ 1'b0 ;
  assign n1981 = n1980 ^ n1655 ^ 1'b0 ;
  assign n1982 = n1472 | n1877 ;
  assign n1983 = n337 & n1122 ;
  assign n1984 = x93 & n947 ;
  assign n1985 = n1984 ^ n1136 ^ 1'b0 ;
  assign n1986 = n1436 & ~n1985 ;
  assign n1987 = ~n370 & n1986 ;
  assign n1988 = n1528 & ~n1786 ;
  assign n1989 = n1987 & n1988 ;
  assign n1990 = n234 | n1067 ;
  assign n1991 = ~n478 & n1217 ;
  assign n1992 = n914 & n1991 ;
  assign n1993 = n507 & n857 ;
  assign n1994 = n707 & n1993 ;
  assign n1995 = ( n719 & n1566 ) | ( n719 & n1994 ) | ( n1566 & n1994 ) ;
  assign n1996 = n1995 ^ n478 ^ x12 ;
  assign n1997 = n1996 ^ n259 ^ x125 ;
  assign n1998 = x21 & x104 ;
  assign n1999 = n592 & n1998 ;
  assign n2001 = ~x2 & n461 ;
  assign n2002 = n2001 ^ n671 ^ n199 ;
  assign n2000 = n1861 ^ n200 ^ 1'b0 ;
  assign n2003 = n2002 ^ n2000 ^ 1'b0 ;
  assign n2005 = n239 | n1212 ;
  assign n2004 = x13 & ~n806 ;
  assign n2006 = n2005 ^ n2004 ^ 1'b0 ;
  assign n2007 = n1633 ^ n553 ^ 1'b0 ;
  assign n2008 = ( ~x3 & x10 ) | ( ~x3 & n1871 ) | ( x10 & n1871 ) ;
  assign n2009 = n143 & n1927 ;
  assign n2010 = n2009 ^ n872 ^ 1'b0 ;
  assign n2011 = ~x11 & n2010 ;
  assign n2012 = n621 & n1928 ;
  assign n2013 = n2012 ^ n1257 ^ 1'b0 ;
  assign n2014 = n631 & n2013 ;
  assign n2015 = n1010 & n1663 ;
  assign n2018 = n385 | n940 ;
  assign n2016 = n1566 ^ n171 ^ 1'b0 ;
  assign n2017 = n487 | n2016 ;
  assign n2019 = n2018 ^ n2017 ^ 1'b0 ;
  assign n2020 = ~x104 & n276 ;
  assign n2021 = n2020 ^ n1261 ^ n1230 ;
  assign n2022 = n1127 ^ n435 ^ 1'b0 ;
  assign n2023 = n1100 & n1407 ;
  assign n2024 = ( n821 & n1022 ) | ( n821 & ~n1155 ) | ( n1022 & ~n1155 ) ;
  assign n2025 = n808 | n2024 ;
  assign n2026 = n2025 ^ x29 ^ 1'b0 ;
  assign n2027 = ( x33 & ~n703 ) | ( x33 & n1854 ) | ( ~n703 & n1854 ) ;
  assign n2028 = n1877 ^ n1010 ^ n893 ;
  assign n2029 = x82 ^ x8 ^ 1'b0 ;
  assign n2030 = x81 & n2029 ;
  assign n2031 = ~n536 & n1587 ;
  assign n2032 = ~n2030 & n2031 ;
  assign n2033 = n2032 ^ n872 ^ 1'b0 ;
  assign n2034 = n2033 ^ n1461 ^ 1'b0 ;
  assign n2035 = n2034 ^ n156 ^ 1'b0 ;
  assign n2036 = n1347 ^ n801 ^ 1'b0 ;
  assign n2037 = n1526 ^ n1343 ^ 1'b0 ;
  assign n2038 = n1940 & n2037 ;
  assign n2039 = n2038 ^ n1493 ^ n965 ;
  assign n2040 = n928 ^ x3 ^ 1'b0 ;
  assign n2042 = x101 & n778 ;
  assign n2043 = n2042 ^ n373 ^ 1'b0 ;
  assign n2041 = n1082 ^ n359 ^ 1'b0 ;
  assign n2044 = n2043 ^ n2041 ^ 1'b0 ;
  assign n2045 = n333 | n2044 ;
  assign n2046 = ( x76 & n189 ) | ( x76 & n1139 ) | ( n189 & n1139 ) ;
  assign n2047 = x54 & n2046 ;
  assign n2048 = n2047 ^ n1820 ^ 1'b0 ;
  assign n2049 = x4 | n1014 ;
  assign n2058 = n1175 ^ n947 ^ n275 ;
  assign n2059 = ( n1432 & n1905 ) | ( n1432 & ~n2058 ) | ( n1905 & ~n2058 ) ;
  assign n2050 = ~n616 & n1125 ;
  assign n2051 = n260 & n2050 ;
  assign n2052 = n447 | n718 ;
  assign n2053 = n2052 ^ n153 ^ 1'b0 ;
  assign n2054 = n2053 ^ n593 ^ 1'b0 ;
  assign n2055 = n781 & n2054 ;
  assign n2056 = ~n920 & n2055 ;
  assign n2057 = n2051 & n2056 ;
  assign n2060 = n2059 ^ n2057 ^ n1251 ;
  assign n2061 = n2060 ^ n1046 ^ 1'b0 ;
  assign n2062 = n2061 ^ n1861 ^ n688 ;
  assign n2063 = n869 & n1639 ;
  assign n2064 = n521 | n1611 ;
  assign n2065 = n1250 & ~n2064 ;
  assign n2066 = x100 & n2002 ;
  assign n2067 = ( n390 & n934 ) | ( n390 & ~n1177 ) | ( n934 & ~n1177 ) ;
  assign n2068 = n1286 ^ n1279 ^ 1'b0 ;
  assign n2069 = n2067 & ~n2068 ;
  assign n2072 = n487 & ~n664 ;
  assign n2073 = n2072 ^ x65 ^ 1'b0 ;
  assign n2071 = n435 & n1868 ;
  assign n2070 = x87 & ~n524 ;
  assign n2074 = n2073 ^ n2071 ^ n2070 ;
  assign n2075 = n1610 | n1901 ;
  assign n2076 = n2074 | n2075 ;
  assign n2086 = n332 ^ x17 ^ 1'b0 ;
  assign n2087 = n691 & n2086 ;
  assign n2088 = ~n562 & n2087 ;
  assign n2089 = n2088 ^ n1933 ^ 1'b0 ;
  assign n2077 = x88 ^ x28 ^ 1'b0 ;
  assign n2078 = x126 ^ x85 ^ 1'b0 ;
  assign n2079 = ~n534 & n2078 ;
  assign n2080 = n461 & n2079 ;
  assign n2081 = n2077 & n2080 ;
  assign n2082 = n1231 & ~n2081 ;
  assign n2083 = n2082 ^ n1025 ^ 1'b0 ;
  assign n2084 = n2083 ^ n790 ^ 1'b0 ;
  assign n2085 = n1120 & n2084 ;
  assign n2090 = n2089 ^ n2085 ^ 1'b0 ;
  assign n2091 = n206 | n488 ;
  assign n2092 = n2091 ^ n469 ^ 1'b0 ;
  assign n2093 = n667 | n2092 ;
  assign n2094 = n1135 & ~n2093 ;
  assign n2095 = n716 & ~n2094 ;
  assign n2096 = n2095 ^ n260 ^ 1'b0 ;
  assign n2097 = n138 & n2096 ;
  assign n2098 = n2097 ^ n1133 ^ 1'b0 ;
  assign n2099 = x101 & ~n309 ;
  assign n2100 = ~n1677 & n2099 ;
  assign n2101 = n319 & n2100 ;
  assign n2102 = ~n1480 & n2101 ;
  assign n2103 = x116 | n2102 ;
  assign n2104 = n1003 | n1922 ;
  assign n2105 = n935 & n2104 ;
  assign n2106 = n655 ^ n645 ^ x31 ;
  assign n2107 = n2106 ^ n539 ^ n533 ;
  assign n2108 = n2107 ^ n150 ^ 1'b0 ;
  assign n2109 = n1006 & ~n2022 ;
  assign n2110 = n984 ^ n799 ^ 1'b0 ;
  assign n2111 = n1209 | n2110 ;
  assign n2112 = n1557 ^ x97 ^ x64 ;
  assign n2113 = n2112 ^ n341 ^ 1'b0 ;
  assign n2114 = ~n1403 & n1765 ;
  assign n2115 = n369 & n2114 ;
  assign n2116 = n1034 | n2115 ;
  assign n2117 = n2116 ^ n1399 ^ 1'b0 ;
  assign n2118 = n2052 ^ n1728 ^ n953 ;
  assign n2119 = n2118 ^ n2061 ^ n311 ;
  assign n2120 = ~n730 & n1564 ;
  assign n2121 = n2120 ^ n840 ^ 1'b0 ;
  assign n2122 = n988 | n2121 ;
  assign n2124 = n1022 ^ n927 ^ 1'b0 ;
  assign n2125 = n355 | n2124 ;
  assign n2123 = n342 | n485 ;
  assign n2126 = n2125 ^ n2123 ^ 1'b0 ;
  assign n2127 = n229 | n1031 ;
  assign n2128 = n369 & ~n2127 ;
  assign n2129 = n439 | n2128 ;
  assign n2130 = n2129 ^ n393 ^ 1'b0 ;
  assign n2131 = n886 & ~n1718 ;
  assign n2132 = n2130 & n2131 ;
  assign n2133 = n1393 & ~n1428 ;
  assign n2134 = ~n731 & n897 ;
  assign n2135 = n282 & n2134 ;
  assign n2136 = n1936 & ~n2135 ;
  assign n2137 = n2136 ^ n651 ^ 1'b0 ;
  assign n2138 = n1708 & ~n1728 ;
  assign n2139 = ~n638 & n1958 ;
  assign n2140 = ~n1235 & n2139 ;
  assign n2141 = n2140 ^ n1033 ^ 1'b0 ;
  assign n2142 = n308 & n2141 ;
  assign n2143 = n210 | n214 ;
  assign n2144 = ~n466 & n1884 ;
  assign n2145 = n2144 ^ n567 ^ 1'b0 ;
  assign n2146 = ~n2143 & n2145 ;
  assign n2147 = n1498 ^ n494 ^ 1'b0 ;
  assign n2148 = ~n748 & n1050 ;
  assign n2149 = n1496 ^ n730 ^ 1'b0 ;
  assign n2150 = n229 | n231 ;
  assign n2151 = n2149 | n2150 ;
  assign n2152 = ( ~n405 & n1851 ) | ( ~n405 & n1854 ) | ( n1851 & n1854 ) ;
  assign n2153 = n562 ^ n486 ^ 1'b0 ;
  assign n2154 = n1520 & n2153 ;
  assign n2155 = ~n1388 & n2154 ;
  assign n2156 = n497 & n1089 ;
  assign n2157 = ~n603 & n2156 ;
  assign n2158 = x88 & ~n744 ;
  assign n2159 = ~x16 & n2158 ;
  assign n2160 = n1724 & n2159 ;
  assign n2161 = n2112 ^ x50 ^ 1'b0 ;
  assign n2162 = n245 & ~n2161 ;
  assign n2163 = n1206 & ~n1269 ;
  assign n2164 = n2163 ^ n482 ^ 1'b0 ;
  assign n2165 = n1130 & ~n1919 ;
  assign n2166 = ~n2015 & n2165 ;
  assign n2167 = n1675 ^ x72 ^ 1'b0 ;
  assign n2168 = n1513 ^ n210 ^ 1'b0 ;
  assign n2169 = n2167 | n2168 ;
  assign n2170 = n969 & ~n2169 ;
  assign n2171 = n1099 ^ n314 ^ 1'b0 ;
  assign n2172 = n1571 & ~n2171 ;
  assign n2173 = ( n319 & n1580 ) | ( n319 & n2172 ) | ( n1580 & n2172 ) ;
  assign n2177 = n2020 ^ n421 ^ 1'b0 ;
  assign n2178 = x12 & ~n2177 ;
  assign n2174 = n1498 ^ x2 ^ 1'b0 ;
  assign n2175 = n817 & ~n2174 ;
  assign n2176 = n830 | n2175 ;
  assign n2179 = n2178 ^ n2176 ^ 1'b0 ;
  assign n2180 = n2173 & ~n2179 ;
  assign n2181 = x42 & n345 ;
  assign n2182 = n1514 & n2181 ;
  assign n2183 = n2106 ^ n612 ^ 1'b0 ;
  assign n2184 = n2182 | n2183 ;
  assign n2185 = n592 & n1791 ;
  assign n2186 = n2185 ^ n1800 ^ 1'b0 ;
  assign n2187 = n1337 | n2186 ;
  assign n2188 = ~n288 & n1217 ;
  assign n2189 = n237 & n2188 ;
  assign n2190 = n353 ^ x94 ^ 1'b0 ;
  assign n2191 = n2190 ^ n744 ^ 1'b0 ;
  assign n2192 = ~n2189 & n2191 ;
  assign n2193 = n1679 ^ n582 ^ n449 ;
  assign n2194 = ~n2192 & n2193 ;
  assign n2198 = n1492 ^ n633 ^ 1'b0 ;
  assign n2195 = n694 | n1761 ;
  assign n2196 = n2195 ^ n536 ^ 1'b0 ;
  assign n2197 = ~n1425 & n2196 ;
  assign n2199 = n2198 ^ n2197 ^ 1'b0 ;
  assign n2203 = n603 | n785 ;
  assign n2200 = ~n141 & n1248 ;
  assign n2201 = ( n352 & n754 ) | ( n352 & n2200 ) | ( n754 & n2200 ) ;
  assign n2202 = n2201 ^ n1504 ^ n149 ;
  assign n2204 = n2203 ^ n2202 ^ n1352 ;
  assign n2205 = n1607 | n2101 ;
  assign n2206 = n901 ^ n849 ^ n664 ;
  assign n2207 = n2206 ^ n1123 ^ 1'b0 ;
  assign n2211 = n1690 ^ x57 ^ 1'b0 ;
  assign n2212 = n1420 | n2211 ;
  assign n2213 = n2212 ^ x75 ^ 1'b0 ;
  assign n2214 = x28 & ~n2213 ;
  assign n2215 = n2214 ^ n639 ^ 1'b0 ;
  assign n2216 = n1321 & ~n2215 ;
  assign n2208 = ~n190 & n620 ;
  assign n2209 = n2208 ^ n1031 ^ 1'b0 ;
  assign n2210 = ~n581 & n2209 ;
  assign n2217 = n2216 ^ n2210 ^ 1'b0 ;
  assign n2218 = n1070 ^ n252 ^ 1'b0 ;
  assign n2219 = n1930 ^ n593 ^ 1'b0 ;
  assign n2220 = ( n197 & n802 ) | ( n197 & n1694 ) | ( n802 & n1694 ) ;
  assign n2221 = n2193 ^ n1663 ^ n912 ;
  assign n2222 = n186 | n454 ;
  assign n2223 = ( x115 & n366 ) | ( x115 & n922 ) | ( n366 & n922 ) ;
  assign n2224 = x66 & n561 ;
  assign n2225 = n2223 & n2224 ;
  assign n2233 = ( x53 & n189 ) | ( x53 & ~n1624 ) | ( n189 & ~n1624 ) ;
  assign n2232 = n470 & ~n740 ;
  assign n2234 = n2233 ^ n2232 ^ 1'b0 ;
  assign n2235 = n2234 ^ n419 ^ 1'b0 ;
  assign n2236 = ~n212 & n2235 ;
  assign n2228 = n801 & ~n808 ;
  assign n2229 = n2228 ^ n648 ^ 1'b0 ;
  assign n2230 = n1449 ^ n534 ^ 1'b0 ;
  assign n2231 = n2229 & ~n2230 ;
  assign n2237 = n2236 ^ n2231 ^ n840 ;
  assign n2226 = x12 & ~n1742 ;
  assign n2227 = ~n982 & n2226 ;
  assign n2238 = n2237 ^ n2227 ^ 1'b0 ;
  assign n2239 = ~n930 & n1454 ;
  assign n2240 = n2239 ^ n1798 ^ 1'b0 ;
  assign n2241 = n2238 & ~n2240 ;
  assign n2242 = n631 & n2241 ;
  assign n2243 = n2242 ^ n1842 ^ 1'b0 ;
  assign n2244 = ( n2222 & ~n2225 ) | ( n2222 & n2243 ) | ( ~n2225 & n2243 ) ;
  assign n2245 = n850 ^ x100 ^ 1'b0 ;
  assign n2246 = n218 & ~n2245 ;
  assign n2247 = n1732 & n2246 ;
  assign n2248 = n445 & n2247 ;
  assign n2249 = n2248 ^ n904 ^ 1'b0 ;
  assign n2250 = n309 & n570 ;
  assign n2251 = n1607 & ~n1753 ;
  assign n2252 = n2251 ^ n1994 ^ 1'b0 ;
  assign n2253 = n1041 ^ n376 ^ n290 ;
  assign n2254 = ~n2125 & n2253 ;
  assign n2256 = n422 & ~n605 ;
  assign n2257 = ~n1920 & n2256 ;
  assign n2255 = n355 ^ n247 ^ x75 ;
  assign n2258 = n2257 ^ n2255 ^ 1'b0 ;
  assign n2259 = n829 & ~n2258 ;
  assign n2260 = n421 & n463 ;
  assign n2261 = n1002 | n1099 ;
  assign n2262 = n884 & ~n2261 ;
  assign n2263 = x33 & ~n2262 ;
  assign n2264 = ~n1788 & n2263 ;
  assign n2265 = n1741 & n1958 ;
  assign n2266 = n2264 & n2265 ;
  assign n2269 = x75 & n502 ;
  assign n2270 = n2269 ^ n1829 ^ 1'b0 ;
  assign n2267 = x27 | n2043 ;
  assign n2268 = n2267 ^ n408 ^ 1'b0 ;
  assign n2271 = n2270 ^ n2268 ^ 1'b0 ;
  assign n2272 = n474 | n1700 ;
  assign n2274 = ~n471 & n620 ;
  assign n2275 = n2274 ^ n194 ^ 1'b0 ;
  assign n2276 = n1059 ^ n526 ^ 1'b0 ;
  assign n2277 = n2275 & ~n2276 ;
  assign n2273 = ~n742 & n1972 ;
  assign n2278 = n2277 ^ n2273 ^ 1'b0 ;
  assign n2279 = n1195 ^ x116 ^ 1'b0 ;
  assign n2280 = n2279 ^ n1600 ^ 1'b0 ;
  assign n2281 = n2280 ^ n1757 ^ 1'b0 ;
  assign n2282 = ~n738 & n2281 ;
  assign n2283 = ( n254 & n1085 ) | ( n254 & n2239 ) | ( n1085 & n2239 ) ;
  assign n2284 = n2283 ^ n952 ^ 1'b0 ;
  assign n2285 = n1077 | n2284 ;
  assign n2289 = n396 & n1246 ;
  assign n2286 = n872 & ~n1923 ;
  assign n2287 = ~n2214 & n2286 ;
  assign n2288 = n450 & ~n2287 ;
  assign n2290 = n2289 ^ n2288 ^ 1'b0 ;
  assign n2291 = n1603 | n2290 ;
  assign n2292 = ( n563 & n2285 ) | ( n563 & ~n2291 ) | ( n2285 & ~n2291 ) ;
  assign n2293 = n1499 ^ n654 ^ 1'b0 ;
  assign n2294 = n176 ^ x110 ^ 1'b0 ;
  assign n2295 = n398 & n2294 ;
  assign n2296 = n2295 ^ x80 ^ 1'b0 ;
  assign n2297 = ( n1705 & ~n2102 ) | ( n1705 & n2296 ) | ( ~n2102 & n2296 ) ;
  assign n2298 = n277 | n1172 ;
  assign n2299 = n368 & ~n2298 ;
  assign n2300 = n2160 | n2299 ;
  assign n2301 = n1268 ^ n310 ^ 1'b0 ;
  assign n2302 = n1815 & ~n2301 ;
  assign n2303 = x16 & n2282 ;
  assign n2304 = n2303 ^ n1002 ^ 1'b0 ;
  assign n2305 = n1455 ^ n1387 ^ 1'b0 ;
  assign n2306 = n2305 ^ n686 ^ 1'b0 ;
  assign n2307 = n1306 ^ n1135 ^ 1'b0 ;
  assign n2308 = n2307 ^ n1065 ^ 1'b0 ;
  assign n2309 = n1851 & ~n2308 ;
  assign n2310 = n1034 ^ x18 ^ 1'b0 ;
  assign n2311 = n2310 ^ n1364 ^ 1'b0 ;
  assign n2312 = n778 & n2311 ;
  assign n2313 = ~n214 & n692 ;
  assign n2314 = n129 & n1534 ;
  assign n2315 = n2314 ^ n1540 ^ 1'b0 ;
  assign n2316 = n1650 ^ n919 ^ n848 ;
  assign n2317 = n1443 | n2316 ;
  assign n2318 = n1192 ^ n508 ^ 1'b0 ;
  assign n2320 = n690 & n1299 ;
  assign n2321 = n2320 ^ n1853 ^ 1'b0 ;
  assign n2322 = n1197 & ~n2321 ;
  assign n2319 = n234 & n1669 ;
  assign n2323 = n2322 ^ n2319 ^ 1'b0 ;
  assign n2324 = n2146 | n2323 ;
  assign n2325 = n2318 | n2324 ;
  assign n2326 = n1286 ^ n547 ^ 1'b0 ;
  assign n2327 = n636 & n1626 ;
  assign n2328 = n2327 ^ n1390 ^ 1'b0 ;
  assign n2329 = n2328 ^ n1894 ^ 1'b0 ;
  assign n2330 = n2329 ^ n1594 ^ 1'b0 ;
  assign n2331 = x111 & ~n312 ;
  assign n2332 = x71 & n2331 ;
  assign n2333 = n2332 ^ n873 ^ 1'b0 ;
  assign n2334 = n2333 ^ n1264 ^ x105 ;
  assign n2335 = n457 & n943 ;
  assign n2336 = n770 ^ x42 ^ 1'b0 ;
  assign n2337 = n395 & n2336 ;
  assign n2338 = n422 & ~n1795 ;
  assign n2339 = ~n2337 & n2338 ;
  assign n2340 = n179 ^ n158 ^ 1'b0 ;
  assign n2341 = n1554 & n2340 ;
  assign n2342 = n2197 ^ n1745 ^ 1'b0 ;
  assign n2343 = n2012 ^ n1492 ^ n590 ;
  assign n2344 = n946 & ~n2343 ;
  assign n2345 = n2237 & n2344 ;
  assign n2346 = ~n1869 & n1989 ;
  assign n2349 = ( n811 & n1195 ) | ( n811 & n2331 ) | ( n1195 & n2331 ) ;
  assign n2350 = n2349 ^ n632 ^ 1'b0 ;
  assign n2347 = n1261 ^ n388 ^ 1'b0 ;
  assign n2348 = ~n1765 & n2347 ;
  assign n2351 = n2350 ^ n2348 ^ 1'b0 ;
  assign n2352 = x38 & ~n1408 ;
  assign n2353 = n2352 ^ n852 ^ 1'b0 ;
  assign n2354 = ( ~n150 & n1530 ) | ( ~n150 & n2353 ) | ( n1530 & n2353 ) ;
  assign n2355 = ( x93 & ~n517 ) | ( x93 & n1203 ) | ( ~n517 & n1203 ) ;
  assign n2356 = n2355 ^ n535 ^ n431 ;
  assign n2357 = n2354 & ~n2356 ;
  assign n2358 = n1716 ^ n950 ^ 1'b0 ;
  assign n2359 = n2112 & ~n2358 ;
  assign n2360 = n1072 ^ x25 ^ 1'b0 ;
  assign n2361 = n473 | n2360 ;
  assign n2362 = n877 & ~n1761 ;
  assign n2363 = n830 ^ n267 ^ 1'b0 ;
  assign n2364 = ~n2122 & n2363 ;
  assign n2365 = n2337 ^ n1184 ^ 1'b0 ;
  assign n2366 = n728 & ~n1700 ;
  assign n2367 = n1677 ^ n445 ^ 1'b0 ;
  assign n2368 = n2366 & n2367 ;
  assign n2370 = n454 & ~n558 ;
  assign n2371 = n2370 ^ n386 ^ 1'b0 ;
  assign n2372 = n1198 ^ n707 ^ 1'b0 ;
  assign n2373 = n1140 & n2372 ;
  assign n2374 = n2373 ^ n1810 ^ 1'b0 ;
  assign n2375 = n928 | n2374 ;
  assign n2376 = ( n166 & ~n2371 ) | ( n166 & n2375 ) | ( ~n2371 & n2375 ) ;
  assign n2369 = n1159 ^ n838 ^ 1'b0 ;
  assign n2377 = n2376 ^ n2369 ^ n848 ;
  assign n2378 = n2377 ^ n1244 ^ 1'b0 ;
  assign n2379 = n1868 | n2378 ;
  assign n2380 = n1212 ^ n798 ^ 1'b0 ;
  assign n2381 = n703 & ~n2380 ;
  assign n2382 = n1375 & n2381 ;
  assign n2383 = n2382 ^ n204 ^ x68 ;
  assign n2384 = n508 | n1370 ;
  assign n2385 = ~n1197 & n2384 ;
  assign n2386 = ~n1997 & n2385 ;
  assign n2387 = n1680 ^ n791 ^ 1'b0 ;
  assign n2388 = n890 & n2387 ;
  assign n2389 = n2388 ^ n348 ^ 1'b0 ;
  assign n2390 = n1329 ^ n338 ^ 1'b0 ;
  assign n2391 = n2390 ^ x113 ^ 1'b0 ;
  assign n2392 = n785 ^ n645 ^ 1'b0 ;
  assign n2393 = n2391 & n2392 ;
  assign n2394 = n1168 & ~n1193 ;
  assign n2395 = ~n2053 & n2394 ;
  assign n2396 = n1140 | n2094 ;
  assign n2397 = n2396 ^ n1115 ^ 1'b0 ;
  assign n2398 = n1031 ^ n722 ^ 1'b0 ;
  assign n2399 = ~n215 & n1567 ;
  assign n2400 = n2398 | n2399 ;
  assign n2401 = n1319 | n2400 ;
  assign n2402 = x23 & ~n1059 ;
  assign n2403 = n503 & n2402 ;
  assign n2404 = n730 & n2403 ;
  assign n2405 = n138 ^ x28 ^ 1'b0 ;
  assign n2406 = n681 & n2405 ;
  assign n2407 = n220 | n1408 ;
  assign n2408 = n2406 | n2407 ;
  assign n2409 = n2408 ^ n2222 ^ 1'b0 ;
  assign n2410 = n578 ^ x80 ^ 1'b0 ;
  assign n2411 = n1746 & ~n2410 ;
  assign n2412 = ~n149 & n2411 ;
  assign n2413 = n2412 ^ n671 ^ 1'b0 ;
  assign n2414 = n2005 ^ n969 ^ n445 ;
  assign n2415 = n361 & ~n2414 ;
  assign n2416 = n1213 & ~n1757 ;
  assign n2417 = n2416 ^ n450 ^ 1'b0 ;
  assign n2418 = n189 | n2417 ;
  assign n2419 = n2418 ^ n1424 ^ 1'b0 ;
  assign n2420 = n2419 ^ n490 ^ 1'b0 ;
  assign n2421 = ( n380 & ~n2415 ) | ( n380 & n2420 ) | ( ~n2415 & n2420 ) ;
  assign n2422 = ( x0 & x121 ) | ( x0 & ~n156 ) | ( x121 & ~n156 ) ;
  assign n2423 = n2422 ^ n2384 ^ 1'b0 ;
  assign n2424 = n212 | n578 ;
  assign n2425 = n1292 & ~n2424 ;
  assign n2426 = n2425 ^ n1412 ^ n1075 ;
  assign n2427 = ~n673 & n962 ;
  assign n2428 = n2426 & n2427 ;
  assign n2429 = n748 & ~n1950 ;
  assign n2430 = ( n746 & n942 ) | ( n746 & ~n988 ) | ( n942 & ~n988 ) ;
  assign n2431 = ~n2429 & n2430 ;
  assign n2432 = n2431 ^ n786 ^ 1'b0 ;
  assign n2433 = n1397 ^ n149 ^ 1'b0 ;
  assign n2434 = n1006 & ~n1041 ;
  assign n2435 = n2420 & n2434 ;
  assign n2436 = n1641 ^ n1004 ^ 1'b0 ;
  assign n2437 = n2436 ^ n728 ^ 1'b0 ;
  assign n2438 = n2437 ^ n1079 ^ n411 ;
  assign n2439 = x95 & n1884 ;
  assign n2440 = ~n1428 & n2439 ;
  assign n2441 = n2440 ^ x113 ^ 1'b0 ;
  assign n2442 = n2441 ^ n2102 ^ n136 ;
  assign n2443 = n2442 ^ n1535 ^ 1'b0 ;
  assign n2444 = ( x120 & n264 ) | ( x120 & n700 ) | ( n264 & n700 ) ;
  assign n2445 = n1442 & ~n2444 ;
  assign n2446 = n935 & n1218 ;
  assign n2447 = ~n1195 & n2446 ;
  assign n2448 = ( n191 & n443 ) | ( n191 & n1041 ) | ( n443 & n1041 ) ;
  assign n2449 = x76 & n2448 ;
  assign n2450 = n1124 ^ n691 ^ 1'b0 ;
  assign n2451 = n2408 & n2450 ;
  assign n2452 = n2449 | n2451 ;
  assign n2453 = n2447 & ~n2452 ;
  assign n2454 = n449 | n1440 ;
  assign n2455 = n2454 ^ x26 ^ 1'b0 ;
  assign n2456 = n2455 ^ n617 ^ n216 ;
  assign n2457 = n910 ^ n632 ^ 1'b0 ;
  assign n2458 = ~n625 & n2096 ;
  assign n2459 = ~n1572 & n2458 ;
  assign n2463 = ( ~n375 & n674 ) | ( ~n375 & n1163 ) | ( n674 & n1163 ) ;
  assign n2464 = ( n642 & n2059 ) | ( n642 & n2463 ) | ( n2059 & n2463 ) ;
  assign n2465 = n1490 | n2464 ;
  assign n2460 = n1940 ^ n619 ^ 1'b0 ;
  assign n2461 = ~n932 & n2460 ;
  assign n2462 = n2461 ^ n708 ^ 1'b0 ;
  assign n2466 = n2465 ^ n2462 ^ 1'b0 ;
  assign n2467 = x92 & ~n801 ;
  assign n2468 = n549 & ~n2467 ;
  assign n2469 = n2468 ^ n1791 ^ 1'b0 ;
  assign n2470 = n2451 ^ n1594 ^ 1'b0 ;
  assign n2471 = n2469 | n2470 ;
  assign n2472 = n1644 ^ n332 ^ 1'b0 ;
  assign n2473 = n2472 ^ n1405 ^ 1'b0 ;
  assign n2474 = x78 | x121 ;
  assign n2481 = n1953 & ~n2094 ;
  assign n2482 = n2481 ^ n1279 ^ 1'b0 ;
  assign n2483 = n597 | n2482 ;
  assign n2475 = x94 ^ x3 ^ 1'b0 ;
  assign n2476 = ~n202 & n2475 ;
  assign n2477 = n1680 ^ n760 ^ 1'b0 ;
  assign n2478 = n1079 & n2477 ;
  assign n2479 = n2478 ^ x59 ^ 1'b0 ;
  assign n2480 = n2476 & ~n2479 ;
  assign n2484 = n2483 ^ n2480 ^ 1'b0 ;
  assign n2488 = n376 & ~n627 ;
  assign n2489 = n225 & n2488 ;
  assign n2490 = n2489 ^ n1555 ^ n970 ;
  assign n2485 = n398 | n2099 ;
  assign n2486 = n594 & n2485 ;
  assign n2487 = n2486 ^ n876 ^ 1'b0 ;
  assign n2491 = n2490 ^ n2487 ^ 1'b0 ;
  assign n2492 = n1535 | n2491 ;
  assign n2493 = n2492 ^ n582 ^ 1'b0 ;
  assign n2494 = n341 ^ x55 ^ 1'b0 ;
  assign n2495 = n2494 ^ n686 ^ n646 ;
  assign n2496 = n2495 ^ n1095 ^ 1'b0 ;
  assign n2497 = n2244 ^ n2130 ^ 1'b0 ;
  assign n2498 = n808 | n2497 ;
  assign n2499 = n1358 & n1442 ;
  assign n2500 = n2499 ^ n1368 ^ 1'b0 ;
  assign n2501 = n2341 ^ x37 ^ 1'b0 ;
  assign n2502 = n2371 ^ n1050 ^ 1'b0 ;
  assign n2503 = n1192 & ~n2502 ;
  assign n2504 = n2111 ^ n373 ^ 1'b0 ;
  assign n2505 = n2503 & ~n2504 ;
  assign n2506 = n962 | n2277 ;
  assign n2507 = x97 ^ x33 ^ 1'b0 ;
  assign n2508 = n1868 ^ n686 ^ x46 ;
  assign n2509 = ( n1168 & ~n1948 ) | ( n1168 & n2508 ) | ( ~n1948 & n2508 ) ;
  assign n2510 = ~n563 & n996 ;
  assign n2511 = n2510 ^ n1055 ^ n969 ;
  assign n2512 = n1710 ^ n225 ^ 1'b0 ;
  assign n2513 = n2511 | n2512 ;
  assign n2514 = ~n886 & n1580 ;
  assign n2515 = n2514 ^ n2275 ^ n562 ;
  assign n2516 = n2515 ^ n2494 ^ 1'b0 ;
  assign n2517 = n2371 | n2516 ;
  assign n2518 = ~n319 & n1166 ;
  assign n2519 = n2518 ^ n1706 ^ 1'b0 ;
  assign n2520 = n150 & n332 ;
  assign n2521 = ~n1481 & n2520 ;
  assign n2522 = n1324 ^ n642 ^ 1'b0 ;
  assign n2523 = n2522 ^ n707 ^ 1'b0 ;
  assign n2524 = n2523 ^ n2254 ^ 1'b0 ;
  assign n2525 = n1352 & ~n2524 ;
  assign n2526 = n1637 ^ n1272 ^ 1'b0 ;
  assign n2527 = n1728 & n2526 ;
  assign n2528 = ~n1842 & n2527 ;
  assign n2529 = n2125 ^ n193 ^ 1'b0 ;
  assign n2530 = n1644 & ~n1786 ;
  assign n2531 = n369 & n2530 ;
  assign n2532 = ( n480 & n1088 ) | ( n480 & ~n1235 ) | ( n1088 & ~n1235 ) ;
  assign n2533 = n1435 ^ x100 ^ 1'b0 ;
  assign n2534 = n362 & n2533 ;
  assign n2535 = n1693 ^ n1451 ^ n1300 ;
  assign n2536 = n2534 & ~n2535 ;
  assign n2537 = ~n1030 & n2536 ;
  assign n2538 = ( ~n2089 & n2133 ) | ( ~n2089 & n2244 ) | ( n2133 & n2244 ) ;
  assign n2547 = n889 ^ n248 ^ x10 ;
  assign n2548 = n2547 ^ n854 ^ 1'b0 ;
  assign n2549 = n341 & n2548 ;
  assign n2542 = n683 ^ n267 ^ 1'b0 ;
  assign n2543 = x92 & ~n2542 ;
  assign n2544 = n2543 ^ x77 ^ 1'b0 ;
  assign n2545 = n1195 & ~n2544 ;
  assign n2546 = n2545 ^ n1973 ^ 1'b0 ;
  assign n2539 = n398 | n475 ;
  assign n2540 = n980 | n2539 ;
  assign n2541 = n2540 ^ n2353 ^ 1'b0 ;
  assign n2550 = n2549 ^ n2546 ^ n2541 ;
  assign n2551 = n1232 ^ n652 ^ 1'b0 ;
  assign n2552 = n2551 ^ n1690 ^ n450 ;
  assign n2553 = n2552 ^ n2406 ^ n1853 ;
  assign n2554 = n673 & ~n2553 ;
  assign n2555 = x19 & x62 ;
  assign n2556 = n2440 & n2555 ;
  assign n2559 = x121 & ~n2239 ;
  assign n2560 = n969 & n2559 ;
  assign n2561 = n436 & n1313 ;
  assign n2562 = n2561 ^ n2226 ^ 1'b0 ;
  assign n2563 = n2562 ^ n599 ^ 1'b0 ;
  assign n2564 = ~n2560 & n2563 ;
  assign n2557 = n1283 & n1568 ;
  assign n2558 = n2557 ^ n1952 ^ 1'b0 ;
  assign n2565 = n2564 ^ n2558 ^ 1'b0 ;
  assign n2566 = ~n1994 & n2565 ;
  assign n2568 = x57 & n381 ;
  assign n2567 = ~n1150 & n1775 ;
  assign n2569 = n2568 ^ n2567 ^ 1'b0 ;
  assign n2570 = ~n895 & n2059 ;
  assign n2571 = n1977 ^ n175 ^ 1'b0 ;
  assign n2572 = n1769 & n2017 ;
  assign n2573 = ~n349 & n2572 ;
  assign n2574 = n1597 & n2573 ;
  assign n2575 = n1088 & n2574 ;
  assign n2576 = n1581 ^ n320 ^ 1'b0 ;
  assign n2577 = n1237 & ~n2576 ;
  assign n2578 = n2546 ^ n1511 ^ 1'b0 ;
  assign n2579 = n2194 | n2578 ;
  assign n2580 = ~n1008 & n2028 ;
  assign n2581 = n2580 ^ n726 ^ 1'b0 ;
  assign n2582 = n2581 ^ n2113 ^ 1'b0 ;
  assign n2583 = n197 & ~n543 ;
  assign n2584 = n2583 ^ n2511 ^ 1'b0 ;
  assign n2585 = ~n868 & n2584 ;
  assign n2586 = n1275 ^ n1074 ^ 1'b0 ;
  assign n2587 = ~n265 & n1407 ;
  assign n2588 = ~n389 & n2587 ;
  assign n2589 = n683 | n2588 ;
  assign n2590 = ~n381 & n2589 ;
  assign n2591 = ( n279 & ~n1476 ) | ( n279 & n2414 ) | ( ~n1476 & n2414 ) ;
  assign n2592 = x36 | n859 ;
  assign n2593 = ( ~x60 & n2154 ) | ( ~x60 & n2592 ) | ( n2154 & n2592 ) ;
  assign n2594 = ( n177 & ~n1230 ) | ( n177 & n2593 ) | ( ~n1230 & n2593 ) ;
  assign n2595 = n1721 ^ n1143 ^ 1'b0 ;
  assign n2596 = x7 & ~n594 ;
  assign n2597 = ( ~x52 & n652 ) | ( ~x52 & n2162 ) | ( n652 & n2162 ) ;
  assign n2598 = n1721 ^ n661 ^ 1'b0 ;
  assign n2599 = n2178 & ~n2598 ;
  assign n2600 = ( ~n910 & n2155 ) | ( ~n910 & n2444 ) | ( n2155 & n2444 ) ;
  assign n2601 = x91 & n130 ;
  assign n2602 = n2601 ^ x38 ^ 1'b0 ;
  assign n2603 = n2340 | n2602 ;
  assign n2604 = n2603 ^ n1629 ^ 1'b0 ;
  assign n2605 = n2275 | n2604 ;
  assign n2606 = ~n487 & n2326 ;
  assign n2607 = n818 & n1403 ;
  assign n2608 = n493 ^ x1 ^ 1'b0 ;
  assign n2609 = n1549 | n2608 ;
  assign n2610 = n1506 ^ n1012 ^ 1'b0 ;
  assign n2611 = n2610 ^ n2472 ^ 1'b0 ;
  assign n2613 = n2295 ^ n1809 ^ 1'b0 ;
  assign n2614 = n1117 & n2033 ;
  assign n2615 = ~n2613 & n2614 ;
  assign n2612 = n2259 ^ n1529 ^ 1'b0 ;
  assign n2616 = n2615 ^ n2612 ^ 1'b0 ;
  assign n2617 = n1950 & n2616 ;
  assign n2618 = n425 & n1920 ;
  assign n2619 = n1173 ^ n586 ^ 1'b0 ;
  assign n2620 = n1191 ^ n1141 ^ 1'b0 ;
  assign n2621 = n1324 ^ n478 ^ x12 ;
  assign n2622 = n1771 ^ n1742 ^ 1'b0 ;
  assign n2623 = n1655 & ~n2622 ;
  assign n2624 = n1953 & n2623 ;
  assign n2625 = ~n2108 & n2624 ;
  assign n2626 = x28 & n2463 ;
  assign n2627 = ~n161 & n2626 ;
  assign n2628 = n2546 & ~n2627 ;
  assign n2629 = n2625 & n2628 ;
  assign n2630 = x44 & x72 ;
  assign n2631 = n2630 ^ n805 ^ 1'b0 ;
  assign n2632 = n838 | n2631 ;
  assign n2633 = n739 & ~n2632 ;
  assign n2634 = ~x124 & n2633 ;
  assign n2635 = n2634 ^ n1070 ^ 1'b0 ;
  assign n2636 = n366 | n2635 ;
  assign n2637 = ~n381 & n2636 ;
  assign n2638 = x91 & n210 ;
  assign n2639 = n1679 ^ n988 ^ 1'b0 ;
  assign n2640 = n2638 | n2639 ;
  assign n2641 = x93 & n2640 ;
  assign n2642 = n2637 & n2641 ;
  assign n2643 = n733 ^ n319 ^ 1'b0 ;
  assign n2644 = x50 & n2643 ;
  assign n2645 = n2644 ^ n454 ^ 1'b0 ;
  assign n2646 = x50 & ~n1362 ;
  assign n2647 = n2645 & n2646 ;
  assign n2648 = n1123 & n2647 ;
  assign n2649 = ~x13 & n2648 ;
  assign n2650 = x20 & n419 ;
  assign n2651 = n2650 ^ n2638 ^ 1'b0 ;
  assign n2652 = n2651 ^ x121 ^ 1'b0 ;
  assign n2653 = n872 | n2027 ;
  assign n2654 = n1374 & ~n2653 ;
  assign n2655 = ~n1382 & n2605 ;
  assign n2656 = ~n848 & n2655 ;
  assign n2659 = n746 & ~n986 ;
  assign n2660 = n2659 ^ n2197 ^ 1'b0 ;
  assign n2661 = ( n179 & ~n190 ) | ( n179 & n2660 ) | ( ~n190 & n2660 ) ;
  assign n2657 = ( n760 & ~n1069 ) | ( n760 & n1765 ) | ( ~n1069 & n1765 ) ;
  assign n2658 = ( n882 & ~n1352 ) | ( n882 & n2657 ) | ( ~n1352 & n2657 ) ;
  assign n2662 = n2661 ^ n2658 ^ 1'b0 ;
  assign n2663 = ( n236 & ~n605 ) | ( n236 & n1288 ) | ( ~n605 & n1288 ) ;
  assign n2664 = n2663 ^ n1680 ^ 1'b0 ;
  assign n2665 = ~n2660 & n2664 ;
  assign n2666 = n2665 ^ n2299 ^ n1624 ;
  assign n2667 = n231 & n1312 ;
  assign n2668 = n891 | n2455 ;
  assign n2669 = ~n654 & n2668 ;
  assign n2670 = n2669 ^ n235 ^ 1'b0 ;
  assign n2671 = n1533 & ~n2640 ;
  assign n2672 = n752 & n2234 ;
  assign n2673 = n503 & n2030 ;
  assign n2674 = n1034 & ~n2673 ;
  assign n2675 = n2674 ^ n1815 ^ 1'b0 ;
  assign n2676 = ( ~n2101 & n2672 ) | ( ~n2101 & n2675 ) | ( n2672 & n2675 ) ;
  assign n2686 = n904 ^ n407 ^ 1'b0 ;
  assign n2687 = n1261 & ~n2686 ;
  assign n2688 = n265 | n2687 ;
  assign n2689 = n2688 ^ x74 ^ 1'b0 ;
  assign n2690 = n2527 & n2689 ;
  assign n2691 = n2690 ^ n1654 ^ 1'b0 ;
  assign n2677 = n135 ^ x32 ^ 1'b0 ;
  assign n2678 = n635 & ~n2677 ;
  assign n2679 = n1688 | n2678 ;
  assign n2680 = n1324 ^ n132 ^ 1'b0 ;
  assign n2681 = n2679 | n2680 ;
  assign n2682 = n189 & n1062 ;
  assign n2683 = n2682 ^ n1800 ^ 1'b0 ;
  assign n2684 = n2681 | n2683 ;
  assign n2685 = x58 & ~n2684 ;
  assign n2692 = n2691 ^ n2685 ^ 1'b0 ;
  assign n2693 = n642 | n953 ;
  assign n2694 = n2600 ^ n790 ^ n215 ;
  assign n2695 = n978 ^ n716 ^ 1'b0 ;
  assign n2696 = ( n536 & n544 ) | ( n536 & ~n1220 ) | ( n544 & ~n1220 ) ;
  assign n2697 = n2696 ^ n1760 ^ x71 ;
  assign n2698 = n2527 & n2697 ;
  assign n2699 = n2698 ^ x126 ^ 1'b0 ;
  assign n2700 = x66 | n1172 ;
  assign n2701 = n2700 ^ n2538 ^ 1'b0 ;
  assign n2702 = x91 & n700 ;
  assign n2703 = ( x120 & ~n1473 ) | ( x120 & n2702 ) | ( ~n1473 & n2702 ) ;
  assign n2705 = n1567 ^ n677 ^ n422 ;
  assign n2704 = n876 | n1949 ;
  assign n2706 = n2705 ^ n2704 ^ 1'b0 ;
  assign n2707 = ~n1172 & n1552 ;
  assign n2708 = n2706 & n2707 ;
  assign n2709 = ~n791 & n1257 ;
  assign n2710 = n2709 ^ n1366 ^ 1'b0 ;
  assign n2711 = x102 ^ x1 ^ 1'b0 ;
  assign n2712 = n683 & ~n2711 ;
  assign n2713 = n1962 | n2712 ;
  assign n2714 = ~n909 & n2713 ;
  assign n2715 = ~n992 & n2714 ;
  assign n2716 = ~n533 & n544 ;
  assign n2717 = n2715 & n2716 ;
  assign n2718 = n415 & ~n1418 ;
  assign n2719 = n2718 ^ n1559 ^ 1'b0 ;
  assign n2720 = n273 | n2010 ;
  assign n2721 = n2720 ^ x106 ^ 1'b0 ;
  assign n2722 = n2721 ^ n1521 ^ 1'b0 ;
  assign n2723 = ~n2719 & n2722 ;
  assign n2724 = ~n961 & n1040 ;
  assign n2725 = n2724 ^ n977 ^ 1'b0 ;
  assign n2726 = n2725 ^ n706 ^ 1'b0 ;
  assign n2727 = ( n319 & n449 ) | ( n319 & ~n1850 ) | ( n449 & ~n1850 ) ;
  assign n2728 = ( n939 & n2254 ) | ( n939 & ~n2727 ) | ( n2254 & ~n2727 ) ;
  assign n2734 = n1100 & ~n2112 ;
  assign n2735 = n2734 ^ n1025 ^ 1'b0 ;
  assign n2732 = n1290 ^ n326 ^ 1'b0 ;
  assign n2733 = n2732 ^ n174 ^ 1'b0 ;
  assign n2736 = n2735 ^ n2733 ^ n588 ;
  assign n2729 = n417 & n560 ;
  assign n2730 = n1948 | n2729 ;
  assign n2731 = n1652 & n2730 ;
  assign n2737 = n2736 ^ n2731 ^ 1'b0 ;
  assign n2738 = n273 | n341 ;
  assign n2739 = n614 & ~n2738 ;
  assign n2740 = n1766 & n2739 ;
  assign n2741 = ~n650 & n1433 ;
  assign n2742 = n1480 ^ n165 ^ 1'b0 ;
  assign n2743 = ~n1929 & n2742 ;
  assign n2744 = n2743 ^ n2594 ^ 1'b0 ;
  assign n2745 = ~n273 & n1594 ;
  assign n2746 = n2745 ^ n413 ^ 1'b0 ;
  assign n2748 = n1054 ^ n308 ^ 1'b0 ;
  assign n2747 = n2498 ^ n1887 ^ n443 ;
  assign n2749 = n2748 ^ n2747 ^ 1'b0 ;
  assign n2750 = x16 | n2479 ;
  assign n2751 = ( x52 & ~n435 ) | ( x52 & n2750 ) | ( ~n435 & n2750 ) ;
  assign n2752 = n840 & ~n2252 ;
  assign n2755 = n429 & n1116 ;
  assign n2756 = ~n980 & n2755 ;
  assign n2753 = ~n179 & n1312 ;
  assign n2754 = ~n2098 & n2753 ;
  assign n2757 = n2756 ^ n2754 ^ 1'b0 ;
  assign n2758 = x68 & ~n2757 ;
  assign n2759 = n2732 ^ n1537 ^ 1'b0 ;
  assign n2760 = n370 & ~n521 ;
  assign n2761 = ( ~n1295 & n1449 ) | ( ~n1295 & n1730 ) | ( n1449 & n1730 ) ;
  assign n2764 = n1130 ^ n396 ^ 1'b0 ;
  assign n2765 = n1329 | n2764 ;
  assign n2762 = n1913 ^ n1321 ^ n651 ;
  assign n2763 = x118 & n2762 ;
  assign n2766 = n2765 ^ n2763 ^ 1'b0 ;
  assign n2767 = n1752 & ~n2766 ;
  assign n2768 = n229 & n285 ;
  assign n2769 = n827 | n2768 ;
  assign n2770 = n612 & ~n2769 ;
  assign n2771 = n973 ^ n663 ^ 1'b0 ;
  assign n2772 = n2758 & ~n2771 ;
  assign n2776 = ~n254 & n619 ;
  assign n2777 = ~n813 & n2776 ;
  assign n2773 = n1684 | n2051 ;
  assign n2774 = n1583 & ~n2773 ;
  assign n2775 = n1832 & ~n2774 ;
  assign n2778 = n2777 ^ n2775 ^ 1'b0 ;
  assign n2779 = n1851 & ~n2778 ;
  assign n2780 = n2779 ^ n1182 ^ n872 ;
  assign n2781 = ~n379 & n1675 ;
  assign n2782 = n469 & n2781 ;
  assign n2783 = n151 & ~n811 ;
  assign n2784 = n2783 ^ x76 ^ 1'b0 ;
  assign n2785 = n2782 | n2784 ;
  assign n2786 = n345 & ~n1143 ;
  assign n2787 = x67 | n1955 ;
  assign n2788 = n2712 & n2760 ;
  assign n2789 = ( n416 & n1409 ) | ( n416 & ~n1670 ) | ( n1409 & ~n1670 ) ;
  assign n2790 = ~n2450 & n2789 ;
  assign n2791 = n2790 ^ n1649 ^ n618 ;
  assign n2792 = n549 & n2175 ;
  assign n2793 = n2791 & n2792 ;
  assign n2795 = n603 ^ n306 ^ 1'b0 ;
  assign n2794 = ~n945 & n1062 ;
  assign n2796 = n2795 ^ n2794 ^ 1'b0 ;
  assign n2797 = n1330 & n2796 ;
  assign n2798 = n576 & n2797 ;
  assign n2799 = n199 | n2798 ;
  assign n2800 = n2799 ^ n1846 ^ 1'b0 ;
  assign n2801 = ~n2030 & n2800 ;
  assign n2802 = n1821 ^ n210 ^ 1'b0 ;
  assign n2803 = n449 ^ x16 ^ 1'b0 ;
  assign n2804 = ~n2802 & n2803 ;
  assign n2805 = n2048 & n2428 ;
  assign n2806 = n844 & ~n2199 ;
  assign n2807 = n485 & n654 ;
  assign n2808 = n1147 ^ n620 ^ 1'b0 ;
  assign n2809 = ~n2807 & n2808 ;
  assign n2810 = n1752 ^ n997 ^ 1'b0 ;
  assign n2811 = n2810 ^ n2085 ^ 1'b0 ;
  assign n2813 = n2479 ^ n1056 ^ 1'b0 ;
  assign n2814 = n1163 | n2813 ;
  assign n2812 = n738 & n1630 ;
  assign n2815 = n2814 ^ n2812 ^ n2426 ;
  assign n2816 = n408 & n2154 ;
  assign n2817 = ~n892 & n2816 ;
  assign n2818 = n530 ^ n150 ^ 1'b0 ;
  assign n2819 = n2818 ^ n1765 ^ n1246 ;
  assign n2820 = ~n2817 & n2819 ;
  assign n2821 = n2820 ^ n1079 ^ 1'b0 ;
  assign n2822 = n1485 ^ x103 ^ 1'b0 ;
  assign n2823 = ~n2092 & n2822 ;
  assign n2824 = n2823 ^ n2379 ^ n994 ;
  assign n2825 = n310 ^ x98 ^ 1'b0 ;
  assign n2826 = n614 ^ n359 ^ x0 ;
  assign n2827 = ( n733 & n1621 ) | ( n733 & n2826 ) | ( n1621 & n2826 ) ;
  assign n2828 = ~n2292 & n2827 ;
  assign n2829 = n2828 ^ n1666 ^ 1'b0 ;
  assign n2830 = ( n2462 & ~n2825 ) | ( n2462 & n2829 ) | ( ~n2825 & n2829 ) ;
  assign n2831 = n1946 ^ n1670 ^ 1'b0 ;
  assign n2832 = ~n340 & n907 ;
  assign n2833 = n363 & n2832 ;
  assign n2834 = n1059 | n2833 ;
  assign n2835 = n2834 ^ n1795 ^ 1'b0 ;
  assign n2836 = n562 & ~n1991 ;
  assign n2837 = n2835 & ~n2836 ;
  assign n2838 = n567 ^ n431 ^ 1'b0 ;
  assign n2839 = n2461 & n2838 ;
  assign n2840 = n2839 ^ n2133 ^ 1'b0 ;
  assign n2841 = x40 & n1818 ;
  assign n2842 = n459 ^ n235 ^ 1'b0 ;
  assign n2843 = n718 & ~n2842 ;
  assign n2844 = n910 & ~n2843 ;
  assign n2845 = n1169 | n2844 ;
  assign n2846 = n1995 ^ n174 ^ 1'b0 ;
  assign n2847 = n340 | n2846 ;
  assign n2848 = n1154 & ~n2847 ;
  assign n2849 = n2848 ^ n1205 ^ 1'b0 ;
  assign n2850 = n868 ^ n619 ^ 1'b0 ;
  assign n2851 = n2850 ^ n2060 ^ n1506 ;
  assign n2852 = x52 & ~n2851 ;
  assign n2853 = n1307 ^ n769 ^ n575 ;
  assign n2854 = n1123 & ~n2853 ;
  assign n2855 = n619 & n2854 ;
  assign n2856 = n1305 ^ n957 ^ 1'b0 ;
  assign n2857 = ~n745 & n2856 ;
  assign n2858 = ~n2436 & n2857 ;
  assign n2859 = n1554 ^ n826 ^ 1'b0 ;
  assign n2860 = ~n2014 & n2859 ;
  assign n2861 = n560 & ~n673 ;
  assign n2862 = n2305 & n2861 ;
  assign n2863 = n2862 ^ n447 ^ 1'b0 ;
  assign n2864 = ( n636 & n1385 ) | ( n636 & n2863 ) | ( n1385 & n2863 ) ;
  assign n2865 = n2307 ^ n1633 ^ 1'b0 ;
  assign n2866 = n706 & n2865 ;
  assign n2867 = n1104 & ~n2482 ;
  assign n2868 = n2867 ^ n1222 ^ 1'b0 ;
  assign n2869 = n2450 ^ n1479 ^ 1'b0 ;
  assign n2870 = ~n254 & n2869 ;
  assign n2871 = n1835 | n1922 ;
  assign n2872 = n369 | n562 ;
  assign n2873 = n1471 | n2872 ;
  assign n2874 = n654 & n2873 ;
  assign n2875 = n2874 ^ n1448 ^ 1'b0 ;
  assign n2877 = ~n381 & n2104 ;
  assign n2876 = n582 & ~n1418 ;
  assign n2878 = n2877 ^ n2876 ^ 1'b0 ;
  assign n2879 = ~n2812 & n2878 ;
  assign n2880 = n2532 & n2879 ;
  assign n2881 = n875 & ~n2768 ;
  assign n2882 = ~n517 & n2881 ;
  assign n2883 = n954 | n1051 ;
  assign n2884 = n1990 | n2785 ;
  assign n2885 = n2884 ^ n567 ^ 1'b0 ;
  assign n2889 = n2195 ^ n615 ^ 1'b0 ;
  assign n2890 = n186 | n2889 ;
  assign n2886 = n1189 | n1765 ;
  assign n2887 = n2886 ^ n1401 ^ 1'b0 ;
  assign n2888 = n1693 & ~n2887 ;
  assign n2891 = n2890 ^ n2888 ^ 1'b0 ;
  assign n2892 = x41 & n2891 ;
  assign n2893 = n1718 ^ n1375 ^ 1'b0 ;
  assign n2894 = n1197 | n2893 ;
  assign n2895 = n640 ^ n628 ^ 1'b0 ;
  assign n2896 = x66 & n2895 ;
  assign n2897 = n681 ^ n153 ^ x64 ;
  assign n2898 = n2897 ^ n231 ^ 1'b0 ;
  assign n2899 = n457 & ~n2898 ;
  assign n2900 = ~n2896 & n2899 ;
  assign n2901 = n1147 | n1234 ;
  assign n2902 = n395 & n2901 ;
  assign n2903 = n2900 & n2902 ;
  assign n2904 = n1686 & ~n1753 ;
  assign n2905 = ~n403 & n2904 ;
  assign n2906 = ( ~n1479 & n2226 ) | ( ~n1479 & n2905 ) | ( n2226 & n2905 ) ;
  assign n2907 = n2906 ^ n1858 ^ n1509 ;
  assign n2908 = ~n169 & n1582 ;
  assign n2909 = n1220 & ~n2908 ;
  assign n2910 = n1061 & n1471 ;
  assign n2911 = ~n166 & n801 ;
  assign n2912 = ~n630 & n2911 ;
  assign n2913 = n2912 ^ n2652 ^ 1'b0 ;
  assign n2914 = n2910 & n2913 ;
  assign n2915 = n631 | n1687 ;
  assign n2916 = n606 | n1033 ;
  assign n2917 = n532 & ~n2916 ;
  assign n2918 = n2289 ^ n1888 ^ n1056 ;
  assign n2919 = n1991 | n2918 ;
  assign n2920 = n2917 & ~n2919 ;
  assign n2921 = ( n1004 & n2415 ) | ( n1004 & ~n2920 ) | ( n2415 & ~n2920 ) ;
  assign n2922 = n1234 ^ n730 ^ 1'b0 ;
  assign n2923 = n2855 ^ n236 ^ 1'b0 ;
  assign n2924 = ( x36 & n262 ) | ( x36 & ~n1566 ) | ( n262 & ~n1566 ) ;
  assign n2925 = ~n349 & n1980 ;
  assign n2926 = ( ~x30 & x68 ) | ( ~x30 & n1218 ) | ( x68 & n1218 ) ;
  assign n2927 = n930 ^ n918 ^ 1'b0 ;
  assign n2928 = n141 | n2927 ;
  assign n2929 = n2033 ^ n1669 ^ x64 ;
  assign n2930 = ( n1378 & ~n2386 ) | ( n1378 & n2403 ) | ( ~n2386 & n2403 ) ;
  assign n2931 = n884 | n1106 ;
  assign n2932 = n2931 ^ n1494 ^ 1'b0 ;
  assign n2933 = ( ~n1375 & n2432 ) | ( ~n1375 & n2932 ) | ( n2432 & n2932 ) ;
  assign n2934 = ( ~n2172 & n2865 ) | ( ~n2172 & n2933 ) | ( n2865 & n2933 ) ;
  assign n2935 = n2055 | n2721 ;
  assign n2936 = n1867 ^ n978 ^ 1'b0 ;
  assign n2937 = n2462 & ~n2936 ;
  assign n2938 = n1051 & n2937 ;
  assign n2939 = n2938 ^ n808 ^ 1'b0 ;
  assign n2940 = n1335 & n2939 ;
  assign n2941 = n964 & ~n1013 ;
  assign n2942 = n2941 ^ n492 ^ 1'b0 ;
  assign n2943 = ~n2612 & n2800 ;
  assign n2944 = n2942 & n2943 ;
  assign n2945 = n1972 ^ n694 ^ n308 ;
  assign n2946 = n297 & n2945 ;
  assign n2947 = n2946 ^ n1721 ^ 1'b0 ;
  assign n2948 = n308 & n1938 ;
  assign n2949 = n2948 ^ n1195 ^ 1'b0 ;
  assign n2950 = n791 | n2441 ;
  assign n2951 = n2950 ^ n1561 ^ 1'b0 ;
  assign n2952 = n1684 ^ n1120 ^ n565 ;
  assign n2953 = n1449 | n2345 ;
  assign n2954 = ~n422 & n2953 ;
  assign n2955 = n1979 ^ n261 ^ 1'b0 ;
  assign n2956 = n625 | n2955 ;
  assign n2957 = n1347 & ~n2956 ;
  assign n2958 = n1230 ^ n742 ^ 1'b0 ;
  assign n2959 = n2958 ^ n811 ^ n654 ;
  assign n2960 = ~n555 & n2959 ;
  assign n2961 = n2957 & n2960 ;
  assign n2962 = n944 & n2414 ;
  assign n2964 = n336 ^ x33 ^ 1'b0 ;
  assign n2965 = n990 & ~n2964 ;
  assign n2963 = n262 & ~n785 ;
  assign n2966 = n2965 ^ n2963 ^ 1'b0 ;
  assign n2967 = ~n2962 & n2966 ;
  assign n2968 = n2128 & n2967 ;
  assign n2969 = n1503 ^ n1445 ^ 1'b0 ;
  assign n2970 = ~n893 & n1499 ;
  assign n2971 = n859 | n1209 ;
  assign n2972 = n2970 & ~n2971 ;
  assign n2973 = n642 ^ x107 ^ 1'b0 ;
  assign n2974 = n2038 & n2973 ;
  assign n2975 = n2974 ^ n1070 ^ 1'b0 ;
  assign n2976 = n2972 | n2975 ;
  assign n2977 = n980 & n1159 ;
  assign n2978 = n2977 ^ n191 ^ 1'b0 ;
  assign n2979 = n2978 ^ n2057 ^ 1'b0 ;
  assign n2984 = n623 ^ n267 ^ 1'b0 ;
  assign n2985 = n143 & n2984 ;
  assign n2986 = x64 & n2687 ;
  assign n2987 = ~n2985 & n2986 ;
  assign n2980 = n454 | n1511 ;
  assign n2981 = ( n696 & ~n1242 ) | ( n696 & n2980 ) | ( ~n1242 & n2980 ) ;
  assign n2982 = n383 & ~n1090 ;
  assign n2983 = ~n2981 & n2982 ;
  assign n2988 = n2987 ^ n2983 ^ 1'b0 ;
  assign n2989 = n2388 ^ n1461 ^ 1'b0 ;
  assign n2990 = n1967 & ~n2989 ;
  assign n2991 = n2990 ^ n2562 ^ 1'b0 ;
  assign n2992 = n487 | n2991 ;
  assign n2993 = x98 & n1266 ;
  assign n2994 = ~n592 & n2993 ;
  assign n2995 = ~n2333 & n2527 ;
  assign n2996 = n2994 & n2995 ;
  assign n2997 = n2992 & ~n2996 ;
  assign n2998 = ~n290 & n1086 ;
  assign n2999 = n2998 ^ n1476 ^ 1'b0 ;
  assign n3000 = x8 & ~n194 ;
  assign n3001 = ~n824 & n3000 ;
  assign n3002 = n764 & ~n3001 ;
  assign n3003 = n3002 ^ n1654 ^ 1'b0 ;
  assign n3004 = n3003 ^ n2401 ^ 1'b0 ;
  assign n3005 = n1950 & n3004 ;
  assign n3006 = ~n169 & n2540 ;
  assign n3007 = n252 & ~n1451 ;
  assign n3008 = ~n3006 & n3007 ;
  assign n3009 = n3008 ^ n2677 ^ 1'b0 ;
  assign n3010 = n2408 ^ n893 ^ 1'b0 ;
  assign n3011 = n3010 ^ n2996 ^ 1'b0 ;
  assign n3012 = n2001 ^ n293 ^ n142 ;
  assign n3013 = n891 | n3012 ;
  assign n3014 = n932 & ~n3013 ;
  assign n3015 = n2634 ^ n1195 ^ n363 ;
  assign n3016 = n306 | n3015 ;
  assign n3017 = n3016 ^ n2538 ^ 1'b0 ;
  assign n3018 = n2178 ^ n456 ^ 1'b0 ;
  assign n3019 = n1239 & ~n3018 ;
  assign n3020 = n929 ^ n420 ^ 1'b0 ;
  assign n3021 = n3020 ^ n1215 ^ 1'b0 ;
  assign n3022 = ( x62 & ~n891 ) | ( x62 & n3021 ) | ( ~n891 & n3021 ) ;
  assign n3023 = n3022 ^ n725 ^ 1'b0 ;
  assign n3024 = n3023 ^ n2591 ^ 1'b0 ;
  assign n3025 = ( n621 & n731 ) | ( n621 & n2027 ) | ( n731 & n2027 ) ;
  assign n3026 = n3025 ^ n1938 ^ n1854 ;
  assign n3027 = n262 | n2280 ;
  assign n3028 = n1408 ^ n1079 ^ n1009 ;
  assign n3029 = ~n1133 & n1584 ;
  assign n3030 = ~n3028 & n3029 ;
  assign n3031 = n1537 | n3030 ;
  assign n3032 = n671 & n2866 ;
  assign n3033 = ~n1892 & n3032 ;
  assign n3034 = n769 | n1261 ;
  assign n3035 = n3034 ^ n2800 ^ n683 ;
  assign n3036 = ~x11 & x54 ;
  assign n3037 = n1001 & n2498 ;
  assign n3038 = n3037 ^ x3 ^ 1'b0 ;
  assign n3039 = n3038 ^ n389 ^ 1'b0 ;
  assign n3040 = n3036 & n3039 ;
  assign n3041 = ~n2599 & n3040 ;
  assign n3042 = n1700 ^ n978 ^ 1'b0 ;
  assign n3043 = ~n1603 & n3042 ;
  assign n3044 = n969 ^ n934 ^ n576 ;
  assign n3045 = n3044 ^ n2864 ^ 1'b0 ;
  assign n3046 = n3043 & ~n3045 ;
  assign n3047 = n2467 ^ n1198 ^ 1'b0 ;
  assign n3048 = ( x2 & x42 ) | ( x2 & ~n3047 ) | ( x42 & ~n3047 ) ;
  assign n3049 = n1788 & n3048 ;
  assign n3050 = n151 & n3049 ;
  assign n3051 = n813 ^ n323 ^ 1'b0 ;
  assign n3052 = n350 | n760 ;
  assign n3053 = n3052 ^ n399 ^ 1'b0 ;
  assign n3054 = n486 | n3053 ;
  assign n3055 = n1030 | n3054 ;
  assign n3056 = n388 & ~n2276 ;
  assign n3057 = n3024 ^ n177 ^ 1'b0 ;
  assign n3058 = ~n616 & n1576 ;
  assign n3059 = ~n2547 & n3058 ;
  assign n3060 = n2083 ^ n2015 ^ 1'b0 ;
  assign n3061 = n3059 & n3060 ;
  assign n3062 = n487 & ~n1269 ;
  assign n3063 = ( n2388 & ~n2608 ) | ( n2388 & n2684 ) | ( ~n2608 & n2684 ) ;
  assign n3066 = n484 ^ x7 ^ 1'b0 ;
  assign n3064 = n763 ^ n470 ^ 1'b0 ;
  assign n3065 = n1130 & n3064 ;
  assign n3067 = n3066 ^ n3065 ^ n508 ;
  assign n3068 = n3067 ^ n1764 ^ 1'b0 ;
  assign n3069 = n3063 & n3068 ;
  assign n3070 = n3069 ^ n1397 ^ 1'b0 ;
  assign n3071 = n161 & ~n2346 ;
  assign n3072 = n2417 ^ n2023 ^ 1'b0 ;
  assign n3073 = n2531 | n3072 ;
  assign n3076 = n859 ^ n381 ^ 1'b0 ;
  assign n3074 = n906 & ~n1471 ;
  assign n3075 = ~n3037 & n3074 ;
  assign n3077 = n3076 ^ n3075 ^ 1'b0 ;
  assign n3078 = n2217 ^ n1583 ^ 1'b0 ;
  assign n3079 = n308 & n3078 ;
  assign n3080 = n2490 & n2725 ;
  assign n3082 = ( ~n1376 & n2248 ) | ( ~n1376 & n2918 ) | ( n2248 & n2918 ) ;
  assign n3081 = n1390 & n2826 ;
  assign n3083 = n3082 ^ n3081 ^ 1'b0 ;
  assign n3084 = n2000 | n2597 ;
  assign n3085 = n1746 ^ n231 ^ 1'b0 ;
  assign n3086 = n473 | n3085 ;
  assign n3087 = n654 | n3086 ;
  assign n3088 = n1587 & n2246 ;
  assign n3089 = n3088 ^ n161 ^ 1'b0 ;
  assign n3090 = n3089 ^ n1927 ^ 1'b0 ;
  assign n3091 = n1627 & ~n3090 ;
  assign n3092 = n3091 ^ n794 ^ 1'b0 ;
  assign n3093 = n3087 & ~n3092 ;
  assign n3094 = n2018 & n3093 ;
  assign n3095 = ~n1722 & n3094 ;
  assign n3096 = n3095 ^ n886 ^ x98 ;
  assign n3097 = n1954 ^ x44 ^ 1'b0 ;
  assign n3098 = n2608 | n3097 ;
  assign n3099 = n962 & ~n2449 ;
  assign n3100 = n3098 & n3099 ;
  assign n3101 = n2932 ^ n323 ^ 1'b0 ;
  assign n3102 = n2035 & ~n3101 ;
  assign n3103 = x2 & ~n3102 ;
  assign n3104 = ( n1229 & ~n1713 ) | ( n1229 & n2173 ) | ( ~n1713 & n2173 ) ;
  assign n3105 = n3104 ^ n156 ^ 1'b0 ;
  assign n3106 = x16 | n2022 ;
  assign n3107 = n310 & ~n3106 ;
  assign n3108 = n2496 & n2703 ;
  assign n3109 = ( n934 & n2254 ) | ( n934 & n3108 ) | ( n2254 & n3108 ) ;
  assign n3110 = n1031 ^ n355 ^ n350 ;
  assign n3111 = n940 & n3110 ;
  assign n3112 = n918 & ~n3111 ;
  assign n3113 = n3112 ^ n267 ^ 1'b0 ;
  assign n3114 = n2302 & n3113 ;
  assign n3115 = n781 & n2875 ;
  assign n3116 = n3115 ^ n1159 ^ 1'b0 ;
  assign n3117 = n986 & n1897 ;
  assign n3118 = ~n186 & n964 ;
  assign n3119 = ~n2519 & n3118 ;
  assign n3120 = n487 ^ x14 ^ 1'b0 ;
  assign n3121 = x13 | n3120 ;
  assign n3122 = n518 | n635 ;
  assign n3123 = n3122 ^ x40 ^ 1'b0 ;
  assign n3124 = n3123 ^ n713 ^ 1'b0 ;
  assign n3125 = n3124 ^ n2022 ^ 1'b0 ;
  assign n3126 = ( n1582 & n3121 ) | ( n1582 & n3125 ) | ( n3121 & n3125 ) ;
  assign n3127 = n796 | n997 ;
  assign n3128 = n512 & ~n2798 ;
  assign n3129 = n3128 ^ n199 ^ 1'b0 ;
  assign n3130 = n3127 & n3129 ;
  assign n3131 = n2216 & ~n2673 ;
  assign n3132 = n3131 ^ n1730 ^ 1'b0 ;
  assign n3133 = n1059 ^ n716 ^ 1'b0 ;
  assign n3134 = n3059 & ~n3133 ;
  assign n3135 = ( ~x121 & n2285 ) | ( ~x121 & n3134 ) | ( n2285 & n3134 ) ;
  assign n3136 = n786 ^ x66 ^ 1'b0 ;
  assign n3137 = n482 & ~n3136 ;
  assign n3138 = n2748 & n3137 ;
  assign n3139 = n3138 ^ x100 ^ 1'b0 ;
  assign n3140 = n2978 & n3139 ;
  assign n3141 = n674 & ~n1576 ;
  assign n3142 = n3141 ^ n1166 ^ 1'b0 ;
  assign n3143 = n1337 | n3142 ;
  assign n3144 = n1711 & n1941 ;
  assign n3145 = n3144 ^ n1971 ^ 1'b0 ;
  assign n3146 = ~n1570 & n3145 ;
  assign n3147 = n601 & n3146 ;
  assign n3148 = n326 | n2706 ;
  assign n3149 = ~n295 & n1229 ;
  assign n3150 = ~n2371 & n3149 ;
  assign n3151 = n3150 ^ n1034 ^ 1'b0 ;
  assign n3152 = ( n2954 & n3148 ) | ( n2954 & ~n3151 ) | ( n3148 & ~n3151 ) ;
  assign n3153 = n3087 ^ n2696 ^ n1959 ;
  assign n3154 = n1236 & ~n2146 ;
  assign n3155 = n2043 & n3154 ;
  assign n3156 = ( n1307 & n3153 ) | ( n1307 & ~n3155 ) | ( n3153 & ~n3155 ) ;
  assign n3157 = n508 | n3156 ;
  assign n3158 = n1175 ^ n245 ^ x17 ;
  assign n3159 = n204 | n1706 ;
  assign n3160 = ~n3158 & n3159 ;
  assign n3161 = n3160 ^ n346 ^ 1'b0 ;
  assign n3162 = n191 & n602 ;
  assign n3163 = n895 & n3162 ;
  assign n3164 = n1273 | n2371 ;
  assign n3165 = n3164 ^ n515 ^ 1'b0 ;
  assign n3166 = n2356 ^ n1413 ^ n322 ;
  assign n3167 = ( n487 & ~n1390 ) | ( n487 & n2473 ) | ( ~n1390 & n2473 ) ;
  assign n3168 = n1667 | n3167 ;
  assign n3169 = n177 & ~n3168 ;
  assign n3170 = n844 | n1810 ;
  assign n3171 = n2661 & n3170 ;
  assign n3172 = n561 & ~n1499 ;
  assign n3173 = n947 & n1189 ;
  assign n3174 = n507 & n519 ;
  assign n3175 = n2618 & n3174 ;
  assign n3176 = n1761 ^ n548 ^ 1'b0 ;
  assign n3178 = n2341 ^ n247 ^ 1'b0 ;
  assign n3177 = n208 & ~n1038 ;
  assign n3179 = n3178 ^ n3177 ^ 1'b0 ;
  assign n3180 = n2357 ^ n1418 ^ 1'b0 ;
  assign n3181 = n1364 & ~n3180 ;
  assign n3183 = n1027 ^ n503 ^ 1'b0 ;
  assign n3184 = n276 & n3183 ;
  assign n3185 = ( ~n1143 & n1842 ) | ( ~n1143 & n3184 ) | ( n1842 & n3184 ) ;
  assign n3182 = n2932 ^ n678 ^ 1'b0 ;
  assign n3186 = n3185 ^ n3182 ^ 1'b0 ;
  assign n3187 = n3027 | n3186 ;
  assign n3188 = n1805 & ~n3187 ;
  assign n3189 = n2001 ^ n959 ^ n134 ;
  assign n3190 = n1860 & n3189 ;
  assign n3191 = n3190 ^ n248 ^ 1'b0 ;
  assign n3192 = n241 & ~n335 ;
  assign n3193 = ~n2859 & n3192 ;
  assign n3194 = n3193 ^ n2636 ^ 1'b0 ;
  assign n3195 = ~n2157 & n3194 ;
  assign n3196 = n3195 ^ n1519 ^ 1'b0 ;
  assign n3197 = n858 & ~n3196 ;
  assign n3198 = n3197 ^ n2431 ^ 1'b0 ;
  assign n3199 = ( n812 & n906 ) | ( n812 & ~n1940 ) | ( n906 & ~n1940 ) ;
  assign n3200 = n494 & n671 ;
  assign n3201 = ~n3199 & n3200 ;
  assign n3202 = n2699 & n3201 ;
  assign n3203 = n346 ^ n214 ^ 1'b0 ;
  assign n3204 = n2032 & ~n3203 ;
  assign n3205 = n868 ^ n379 ^ 1'b0 ;
  assign n3206 = n3205 ^ n1954 ^ 1'b0 ;
  assign n3207 = ~n350 & n646 ;
  assign n3208 = n3207 ^ n505 ^ 1'b0 ;
  assign n3209 = ~n769 & n3208 ;
  assign n3210 = ( n2793 & ~n3165 ) | ( n2793 & n3209 ) | ( ~n3165 & n3209 ) ;
  assign n3211 = n2631 ^ n2109 ^ 1'b0 ;
  assign n3212 = n2323 ^ n2253 ^ 1'b0 ;
  assign n3213 = ( n876 & ~n3172 ) | ( n876 & n3212 ) | ( ~n3172 & n3212 ) ;
  assign n3214 = n1819 & ~n3124 ;
  assign n3215 = n1677 ^ n977 ^ 1'b0 ;
  assign n3216 = n3214 & n3215 ;
  assign n3217 = n619 | n1276 ;
  assign n3218 = n130 & ~n2135 ;
  assign n3219 = n1490 & n3218 ;
  assign n3220 = n3219 ^ n479 ^ 1'b0 ;
  assign n3221 = ~n2413 & n3220 ;
  assign n3222 = n275 ^ x29 ^ 1'b0 ;
  assign n3223 = x12 & ~n3222 ;
  assign n3224 = n3223 ^ n1655 ^ 1'b0 ;
  assign n3225 = n1067 ^ n845 ^ 1'b0 ;
  assign n3226 = n3224 | n3225 ;
  assign n3227 = n2625 | n3226 ;
  assign n3228 = n756 & ~n3227 ;
  assign n3229 = n420 & ~n1771 ;
  assign n3230 = n3229 ^ n2406 ^ n783 ;
  assign n3231 = ~n1012 & n3230 ;
  assign n3232 = n2663 & n3231 ;
  assign n3233 = n2335 & ~n2811 ;
  assign n3234 = ~x72 & n3233 ;
  assign n3235 = n2101 ^ n190 ^ 1'b0 ;
  assign n3236 = ( n644 & n1448 ) | ( n644 & n2223 ) | ( n1448 & n2223 ) ;
  assign n3237 = n2264 | n3236 ;
  assign n3238 = n3235 | n3237 ;
  assign n3239 = n3234 & ~n3238 ;
  assign n3240 = ~n570 & n1913 ;
  assign n3241 = n1004 | n2225 ;
  assign n3242 = n3240 | n3241 ;
  assign n3243 = ( n729 & n773 ) | ( n729 & n3242 ) | ( n773 & n3242 ) ;
  assign n3244 = ( n1418 & n2798 ) | ( n1418 & ~n2853 ) | ( n2798 & ~n2853 ) ;
  assign n3245 = n3244 ^ n2048 ^ 1'b0 ;
  assign n3246 = x49 & ~n791 ;
  assign n3247 = ~n1088 & n3246 ;
  assign n3248 = n3158 | n3203 ;
  assign n3249 = n3247 & ~n3248 ;
  assign n3250 = ( n1212 & n2471 ) | ( n1212 & n3249 ) | ( n2471 & n3249 ) ;
  assign n3251 = n1067 | n1917 ;
  assign n3252 = n3250 & ~n3251 ;
  assign n3253 = n2070 & ~n2231 ;
  assign n3254 = n938 | n3034 ;
  assign n3255 = ~n2864 & n3254 ;
  assign n3256 = n2603 ^ n2331 ^ n2003 ;
  assign n3257 = ~n1874 & n3256 ;
  assign n3258 = ~n2329 & n3257 ;
  assign n3263 = n1116 ^ n171 ^ 1'b0 ;
  assign n3264 = n1892 & n3263 ;
  assign n3259 = x58 & n1077 ;
  assign n3260 = ~n849 & n3259 ;
  assign n3261 = n3260 ^ n1511 ^ 1'b0 ;
  assign n3262 = n2875 & n3261 ;
  assign n3265 = n3264 ^ n3262 ^ 1'b0 ;
  assign n3266 = ( ~n510 & n1330 ) | ( ~n510 & n2206 ) | ( n1330 & n2206 ) ;
  assign n3267 = n1808 ^ n1684 ^ 1'b0 ;
  assign n3268 = n3126 ^ n2574 ^ n812 ;
  assign n3269 = n216 ^ x28 ^ 1'b0 ;
  assign n3270 = n3269 ^ n697 ^ 1'b0 ;
  assign n3271 = n323 & ~n2092 ;
  assign n3272 = n842 & n3271 ;
  assign n3273 = n2758 & ~n3272 ;
  assign n3274 = n3273 ^ n1405 ^ 1'b0 ;
  assign n3275 = x58 & ~n582 ;
  assign n3276 = ( n939 & n1238 ) | ( n939 & n1603 ) | ( n1238 & n1603 ) ;
  assign n3277 = n380 & n3276 ;
  assign n3278 = n1271 ^ x17 ^ 1'b0 ;
  assign n3279 = n3277 & n3278 ;
  assign n3285 = n651 ^ n149 ^ 1'b0 ;
  assign n3280 = n1084 & ~n3066 ;
  assign n3281 = n3280 ^ n1692 ^ 1'b0 ;
  assign n3282 = n956 & n3281 ;
  assign n3283 = n3208 ^ n261 ^ 1'b0 ;
  assign n3284 = n3282 & ~n3283 ;
  assign n3286 = n3285 ^ n3284 ^ 1'b0 ;
  assign n3287 = n1732 ^ n828 ^ x6 ;
  assign n3288 = x12 | n1994 ;
  assign n3289 = n2219 ^ n2055 ^ 1'b0 ;
  assign n3290 = n2001 ^ n1976 ^ 1'b0 ;
  assign n3291 = ( x23 & n1323 ) | ( x23 & n3290 ) | ( n1323 & n3290 ) ;
  assign n3292 = n1045 | n3291 ;
  assign n3293 = n1855 | n3292 ;
  assign n3294 = n1539 & ~n3293 ;
  assign n3296 = ~n442 & n2514 ;
  assign n3297 = n3296 ^ n2462 ^ n1461 ;
  assign n3295 = n967 & ~n2956 ;
  assign n3298 = n3297 ^ n3295 ^ 1'b0 ;
  assign n3299 = x80 & ~n2711 ;
  assign n3300 = n2106 & ~n3299 ;
  assign n3301 = n3300 ^ n1347 ^ 1'b0 ;
  assign n3302 = ( n833 & n2620 ) | ( n833 & n3301 ) | ( n2620 & n3301 ) ;
  assign n3303 = n376 & n1197 ;
  assign n3304 = n909 & n3303 ;
  assign n3306 = n2938 ^ n2451 ^ 1'b0 ;
  assign n3305 = x32 & ~n1656 ;
  assign n3307 = n3306 ^ n3305 ^ 1'b0 ;
  assign n3308 = n2735 ^ n1703 ^ 1'b0 ;
  assign n3309 = n297 & ~n3308 ;
  assign n3310 = ~n1056 & n3309 ;
  assign n3311 = n2393 ^ n317 ^ 1'b0 ;
  assign n3312 = n612 & ~n3311 ;
  assign n3314 = n1743 ^ n498 ^ 1'b0 ;
  assign n3315 = ~n642 & n3314 ;
  assign n3316 = n3315 ^ n1122 ^ n227 ;
  assign n3313 = n696 & ~n832 ;
  assign n3317 = n3316 ^ n3313 ^ 1'b0 ;
  assign n3318 = ~n2027 & n2566 ;
  assign n3319 = n3318 ^ x46 ^ 1'b0 ;
  assign n3320 = n961 | n2777 ;
  assign n3321 = ~x58 & n276 ;
  assign n3322 = n2329 & ~n3321 ;
  assign n3323 = n3322 ^ n2496 ^ 1'b0 ;
  assign n3324 = n1108 | n1746 ;
  assign n3325 = n3323 & ~n3324 ;
  assign n3326 = n1713 ^ n1387 ^ 1'b0 ;
  assign n3327 = n1154 & ~n2791 ;
  assign n3328 = ~n3326 & n3327 ;
  assign n3329 = ~n3237 & n3328 ;
  assign n3330 = n2662 ^ x76 ^ 1'b0 ;
  assign n3331 = x84 & ~n411 ;
  assign n3332 = ~n408 & n3331 ;
  assign n3333 = n3332 ^ n956 ^ 1'b0 ;
  assign n3334 = n519 & n3333 ;
  assign n3335 = n2341 & ~n3009 ;
  assign n3336 = n1685 | n3304 ;
  assign n3341 = x45 & ~n494 ;
  assign n3342 = n3341 ^ n1097 ^ 1'b0 ;
  assign n3338 = ~n555 & n783 ;
  assign n3339 = ~n2603 & n3338 ;
  assign n3340 = ~n1809 & n3339 ;
  assign n3343 = n3342 ^ n3340 ^ 1'b0 ;
  assign n3337 = ~n1261 & n1771 ;
  assign n3344 = n3343 ^ n3337 ^ 1'b0 ;
  assign n3345 = n3208 ^ n1366 ^ n1320 ;
  assign n3346 = n194 & ~n3345 ;
  assign n3347 = n443 & n3346 ;
  assign n3348 = n479 & n2873 ;
  assign n3352 = n2166 ^ n1936 ^ 1'b0 ;
  assign n3350 = ~n740 & n1433 ;
  assign n3351 = n3350 ^ n2282 ^ x110 ;
  assign n3349 = n1897 ^ n978 ^ 1'b0 ;
  assign n3353 = n3352 ^ n3351 ^ n3349 ;
  assign n3354 = n223 & n2589 ;
  assign n3355 = ( n1222 & ~n3317 ) | ( n1222 & n3354 ) | ( ~n3317 & n3354 ) ;
  assign n3357 = ( x66 & n479 ) | ( x66 & n1874 ) | ( n479 & n1874 ) ;
  assign n3356 = n690 & n804 ;
  assign n3358 = n3357 ^ n3356 ^ 1'b0 ;
  assign n3359 = n2817 ^ n549 ^ 1'b0 ;
  assign n3360 = ~n891 & n3359 ;
  assign n3361 = ~n1844 & n3360 ;
  assign n3362 = n3361 ^ n2348 ^ n1842 ;
  assign n3363 = n1796 ^ n323 ^ 1'b0 ;
  assign n3364 = n3028 ^ n1740 ^ 1'b0 ;
  assign n3365 = n3363 & n3364 ;
  assign n3366 = n3362 & n3365 ;
  assign n3367 = n1141 & n2222 ;
  assign n3368 = n290 | n377 ;
  assign n3369 = n3368 ^ n1014 ^ 1'b0 ;
  assign n3370 = n343 & n529 ;
  assign n3371 = n3369 & n3370 ;
  assign n3372 = n1977 & n3371 ;
  assign n3373 = n1177 | n1520 ;
  assign n3374 = ( n2326 & ~n2671 ) | ( n2326 & n3373 ) | ( ~n2671 & n3373 ) ;
  assign n3375 = ~n1841 & n3374 ;
  assign n3376 = n3375 ^ n692 ^ 1'b0 ;
  assign n3377 = n3376 ^ n2600 ^ 1'b0 ;
  assign n3378 = x3 & x65 ;
  assign n3379 = n3378 ^ n1765 ^ 1'b0 ;
  assign n3380 = n671 & ~n3379 ;
  assign n3381 = n730 | n2157 ;
  assign n3382 = n3259 & ~n3381 ;
  assign n3383 = ( ~n577 & n2085 ) | ( ~n577 & n2517 ) | ( n2085 & n2517 ) ;
  assign n3384 = n1863 ^ n1339 ^ n1231 ;
  assign n3385 = n1828 ^ n889 ^ 1'b0 ;
  assign n3386 = n1457 | n1933 ;
  assign n3387 = n3386 ^ n2795 ^ 1'b0 ;
  assign n3388 = n1175 & ~n2222 ;
  assign n3389 = ~n3387 & n3388 ;
  assign n3390 = n954 & ~n3389 ;
  assign n3391 = n3390 ^ n2142 ^ 1'b0 ;
  assign n3392 = n2166 & ~n3325 ;
  assign n3393 = ~n671 & n3392 ;
  assign n3394 = n872 | n1375 ;
  assign n3395 = n3394 ^ n415 ^ 1'b0 ;
  assign n3399 = n897 ^ x19 ^ 1'b0 ;
  assign n3396 = x119 & n1512 ;
  assign n3397 = n3396 ^ n3324 ^ 1'b0 ;
  assign n3398 = ~n413 & n3397 ;
  assign n3400 = n3399 ^ n3398 ^ 1'b0 ;
  assign n3401 = n2120 | n3400 ;
  assign n3402 = n1080 & ~n1312 ;
  assign n3403 = n3048 ^ n1271 ^ n691 ;
  assign n3404 = n3403 ^ n2818 ^ 1'b0 ;
  assign n3405 = n1472 ^ n997 ^ 1'b0 ;
  assign n3406 = n241 & n3405 ;
  assign n3407 = n3290 ^ n707 ^ 1'b0 ;
  assign n3408 = n3406 & n3407 ;
  assign n3409 = ( n359 & ~n623 ) | ( n359 & n3175 ) | ( ~n623 & n3175 ) ;
  assign n3410 = n1472 & ~n2073 ;
  assign n3411 = ~n280 & n3410 ;
  assign n3414 = n214 ^ x102 ^ 1'b0 ;
  assign n3413 = n1277 ^ n346 ^ 1'b0 ;
  assign n3412 = n1013 ^ n1000 ^ 1'b0 ;
  assign n3415 = n3414 ^ n3413 ^ n3412 ;
  assign n3416 = n3415 ^ n517 ^ 1'b0 ;
  assign n3417 = ~n3411 & n3416 ;
  assign n3418 = n1192 & ~n3409 ;
  assign n3419 = n1023 ^ n668 ^ 1'b0 ;
  assign n3420 = n3205 ^ n2003 ^ 1'b0 ;
  assign n3421 = n3420 ^ n442 ^ 1'b0 ;
  assign n3422 = ~n3419 & n3421 ;
  assign n3423 = n352 & ~n2733 ;
  assign n3424 = ~n3422 & n3423 ;
  assign n3425 = x57 & n166 ;
  assign n3426 = n3425 ^ n1680 ^ 1'b0 ;
  assign n3427 = ~n319 & n3426 ;
  assign n3428 = n3427 ^ n2723 ^ 1'b0 ;
  assign n3429 = ( x70 & ~n1545 ) | ( x70 & n3428 ) | ( ~n1545 & n3428 ) ;
  assign n3430 = ~n167 & n383 ;
  assign n3431 = n3429 & n3430 ;
  assign n3432 = n1238 | n2399 ;
  assign n3434 = n3321 ^ n954 ^ x75 ;
  assign n3433 = n516 & ~n1364 ;
  assign n3435 = n3434 ^ n3433 ^ n2334 ;
  assign n3436 = n1550 & ~n1627 ;
  assign n3437 = n1376 ^ n983 ^ 1'b0 ;
  assign n3438 = n243 & ~n3342 ;
  assign n3439 = n3030 ^ n431 ^ 1'b0 ;
  assign n3440 = n2632 ^ n200 ^ 1'b0 ;
  assign n3441 = ~n138 & n3440 ;
  assign n3442 = n3441 ^ n2489 ^ 1'b0 ;
  assign n3443 = n873 & n1561 ;
  assign n3444 = n3443 ^ n3077 ^ 1'b0 ;
  assign n3445 = x54 & n1192 ;
  assign n3446 = ~n216 & n3445 ;
  assign n3447 = ( n1013 & ~n1736 ) | ( n1013 & n1775 ) | ( ~n1736 & n1775 ) ;
  assign n3448 = ( n1886 & ~n2333 ) | ( n1886 & n3447 ) | ( ~n2333 & n3447 ) ;
  assign n3449 = n1171 | n3448 ;
  assign n3450 = n3449 ^ n1095 ^ 1'b0 ;
  assign n3459 = n1664 ^ n881 ^ 1'b0 ;
  assign n3460 = ~n536 & n3459 ;
  assign n3455 = ( n1064 & n1197 ) | ( n1064 & n2216 ) | ( n1197 & n2216 ) ;
  assign n3456 = ( n1856 & n2380 ) | ( n1856 & ~n3455 ) | ( n2380 & ~n3455 ) ;
  assign n3451 = n918 & n1070 ;
  assign n3452 = ~n208 & n3451 ;
  assign n3453 = n621 & ~n3452 ;
  assign n3454 = ~n2957 & n3453 ;
  assign n3457 = n3456 ^ n3454 ^ 1'b0 ;
  assign n3458 = ~n2817 & n3457 ;
  assign n3461 = n3460 ^ n3458 ^ 1'b0 ;
  assign n3462 = n2531 ^ n2376 ^ 1'b0 ;
  assign n3463 = ~n2255 & n3462 ;
  assign n3464 = n3463 ^ n1529 ^ 1'b0 ;
  assign n3465 = n1157 ^ n138 ^ 1'b0 ;
  assign n3466 = n3465 ^ n2506 ^ n341 ;
  assign n3467 = n2293 ^ n478 ^ 1'b0 ;
  assign n3472 = n214 | n651 ;
  assign n3468 = n1358 | n2043 ;
  assign n3469 = n1566 & n3468 ;
  assign n3470 = n1487 & n3469 ;
  assign n3471 = ( n210 & ~n3386 ) | ( n210 & n3470 ) | ( ~n3386 & n3470 ) ;
  assign n3473 = n3472 ^ n3471 ^ 1'b0 ;
  assign n3474 = ~x97 & n3473 ;
  assign n3475 = ~n2732 & n3474 ;
  assign n3476 = n3447 ^ n977 ^ 1'b0 ;
  assign n3477 = n2756 & ~n3476 ;
  assign n3478 = n409 & n3477 ;
  assign n3479 = n273 ^ x116 ^ 1'b0 ;
  assign n3480 = n3479 ^ n3429 ^ 1'b0 ;
  assign n3481 = ~n812 & n3281 ;
  assign n3482 = n3481 ^ n512 ^ 1'b0 ;
  assign n3483 = n3482 ^ n2024 ^ 1'b0 ;
  assign n3484 = n3166 & ~n3483 ;
  assign n3486 = n744 | n2964 ;
  assign n3487 = n3486 ^ n421 ^ 1'b0 ;
  assign n3488 = n703 & ~n3487 ;
  assign n3485 = n2534 ^ x2 ^ 1'b0 ;
  assign n3489 = n3488 ^ n3485 ^ 1'b0 ;
  assign n3490 = n2226 & n3489 ;
  assign n3491 = ~n1100 & n3490 ;
  assign n3492 = n1840 | n2178 ;
  assign n3493 = ~n346 & n3055 ;
  assign n3494 = n3493 ^ n838 ^ 1'b0 ;
  assign n3495 = n3494 ^ x123 ^ 1'b0 ;
  assign n3496 = ~n3492 & n3495 ;
  assign n3497 = ( n145 & n494 ) | ( n145 & n1130 ) | ( n494 & n1130 ) ;
  assign n3498 = n592 ^ x13 ^ 1'b0 ;
  assign n3499 = n3497 & ~n3498 ;
  assign n3500 = n597 & n3499 ;
  assign n3501 = ~n597 & n3500 ;
  assign n3502 = n1061 ^ n343 ^ 1'b0 ;
  assign n3503 = ~n254 & n3502 ;
  assign n3504 = n1072 | n2112 ;
  assign n3505 = n1072 & ~n3504 ;
  assign n3506 = n3503 & ~n3505 ;
  assign n3507 = ~n3503 & n3506 ;
  assign n3508 = n977 | n3507 ;
  assign n3509 = n1809 ^ n1693 ^ 1'b0 ;
  assign n3510 = ( n1269 & n1758 ) | ( n1269 & ~n1796 ) | ( n1758 & ~n1796 ) ;
  assign n3511 = ~n3509 & n3510 ;
  assign n3512 = ( ~n3501 & n3508 ) | ( ~n3501 & n3511 ) | ( n3508 & n3511 ) ;
  assign n3513 = n1416 ^ x12 ^ 1'b0 ;
  assign n3514 = ~n3217 & n3279 ;
  assign n3515 = ~n3513 & n3514 ;
  assign n3517 = x19 & n861 ;
  assign n3518 = ~n1046 & n3517 ;
  assign n3516 = ( x1 & ~n803 ) | ( x1 & n1203 ) | ( ~n803 & n1203 ) ;
  assign n3519 = n3518 ^ n3516 ^ n1481 ;
  assign n3520 = x23 | n850 ;
  assign n3521 = n2033 | n3520 ;
  assign n3522 = ~n1553 & n1578 ;
  assign n3523 = ~n3195 & n3522 ;
  assign n3524 = n1726 & ~n3091 ;
  assign n3525 = ( ~n1435 & n1860 ) | ( ~n1435 & n1959 ) | ( n1860 & n1959 ) ;
  assign n3526 = n2335 & n3525 ;
  assign n3527 = n271 ^ n199 ^ 1'b0 ;
  assign n3528 = n1718 | n3527 ;
  assign n3529 = n2195 ^ n1666 ^ 1'b0 ;
  assign n3530 = n2802 | n3529 ;
  assign n3531 = n3528 & ~n3530 ;
  assign n3532 = ~n1257 & n1698 ;
  assign n3535 = ( n891 & n1379 ) | ( n891 & n3277 ) | ( n1379 & n3277 ) ;
  assign n3533 = n161 | n1888 ;
  assign n3534 = n2349 & ~n3533 ;
  assign n3536 = n3535 ^ n3534 ^ 1'b0 ;
  assign n3537 = n129 & ~n2639 ;
  assign n3538 = ( n314 & n1088 ) | ( n314 & ~n3537 ) | ( n1088 & ~n3537 ) ;
  assign n3539 = n513 & ~n1989 ;
  assign n3540 = n3539 ^ n1565 ^ 1'b0 ;
  assign n3541 = n2200 | n3540 ;
  assign n3542 = n3541 ^ n145 ^ 1'b0 ;
  assign n3543 = n3538 & n3542 ;
  assign n3544 = n3543 ^ n2638 ^ 1'b0 ;
  assign n3545 = n2538 & ~n2622 ;
  assign n3546 = n671 & n3545 ;
  assign n3549 = n419 ^ x48 ^ 1'b0 ;
  assign n3550 = ~n396 & n3549 ;
  assign n3551 = n3550 ^ n1940 ^ x67 ;
  assign n3552 = n3551 ^ n327 ^ 1'b0 ;
  assign n3547 = ( ~x78 & n210 ) | ( ~x78 & n220 ) | ( n210 & n220 ) ;
  assign n3548 = n2258 & ~n3547 ;
  assign n3553 = n3552 ^ n3548 ^ 1'b0 ;
  assign n3556 = n726 ^ n370 ^ 1'b0 ;
  assign n3557 = n2255 ^ n1839 ^ x58 ;
  assign n3558 = ( ~n858 & n3556 ) | ( ~n858 & n3557 ) | ( n3556 & n3557 ) ;
  assign n3554 = n1291 & ~n1619 ;
  assign n3555 = n2740 & n3554 ;
  assign n3559 = n3558 ^ n3555 ^ 1'b0 ;
  assign n3560 = n912 ^ n431 ^ 1'b0 ;
  assign n3561 = n3560 ^ n1588 ^ x71 ;
  assign n3562 = ( n686 & n1809 ) | ( n686 & n3022 ) | ( n1809 & n3022 ) ;
  assign n3563 = n2406 & n3562 ;
  assign n3564 = n3561 & n3563 ;
  assign n3565 = n574 | n3367 ;
  assign n3566 = n3357 ^ n3157 ^ 1'b0 ;
  assign n3567 = n2908 & n3566 ;
  assign n3568 = ~x78 & n653 ;
  assign n3569 = n373 | n3568 ;
  assign n3570 = n1669 & n3569 ;
  assign n3571 = ~n380 & n3570 ;
  assign n3572 = n762 | n1067 ;
  assign n3573 = n957 & ~n3572 ;
  assign n3574 = n3573 ^ n1690 ^ 1'b0 ;
  assign n3575 = n398 & ~n3574 ;
  assign n3579 = n1059 | n1747 ;
  assign n3580 = n3579 ^ n2063 ^ 1'b0 ;
  assign n3576 = n1791 ^ n750 ^ 1'b0 ;
  assign n3577 = n3576 ^ n2198 ^ 1'b0 ;
  assign n3578 = n1619 | n3577 ;
  assign n3581 = n3580 ^ n3578 ^ n3211 ;
  assign n3583 = n473 | n909 ;
  assign n3582 = n2687 ^ n760 ^ 1'b0 ;
  assign n3584 = n3583 ^ n3582 ^ 1'b0 ;
  assign n3585 = n1884 ^ n786 ^ 1'b0 ;
  assign n3589 = n1042 ^ n892 ^ n586 ;
  assign n3587 = ( ~n361 & n1082 ) | ( ~n361 & n2328 ) | ( n1082 & n2328 ) ;
  assign n3588 = n454 & n3587 ;
  assign n3590 = n3589 ^ n3588 ^ 1'b0 ;
  assign n3586 = n1374 ^ n332 ^ 1'b0 ;
  assign n3591 = n3590 ^ n3586 ^ n2317 ;
  assign n3592 = n2252 & n3591 ;
  assign n3593 = ~n2107 & n3592 ;
  assign n3594 = n2433 & ~n3593 ;
  assign n3595 = ~n824 & n1894 ;
  assign n3596 = n3595 ^ n2906 ^ 1'b0 ;
  assign n3597 = n1780 ^ n1512 ^ n636 ;
  assign n3598 = n2146 | n3597 ;
  assign n3599 = n3598 ^ n2958 ^ 1'b0 ;
  assign n3600 = ~n2988 & n3599 ;
  assign n3601 = n236 | n353 ;
  assign n3602 = n3601 ^ n3125 ^ 1'b0 ;
  assign n3603 = ~n1297 & n3602 ;
  assign n3604 = n2845 & n3603 ;
  assign n3616 = ~n791 & n1586 ;
  assign n3617 = n3616 ^ n671 ^ 1'b0 ;
  assign n3605 = n1234 ^ n179 ^ 1'b0 ;
  assign n3608 = n1378 ^ n1284 ^ n1036 ;
  assign n3606 = ~n479 & n863 ;
  assign n3607 = n3606 ^ x4 ^ 1'b0 ;
  assign n3609 = n3608 ^ n3607 ^ n959 ;
  assign n3610 = n3609 ^ n220 ^ 1'b0 ;
  assign n3611 = n3610 ^ n883 ^ 1'b0 ;
  assign n3612 = ~n3605 & n3611 ;
  assign n3613 = ~n1135 & n1413 ;
  assign n3614 = n3613 ^ n2197 ^ 1'b0 ;
  assign n3615 = n3612 & n3614 ;
  assign n3618 = n3617 ^ n3615 ^ 1'b0 ;
  assign n3619 = ~x95 & n3440 ;
  assign n3620 = ( n1463 & ~n1582 ) | ( n1463 & n1893 ) | ( ~n1582 & n1893 ) ;
  assign n3621 = n461 & ~n1484 ;
  assign n3622 = n3620 & n3621 ;
  assign n3623 = x125 & n612 ;
  assign n3624 = ( ~n502 & n1461 ) | ( ~n502 & n3623 ) | ( n1461 & n3623 ) ;
  assign n3625 = n1920 ^ n1854 ^ 1'b0 ;
  assign n3626 = n645 & n1235 ;
  assign n3627 = ~n3424 & n3626 ;
  assign n3628 = n1156 & n3627 ;
  assign n3629 = ~n933 & n2928 ;
  assign n3630 = ~n1741 & n3629 ;
  assign n3631 = n1237 ^ n399 ^ x114 ;
  assign n3632 = n581 | n2696 ;
  assign n3633 = n3632 ^ n1371 ^ 1'b0 ;
  assign n3634 = n3633 ^ n2505 ^ n2239 ;
  assign n3635 = ~n3631 & n3634 ;
  assign n3636 = ~n1600 & n2747 ;
  assign n3637 = n977 | n1562 ;
  assign n3638 = n1031 ^ n671 ^ 1'b0 ;
  assign n3639 = ( n1267 & n1638 ) | ( n1267 & n2985 ) | ( n1638 & n2985 ) ;
  assign n3640 = n2322 ^ n1667 ^ 1'b0 ;
  assign n3641 = n262 & n3640 ;
  assign n3643 = n934 & ~n969 ;
  assign n3642 = n1434 & n3130 ;
  assign n3644 = n3643 ^ n3642 ^ 1'b0 ;
  assign n3645 = n3462 & n3644 ;
  assign n3646 = n3645 ^ n3474 ^ 1'b0 ;
  assign n3647 = n1973 ^ n742 ^ n639 ;
  assign n3648 = n3509 & n3647 ;
  assign n3649 = ( ~n405 & n895 ) | ( ~n405 & n3648 ) | ( n895 & n3648 ) ;
  assign n3650 = n3649 ^ n474 ^ 1'b0 ;
  assign n3651 = ~n1780 & n3650 ;
  assign n3652 = n688 & ~n785 ;
  assign n3653 = n3290 ^ n612 ^ 1'b0 ;
  assign n3654 = n1955 ^ n1345 ^ n260 ;
  assign n3655 = ( n752 & n1684 ) | ( n752 & n3654 ) | ( n1684 & n3654 ) ;
  assign n3656 = n445 & n3153 ;
  assign n3657 = n370 | n3001 ;
  assign n3659 = n487 & n1267 ;
  assign n3660 = n3659 ^ n2271 ^ 1'b0 ;
  assign n3658 = n935 & n1864 ;
  assign n3661 = n3660 ^ n3658 ^ 1'b0 ;
  assign n3662 = n1083 & ~n3661 ;
  assign n3663 = n3657 & n3662 ;
  assign n3664 = ( n605 & ~n840 ) | ( n605 & n2742 ) | ( ~n840 & n2742 ) ;
  assign n3665 = x123 & ~n3664 ;
  assign n3666 = n3665 ^ x52 ^ 1'b0 ;
  assign n3667 = n3533 ^ n2515 ^ 1'b0 ;
  assign n3668 = ~n3666 & n3667 ;
  assign n3669 = n3668 ^ n2888 ^ n712 ;
  assign n3670 = n3515 ^ n869 ^ 1'b0 ;
  assign n3671 = n949 & ~n2835 ;
  assign n3672 = n1226 & n3671 ;
  assign n3673 = ( n1168 & n1479 ) | ( n1168 & ~n2285 ) | ( n1479 & ~n2285 ) ;
  assign n3674 = n1003 & n3673 ;
  assign n3675 = n627 & ~n2610 ;
  assign n3676 = n541 | n1938 ;
  assign n3677 = n1086 | n1506 ;
  assign n3678 = n324 & ~n3677 ;
  assign n3679 = n3678 ^ n1217 ^ 1'b0 ;
  assign n3680 = ( n1477 & n1860 ) | ( n1477 & n3679 ) | ( n1860 & n3679 ) ;
  assign n3681 = ~n2248 & n3680 ;
  assign n3682 = ( ~n499 & n1780 ) | ( ~n499 & n2668 ) | ( n1780 & n2668 ) ;
  assign n3683 = n756 | n3682 ;
  assign n3684 = n1162 | n3683 ;
  assign n3685 = ~n494 & n3684 ;
  assign n3686 = ~n3496 & n3685 ;
  assign n3687 = ( ~x57 & n1675 ) | ( ~x57 & n2829 ) | ( n1675 & n2829 ) ;
  assign n3688 = ( n398 & ~n1267 ) | ( n398 & n1505 ) | ( ~n1267 & n1505 ) ;
  assign n3689 = n3688 ^ n2583 ^ 1'b0 ;
  assign n3690 = ~n1149 & n3689 ;
  assign n3691 = n3690 ^ n2983 ^ 1'b0 ;
  assign n3692 = ~n403 & n3691 ;
  assign n3693 = ~n388 & n3692 ;
  assign n3694 = n1990 & ~n2579 ;
  assign n3695 = ~n558 & n2495 ;
  assign n3696 = n3694 & n3695 ;
  assign n3697 = n1820 | n3696 ;
  assign n3698 = ( n478 & ~n950 ) | ( n478 & n1200 ) | ( ~n950 & n1200 ) ;
  assign n3699 = n3698 ^ n237 ^ 1'b0 ;
  assign n3700 = n946 & n2058 ;
  assign n3701 = n3700 ^ n3633 ^ 1'b0 ;
  assign n3702 = n3240 & ~n3701 ;
  assign n3703 = n1106 ^ x98 ^ 1'b0 ;
  assign n3704 = n519 & ~n3703 ;
  assign n3705 = ~n1670 & n3704 ;
  assign n3706 = n3705 ^ n566 ^ 1'b0 ;
  assign n3707 = n3706 ^ n2789 ^ 1'b0 ;
  assign n3708 = n2290 & n3707 ;
  assign n3709 = ~n1042 & n1858 ;
  assign n3710 = ( n254 & n362 ) | ( n254 & n2814 ) | ( n362 & n2814 ) ;
  assign n3711 = n1683 | n1767 ;
  assign n3712 = n1520 | n3711 ;
  assign n3713 = ~n1971 & n3712 ;
  assign n3714 = n3713 ^ n781 ^ 1'b0 ;
  assign n3715 = n3710 | n3714 ;
  assign n3716 = n3476 & ~n3715 ;
  assign n3717 = n3716 ^ n150 ^ 1'b0 ;
  assign n3718 = x87 & n1229 ;
  assign n3719 = n2647 & ~n3718 ;
  assign n3720 = n3085 ^ n2719 ^ 1'b0 ;
  assign n3721 = n510 & n3720 ;
  assign n3722 = n2041 & n3721 ;
  assign n3723 = n3000 & n3722 ;
  assign n3724 = n1448 ^ n1088 ^ 1'b0 ;
  assign n3725 = n1428 & ~n1545 ;
  assign n3726 = n3725 ^ n2951 ^ 1'b0 ;
  assign n3727 = ~n3696 & n3726 ;
  assign n3728 = n2106 ^ n2003 ^ n1784 ;
  assign n3729 = n2817 ^ n1736 ^ 1'b0 ;
  assign n3730 = n3487 & ~n3729 ;
  assign n3731 = n3730 ^ n1291 ^ 1'b0 ;
  assign n3734 = n586 ^ n380 ^ 1'b0 ;
  assign n3732 = n2353 ^ n1228 ^ 1'b0 ;
  assign n3733 = ~n854 & n3732 ;
  assign n3735 = n3734 ^ n3733 ^ 1'b0 ;
  assign n3736 = n3371 ^ n231 ^ 1'b0 ;
  assign n3737 = n796 & n3736 ;
  assign n3738 = n380 & n3737 ;
  assign n3739 = n3735 | n3738 ;
  assign n3740 = x51 & n2678 ;
  assign n3741 = n1189 ^ n886 ^ 1'b0 ;
  assign n3742 = n939 ^ n273 ^ 1'b0 ;
  assign n3743 = ~n2045 & n3742 ;
  assign n3744 = ~n1166 & n3743 ;
  assign n3745 = n925 ^ n692 ^ 1'b0 ;
  assign n3746 = ~n1113 & n3745 ;
  assign n3747 = n275 | n3746 ;
  assign n3748 = n2112 & n3747 ;
  assign n3749 = ~x48 & n3748 ;
  assign n3750 = n1689 & n2058 ;
  assign n3751 = n3750 ^ n969 ^ 1'b0 ;
  assign n3752 = ~n1765 & n3751 ;
  assign n3753 = n1671 & ~n3752 ;
  assign n3754 = n3192 ^ x52 ^ 1'b0 ;
  assign n3755 = n2777 ^ n1281 ^ 1'b0 ;
  assign n3756 = n3755 ^ n2249 ^ n227 ;
  assign n3757 = n1236 ^ n148 ^ 1'b0 ;
  assign n3758 = ( ~n2104 & n3756 ) | ( ~n2104 & n3757 ) | ( n3756 & n3757 ) ;
  assign n3759 = ( n1219 & n2826 ) | ( n1219 & ~n3001 ) | ( n2826 & ~n3001 ) ;
  assign n3760 = n3759 ^ n474 ^ 1'b0 ;
  assign n3761 = ~n2594 & n2839 ;
  assign n3764 = n2964 ^ n1231 ^ 1'b0 ;
  assign n3765 = n1920 | n3764 ;
  assign n3766 = ~n1288 & n3765 ;
  assign n3767 = ~n478 & n3766 ;
  assign n3762 = ~n1840 & n3751 ;
  assign n3763 = n3762 ^ n2608 ^ 1'b0 ;
  assign n3768 = n3767 ^ n3763 ^ 1'b0 ;
  assign n3772 = n986 ^ n149 ^ 1'b0 ;
  assign n3773 = ~n605 & n3772 ;
  assign n3774 = ~n1654 & n3773 ;
  assign n3775 = n3774 ^ n1432 ^ 1'b0 ;
  assign n3769 = ~n381 & n706 ;
  assign n3770 = n3769 ^ n141 ^ 1'b0 ;
  assign n3771 = n2343 | n3770 ;
  assign n3776 = n3775 ^ n3771 ^ 1'b0 ;
  assign n3777 = ( ~n1219 & n1479 ) | ( ~n1219 & n3440 ) | ( n1479 & n3440 ) ;
  assign n3778 = n3460 ^ n1762 ^ 1'b0 ;
  assign n3779 = n3777 & n3778 ;
  assign n3780 = n2313 & n3779 ;
  assign n3781 = n3780 ^ n586 ^ 1'b0 ;
  assign n3782 = n2376 ^ n794 ^ 1'b0 ;
  assign n3783 = n261 & n3782 ;
  assign n3784 = n2711 & n3783 ;
  assign n3785 = n3784 ^ n422 ^ 1'b0 ;
  assign n3786 = n3785 ^ n3080 ^ 1'b0 ;
  assign n3787 = n1594 & ~n2182 ;
  assign n3788 = n3787 ^ n2070 ^ 1'b0 ;
  assign n3789 = n3788 ^ n3644 ^ 1'b0 ;
  assign n3790 = n3529 ^ n2623 ^ 1'b0 ;
  assign n3791 = n1722 & ~n3790 ;
  assign n3792 = n671 ^ n533 ^ 1'b0 ;
  assign n3793 = n3792 ^ n3434 ^ 1'b0 ;
  assign n3796 = n1648 ^ n530 ^ 1'b0 ;
  assign n3797 = n2818 & ~n3796 ;
  assign n3794 = ( n982 & n2115 ) | ( n982 & ~n3525 ) | ( n2115 & ~n3525 ) ;
  assign n3795 = n2302 | n3794 ;
  assign n3798 = n3797 ^ n3795 ^ 1'b0 ;
  assign n3799 = n2985 & n3798 ;
  assign n3800 = ( n1718 & ~n2067 ) | ( n1718 & n3799 ) | ( ~n2067 & n3799 ) ;
  assign n3801 = n2375 | n2482 ;
  assign n3802 = n3801 ^ n681 ^ 1'b0 ;
  assign n3803 = ( n754 & n986 ) | ( n754 & n1594 ) | ( n986 & n1594 ) ;
  assign n3804 = x65 & ~n3803 ;
  assign n3805 = n3804 ^ n1408 ^ 1'b0 ;
  assign n3806 = n3615 & n3805 ;
  assign n3807 = n3806 ^ n3628 ^ 1'b0 ;
  assign n3808 = n2373 & ~n3158 ;
  assign n3809 = n2765 ^ n901 ^ 1'b0 ;
  assign n3810 = n1288 | n3809 ;
  assign n3811 = n3810 ^ n3740 ^ n301 ;
  assign n3812 = n655 & n672 ;
  assign n3813 = n575 & n1257 ;
  assign n3814 = ~n1416 & n3813 ;
  assign n3815 = n3814 ^ n974 ^ 1'b0 ;
  assign n3816 = ( n259 & n1072 ) | ( n259 & ~n2956 ) | ( n1072 & ~n2956 ) ;
  assign n3817 = n3229 | n3816 ;
  assign n3818 = n2111 & ~n3817 ;
  assign n3819 = n337 & n1123 ;
  assign n3820 = n3819 ^ n1892 ^ 1'b0 ;
  assign n3821 = n2839 & ~n3476 ;
  assign n3823 = n1139 ^ n945 ^ 1'b0 ;
  assign n3824 = n3823 ^ n1333 ^ 1'b0 ;
  assign n3825 = n345 & ~n3824 ;
  assign n3822 = n760 | n2905 ;
  assign n3826 = n3825 ^ n3822 ^ 1'b0 ;
  assign n3827 = n2517 & n2775 ;
  assign n3828 = n3827 ^ n3491 ^ 1'b0 ;
  assign n3829 = ~n1917 & n2399 ;
  assign n3830 = ~n418 & n3829 ;
  assign n3831 = ~n2864 & n3830 ;
  assign n3832 = ( n1791 & n2330 ) | ( n1791 & ~n3358 ) | ( n2330 & ~n3358 ) ;
  assign n3833 = n576 ^ n479 ^ 1'b0 ;
  assign n3834 = ~n616 & n3833 ;
  assign n3835 = ( n1117 & n1439 ) | ( n1117 & n3834 ) | ( n1439 & n3834 ) ;
  assign n3836 = n3766 ^ n3509 ^ n517 ;
  assign n3837 = n1286 | n3626 ;
  assign n3838 = n1106 & ~n3837 ;
  assign n3839 = n3838 ^ n1480 ^ 1'b0 ;
  assign n3840 = n1238 & n3839 ;
  assign n3841 = ~x27 & n801 ;
  assign n3842 = ~n3840 & n3841 ;
  assign n3843 = n3836 ^ n379 ^ 1'b0 ;
  assign n3844 = n744 | n3843 ;
  assign n3845 = n3038 ^ n1238 ^ 1'b0 ;
  assign n3846 = n3845 ^ n1907 ^ 1'b0 ;
  assign n3847 = n2036 ^ n912 ^ 1'b0 ;
  assign n3848 = n143 & n692 ;
  assign n3849 = n3848 ^ n405 ^ 1'b0 ;
  assign n3850 = n271 & ~n3373 ;
  assign n3851 = n3850 ^ n2008 ^ 1'b0 ;
  assign n3852 = n1306 | n3851 ;
  assign n3853 = n3849 | n3852 ;
  assign n3854 = n712 & n3853 ;
  assign n3855 = ~n3847 & n3854 ;
  assign n3856 = ~n3846 & n3855 ;
  assign n3857 = ~n148 & n3089 ;
  assign n3858 = n3857 ^ n2087 ^ n1455 ;
  assign n3859 = n2678 | n3055 ;
  assign n3860 = n3859 ^ n1936 ^ 1'b0 ;
  assign n3861 = n1545 & ~n1953 ;
  assign n3862 = n3861 ^ n3170 ^ n1045 ;
  assign n3863 = n3862 ^ n3156 ^ 1'b0 ;
  assign n3864 = x91 & n3863 ;
  assign n3865 = n3041 ^ n254 ^ 1'b0 ;
  assign n3866 = n3864 & ~n3865 ;
  assign n3867 = n821 | n1835 ;
  assign n3868 = n3867 ^ n584 ^ 1'b0 ;
  assign n3869 = n3468 ^ n2026 ^ n593 ;
  assign n3870 = ( n651 & n888 ) | ( n651 & n3869 ) | ( n888 & n3869 ) ;
  assign n3871 = n3870 ^ n2169 ^ n1532 ;
  assign n3872 = n3871 ^ n773 ^ 1'b0 ;
  assign n3873 = n1308 ^ n371 ^ 1'b0 ;
  assign n3874 = n463 & ~n3873 ;
  assign n3879 = ( n1009 & n1123 ) | ( n1009 & ~n1682 ) | ( n1123 & ~n1682 ) ;
  assign n3875 = n1293 & ~n2366 ;
  assign n3876 = n3875 ^ n1321 ^ 1'b0 ;
  assign n3877 = n1074 & ~n3876 ;
  assign n3878 = n215 & n3877 ;
  assign n3880 = n3879 ^ n3878 ^ 1'b0 ;
  assign n3881 = n3874 & ~n3880 ;
  assign n3882 = ~x3 & n248 ;
  assign n3891 = n1061 ^ n960 ^ 1'b0 ;
  assign n3892 = n657 | n3891 ;
  assign n3893 = ~n1610 & n1721 ;
  assign n3894 = n3893 ^ n1350 ^ 1'b0 ;
  assign n3895 = ~n3892 & n3894 ;
  assign n3896 = n1607 & ~n3895 ;
  assign n3885 = n1075 & n2195 ;
  assign n3883 = n1876 ^ n729 ^ 1'b0 ;
  assign n3884 = n370 & ~n3883 ;
  assign n3886 = n3885 ^ n3884 ^ 1'b0 ;
  assign n3887 = ( n2022 & n2441 ) | ( n2022 & n3886 ) | ( n2441 & n3886 ) ;
  assign n3888 = n2111 | n2574 ;
  assign n3889 = n2187 & ~n3888 ;
  assign n3890 = n3887 | n3889 ;
  assign n3897 = n3896 ^ n3890 ^ 1'b0 ;
  assign n3898 = n605 | n1059 ;
  assign n3899 = n148 & ~n3898 ;
  assign n3900 = ( n1849 & n2253 ) | ( n1849 & ~n3899 ) | ( n2253 & ~n3899 ) ;
  assign n3901 = ( n532 & n2190 ) | ( n532 & n3900 ) | ( n2190 & n3900 ) ;
  assign n3902 = n2112 & n2300 ;
  assign n3903 = n1505 & n3902 ;
  assign n3904 = ~n3901 & n3903 ;
  assign n3905 = n262 & n3904 ;
  assign n3906 = n3897 & n3905 ;
  assign n3907 = ~n2254 & n3153 ;
  assign n3908 = n3907 ^ n2252 ^ 1'b0 ;
  assign n3909 = n411 | n3908 ;
  assign n3910 = n3909 ^ n1062 ^ 1'b0 ;
  assign n3911 = n1000 | n1913 ;
  assign n3913 = ~n1023 & n1062 ;
  assign n3914 = x97 & n3913 ;
  assign n3912 = ~n1768 & n2257 ;
  assign n3915 = n3914 ^ n3912 ^ 1'b0 ;
  assign n3916 = n486 & n3915 ;
  assign n3917 = n475 ^ n361 ^ 1'b0 ;
  assign n3918 = ~n677 & n3917 ;
  assign n3919 = n3918 ^ n3182 ^ n1079 ;
  assign n3920 = n3919 ^ n3893 ^ n3159 ;
  assign n3921 = n3920 ^ n1722 ^ 1'b0 ;
  assign n3922 = n1864 & ~n3921 ;
  assign n3923 = n832 | n2767 ;
  assign n3924 = n2827 | n3923 ;
  assign n3925 = n997 & n3732 ;
  assign n3926 = ~n944 & n3925 ;
  assign n3927 = n3926 ^ n3441 ^ n3351 ;
  assign n3928 = n1585 & n2355 ;
  assign n3929 = n3928 ^ n1492 ^ 1'b0 ;
  assign n3930 = n470 ^ n346 ^ n338 ;
  assign n3931 = n3929 | n3930 ;
  assign n3932 = n173 & ~n1805 ;
  assign n3933 = ~n483 & n3932 ;
  assign n3934 = n3933 ^ n791 ^ 1'b0 ;
  assign n3935 = n1895 ^ x16 ^ 1'b0 ;
  assign n3936 = ~n403 & n1345 ;
  assign n3937 = n3935 & n3936 ;
  assign n3938 = n1840 ^ n1284 ^ 1'b0 ;
  assign n3939 = n3938 ^ n2060 ^ x79 ;
  assign n3940 = ~n3249 & n3939 ;
  assign n3943 = n2749 ^ n216 ^ 1'b0 ;
  assign n3944 = n1374 | n3943 ;
  assign n3945 = n1858 | n3944 ;
  assign n3941 = n3050 ^ n411 ^ 1'b0 ;
  assign n3942 = ~n2706 & n3941 ;
  assign n3946 = n3945 ^ n3942 ^ n3688 ;
  assign n3947 = n1162 ^ n305 ^ x115 ;
  assign n3948 = n319 & ~n3947 ;
  assign n3949 = n1974 ^ x67 ^ 1'b0 ;
  assign n3950 = n2130 | n3949 ;
  assign n3951 = n2602 | n3950 ;
  assign n3952 = n3951 ^ n2399 ^ 1'b0 ;
  assign n3953 = x81 & n1771 ;
  assign n3954 = x16 | n723 ;
  assign n3955 = n1370 ^ n129 ^ 1'b0 ;
  assign n3956 = ( n3953 & n3954 ) | ( n3953 & ~n3955 ) | ( n3954 & ~n3955 ) ;
  assign n3957 = n529 & n2621 ;
  assign n3958 = n3287 ^ n854 ^ 1'b0 ;
  assign n3959 = n2019 | n2027 ;
  assign n3960 = ~n875 & n3959 ;
  assign n3961 = n3492 ^ n1138 ^ 1'b0 ;
  assign n3962 = n1669 & n2864 ;
  assign n3965 = n190 | n2634 ;
  assign n3966 = n3965 ^ n1380 ^ 1'b0 ;
  assign n3967 = n3966 ^ n398 ^ 1'b0 ;
  assign n3968 = n3967 ^ n2640 ^ 1'b0 ;
  assign n3969 = n3643 | n3968 ;
  assign n3963 = n863 | n3766 ;
  assign n3964 = ( n1191 & n2159 ) | ( n1191 & ~n3963 ) | ( n2159 & ~n3963 ) ;
  assign n3970 = n3969 ^ n3964 ^ n1784 ;
  assign n3971 = n388 & n927 ;
  assign n3972 = n3971 ^ n1656 ^ 1'b0 ;
  assign n3973 = n3970 & n3972 ;
  assign n3974 = n1654 & n3973 ;
  assign n3975 = n3583 ^ n1566 ^ n1436 ;
  assign n3976 = x93 | n1360 ;
  assign n3977 = n3976 ^ n3354 ^ 1'b0 ;
  assign n3978 = ~n2725 & n3751 ;
  assign n3979 = n3978 ^ n319 ^ 1'b0 ;
  assign n3980 = x13 & ~n2952 ;
  assign n3981 = ~n1559 & n3143 ;
  assign n3982 = ( ~n190 & n3128 ) | ( ~n190 & n3247 ) | ( n3128 & n3247 ) ;
  assign n3983 = x32 & n2231 ;
  assign n3984 = ~n1300 & n3983 ;
  assign n3985 = n150 ^ x15 ^ 1'b0 ;
  assign n3986 = n1258 | n3985 ;
  assign n3987 = n3664 ^ n3455 ^ 1'b0 ;
  assign n3988 = x62 & n3987 ;
  assign n3989 = n3988 ^ n2291 ^ 1'b0 ;
  assign n3990 = n2853 ^ n740 ^ 1'b0 ;
  assign n3991 = n3990 ^ n3447 ^ 1'b0 ;
  assign n3992 = ~n1821 & n2617 ;
  assign n3993 = n2639 & n3992 ;
  assign n3994 = ( n188 & n1145 ) | ( n188 & ~n3608 ) | ( n1145 & ~n3608 ) ;
  assign n3995 = n3185 ^ n2214 ^ n980 ;
  assign n3996 = n3995 ^ n2419 ^ 1'b0 ;
  assign n3997 = n3996 ^ n3025 ^ n2041 ;
  assign n3998 = n1231 & n2706 ;
  assign n3999 = n1948 ^ n635 ^ n371 ;
  assign n4000 = n1100 | n3999 ;
  assign n4001 = n2964 ^ n1173 ^ 1'b0 ;
  assign n4002 = ~n1776 & n4001 ;
  assign n4003 = n530 ^ n461 ^ 1'b0 ;
  assign n4004 = ~n1000 & n4003 ;
  assign n4005 = ~n723 & n3572 ;
  assign n4006 = x68 & ~n4005 ;
  assign n4007 = n4004 & n4006 ;
  assign n4008 = ~x28 & n4007 ;
  assign n4009 = n529 & n1394 ;
  assign n4010 = n4009 ^ n237 ^ 1'b0 ;
  assign n4011 = n990 & n3066 ;
  assign n4012 = ( ~n324 & n2795 ) | ( ~n324 & n3980 ) | ( n2795 & n3980 ) ;
  assign n4013 = n946 & ~n1636 ;
  assign n4014 = n4013 ^ x70 ^ 1'b0 ;
  assign n4015 = n908 & n1815 ;
  assign n4016 = n4014 & n4015 ;
  assign n4017 = n1981 & n3547 ;
  assign n4018 = n578 & ~n4017 ;
  assign n4019 = n823 ^ n200 ^ 1'b0 ;
  assign n4020 = ( ~n909 & n2140 ) | ( ~n909 & n4019 ) | ( n2140 & n4019 ) ;
  assign n4021 = ~n1654 & n4020 ;
  assign n4022 = ~n671 & n4021 ;
  assign n4023 = n4022 ^ n623 ^ 1'b0 ;
  assign n4024 = n235 & n3940 ;
  assign n4026 = n701 ^ n429 ^ 1'b0 ;
  assign n4025 = n1265 ^ n753 ^ 1'b0 ;
  assign n4027 = n4026 ^ n4025 ^ 1'b0 ;
  assign n4028 = n141 | n4027 ;
  assign n4029 = n1450 | n1627 ;
  assign n4030 = n3793 & n4029 ;
  assign n4031 = n261 & n2238 ;
  assign n4032 = n4031 ^ n2219 ^ 1'b0 ;
  assign n4033 = n654 ^ n597 ^ n403 ;
  assign n4034 = n1529 | n4033 ;
  assign n4035 = n2291 ^ x97 ^ 1'b0 ;
  assign n4036 = n1754 & ~n4035 ;
  assign n4037 = n4034 & n4036 ;
  assign n4038 = n1671 ^ n469 ^ 1'b0 ;
  assign n4039 = n1892 ^ n1181 ^ n271 ;
  assign n4040 = n3438 ^ n2595 ^ 1'b0 ;
  assign n4041 = n4039 & ~n4040 ;
  assign n4042 = n2176 | n3657 ;
  assign n4043 = n813 & ~n4042 ;
  assign n4048 = x7 | n363 ;
  assign n4049 = n4048 ^ n2180 ^ 1'b0 ;
  assign n4044 = n1373 & ~n1730 ;
  assign n4045 = n1388 ^ n421 ^ 1'b0 ;
  assign n4046 = ~n852 & n4045 ;
  assign n4047 = ( ~n3878 & n4044 ) | ( ~n3878 & n4046 ) | ( n4044 & n4046 ) ;
  assign n4050 = n4049 ^ n4047 ^ n1370 ;
  assign n4052 = n1698 ^ n1588 ^ 1'b0 ;
  assign n4051 = n256 & ~n2143 ;
  assign n4053 = n4052 ^ n4051 ^ 1'b0 ;
  assign n4054 = n2180 ^ n1922 ^ n1650 ;
  assign n4055 = n4054 ^ n3269 ^ n2793 ;
  assign n4056 = n529 & n2787 ;
  assign n4057 = n4056 ^ n239 ^ 1'b0 ;
  assign n4058 = n2958 ^ n2155 ^ 1'b0 ;
  assign n4059 = n673 & n865 ;
  assign n4060 = ~n466 & n4059 ;
  assign n4061 = n4060 ^ n2546 ^ 1'b0 ;
  assign n4062 = x58 & ~n833 ;
  assign n4063 = n1307 | n2102 ;
  assign n4064 = n156 | n4063 ;
  assign n4065 = ( ~n3494 & n4062 ) | ( ~n3494 & n4064 ) | ( n4062 & n4064 ) ;
  assign n4066 = n161 & ~n4065 ;
  assign n4067 = ~n2649 & n4066 ;
  assign n4068 = n950 & n2201 ;
  assign n4069 = n1596 ^ n942 ^ 1'b0 ;
  assign n4070 = n2077 | n4069 ;
  assign n4071 = ( ~n1309 & n4068 ) | ( ~n1309 & n4070 ) | ( n4068 & n4070 ) ;
  assign n4072 = ~n4067 & n4071 ;
  assign n4073 = n3111 & n4072 ;
  assign n4074 = n4073 ^ n884 ^ 1'b0 ;
  assign n4075 = ~n4061 & n4074 ;
  assign n4076 = n653 ^ x22 ^ 1'b0 ;
  assign n4078 = ( ~n380 & n461 ) | ( ~n380 & n1034 ) | ( n461 & n1034 ) ;
  assign n4077 = n2444 & ~n2912 ;
  assign n4079 = n4078 ^ n4077 ^ 1'b0 ;
  assign n4080 = x58 & n4079 ;
  assign n4081 = n4080 ^ n1684 ^ 1'b0 ;
  assign n4082 = n3139 ^ n2285 ^ n129 ;
  assign n4083 = ~n584 & n1560 ;
  assign n4084 = n4083 ^ n3290 ^ 1'b0 ;
  assign n4085 = n1387 & ~n4084 ;
  assign n4086 = n1605 | n3551 ;
  assign n4087 = n4086 ^ n2817 ^ 1'b0 ;
  assign n4088 = n4087 ^ n3134 ^ 1'b0 ;
  assign n4089 = n4085 | n4088 ;
  assign n4090 = n4089 ^ n1465 ^ 1'b0 ;
  assign n4091 = ( n381 & n1764 ) | ( n381 & ~n2831 ) | ( n1764 & ~n2831 ) ;
  assign n4092 = ~n271 & n4091 ;
  assign n4093 = x7 & n3137 ;
  assign n4094 = n3084 & n4093 ;
  assign n4095 = n2638 ^ n1963 ^ x123 ;
  assign n4096 = n4094 | n4095 ;
  assign n4097 = n2111 ^ n1890 ^ 1'b0 ;
  assign n4098 = n1370 | n3954 ;
  assign n4099 = n4098 ^ n3802 ^ 1'b0 ;
  assign n4100 = n3158 ^ n1843 ^ 1'b0 ;
  assign n4101 = ~n3193 & n4100 ;
  assign n4102 = ~n3834 & n4101 ;
  assign n4103 = n2237 | n4102 ;
  assign n4104 = n312 | n4103 ;
  assign n4105 = n1487 & ~n2696 ;
  assign n4106 = n2262 & ~n3435 ;
  assign n4111 = n3857 ^ n293 ^ 1'b0 ;
  assign n4107 = n1590 & n3525 ;
  assign n4108 = n4107 ^ n1261 ^ n1067 ;
  assign n4109 = n1943 & ~n4108 ;
  assign n4110 = n872 & n4109 ;
  assign n4112 = n4111 ^ n4110 ^ 1'b0 ;
  assign n4113 = ~n1584 & n4112 ;
  assign n4114 = n2589 & n3503 ;
  assign n4115 = n4114 ^ n3947 ^ 1'b0 ;
  assign n4116 = n204 & ~n2694 ;
  assign n4117 = n4115 & n4116 ;
  assign n4118 = n4117 ^ n3411 ^ 1'b0 ;
  assign n4119 = n3499 ^ n2202 ^ n1771 ;
  assign n4120 = ( n1163 & n1528 ) | ( n1163 & ~n4119 ) | ( n1528 & ~n4119 ) ;
  assign n4121 = n3402 ^ n202 ^ 1'b0 ;
  assign n4122 = n4121 ^ n1953 ^ 1'b0 ;
  assign n4123 = ( ~n1213 & n1244 ) | ( ~n1213 & n4107 ) | ( n1244 & n4107 ) ;
  assign n4124 = ~n510 & n3482 ;
  assign n4125 = x22 & ~n467 ;
  assign n4126 = n4125 ^ n3788 ^ 1'b0 ;
  assign n4127 = n577 & ~n4126 ;
  assign n4128 = ~n4124 & n4127 ;
  assign n4129 = ~n1276 & n4128 ;
  assign n4130 = n2733 & n3948 ;
  assign n4131 = n1212 & ~n1364 ;
  assign n4132 = n2435 ^ n1847 ^ 1'b0 ;
  assign n4133 = n2309 & n4132 ;
  assign n4134 = n3586 & ~n4133 ;
  assign n4135 = n4134 ^ n1197 ^ 1'b0 ;
  assign n4136 = n2688 & ~n3098 ;
  assign n4137 = n1626 ^ n1305 ^ 1'b0 ;
  assign n4138 = ~n3323 & n4137 ;
  assign n4139 = n1863 & n4136 ;
  assign n4140 = ~n4138 & n4139 ;
  assign n4141 = n1376 & ~n1973 ;
  assign n4142 = x35 & ~n4141 ;
  assign n4143 = n4142 ^ n954 ^ 1'b0 ;
  assign n4144 = n250 ^ n191 ^ 1'b0 ;
  assign n4145 = n2485 ^ n548 ^ x100 ;
  assign n4146 = n4145 ^ n3367 ^ 1'b0 ;
  assign n4147 = ~n225 & n4146 ;
  assign n4148 = n1279 & n1693 ;
  assign n4149 = n4132 & n4148 ;
  assign n4150 = ~x39 & n283 ;
  assign n4151 = n1697 & n4150 ;
  assign n4152 = ~n854 & n2142 ;
  assign n4153 = ~n3134 & n4152 ;
  assign n4154 = n1999 & n4122 ;
  assign n4155 = ( n1088 & n1193 ) | ( n1088 & n1632 ) | ( n1193 & n1632 ) ;
  assign n4156 = n1867 & ~n4155 ;
  assign n4157 = n429 & ~n1074 ;
  assign n4158 = n380 & n2495 ;
  assign n4159 = n4157 & n4158 ;
  assign n4160 = n1452 & ~n4159 ;
  assign n4161 = n975 & n4160 ;
  assign n4162 = ~n471 & n2782 ;
  assign n4165 = n2721 ^ n919 ^ 1'b0 ;
  assign n4163 = ~x61 & n1766 ;
  assign n4164 = n1806 & ~n4163 ;
  assign n4166 = n4165 ^ n4164 ^ 1'b0 ;
  assign n4167 = n1513 & n4166 ;
  assign n4168 = ~n4162 & n4167 ;
  assign n4169 = n4168 ^ n2027 ^ 1'b0 ;
  assign n4170 = n1871 & n4169 ;
  assign n4171 = n4170 ^ n1894 ^ 1'b0 ;
  assign n4172 = n990 & n1217 ;
  assign n4173 = ~n2353 & n4172 ;
  assign n4174 = n1286 | n4173 ;
  assign n4175 = ~n1347 & n2796 ;
  assign n4176 = n4175 ^ n1039 ^ 1'b0 ;
  assign n4177 = n1320 & n4176 ;
  assign n4178 = n4177 ^ n3802 ^ 1'b0 ;
  assign n4179 = n523 | n630 ;
  assign n4180 = n4179 ^ n982 ^ 1'b0 ;
  assign n4181 = n2830 & n4180 ;
  assign n4182 = ~n3229 & n4181 ;
  assign n4183 = n4182 ^ n3760 ^ 1'b0 ;
  assign n4184 = n2898 ^ n1918 ^ n630 ;
  assign n4185 = n1033 ^ n791 ^ x110 ;
  assign n4186 = ( n2041 & ~n2523 ) | ( n2041 & n4185 ) | ( ~n2523 & n4185 ) ;
  assign n4187 = n1815 ^ n1267 ^ n998 ;
  assign n4188 = ~n4186 & n4187 ;
  assign n4189 = x64 & n176 ;
  assign n4190 = ~n1347 & n4189 ;
  assign n4191 = ~n381 & n4190 ;
  assign n4192 = ~n2972 & n4191 ;
  assign n4193 = n1406 & n1467 ;
  assign n4194 = n4193 ^ x107 ^ 1'b0 ;
  assign n4195 = n2866 | n4194 ;
  assign n4196 = ~n884 & n1454 ;
  assign n4197 = n4196 ^ n1907 ^ 1'b0 ;
  assign n4201 = x54 & ~n348 ;
  assign n4202 = ~n286 & n4201 ;
  assign n4203 = n417 & n796 ;
  assign n4204 = n4202 & n4203 ;
  assign n4205 = n901 & ~n4204 ;
  assign n4206 = x76 & n4205 ;
  assign n4207 = ~n373 & n4206 ;
  assign n4198 = x87 & n3205 ;
  assign n4199 = n4198 ^ n2422 ^ 1'b0 ;
  assign n4200 = n3710 | n4199 ;
  assign n4208 = n4207 ^ n4200 ^ 1'b0 ;
  assign n4209 = ~n752 & n944 ;
  assign n4210 = x121 & n4209 ;
  assign n4211 = n4210 ^ n210 ^ 1'b0 ;
  assign n4212 = n4211 ^ n615 ^ 1'b0 ;
  assign n4213 = n3472 & ~n4212 ;
  assign n4214 = n1387 & n1458 ;
  assign n4215 = n1976 ^ x16 ^ 1'b0 ;
  assign n4216 = n1583 | n4215 ;
  assign n4217 = n3176 | n3199 ;
  assign n4218 = n1198 | n4217 ;
  assign n4219 = n1634 & ~n4218 ;
  assign n4220 = n3163 | n4219 ;
  assign n4221 = n3529 ^ n2373 ^ n1747 ;
  assign n4222 = n4221 ^ n1017 ^ 1'b0 ;
  assign n4223 = n1222 & n2607 ;
  assign n4224 = ~n3247 & n4088 ;
  assign n4225 = n804 ^ n691 ^ 1'b0 ;
  assign n4226 = ~n4224 & n4225 ;
  assign n4227 = n4226 ^ n2629 ^ 1'b0 ;
  assign n4228 = n1293 & ~n2890 ;
  assign n4229 = n4228 ^ n2406 ^ 1'b0 ;
  assign n4230 = n707 & n1151 ;
  assign n4231 = n4230 ^ n2597 ^ 1'b0 ;
  assign n4232 = x113 & ~n530 ;
  assign n4233 = n3985 ^ n3006 ^ 1'b0 ;
  assign n4234 = x94 & ~n842 ;
  assign n4235 = n4234 ^ n764 ^ 1'b0 ;
  assign n4236 = n2693 ^ n331 ^ 1'b0 ;
  assign n4237 = ~n3969 & n4236 ;
  assign n4238 = ( n987 & n4235 ) | ( n987 & ~n4237 ) | ( n4235 & ~n4237 ) ;
  assign n4239 = ( n603 & n628 ) | ( n603 & ~n1648 ) | ( n628 & ~n1648 ) ;
  assign n4240 = ~x126 & n4239 ;
  assign n4241 = n4240 ^ n507 ^ 1'b0 ;
  assign n4242 = n661 | n2782 ;
  assign n4243 = n4242 ^ n442 ^ 1'b0 ;
  assign n4244 = ~n1048 & n4205 ;
  assign n4245 = n4244 ^ n1785 ^ 1'b0 ;
  assign n4246 = n4245 ^ n978 ^ 1'b0 ;
  assign n4247 = n4246 ^ n3434 ^ n1303 ;
  assign n4248 = n4243 | n4247 ;
  assign n4249 = n994 | n4248 ;
  assign n4250 = n214 | n218 ;
  assign n4251 = n961 | n1297 ;
  assign n4252 = n2016 | n4251 ;
  assign n4253 = n4252 ^ n2988 ^ 1'b0 ;
  assign n4254 = n1494 ^ n980 ^ n755 ;
  assign n4255 = n630 & ~n1118 ;
  assign n4256 = n2705 | n3067 ;
  assign n4257 = n711 | n4256 ;
  assign n4258 = n2444 & n4257 ;
  assign n4259 = n1240 & n4258 ;
  assign n4260 = x18 & ~n2708 ;
  assign n4261 = n4260 ^ n2845 ^ 1'b0 ;
  assign n4262 = ( n4255 & n4259 ) | ( n4255 & n4261 ) | ( n4259 & n4261 ) ;
  assign n4263 = n2018 ^ n1053 ^ 1'b0 ;
  assign n4264 = ~n2377 & n4263 ;
  assign n4266 = ( n2109 & ~n2390 ) | ( n2109 & n3282 ) | ( ~n2390 & n3282 ) ;
  assign n4265 = n2260 & ~n2323 ;
  assign n4267 = n4266 ^ n4265 ^ 1'b0 ;
  assign n4268 = x110 & n1136 ;
  assign n4269 = n415 & n2568 ;
  assign n4270 = n4269 ^ n1169 ^ 1'b0 ;
  assign n4271 = ~n4224 & n4270 ;
  assign n4272 = n4271 ^ n3783 ^ n2795 ;
  assign n4273 = ( n1605 & n4268 ) | ( n1605 & ~n4272 ) | ( n4268 & ~n4272 ) ;
  assign n4274 = n4273 ^ n1041 ^ 1'b0 ;
  assign n4275 = ~n4267 & n4274 ;
  assign n4276 = n1939 ^ n599 ^ 1'b0 ;
  assign n4277 = n4276 ^ n519 ^ 1'b0 ;
  assign n4278 = n305 & ~n1718 ;
  assign n4279 = n4199 & n4278 ;
  assign n4280 = n2256 | n4279 ;
  assign n4281 = x107 & n2529 ;
  assign n4283 = ~x7 & n2700 ;
  assign n4284 = ~n1155 & n3503 ;
  assign n4285 = ~n4283 & n4284 ;
  assign n4282 = n4141 ^ n2855 ^ 1'b0 ;
  assign n4286 = n4285 ^ n4282 ^ n1057 ;
  assign n4287 = n283 & n2151 ;
  assign n4288 = n4287 ^ n975 ^ 1'b0 ;
  assign n4289 = ( n3249 & ~n3758 ) | ( n3249 & n4288 ) | ( ~n3758 & n4288 ) ;
  assign n4291 = n3452 ^ x97 ^ 1'b0 ;
  assign n4290 = ~n881 & n3436 ;
  assign n4292 = n4291 ^ n4290 ^ 1'b0 ;
  assign n4293 = n1452 & n1794 ;
  assign n4294 = n2608 & ~n4293 ;
  assign n4295 = ( n1708 & n3656 ) | ( n1708 & n4294 ) | ( n3656 & n4294 ) ;
  assign n4299 = n547 ^ n275 ^ 1'b0 ;
  assign n4300 = n529 & n4299 ;
  assign n4296 = n2728 ^ n1850 ^ 1'b0 ;
  assign n4297 = n1805 | n4296 ;
  assign n4298 = ~n225 & n4297 ;
  assign n4301 = n4300 ^ n4298 ^ n1291 ;
  assign n4302 = n2766 & ~n2932 ;
  assign n4303 = n4302 ^ n1042 ^ 1'b0 ;
  assign n4304 = n1955 | n4303 ;
  assign n4305 = n2907 | n4304 ;
  assign n4306 = n1882 ^ n1573 ^ n688 ;
  assign n4307 = ( n681 & ~n3953 ) | ( n681 & n3969 ) | ( ~n3953 & n3969 ) ;
  assign n4308 = n2814 & n3365 ;
  assign n4309 = n2482 ^ n1433 ^ n1154 ;
  assign n4310 = n1439 | n4309 ;
  assign n4311 = n4310 ^ n2277 ^ 1'b0 ;
  assign n4312 = n2923 ^ n1554 ^ 1'b0 ;
  assign n4313 = ~n370 & n3326 ;
  assign n4314 = n1450 | n4313 ;
  assign n4316 = n1973 ^ n1370 ^ 1'b0 ;
  assign n4317 = ~n1567 & n4316 ;
  assign n4318 = n132 & ~n4317 ;
  assign n4315 = n3302 ^ n3034 ^ n1684 ;
  assign n4319 = n4318 ^ n4315 ^ n2537 ;
  assign n4320 = n2927 ^ n2390 ^ 1'b0 ;
  assign n4321 = n1948 | n4186 ;
  assign n4322 = n4320 | n4321 ;
  assign n4323 = n182 | n4322 ;
  assign n4324 = n1785 ^ n395 ^ 1'b0 ;
  assign n4325 = n691 & n4324 ;
  assign n4326 = n1074 & n3047 ;
  assign n4327 = ~n4325 & n4326 ;
  assign n4329 = n1829 ^ n1219 ^ 1'b0 ;
  assign n4330 = ~n3576 & n4329 ;
  assign n4328 = ~n1506 & n3557 ;
  assign n4331 = n4330 ^ n4328 ^ 1'b0 ;
  assign n4332 = n2582 & ~n4331 ;
  assign n4333 = n2489 & n4332 ;
  assign n4334 = n1835 ^ x100 ^ 1'b0 ;
  assign n4335 = n2687 & ~n4334 ;
  assign n4336 = ( ~n138 & n3317 ) | ( ~n138 & n4335 ) | ( n3317 & n4335 ) ;
  assign n4337 = n1111 ^ x65 ^ 1'b0 ;
  assign n4338 = n462 & n597 ;
  assign n4339 = n4337 & n4338 ;
  assign n4340 = x31 & n1752 ;
  assign n4341 = ~n1517 & n4340 ;
  assign n4342 = n4339 & n4341 ;
  assign n4343 = ( n2453 & n2796 ) | ( n2453 & ~n4342 ) | ( n2796 & ~n4342 ) ;
  assign n4344 = n2222 ^ n1378 ^ n725 ;
  assign n4346 = n824 ^ n775 ^ n312 ;
  assign n4345 = n844 & ~n2128 ;
  assign n4347 = n4346 ^ n4345 ^ 1'b0 ;
  assign n4348 = n4347 ^ n3674 ^ 1'b0 ;
  assign n4353 = n1800 & n3197 ;
  assign n4350 = ~n2321 & n3755 ;
  assign n4351 = n4350 ^ n2710 ^ 1'b0 ;
  assign n4352 = n3292 | n4351 ;
  assign n4354 = n4353 ^ n4352 ^ 1'b0 ;
  assign n4349 = n912 & n3304 ;
  assign n4355 = n4354 ^ n4349 ^ 1'b0 ;
  assign n4356 = n3544 ^ x89 ^ 1'b0 ;
  assign n4357 = n2172 & ~n4356 ;
  assign n4358 = n603 | n3376 ;
  assign n4359 = n3565 ^ n179 ^ 1'b0 ;
  assign n4362 = x81 & ~n1966 ;
  assign n4360 = n1184 & ~n2750 ;
  assign n4361 = n4360 ^ n1766 ^ 1'b0 ;
  assign n4363 = n4362 ^ n4361 ^ 1'b0 ;
  assign n4364 = n4184 ^ n1940 ^ 1'b0 ;
  assign n4365 = n3479 ^ n2066 ^ 1'b0 ;
  assign n4366 = ~n2917 & n4365 ;
  assign n4367 = ~n923 & n1184 ;
  assign n4368 = n4367 ^ n1198 ^ 1'b0 ;
  assign n4369 = n4368 ^ n3497 ^ 1'b0 ;
  assign n4370 = ~n3847 & n3886 ;
  assign n4371 = n4369 & n4370 ;
  assign n4372 = n508 | n2636 ;
  assign n4373 = n4372 ^ n1576 ^ 1'b0 ;
  assign n4374 = n539 & n4373 ;
  assign n4375 = n2437 ^ n788 ^ 1'b0 ;
  assign n4376 = n4375 ^ n2526 ^ 1'b0 ;
  assign n4377 = n671 & ~n4376 ;
  assign n4378 = n3997 & n4377 ;
  assign n4379 = n2935 | n4049 ;
  assign n4380 = n3102 ^ n524 ^ 1'b0 ;
  assign n4381 = n1886 ^ n762 ^ 1'b0 ;
  assign n4382 = n957 & n4381 ;
  assign n4383 = x11 & n4004 ;
  assign n4384 = ~n4382 & n4383 ;
  assign n4385 = ( n876 & ~n1061 ) | ( n876 & n1584 ) | ( ~n1061 & n1584 ) ;
  assign n4386 = n2107 & ~n4385 ;
  assign n4387 = n2880 & n4386 ;
  assign n4388 = ~n3329 & n4387 ;
  assign n4389 = n4384 | n4388 ;
  assign n4390 = n4380 | n4389 ;
  assign n4391 = n2645 ^ n664 ^ x126 ;
  assign n4392 = ( ~n4188 & n4322 ) | ( ~n4188 & n4391 ) | ( n4322 & n4391 ) ;
  assign n4393 = n1798 ^ n1626 ^ 1'b0 ;
  assign n4394 = ( ~n214 & n615 ) | ( ~n214 & n1690 ) | ( n615 & n1690 ) ;
  assign n4395 = n4394 ^ n4346 ^ 1'b0 ;
  assign n4396 = n2865 ^ n534 ^ 1'b0 ;
  assign n4397 = n4395 | n4396 ;
  assign n4398 = n3022 ^ n2747 ^ 1'b0 ;
  assign n4399 = ~n745 & n3414 ;
  assign n4400 = ( n217 & n3631 ) | ( n217 & n4399 ) | ( n3631 & n4399 ) ;
  assign n4401 = n812 & ~n1486 ;
  assign n4402 = n4401 ^ n873 ^ 1'b0 ;
  assign n4403 = x94 & ~n200 ;
  assign n4404 = n4403 ^ n1208 ^ 1'b0 ;
  assign n4405 = ( n582 & n4402 ) | ( n582 & n4404 ) | ( n4402 & n4404 ) ;
  assign n4406 = n1061 & ~n4405 ;
  assign n4407 = ( n3755 & ~n4400 ) | ( n3755 & n4406 ) | ( ~n4400 & n4406 ) ;
  assign n4408 = n3308 ^ n3139 ^ n1314 ;
  assign n4409 = ( n1002 & n1036 ) | ( n1002 & n4085 ) | ( n1036 & n4085 ) ;
  assign n4410 = n4408 & n4409 ;
  assign n4411 = ~n850 & n1061 ;
  assign n4412 = n850 & n4411 ;
  assign n4413 = n594 & ~n4412 ;
  assign n4414 = n4412 & n4413 ;
  assign n4415 = n1421 | n4414 ;
  assign n4416 = n4414 & ~n4415 ;
  assign n4418 = ~n237 & n2340 ;
  assign n4419 = n4418 ^ x14 ^ 1'b0 ;
  assign n4417 = x102 & ~n830 ;
  assign n4420 = n4419 ^ n4417 ^ 1'b0 ;
  assign n4421 = ~n1486 & n4420 ;
  assign n4422 = n4421 ^ n3428 ^ 1'b0 ;
  assign n4423 = ~n4416 & n4422 ;
  assign n4424 = ~n3938 & n4423 ;
  assign n4425 = n3191 ^ n2901 ^ 1'b0 ;
  assign n4426 = n3420 | n4425 ;
  assign n4427 = n701 | n1603 ;
  assign n4428 = n4427 ^ x78 ^ 1'b0 ;
  assign n4430 = n1938 ^ n1880 ^ 1'b0 ;
  assign n4431 = n4430 ^ n2985 ^ 1'b0 ;
  assign n4432 = n1998 & ~n4431 ;
  assign n4429 = ~n1250 & n1320 ;
  assign n4433 = n4432 ^ n4429 ^ 1'b0 ;
  assign n4434 = n4428 & n4433 ;
  assign n4435 = n4434 ^ n933 ^ 1'b0 ;
  assign n4436 = ~n256 & n4435 ;
  assign n4438 = n210 & ~n2356 ;
  assign n4439 = n1718 & n4438 ;
  assign n4437 = n2404 & ~n2451 ;
  assign n4440 = n4439 ^ n4437 ^ 1'b0 ;
  assign n4441 = n348 & n4440 ;
  assign n4444 = n404 & ~n3326 ;
  assign n4442 = n1212 ^ n1193 ^ 1'b0 ;
  assign n4443 = n4442 ^ n1730 ^ 1'b0 ;
  assign n4445 = n4444 ^ n4443 ^ 1'b0 ;
  assign n4446 = n4445 ^ n4121 ^ 1'b0 ;
  assign n4447 = n990 & n2401 ;
  assign n4448 = x51 & ~n794 ;
  assign n4449 = n4443 ^ n3686 ^ 1'b0 ;
  assign n4450 = n4449 ^ n1666 ^ 1'b0 ;
  assign n4451 = n379 | n805 ;
  assign n4452 = n1374 | n4451 ;
  assign n4453 = n479 & n1131 ;
  assign n4454 = n3040 ^ n1041 ^ 1'b0 ;
  assign n4455 = ~n808 & n2376 ;
  assign n4456 = n3589 | n4455 ;
  assign n4457 = n2423 ^ n299 ^ 1'b0 ;
  assign n4458 = n4363 ^ n1149 ^ 1'b0 ;
  assign n4459 = n3468 & ~n4458 ;
  assign n4460 = ( x40 & n1079 ) | ( x40 & n4369 ) | ( n1079 & n4369 ) ;
  assign n4461 = n3124 ^ n1967 ^ 1'b0 ;
  assign n4462 = n3143 | n4461 ;
  assign n4463 = n4462 ^ n3705 ^ 1'b0 ;
  assign n4464 = ~n2608 & n4463 ;
  assign n4465 = n1151 & ~n3710 ;
  assign n4466 = ( n876 & n1116 ) | ( n876 & ~n2455 ) | ( n1116 & ~n2455 ) ;
  assign n4467 = ( n417 & ~n1920 ) | ( n417 & n2143 ) | ( ~n1920 & n2143 ) ;
  assign n4468 = n264 & n4467 ;
  assign n4469 = ( n4225 & n4466 ) | ( n4225 & ~n4468 ) | ( n4466 & ~n4468 ) ;
  assign n4470 = n4469 ^ n1500 ^ n838 ;
  assign n4471 = n403 & n4335 ;
  assign n4472 = n1687 | n1922 ;
  assign n4473 = n4472 ^ n955 ^ 1'b0 ;
  assign n4474 = n3758 | n4473 ;
  assign n4475 = n2318 ^ n654 ^ 1'b0 ;
  assign n4476 = ( n677 & n1236 ) | ( n677 & ~n2026 ) | ( n1236 & ~n2026 ) ;
  assign n4477 = n4476 ^ n4375 ^ n2389 ;
  assign n4478 = n436 ^ n176 ^ 1'b0 ;
  assign n4479 = n3025 ^ n429 ^ 1'b0 ;
  assign n4480 = n3304 ^ n2915 ^ 1'b0 ;
  assign n4481 = n740 | n4480 ;
  assign n4482 = ~n1403 & n1800 ;
  assign n4483 = ~n1706 & n4482 ;
  assign n4484 = n4362 | n4483 ;
  assign n4485 = n2988 & ~n4484 ;
  assign n4486 = n1938 & n2085 ;
  assign n4487 = n1286 & n4486 ;
  assign n4488 = n612 | n2503 ;
  assign n4489 = ~n4487 & n4488 ;
  assign n4490 = n1103 & ~n4489 ;
  assign n4492 = n1933 ^ n1070 ^ n575 ;
  assign n4493 = n1639 | n4492 ;
  assign n4494 = n4493 ^ n2651 ^ 1'b0 ;
  assign n4491 = ( n341 & ~n1983 ) | ( n341 & n2721 ) | ( ~n1983 & n2721 ) ;
  assign n4495 = n4494 ^ n4491 ^ n2094 ;
  assign n4496 = n2976 | n4495 ;
  assign n4497 = n4496 ^ n282 ^ 1'b0 ;
  assign n4498 = n1931 | n2853 ;
  assign n4499 = ~n2279 & n4498 ;
  assign n4500 = n4497 & n4499 ;
  assign n4501 = n726 & ~n3470 ;
  assign n4502 = n2469 & n4501 ;
  assign n4503 = n4502 ^ n1173 ^ 1'b0 ;
  assign n4504 = n1871 ^ n1641 ^ n1008 ;
  assign n4505 = n2052 ^ n953 ^ 1'b0 ;
  assign n4506 = n3206 | n4505 ;
  assign n4507 = n4504 & ~n4506 ;
  assign n4508 = n3998 & n4507 ;
  assign n4509 = ~n443 & n574 ;
  assign n4510 = n4509 ^ n938 ^ 1'b0 ;
  assign n4511 = n478 & ~n4510 ;
  assign n4512 = n4511 ^ n403 ^ x93 ;
  assign n4513 = x16 & n1271 ;
  assign n4514 = n3519 & n4513 ;
  assign n4515 = n439 & n2060 ;
  assign n4516 = n2079 ^ n2073 ^ 1'b0 ;
  assign n4517 = n2032 ^ n630 ^ 1'b0 ;
  assign n4518 = n408 & n4517 ;
  assign n4519 = ~n740 & n4518 ;
  assign n4520 = n4519 ^ n427 ^ 1'b0 ;
  assign n4521 = n130 & n1667 ;
  assign n4522 = n132 & n692 ;
  assign n4523 = n2870 & ~n4522 ;
  assign n4524 = n4521 & n4523 ;
  assign n4525 = n241 & ~n627 ;
  assign n4526 = n4525 ^ n2627 ^ 1'b0 ;
  assign n4527 = n2906 ^ n1086 ^ 1'b0 ;
  assign n4528 = ~n606 & n2746 ;
  assign n4529 = n4527 & n4528 ;
  assign n4530 = n2464 ^ x34 ^ 1'b0 ;
  assign n4531 = n2933 & n4530 ;
  assign n4532 = n3291 ^ n1088 ^ 1'b0 ;
  assign n4533 = n707 ^ n582 ^ 1'b0 ;
  assign n4534 = n4532 | n4533 ;
  assign n4535 = n4531 | n4534 ;
  assign n4537 = n2583 ^ n410 ^ 1'b0 ;
  assign n4536 = n1341 | n4113 ;
  assign n4538 = n4537 ^ n4536 ^ 1'b0 ;
  assign n4539 = n2937 ^ n1077 ^ n372 ;
  assign n4540 = n452 & n1844 ;
  assign n4541 = n4540 ^ x24 ^ 1'b0 ;
  assign n4542 = n1371 & ~n4541 ;
  assign n4543 = n196 & n4542 ;
  assign n4544 = n2126 | n2681 ;
  assign n4545 = n436 | n4544 ;
  assign n4546 = ~n553 & n4545 ;
  assign n4547 = n4546 ^ n3166 ^ 1'b0 ;
  assign n4548 = n1897 & ~n4547 ;
  assign n4549 = n3538 ^ n2443 ^ 1'b0 ;
  assign n4550 = ~n1092 & n4549 ;
  assign n4551 = n277 | n2978 ;
  assign n4552 = n4551 ^ n1632 ^ 1'b0 ;
  assign n4553 = n4550 | n4552 ;
  assign n4554 = n4491 ^ n3743 ^ 1'b0 ;
  assign n4555 = n4245 & n4554 ;
  assign n4558 = n673 | n884 ;
  assign n4559 = n4558 ^ n1069 ^ 1'b0 ;
  assign n4557 = ( ~n2333 & n3175 ) | ( ~n2333 & n4387 ) | ( n3175 & n4387 ) ;
  assign n4560 = n4559 ^ n4557 ^ n3304 ;
  assign n4561 = n3109 | n4560 ;
  assign n4556 = ~n182 & n4044 ;
  assign n4562 = n4561 ^ n4556 ^ 1'b0 ;
  assign n4563 = n783 & ~n1947 ;
  assign n4564 = ( n543 & n1159 ) | ( n543 & ~n4563 ) | ( n1159 & ~n4563 ) ;
  assign n4565 = n1501 ^ n648 ^ 1'b0 ;
  assign n4566 = n4565 ^ n2157 ^ 1'b0 ;
  assign n4567 = n2189 ^ n1390 ^ 1'b0 ;
  assign n4568 = n2112 & n4567 ;
  assign n4569 = ~n1309 & n4568 ;
  assign n4570 = ~n3945 & n4569 ;
  assign n4571 = n3607 | n3664 ;
  assign n4572 = n166 | n4571 ;
  assign n4573 = ~n1265 & n4572 ;
  assign n4574 = n3864 ^ n664 ^ 1'b0 ;
  assign n4575 = n1358 | n4574 ;
  assign n4576 = ( n1265 & n1440 ) | ( n1265 & ~n3803 ) | ( n1440 & ~n3803 ) ;
  assign n4577 = n4576 ^ n4538 ^ 1'b0 ;
  assign n4578 = ~n1286 & n4577 ;
  assign n4579 = n3562 ^ x86 ^ 1'b0 ;
  assign n4580 = n4503 ^ n4085 ^ 1'b0 ;
  assign n4583 = x42 & n716 ;
  assign n4584 = n4583 ^ n3487 ^ 1'b0 ;
  assign n4582 = n273 | n431 ;
  assign n4581 = n992 | n1765 ;
  assign n4585 = n4584 ^ n4582 ^ n4581 ;
  assign n4586 = n2759 ^ n2346 ^ n2184 ;
  assign n4588 = n461 & ~n1854 ;
  assign n4589 = n661 & n4588 ;
  assign n4587 = ~n1048 & n1592 ;
  assign n4590 = n4589 ^ n4587 ^ 1'b0 ;
  assign n4591 = ~n4586 & n4590 ;
  assign n4592 = n1326 & ~n1486 ;
  assign n4593 = ~n530 & n4592 ;
  assign n4594 = n369 & ~n4593 ;
  assign n4595 = ~n785 & n3918 ;
  assign n4596 = n4595 ^ n2631 ^ 1'b0 ;
  assign n4597 = n1153 & n4596 ;
  assign n4598 = n4449 & n4597 ;
  assign n4599 = ~n2737 & n4598 ;
  assign n4600 = ( ~n2194 & n3401 ) | ( ~n2194 & n4599 ) | ( n3401 & n4599 ) ;
  assign n4601 = n1687 & n3775 ;
  assign n4602 = n4601 ^ n1981 ^ 1'b0 ;
  assign n4603 = ~n700 & n1853 ;
  assign n4604 = n1788 & n3846 ;
  assign n4605 = ~n4603 & n4604 ;
  assign n4606 = x63 & ~n1739 ;
  assign n4607 = n4606 ^ n1710 ^ 1'b0 ;
  assign n4608 = n3528 | n4607 ;
  assign n4609 = n4608 ^ n2985 ^ 1'b0 ;
  assign n4610 = n493 & n4609 ;
  assign n4611 = n1237 ^ n526 ^ n380 ;
  assign n4612 = n4611 ^ n2811 ^ n707 ;
  assign n4613 = n992 ^ x24 ^ 1'b0 ;
  assign n4614 = n1740 & n3139 ;
  assign n4615 = n746 & ~n2498 ;
  assign n4616 = ~n4614 & n4615 ;
  assign n4617 = n1494 ^ n1295 ^ 1'b0 ;
  assign n4618 = n3623 & n4617 ;
  assign n4619 = n3334 & n4618 ;
  assign n4620 = n2591 & n4619 ;
  assign n4621 = n4620 ^ n1821 ^ 1'b0 ;
  assign n4622 = ~n3663 & n4621 ;
  assign n4623 = n2433 ^ n1585 ^ n1089 ;
  assign n4624 = ( n1566 & n3950 ) | ( n1566 & n4279 ) | ( n3950 & n4279 ) ;
  assign n4625 = ( ~n4174 & n4623 ) | ( ~n4174 & n4624 ) | ( n4623 & n4624 ) ;
  assign n4626 = n379 | n3220 ;
  assign n4629 = n719 & n1074 ;
  assign n4630 = n4629 ^ n2807 ^ 1'b0 ;
  assign n4627 = ~n657 & n2577 ;
  assign n4628 = n3387 & n4627 ;
  assign n4631 = n4630 ^ n4628 ^ 1'b0 ;
  assign n4632 = ( n1738 & n2596 ) | ( n1738 & ~n4084 ) | ( n2596 & ~n4084 ) ;
  assign n4633 = n4001 & ~n4279 ;
  assign n4634 = ~n4004 & n4633 ;
  assign n4635 = n633 | n1692 ;
  assign n4636 = n3139 | n4635 ;
  assign n4637 = n2958 & n4254 ;
  assign n4638 = n719 & n2112 ;
  assign n4639 = n938 & n4638 ;
  assign n4640 = n4639 ^ n4099 ^ 1'b0 ;
  assign n4641 = n1313 & n3585 ;
  assign n4642 = n4452 & ~n4641 ;
  assign n4643 = ~n326 & n1432 ;
  assign n4644 = ~n3554 & n4643 ;
  assign n4645 = n4644 ^ n2003 ^ 1'b0 ;
  assign n4646 = n2167 | n2821 ;
  assign n4647 = n4646 ^ x97 ^ 1'b0 ;
  assign n4648 = n4647 ^ n2325 ^ n605 ;
  assign n4649 = n1374 | n4162 ;
  assign n4650 = n4509 & ~n4649 ;
  assign n4651 = n370 & ~n979 ;
  assign n4652 = ~n607 & n4651 ;
  assign n4653 = n1582 & n2130 ;
  assign n4654 = ( n4650 & n4652 ) | ( n4650 & ~n4653 ) | ( n4652 & ~n4653 ) ;
  assign n4655 = n3612 ^ n2275 ^ 1'b0 ;
  assign n4656 = ~n1198 & n2406 ;
  assign n4657 = n1293 & n4656 ;
  assign n4658 = ~n3689 & n4657 ;
  assign n4659 = n236 | n467 ;
  assign n4660 = n4659 ^ n1828 ^ 1'b0 ;
  assign n4661 = ~n1877 & n1912 ;
  assign n4662 = n4466 & n4661 ;
  assign n4663 = n2985 | n4662 ;
  assign n4664 = ( n2062 & n3914 ) | ( n2062 & n4663 ) | ( n3914 & n4663 ) ;
  assign n4665 = n4664 ^ n3623 ^ 1'b0 ;
  assign n4667 = n1985 | n2647 ;
  assign n4666 = n301 | n2346 ;
  assign n4668 = n4667 ^ n4666 ^ 1'b0 ;
  assign n4669 = n4668 ^ n1752 ^ 1'b0 ;
  assign n4670 = n1869 | n3468 ;
  assign n4671 = n4669 | n4670 ;
  assign n4672 = n488 & n4671 ;
  assign n4673 = n186 | n3232 ;
  assign n4674 = n2622 | n4673 ;
  assign n4675 = x99 | n1680 ;
  assign n4676 = n4675 ^ n942 ^ 1'b0 ;
  assign n4677 = ~n755 & n4676 ;
  assign n4678 = ~n3363 & n4677 ;
  assign n4679 = n2431 ^ n1703 ^ 1'b0 ;
  assign n4680 = ~n1470 & n2309 ;
  assign n4681 = ~n4479 & n4680 ;
  assign n4682 = n956 ^ n345 ^ 1'b0 ;
  assign n4683 = n3210 & ~n4682 ;
  assign n4684 = n1854 | n4171 ;
  assign n4685 = n3591 ^ n3354 ^ n2662 ;
  assign n4688 = ~n179 & n1479 ;
  assign n4689 = n4688 ^ n760 ^ 1'b0 ;
  assign n4690 = n4689 ^ n3135 ^ n2510 ;
  assign n4686 = ~n1979 & n4084 ;
  assign n4687 = ~n1376 & n4686 ;
  assign n4691 = n4690 ^ n4687 ^ 1'b0 ;
  assign n4692 = n3678 ^ n337 ^ 1'b0 ;
  assign n4693 = n4691 & n4692 ;
  assign n4694 = n503 ^ x26 ^ 1'b0 ;
  assign n4695 = n4618 & ~n4694 ;
  assign n4696 = n3651 ^ n1824 ^ 1'b0 ;
  assign n4697 = ~n640 & n4696 ;
  assign n4698 = n4115 ^ n1766 ^ 1'b0 ;
  assign n4699 = ( ~n2435 & n3491 ) | ( ~n2435 & n4312 ) | ( n3491 & n4312 ) ;
  assign n4700 = n726 & ~n4699 ;
  assign n4701 = x5 & n182 ;
  assign n4702 = ( n206 & n560 ) | ( n206 & ~n1776 ) | ( n560 & ~n1776 ) ;
  assign n4703 = n4059 ^ x33 ^ 1'b0 ;
  assign n4704 = ( n377 & n1947 ) | ( n377 & n1985 ) | ( n1947 & n1985 ) ;
  assign n4705 = n4704 ^ n3954 ^ 1'b0 ;
  assign n4706 = ~n2574 & n3594 ;
  assign n4707 = n4706 ^ n2552 ^ 1'b0 ;
  assign n4708 = n4707 ^ n4059 ^ 1'b0 ;
  assign n4709 = x111 & n1062 ;
  assign n4710 = ~n703 & n4709 ;
  assign n4711 = n3362 | n4710 ;
  assign n4712 = n4711 ^ n809 ^ 1'b0 ;
  assign n4713 = ( n1268 & n1307 ) | ( n1268 & n4712 ) | ( n1307 & n4712 ) ;
  assign n4714 = n3048 ^ n2386 ^ n325 ;
  assign n4715 = n1856 | n3698 ;
  assign n4716 = n3272 ^ n2307 ^ 1'b0 ;
  assign n4717 = n4716 ^ n1575 ^ 1'b0 ;
  assign n4718 = n4263 ^ n2340 ^ n341 ;
  assign n4720 = ( n1327 & n3857 ) | ( n1327 & n4162 ) | ( n3857 & n4162 ) ;
  assign n4719 = n1650 & n3644 ;
  assign n4721 = n4720 ^ n4719 ^ 1'b0 ;
  assign n4722 = n1307 & n4721 ;
  assign n4723 = n3374 & n3572 ;
  assign n4724 = n403 & n1162 ;
  assign n4725 = n4724 ^ n202 ^ 1'b0 ;
  assign n4726 = n4725 ^ n2346 ^ 1'b0 ;
  assign n4727 = n416 & ~n4726 ;
  assign n4728 = n4727 ^ n303 ^ 1'b0 ;
  assign n4729 = n4723 & ~n4728 ;
  assign n4733 = ~n1343 & n2762 ;
  assign n4734 = n2810 & n4733 ;
  assign n4735 = n4734 ^ n149 ^ 1'b0 ;
  assign n4736 = n2476 & n4735 ;
  assign n4731 = n817 & ~n1649 ;
  assign n4732 = n4731 ^ n2255 ^ 1'b0 ;
  assign n4730 = ( n1496 & ~n1920 ) | ( n1496 & n2696 ) | ( ~n1920 & n2696 ) ;
  assign n4737 = n4736 ^ n4732 ^ n4730 ;
  assign n4738 = n1953 ^ n630 ^ 1'b0 ;
  assign n4739 = n4737 | n4738 ;
  assign n4740 = n1283 & ~n2340 ;
  assign n4741 = n4740 ^ n2887 ^ 1'b0 ;
  assign n4742 = n1792 & n4741 ;
  assign n4743 = n837 ^ n373 ^ 1'b0 ;
  assign n4744 = n1266 & n2443 ;
  assign n4745 = n4744 ^ n796 ^ 1'b0 ;
  assign n4746 = ( n1044 & ~n2878 ) | ( n1044 & n4125 ) | ( ~n2878 & n4125 ) ;
  assign n4747 = n2091 & ~n2160 ;
  assign n4748 = n1506 | n4747 ;
  assign n4749 = n1519 | n1624 ;
  assign n4750 = n4749 ^ n3740 ^ 1'b0 ;
  assign n4751 = n4593 ^ n3142 ^ n2104 ;
  assign n4752 = n3093 ^ x32 ^ 1'b0 ;
  assign n4753 = n4751 & n4752 ;
  assign n4754 = n4753 ^ n3994 ^ 1'b0 ;
  assign n4755 = n3701 ^ n1586 ^ 1'b0 ;
  assign n4756 = n4755 ^ n2622 ^ 1'b0 ;
  assign n4757 = n2503 & ~n4756 ;
  assign n4758 = n4076 ^ n3800 ^ 1'b0 ;
  assign n4759 = n3724 ^ n1123 ^ 1'b0 ;
  assign n4760 = n2966 ^ n2787 ^ 1'b0 ;
  assign n4761 = n2582 & ~n3922 ;
  assign n4762 = ~n652 & n725 ;
  assign n4763 = n2364 & n4762 ;
  assign n4764 = n4763 ^ n2135 ^ 1'b0 ;
  assign n4767 = n2905 ^ n2821 ^ n2053 ;
  assign n4765 = n1195 & ~n2112 ;
  assign n4766 = ~n2051 & n4765 ;
  assign n4768 = n4767 ^ n4766 ^ 1'b0 ;
  assign n4769 = n845 | n1109 ;
  assign n4770 = n1212 & n2479 ;
  assign n4771 = n4770 ^ n3277 ^ 1'b0 ;
  assign n4772 = ( n3627 & ~n4769 ) | ( n3627 & n4771 ) | ( ~n4769 & n4771 ) ;
  assign n4773 = n1088 ^ n1085 ^ n129 ;
  assign n4774 = n4773 ^ n2175 ^ 1'b0 ;
  assign n4775 = n1040 & ~n4774 ;
  assign n4776 = ~n2888 & n4205 ;
  assign n4777 = n1451 & ~n2077 ;
  assign n4778 = ( n681 & ~n3139 ) | ( n681 & n4777 ) | ( ~n3139 & n4777 ) ;
  assign n4779 = n3967 | n4778 ;
  assign n4780 = ( ~n1127 & n1318 ) | ( ~n1127 & n4095 ) | ( n1318 & n4095 ) ;
  assign n4781 = x85 & n2505 ;
  assign n4782 = ~n3854 & n4781 ;
  assign n4783 = n798 & n3433 ;
  assign n4784 = ~n3152 & n3631 ;
  assign n4785 = ~n4323 & n4784 ;
  assign n4786 = ( ~n571 & n3230 ) | ( ~n571 & n3785 ) | ( n3230 & n3785 ) ;
  assign n4787 = n4563 & n4786 ;
  assign n4788 = ~n457 & n2444 ;
  assign n4789 = n4161 ^ n2553 ^ 1'b0 ;
  assign n4790 = n2922 ^ n2772 ^ 1'b0 ;
  assign n4791 = n4442 | n4790 ;
  assign n4792 = n3353 & ~n4791 ;
  assign n4793 = n4789 & n4792 ;
  assign n4796 = n2000 & n3172 ;
  assign n4794 = n1057 & ~n1489 ;
  assign n4795 = n1688 & n4794 ;
  assign n4797 = n4796 ^ n4795 ^ 1'b0 ;
  assign n4798 = n1455 & n4429 ;
  assign n4799 = n4798 ^ n1760 ^ 1'b0 ;
  assign n4800 = n4799 ^ n1943 ^ 1'b0 ;
  assign n4801 = n4347 & ~n4800 ;
  assign n4802 = x80 & n4801 ;
  assign n4803 = n1123 ^ n186 ^ 1'b0 ;
  assign n4804 = ~n2569 & n3712 ;
  assign n4805 = ~n4803 & n4804 ;
  assign n4806 = n2549 ^ n2064 ^ n798 ;
  assign n4807 = n4420 & ~n4806 ;
  assign n4808 = n4807 ^ x62 ^ 1'b0 ;
  assign n4809 = n463 & ~n1379 ;
  assign n4810 = n4809 ^ n1786 ^ 1'b0 ;
  assign n4811 = n4810 ^ n1718 ^ n524 ;
  assign n4812 = n1273 ^ n1175 ^ 1'b0 ;
  assign n4820 = n4204 ^ n2663 ^ 1'b0 ;
  assign n4813 = n3324 ^ n2985 ^ 1'b0 ;
  assign n4814 = n965 ^ n651 ^ 1'b0 ;
  assign n4815 = n169 | n4814 ;
  assign n4816 = n2206 & ~n4815 ;
  assign n4817 = n4816 ^ n2249 ^ 1'b0 ;
  assign n4818 = x122 & ~n4817 ;
  assign n4819 = n4813 & n4818 ;
  assign n4821 = n4820 ^ n4819 ^ 1'b0 ;
  assign n4822 = n762 ^ x106 ^ 1'b0 ;
  assign n4823 = n4822 ^ n156 ^ 1'b0 ;
  assign n4824 = n831 & n4823 ;
  assign n4825 = x125 & ~n3193 ;
  assign n4826 = n4825 ^ n875 ^ 1'b0 ;
  assign n4827 = ( n2643 & n4824 ) | ( n2643 & n4826 ) | ( n4824 & n4826 ) ;
  assign n4828 = n3916 ^ n1948 ^ n1636 ;
  assign n4829 = n4827 | n4828 ;
  assign n4831 = ~n1772 & n2843 ;
  assign n4832 = n4831 ^ x107 ^ 1'b0 ;
  assign n4833 = ( x25 & n159 ) | ( x25 & n986 ) | ( n159 & n986 ) ;
  assign n4834 = n584 | n4833 ;
  assign n4835 = n4832 & ~n4834 ;
  assign n4830 = ~n2903 & n4727 ;
  assign n4836 = n4835 ^ n4830 ^ 1'b0 ;
  assign n4837 = n4836 ^ n1525 ^ 1'b0 ;
  assign n4838 = n389 & ~n2840 ;
  assign n4839 = n4838 ^ n4479 ^ 1'b0 ;
  assign n4840 = ~n369 & n1305 ;
  assign n4841 = n4840 ^ n661 ^ 1'b0 ;
  assign n4842 = n4839 & n4841 ;
  assign n4844 = n1401 ^ n708 ^ n524 ;
  assign n4843 = ~n1055 & n3565 ;
  assign n4845 = n4844 ^ n4843 ^ 1'b0 ;
  assign n4846 = n2373 & n3020 ;
  assign n4847 = n2299 & ~n3908 ;
  assign n4848 = n728 & ~n4757 ;
  assign n4849 = x119 & n1050 ;
  assign n4850 = ~n374 & n4849 ;
  assign n4851 = ( x86 & n3373 ) | ( x86 & ~n4850 ) | ( n3373 & ~n4850 ) ;
  assign n4852 = n1566 & n2355 ;
  assign n4853 = ~n4851 & n4852 ;
  assign n4854 = ( n240 & n582 ) | ( n240 & ~n1870 ) | ( n582 & ~n1870 ) ;
  assign n4855 = n3499 ^ n1084 ^ n417 ;
  assign n4856 = n4854 | n4855 ;
  assign n4857 = n4853 & ~n4856 ;
  assign n4858 = n2396 ^ n1907 ^ n1224 ;
  assign n4859 = n4565 | n4858 ;
  assign n4860 = n436 & ~n2940 ;
  assign n4861 = ~n381 & n416 ;
  assign n4862 = n4861 ^ n1629 ^ 1'b0 ;
  assign n4863 = n4154 | n4862 ;
  assign n4864 = n4863 ^ n3739 ^ n1571 ;
  assign n4866 = n2087 ^ x68 ^ 1'b0 ;
  assign n4865 = n4552 ^ n2796 ^ 1'b0 ;
  assign n4867 = n4866 ^ n4865 ^ n1492 ;
  assign n4868 = n2248 & n3590 ;
  assign n4869 = n3020 ^ n892 ^ 1'b0 ;
  assign n4870 = n4869 ^ n2727 ^ 1'b0 ;
  assign n4871 = n1238 & n1946 ;
  assign n4872 = n4870 & n4871 ;
  assign n4873 = n1954 & ~n4872 ;
  assign n4874 = n920 & n4873 ;
  assign n4875 = n1088 & n3377 ;
  assign n4876 = n845 & ~n3399 ;
  assign n4877 = ( n314 & n1869 ) | ( n314 & n4876 ) | ( n1869 & n4876 ) ;
  assign n4878 = n1722 & n2074 ;
  assign n4879 = n449 & n4878 ;
  assign n4880 = n395 & ~n4879 ;
  assign n4881 = n4880 ^ n4820 ^ 1'b0 ;
  assign n4882 = n4877 & n4881 ;
  assign n4883 = ~n4875 & n4882 ;
  assign n4884 = n3395 ^ n261 ^ 1'b0 ;
  assign n4885 = n805 & n4119 ;
  assign n4886 = n4885 ^ n1528 ^ 1'b0 ;
  assign n4887 = n4106 | n4860 ;
  assign n4888 = ~n712 & n2053 ;
  assign n4889 = ~n2053 & n4888 ;
  assign n4890 = n1954 | n4889 ;
  assign n4891 = n4890 ^ n3993 ^ n3289 ;
  assign n4892 = ~n3244 & n3732 ;
  assign n4893 = n4892 ^ n3893 ^ 1'b0 ;
  assign n4894 = x21 & n1821 ;
  assign n4895 = n4894 ^ n3184 ^ 1'b0 ;
  assign n4896 = n1088 & ~n4895 ;
  assign n4897 = n4380 & ~n4876 ;
  assign n4898 = n2456 & n3510 ;
  assign n4899 = n764 & n4686 ;
  assign n4900 = ~n3879 & n4899 ;
  assign n4901 = n883 & n1566 ;
  assign n4902 = n1885 & n4901 ;
  assign n4903 = n1269 & ~n3969 ;
  assign n4904 = n3102 | n4903 ;
  assign n4905 = n4904 ^ n456 ^ 1'b0 ;
  assign n4906 = n4902 | n4905 ;
  assign n4907 = n4906 ^ n4078 ^ n524 ;
  assign n4908 = ~n760 & n2959 ;
  assign n4909 = n4908 ^ n3981 ^ 1'b0 ;
  assign n4910 = n3455 ^ n697 ^ 1'b0 ;
  assign n4911 = n2527 & n4910 ;
  assign n4912 = n4911 ^ n2243 ^ 1'b0 ;
  assign n4913 = n4912 ^ n3249 ^ 1'b0 ;
  assign n4914 = n2954 ^ n2708 ^ 1'b0 ;
  assign n4915 = ~n4913 & n4914 ;
  assign n4916 = n2443 & ~n2945 ;
  assign n4917 = ~n879 & n4916 ;
  assign n4918 = x44 & n424 ;
  assign n4919 = n443 & n4918 ;
  assign n4920 = n3900 ^ n1966 ^ 1'b0 ;
  assign n4921 = n2908 & n4920 ;
  assign n4922 = n4921 ^ n3187 ^ 1'b0 ;
  assign n4923 = n4919 | n4922 ;
  assign n4924 = n1911 & ~n2853 ;
  assign n4925 = n4924 ^ n1048 ^ 1'b0 ;
  assign n4926 = n4057 & n4925 ;
  assign n4927 = n4923 & n4926 ;
  assign n4928 = n3689 & ~n4927 ;
  assign n4929 = n4928 ^ n2726 ^ 1'b0 ;
  assign n4930 = n588 & ~n1959 ;
  assign n4931 = n4459 ^ n1734 ^ 1'b0 ;
  assign n4932 = n3031 ^ n1150 ^ n216 ;
  assign n4933 = ( n150 & n2309 ) | ( n150 & ~n4932 ) | ( n2309 & ~n4932 ) ;
  assign n4934 = ~n2656 & n3130 ;
  assign n4935 = ~n1644 & n4934 ;
  assign n4936 = ( n443 & ~n1354 ) | ( n443 & n1909 ) | ( ~n1354 & n1909 ) ;
  assign n4937 = n4935 & n4936 ;
  assign n4938 = n3275 | n4937 ;
  assign n4943 = n1335 ^ n888 ^ 1'b0 ;
  assign n4944 = ~n277 & n4943 ;
  assign n4940 = n2920 ^ n2382 ^ n276 ;
  assign n4939 = n259 | n4740 ;
  assign n4941 = n4940 ^ n4939 ^ 1'b0 ;
  assign n4942 = ~n1645 & n4941 ;
  assign n4945 = n4944 ^ n4942 ^ 1'b0 ;
  assign n4946 = n527 & ~n2219 ;
  assign n4948 = ( n830 & ~n919 ) | ( n830 & n1147 ) | ( ~n919 & n1147 ) ;
  assign n4949 = n4948 ^ n2668 ^ 1'b0 ;
  assign n4950 = n2910 & n4949 ;
  assign n4947 = n1380 & ~n2863 ;
  assign n4951 = n4950 ^ n4947 ^ 1'b0 ;
  assign n4952 = ( ~n1953 & n4946 ) | ( ~n1953 & n4951 ) | ( n4946 & n4951 ) ;
  assign n4953 = ~n2998 & n4357 ;
  assign n4954 = n1081 & n4953 ;
  assign n4955 = n4156 ^ n1810 ^ 1'b0 ;
  assign n4956 = n619 ^ n427 ^ 1'b0 ;
  assign n4957 = n4956 ^ n1679 ^ 1'b0 ;
  assign n4958 = n1989 ^ n1594 ^ 1'b0 ;
  assign n4959 = n1276 & n4958 ;
  assign n4960 = n4959 ^ n3014 ^ 1'b0 ;
  assign n4961 = n1081 | n4960 ;
  assign n4962 = n2283 ^ n1372 ^ 1'b0 ;
  assign n4963 = n4962 ^ n4932 ^ 1'b0 ;
  assign n4964 = n1652 & ~n2739 ;
  assign n4965 = n3975 & ~n4639 ;
  assign n4966 = n4757 & n4965 ;
  assign n4967 = n1785 | n2741 ;
  assign n4968 = n4967 ^ n4084 ^ 1'b0 ;
  assign n4969 = x23 & n4968 ;
  assign n4970 = n1200 & n4969 ;
  assign n4971 = n4970 ^ n4333 ^ 1'b0 ;
  assign n4972 = n337 & n4971 ;
  assign n4973 = ~n972 & n4972 ;
  assign n4974 = n4973 ^ n2167 ^ 1'b0 ;
  assign n4975 = n3552 ^ n1418 ^ 1'b0 ;
  assign n4976 = n4975 ^ n3882 ^ 1'b0 ;
  assign n4977 = n503 | n4976 ;
  assign n4978 = x121 ^ x99 ^ 1'b0 ;
  assign n4979 = n2755 & ~n4978 ;
  assign n4980 = n406 & n4979 ;
  assign n4981 = ~n539 & n4980 ;
  assign n4982 = n3958 & ~n4981 ;
  assign n4983 = ~x45 & n4982 ;
  assign n4984 = ( n1277 & n4730 ) | ( n1277 & ~n4983 ) | ( n4730 & ~n4983 ) ;
  assign n4985 = n3119 ^ n1591 ^ n1286 ;
  assign n4986 = ~n2157 & n4985 ;
  assign n4987 = n4986 ^ n2888 ^ 1'b0 ;
  assign n4988 = n2012 ^ n538 ^ 1'b0 ;
  assign n4989 = n4988 ^ n1525 ^ 1'b0 ;
  assign n4990 = n2000 & n4989 ;
  assign n4991 = n4990 ^ n2742 ^ n179 ;
  assign n4992 = n4100 ^ n2807 ^ n2692 ;
  assign n4993 = n4992 ^ n1721 ^ 1'b0 ;
  assign n4994 = ~n1081 & n4046 ;
  assign n4995 = n4993 & n4994 ;
  assign n4996 = n4675 | n4725 ;
  assign n4997 = n745 | n959 ;
  assign n4998 = n4997 ^ n577 ^ 1'b0 ;
  assign n4999 = ( n1042 & n4639 ) | ( n1042 & ~n4998 ) | ( n4639 & ~n4998 ) ;
  assign n5000 = n1811 | n4999 ;
  assign n5001 = n2736 & ~n5000 ;
  assign n5002 = x89 & n1166 ;
  assign n5003 = n3625 ^ n490 ^ 1'b0 ;
  assign n5004 = n654 & ~n1193 ;
  assign n5005 = n3547 ^ n383 ^ 1'b0 ;
  assign n5006 = ~n3682 & n5005 ;
  assign n5007 = n5006 ^ n4916 ^ 1'b0 ;
  assign n5008 = n5004 & ~n5007 ;
  assign n5009 = n1069 ^ n830 ^ 1'b0 ;
  assign n5010 = n5009 ^ n2064 ^ 1'b0 ;
  assign n5011 = ~n1172 & n5010 ;
  assign n5012 = n5011 ^ n2535 ^ 1'b0 ;
  assign n5013 = n794 | n5012 ;
  assign n5014 = n4801 ^ n3587 ^ n2981 ;
  assign n5015 = n1155 ^ n254 ^ 1'b0 ;
  assign n5016 = n1026 & n5015 ;
  assign n5017 = n1162 ^ n1013 ^ 1'b0 ;
  assign n5018 = n2549 | n3249 ;
  assign n5019 = n3818 | n5018 ;
  assign n5020 = n1251 | n5019 ;
  assign n5021 = n3382 ^ n1636 ^ 1'b0 ;
  assign n5022 = n1776 ^ x80 ^ 1'b0 ;
  assign n5023 = n2581 ^ n2018 ^ 1'b0 ;
  assign n5024 = n5022 & ~n5023 ;
  assign n5025 = n1131 & n5024 ;
  assign n5026 = n2796 & n3077 ;
  assign n5027 = n5026 ^ n962 ^ 1'b0 ;
  assign n5028 = n3320 ^ n997 ^ 1'b0 ;
  assign n5029 = n5027 | n5028 ;
  assign n5030 = n2479 ^ n2241 ^ 1'b0 ;
  assign n5031 = n5030 ^ n2365 ^ 1'b0 ;
  assign n5032 = ( ~n1229 & n2362 ) | ( ~n1229 & n5031 ) | ( n2362 & n5031 ) ;
  assign n5033 = n2957 ^ n607 ^ 1'b0 ;
  assign n5034 = n750 & n5033 ;
  assign n5035 = n1364 & ~n4667 ;
  assign n5036 = ~n5034 & n5035 ;
  assign n5037 = n179 | n314 ;
  assign n5038 = n395 | n1384 ;
  assign n5039 = n5037 & ~n5038 ;
  assign n5040 = n2334 ^ n1430 ^ 1'b0 ;
  assign n5041 = ( n893 & n3036 ) | ( n893 & n5040 ) | ( n3036 & n5040 ) ;
  assign n5042 = n671 & ~n3126 ;
  assign n5043 = n5042 ^ x40 ^ 1'b0 ;
  assign n5044 = n1445 & ~n5043 ;
  assign n5045 = n5041 & n5044 ;
  assign n5046 = n2019 & ~n4820 ;
  assign n5047 = n4578 ^ n1008 ^ 1'b0 ;
  assign n5048 = n2640 & ~n5047 ;
  assign n5049 = n691 & n1186 ;
  assign n5050 = n2275 & n5049 ;
  assign n5051 = n5050 ^ n3403 ^ 1'b0 ;
  assign n5052 = n2544 ^ n2060 ^ 1'b0 ;
  assign n5053 = n5052 ^ n729 ^ 1'b0 ;
  assign n5055 = n1976 ^ n564 ^ 1'b0 ;
  assign n5056 = n1461 | n5055 ;
  assign n5054 = n876 | n2128 ;
  assign n5057 = n5056 ^ n5054 ^ 1'b0 ;
  assign n5058 = n5057 ^ n3435 ^ n1513 ;
  assign n5059 = ~n362 & n3489 ;
  assign n5060 = ~n1240 & n3494 ;
  assign n5061 = ( n3768 & n5059 ) | ( n3768 & n5060 ) | ( n5059 & n5060 ) ;
  assign n5062 = n1405 | n4532 ;
  assign n5063 = n5062 ^ n895 ^ 1'b0 ;
  assign n5064 = n173 & ~n935 ;
  assign n5065 = n1583 | n5064 ;
  assign n5066 = n4252 | n5065 ;
  assign n5067 = n5063 & n5066 ;
  assign n5068 = n1319 & ~n5067 ;
  assign n5069 = ~n3173 & n5068 ;
  assign n5070 = n3296 ^ n1462 ^ 1'b0 ;
  assign n5071 = n442 | n5070 ;
  assign n5072 = n5071 ^ n2403 ^ 1'b0 ;
  assign n5073 = n267 | n381 ;
  assign n5074 = n5073 ^ n754 ^ 1'b0 ;
  assign n5075 = n4157 ^ n2568 ^ 1'b0 ;
  assign n5076 = n5074 & ~n5075 ;
  assign n5077 = n5076 ^ n959 ^ n474 ;
  assign n5078 = n5077 ^ n1189 ^ 1'b0 ;
  assign n5079 = ~n3993 & n5078 ;
  assign n5080 = n1120 & ~n1663 ;
  assign n5081 = n1721 & n5080 ;
  assign n5082 = n3783 & ~n5081 ;
  assign n5083 = ~n4395 & n5082 ;
  assign n5084 = n668 & n2058 ;
  assign n5085 = n5084 ^ n2966 ^ 1'b0 ;
  assign n5087 = x26 & ~n3999 ;
  assign n5088 = n4521 & n5087 ;
  assign n5089 = n964 | n5088 ;
  assign n5086 = n1711 & n4260 ;
  assign n5090 = n5089 ^ n5086 ^ 1'b0 ;
  assign n5092 = n4186 ^ n930 ^ 1'b0 ;
  assign n5093 = n5092 ^ n2693 ^ 1'b0 ;
  assign n5091 = n3012 ^ n2318 ^ 1'b0 ;
  assign n5094 = n5093 ^ n5091 ^ n1025 ;
  assign n5095 = x23 | n1163 ;
  assign n5096 = n5095 ^ n982 ^ 1'b0 ;
  assign n5097 = n5096 ^ n3763 ^ n2871 ;
  assign n5098 = n1519 & n2388 ;
  assign n5099 = ( n630 & n2798 ) | ( n630 & n4985 ) | ( n2798 & n4985 ) ;
  assign n5100 = n2028 & n2069 ;
  assign n5101 = n5100 ^ n725 ^ 1'b0 ;
  assign n5102 = n2091 & n5101 ;
  assign n5103 = n1644 & ~n1936 ;
  assign n5104 = n2204 & n4931 ;
  assign n5105 = ~n5103 & n5104 ;
  assign n5106 = n3209 ^ n1907 ^ 1'b0 ;
  assign n5107 = n886 ^ x17 ^ 1'b0 ;
  assign n5108 = n3012 ^ n413 ^ 1'b0 ;
  assign n5109 = ~n677 & n5108 ;
  assign n5110 = n5109 ^ n2111 ^ 1'b0 ;
  assign n5111 = n2241 & n5110 ;
  assign n5112 = n1661 & n5111 ;
  assign n5113 = n3304 ^ n773 ^ 1'b0 ;
  assign n5114 = n5113 ^ n4123 ^ 1'b0 ;
  assign n5115 = ~n1077 & n1147 ;
  assign n5116 = n5115 ^ n265 ^ 1'b0 ;
  assign n5117 = ( ~n1072 & n1706 ) | ( ~n1072 & n5116 ) | ( n1706 & n5116 ) ;
  assign n5118 = ~n1905 & n5117 ;
  assign n5119 = n241 | n4939 ;
  assign n5120 = n3185 ^ n990 ^ 1'b0 ;
  assign n5121 = n3137 & n5120 ;
  assign n5122 = n4487 ^ x70 ^ 1'b0 ;
  assign n5125 = n2234 & n4384 ;
  assign n5124 = n480 | n3537 ;
  assign n5123 = ~n369 & n928 ;
  assign n5126 = n5125 ^ n5124 ^ n5123 ;
  assign n5127 = ( n844 & n2906 ) | ( n844 & ~n5126 ) | ( n2906 & ~n5126 ) ;
  assign n5129 = n452 ^ n451 ^ 1'b0 ;
  assign n5128 = n4373 ^ n2755 ^ n2376 ;
  assign n5130 = n5129 ^ n5128 ^ 1'b0 ;
  assign n5132 = ( n824 & n1373 ) | ( n824 & ~n2852 ) | ( n1373 & ~n2852 ) ;
  assign n5131 = n608 & ~n1337 ;
  assign n5133 = n5132 ^ n5131 ^ 1'b0 ;
  assign n5136 = n1953 ^ x18 ^ 1'b0 ;
  assign n5137 = ~n2297 & n5136 ;
  assign n5134 = n3828 ^ n2077 ^ 1'b0 ;
  assign n5135 = ~n2164 & n5134 ;
  assign n5138 = n5137 ^ n5135 ^ 1'b0 ;
  assign n5140 = n2323 ^ n2302 ^ 1'b0 ;
  assign n5141 = n2055 & ~n5140 ;
  assign n5139 = n245 & ~n1226 ;
  assign n5142 = n5141 ^ n5139 ^ 1'b0 ;
  assign n5143 = n188 & n5084 ;
  assign n5144 = n5143 ^ x2 ^ 1'b0 ;
  assign n5145 = n2829 & ~n4879 ;
  assign n5146 = n1016 | n5145 ;
  assign n5147 = n5146 ^ n3763 ^ 1'b0 ;
  assign n5148 = ~n4333 & n5147 ;
  assign n5149 = ~n5144 & n5148 ;
  assign n5150 = n3488 ^ n3209 ^ 1'b0 ;
  assign n5151 = n367 ^ x52 ^ 1'b0 ;
  assign n5152 = n3760 & n5151 ;
  assign n5153 = n507 & ~n828 ;
  assign n5154 = n5153 ^ n804 ^ 1'b0 ;
  assign n5155 = ( n3184 & n4667 ) | ( n3184 & n5154 ) | ( n4667 & n5154 ) ;
  assign n5156 = ( n2898 & n4578 ) | ( n2898 & ~n5155 ) | ( n4578 & ~n5155 ) ;
  assign n5157 = n1316 & ~n1987 ;
  assign n5158 = n635 & n5157 ;
  assign n5159 = n5158 ^ n2727 ^ 1'b0 ;
  assign n5160 = n1284 & n5159 ;
  assign n5161 = n1245 ^ n221 ^ 1'b0 ;
  assign n5162 = n560 & n5010 ;
  assign n5163 = n5162 ^ x53 ^ 1'b0 ;
  assign n5164 = n5163 ^ n2544 ^ 1'b0 ;
  assign n5165 = ~n4455 & n5164 ;
  assign n5166 = ( n2340 & n2484 ) | ( n2340 & ~n5165 ) | ( n2484 & ~n5165 ) ;
  assign n5167 = n1307 | n5166 ;
  assign n5168 = n4359 & ~n5167 ;
  assign n5169 = ( n1540 & n3053 ) | ( n1540 & ~n4243 ) | ( n3053 & ~n4243 ) ;
  assign n5170 = n1486 | n2652 ;
  assign n5171 = n5170 ^ x124 ^ 1'b0 ;
  assign n5172 = n5171 ^ n3474 ^ 1'b0 ;
  assign n5173 = ~n3167 & n5172 ;
  assign n5175 = n4358 ^ n2618 ^ n1624 ;
  assign n5174 = n1843 | n3956 ;
  assign n5176 = n5175 ^ n5174 ^ 1'b0 ;
  assign n5178 = n1311 | n1446 ;
  assign n5179 = n5178 ^ n3900 ^ n3236 ;
  assign n5177 = n805 ^ n293 ^ 1'b0 ;
  assign n5180 = n5179 ^ n5177 ^ 1'b0 ;
  assign n5181 = x102 & n5180 ;
  assign n5182 = n1819 ^ n1218 ^ 1'b0 ;
  assign n5183 = x95 & n5182 ;
  assign n5184 = ~n4485 & n5183 ;
  assign n5185 = n5184 ^ n4737 ^ 1'b0 ;
  assign n5186 = n4796 ^ n2552 ^ 1'b0 ;
  assign n5187 = n950 & n5186 ;
  assign n5188 = ~n947 & n5187 ;
  assign n5189 = ( n1461 & n1644 ) | ( n1461 & n2474 ) | ( n1644 & n2474 ) ;
  assign n5190 = n3565 & n5189 ;
  assign n5191 = n5188 | n5190 ;
  assign n5192 = n1061 & ~n2547 ;
  assign n5193 = n5192 ^ n3005 ^ 1'b0 ;
  assign n5194 = ( ~n1649 & n3746 ) | ( ~n1649 & n5193 ) | ( n3746 & n5193 ) ;
  assign n5195 = n2046 & ~n2277 ;
  assign n5196 = ~n1476 & n5195 ;
  assign n5197 = n570 & ~n4650 ;
  assign n5198 = n707 & n5197 ;
  assign n5199 = n2453 & ~n5198 ;
  assign n5200 = n3285 ^ n1832 ^ 1'b0 ;
  assign n5201 = n2149 & n5200 ;
  assign n5202 = n2914 & n5201 ;
  assign n5203 = n4447 & n5202 ;
  assign n5204 = ~n1200 & n1931 ;
  assign n5205 = n5070 ^ n4091 ^ n1687 ;
  assign n5206 = n5205 ^ n4260 ^ 1'b0 ;
  assign n5207 = ( n998 & n3226 ) | ( n998 & ~n3324 ) | ( n3226 & ~n3324 ) ;
  assign n5208 = n5207 ^ n2112 ^ x113 ;
  assign n5209 = n676 | n1893 ;
  assign n5210 = n5208 | n5209 ;
  assign n5211 = n5210 ^ n1695 ^ 1'b0 ;
  assign n5212 = n5211 ^ n2390 ^ n1475 ;
  assign n5213 = n2681 ^ x121 ^ 1'b0 ;
  assign n5214 = n497 & ~n4895 ;
  assign n5215 = ~n1192 & n5214 ;
  assign n5216 = ( ~n3844 & n5213 ) | ( ~n3844 & n5215 ) | ( n5213 & n5215 ) ;
  assign n5217 = n4320 & n4568 ;
  assign n5218 = n4316 & n5217 ;
  assign n5219 = ( ~n505 & n811 ) | ( ~n505 & n1819 ) | ( n811 & n1819 ) ;
  assign n5220 = n422 & ~n932 ;
  assign n5221 = n5220 ^ n332 ^ 1'b0 ;
  assign n5222 = n2665 ^ n933 ^ 1'b0 ;
  assign n5223 = ( n449 & ~n2070 ) | ( n449 & n2985 ) | ( ~n2070 & n2985 ) ;
  assign n5224 = n2710 ^ n130 ^ 1'b0 ;
  assign n5225 = n4146 | n4725 ;
  assign n5226 = n869 & n4000 ;
  assign n5227 = n954 & n5226 ;
  assign n5228 = n247 ^ n189 ^ 1'b0 ;
  assign n5229 = n1256 | n5228 ;
  assign n5230 = n4199 ^ n1492 ^ 1'b0 ;
  assign n5231 = n848 & n5230 ;
  assign n5232 = n5017 ^ n1278 ^ 1'b0 ;
  assign n5233 = n386 & n5232 ;
  assign n5234 = n3641 ^ n3563 ^ 1'b0 ;
  assign n5235 = n5233 & n5234 ;
  assign n5236 = ( n1313 & n1765 ) | ( n1313 & ~n3827 ) | ( n1765 & ~n3827 ) ;
  assign n5237 = n1324 | n3399 ;
  assign n5238 = n2197 & ~n3657 ;
  assign n5239 = n1584 & ~n5238 ;
  assign n5240 = n5239 ^ n2411 ^ 1'b0 ;
  assign n5241 = n4395 ^ n3869 ^ n2236 ;
  assign n5242 = n301 | n5241 ;
  assign n5243 = ( n159 & n2495 ) | ( n159 & n3716 ) | ( n2495 & n3716 ) ;
  assign n5244 = n3696 ^ n1271 ^ 1'b0 ;
  assign n5245 = ~n1639 & n5244 ;
  assign n5246 = n4053 & n5245 ;
  assign n5247 = n4618 ^ n3439 ^ 1'b0 ;
  assign n5248 = n2534 & ~n3249 ;
  assign n5249 = n5248 ^ n1799 ^ 1'b0 ;
  assign n5250 = ( n739 & n3612 ) | ( n739 & n5249 ) | ( n3612 & n5249 ) ;
  assign n5251 = n3256 | n5250 ;
  assign n5252 = n4149 ^ n4115 ^ 1'b0 ;
  assign n5253 = n4811 & ~n5252 ;
  assign n5254 = ~n3067 & n3125 ;
  assign n5255 = n1853 & n5254 ;
  assign n5256 = n4903 ^ n4870 ^ x77 ;
  assign n5257 = n256 & ~n4375 ;
  assign n5258 = ~n5256 & n5257 ;
  assign n5261 = n4194 ^ n1842 ^ n711 ;
  assign n5259 = ( n179 & n676 ) | ( n179 & ~n1673 ) | ( n676 & ~n1673 ) ;
  assign n5260 = n4439 | n5259 ;
  assign n5262 = n5261 ^ n5260 ^ 1'b0 ;
  assign n5263 = n429 & n607 ;
  assign n5264 = ~n2295 & n5263 ;
  assign n5265 = n5219 ^ n2506 ^ 1'b0 ;
  assign n5266 = n3171 ^ n2660 ^ 1'b0 ;
  assign n5267 = n462 & ~n2382 ;
  assign n5268 = n752 | n5267 ;
  assign n5269 = n5268 ^ n1721 ^ 1'b0 ;
  assign n5270 = ~n1656 & n4478 ;
  assign n5271 = n5270 ^ x36 ^ 1'b0 ;
  assign n5272 = n3025 | n5271 ;
  assign n5273 = n1976 & ~n5272 ;
  assign n5274 = n3572 ^ n1843 ^ 1'b0 ;
  assign n5275 = n4600 & ~n5274 ;
  assign n5276 = n955 & ~n4574 ;
  assign n5277 = n5276 ^ n3952 ^ 1'b0 ;
  assign n5278 = n5277 ^ n536 ^ 1'b0 ;
  assign n5279 = n828 & n3482 ;
  assign n5280 = n519 ^ x32 ^ 1'b0 ;
  assign n5281 = n276 & n5280 ;
  assign n5282 = n5281 ^ n191 ^ 1'b0 ;
  assign n5283 = n1603 ^ n1203 ^ 1'b0 ;
  assign n5284 = n5283 ^ n2910 ^ 1'b0 ;
  assign n5285 = n1571 ^ n328 ^ 1'b0 ;
  assign n5286 = n5056 ^ n2214 ^ 1'b0 ;
  assign n5287 = n4202 ^ n612 ^ 1'b0 ;
  assign n5288 = n1439 | n5287 ;
  assign n5289 = n143 | n2222 ;
  assign n5290 = n5289 ^ n2517 ^ n1589 ;
  assign n5291 = n3158 | n5290 ;
  assign n5292 = n5288 | n5291 ;
  assign n5293 = n1954 | n2397 ;
  assign n5294 = n338 | n5293 ;
  assign n5295 = n5294 ^ n1915 ^ 1'b0 ;
  assign n5296 = n1079 & n3626 ;
  assign n5297 = n5296 ^ n1413 ^ n955 ;
  assign n5298 = ( n327 & ~n387 ) | ( n327 & n3291 ) | ( ~n387 & n3291 ) ;
  assign n5299 = ~n1821 & n3743 ;
  assign n5300 = ~n1025 & n5299 ;
  assign n5302 = x12 & n2302 ;
  assign n5303 = n5302 ^ n2517 ^ 1'b0 ;
  assign n5301 = ~n199 & n1513 ;
  assign n5304 = n5303 ^ n5301 ^ 1'b0 ;
  assign n5305 = n5304 ^ n2906 ^ n2720 ;
  assign n5306 = ( n527 & n1290 ) | ( n527 & n5305 ) | ( n1290 & n5305 ) ;
  assign n5307 = n3513 ^ n2255 ^ 1'b0 ;
  assign n5308 = n1583 & n5307 ;
  assign n5309 = n493 & ~n3589 ;
  assign n5310 = n2754 & n5309 ;
  assign n5311 = n2132 ^ n398 ^ 1'b0 ;
  assign n5312 = n4160 & ~n5311 ;
  assign n5313 = n701 | n3663 ;
  assign n5314 = n4691 | n5313 ;
  assign n5315 = ~n508 & n5314 ;
  assign n5316 = ~n3792 & n5315 ;
  assign n5317 = n306 | n1171 ;
  assign n5318 = n3276 | n5317 ;
  assign n5319 = n1000 ^ x33 ^ 1'b0 ;
  assign n5320 = n5318 & ~n5319 ;
  assign n5321 = ~n1171 & n4693 ;
  assign n5329 = n1938 ^ n945 ^ 1'b0 ;
  assign n5330 = n2779 & ~n5329 ;
  assign n5322 = n3540 | n4207 ;
  assign n5323 = n5322 ^ n2039 ^ 1'b0 ;
  assign n5325 = n498 | n1451 ;
  assign n5326 = n5325 ^ n1095 ^ 1'b0 ;
  assign n5324 = n2972 ^ n723 ^ 1'b0 ;
  assign n5327 = n5326 ^ n5324 ^ x126 ;
  assign n5328 = ( n2172 & n5323 ) | ( n2172 & ~n5327 ) | ( n5323 & ~n5327 ) ;
  assign n5331 = n5330 ^ n5328 ^ n1982 ;
  assign n5332 = n2478 ^ n1025 ^ 1'b0 ;
  assign n5333 = x55 & ~n5332 ;
  assign n5334 = n1341 ^ n319 ^ 1'b0 ;
  assign n5335 = ~n3823 & n5334 ;
  assign n5336 = n5335 ^ n1991 ^ 1'b0 ;
  assign n5337 = n2149 & ~n2767 ;
  assign n5338 = ~n5336 & n5337 ;
  assign n5339 = n2821 & ~n5338 ;
  assign n5340 = n5339 ^ n1668 ^ 1'b0 ;
  assign n5341 = n308 & ~n346 ;
  assign n5342 = n5341 ^ n4239 ^ 1'b0 ;
  assign n5343 = n5278 ^ n5142 ^ 1'b0 ;
  assign n5344 = n5342 | n5343 ;
  assign n5352 = n3389 ^ n1669 ^ x88 ;
  assign n5347 = n575 ^ n395 ^ 1'b0 ;
  assign n5345 = n1794 ^ n1338 ^ 1'b0 ;
  assign n5346 = ~n3478 & n5345 ;
  assign n5348 = n5347 ^ n5346 ^ 1'b0 ;
  assign n5349 = n4669 | n5348 ;
  assign n5350 = n3849 & ~n5349 ;
  assign n5351 = n5350 ^ n5335 ^ 1'b0 ;
  assign n5353 = n5352 ^ n5351 ^ 1'b0 ;
  assign n5354 = n4613 ^ n1077 ^ 1'b0 ;
  assign n5355 = n4699 | n5354 ;
  assign n5359 = n1150 | n1658 ;
  assign n5356 = n3743 ^ n1264 ^ 1'b0 ;
  assign n5357 = n5356 ^ n454 ^ 1'b0 ;
  assign n5358 = ~n4746 & n5357 ;
  assign n5360 = n5359 ^ n5358 ^ 1'b0 ;
  assign n5361 = n1496 ^ n1326 ^ 1'b0 ;
  assign n5362 = ~n740 & n2772 ;
  assign n5363 = n5362 ^ n3362 ^ 1'b0 ;
  assign n5364 = n5361 & n5363 ;
  assign n5365 = ~n2256 & n5364 ;
  assign n5366 = n1810 & n4115 ;
  assign n5367 = n5366 ^ n4704 ^ 1'b0 ;
  assign n5368 = n5144 ^ n3525 ^ 1'b0 ;
  assign n5369 = n1250 & n5368 ;
  assign n5370 = n5369 ^ x81 ^ 1'b0 ;
  assign n5371 = ~n3055 & n5370 ;
  assign n5372 = n631 & n2485 ;
  assign n5373 = n5372 ^ n1736 ^ 1'b0 ;
  assign n5374 = n5373 ^ n1780 ^ 1'b0 ;
  assign n5375 = ~n1150 & n5374 ;
  assign n5376 = ~n4027 & n5375 ;
  assign n5377 = n411 ^ n276 ^ 1'b0 ;
  assign n5378 = n5377 ^ n663 ^ n193 ;
  assign n5379 = n3938 ^ n1239 ^ n379 ;
  assign n5380 = n2355 | n5379 ;
  assign n5381 = n5380 ^ n4806 ^ 1'b0 ;
  assign n5382 = ( ~n1714 & n2738 ) | ( ~n1714 & n5381 ) | ( n2738 & n5381 ) ;
  assign n5383 = n150 & n3077 ;
  assign n5384 = n5382 & n5383 ;
  assign n5385 = ~n3560 & n5384 ;
  assign n5386 = n256 | n3672 ;
  assign n5387 = n1660 & ~n5386 ;
  assign n5388 = n672 ^ n457 ^ 1'b0 ;
  assign n5389 = ~n2253 & n5388 ;
  assign n5390 = n928 | n1124 ;
  assign n5391 = n1219 & ~n5390 ;
  assign n5392 = n5389 | n5391 ;
  assign n5393 = n1911 ^ n932 ^ 1'b0 ;
  assign n5394 = n1267 | n5393 ;
  assign n5395 = ~n2346 & n3847 ;
  assign n5396 = ( n1175 & n1181 ) | ( n1175 & n5395 ) | ( n1181 & n5395 ) ;
  assign n5397 = ( ~n1206 & n5394 ) | ( ~n1206 & n5396 ) | ( n5394 & n5396 ) ;
  assign n5398 = n3961 & n4599 ;
  assign n5399 = n1191 ^ n744 ^ 1'b0 ;
  assign n5400 = ( ~n3181 & n3673 ) | ( ~n3181 & n4827 ) | ( n3673 & n4827 ) ;
  assign n5401 = n1600 ^ n1323 ^ 1'b0 ;
  assign n5402 = ~n3984 & n5401 ;
  assign n5403 = n5400 & n5402 ;
  assign n5404 = n5399 & n5403 ;
  assign n5405 = n2094 | n2836 ;
  assign n5406 = n3614 & ~n5405 ;
  assign n5407 = ( n2681 & n3371 ) | ( n2681 & ~n5406 ) | ( n3371 & ~n5406 ) ;
  assign n5408 = n2625 | n5407 ;
  assign n5409 = n4428 | n5408 ;
  assign n5410 = n4220 ^ n2887 ^ n730 ;
  assign n5411 = n1760 ^ n943 ^ 1'b0 ;
  assign n5412 = n282 & ~n5411 ;
  assign n5413 = ( n2375 & n2508 ) | ( n2375 & ~n3119 ) | ( n2508 & ~n3119 ) ;
  assign n5414 = x34 & n5413 ;
  assign n5415 = ( ~n2271 & n2316 ) | ( ~n2271 & n3192 ) | ( n2316 & n3192 ) ;
  assign n5416 = n4606 ^ n1815 ^ 1'b0 ;
  assign n5417 = n3531 ^ n1854 ^ 1'b0 ;
  assign n5418 = ( n1646 & ~n4406 ) | ( n1646 & n5417 ) | ( ~n4406 & n5417 ) ;
  assign n5419 = n5418 ^ n967 ^ 1'b0 ;
  assign n5420 = n3599 ^ n1414 ^ 1'b0 ;
  assign n5421 = ~n564 & n5420 ;
  assign n5422 = n3414 & ~n4337 ;
  assign n5423 = n2921 & n5422 ;
  assign n5424 = n2678 ^ n1631 ^ 1'b0 ;
  assign n5425 = x8 & ~n5424 ;
  assign n5426 = n5425 ^ n4689 ^ 1'b0 ;
  assign n5427 = ~n375 & n5426 ;
  assign n5428 = ~n829 & n5427 ;
  assign n5429 = n5428 ^ n264 ^ 1'b0 ;
  assign n5430 = n1798 & n4663 ;
  assign n5431 = n4815 & n5430 ;
  assign n5432 = n4019 ^ n322 ^ 1'b0 ;
  assign n5433 = ~n1880 & n5432 ;
  assign n5434 = ( ~n1854 & n5431 ) | ( ~n1854 & n5433 ) | ( n5431 & n5433 ) ;
  assign n5435 = x7 & ~n1592 ;
  assign n5436 = n1083 & n5116 ;
  assign n5437 = ~n5435 & n5436 ;
  assign n5438 = n1026 & ~n2492 ;
  assign n5439 = ~n2823 & n5438 ;
  assign n5440 = n5439 ^ n3680 ^ 1'b0 ;
  assign n5441 = ( n3868 & n4561 ) | ( n3868 & ~n5440 ) | ( n4561 & ~n5440 ) ;
  assign n5442 = ~n485 & n2404 ;
  assign n5443 = n5442 ^ n1473 ^ 1'b0 ;
  assign n5444 = n5326 ^ n3900 ^ 1'b0 ;
  assign n5445 = n5443 & ~n5444 ;
  assign n5446 = n4835 & n5445 ;
  assign n5447 = n3893 ^ n2359 ^ n663 ;
  assign n5448 = n5447 ^ n4410 ^ n3630 ;
  assign n5449 = n5448 ^ n3709 ^ 1'b0 ;
  assign n5450 = n3492 ^ n1938 ^ 1'b0 ;
  assign n5451 = n2897 | n5450 ;
  assign n5452 = n5451 ^ n4276 ^ 1'b0 ;
  assign n5453 = n2861 & ~n5452 ;
  assign n5454 = n5453 ^ n3335 ^ 1'b0 ;
  assign n5455 = n4857 ^ n1624 ^ 1'b0 ;
  assign n5456 = n3942 & ~n5455 ;
  assign n5457 = n4026 ^ n872 ^ x87 ;
  assign n5458 = n5457 ^ n4656 ^ 1'b0 ;
  assign n5459 = ( ~x57 & n603 ) | ( ~x57 & n2588 ) | ( n603 & n2588 ) ;
  assign n5460 = n4237 & ~n5459 ;
  assign n5461 = n5460 ^ n3976 ^ 1'b0 ;
  assign n5462 = ~n2692 & n5461 ;
  assign n5463 = n3934 & n5462 ;
  assign n5464 = n965 ^ n833 ^ n155 ;
  assign n5465 = n1581 & n5464 ;
  assign n5466 = n5463 & n5465 ;
  assign n5470 = ~n1732 & n4614 ;
  assign n5467 = ~n1356 & n1424 ;
  assign n5468 = n5467 ^ x49 ^ 1'b0 ;
  assign n5469 = n3691 & ~n5468 ;
  assign n5471 = n5470 ^ n5469 ^ 1'b0 ;
  assign n5472 = ( n674 & n5371 ) | ( n674 & ~n5471 ) | ( n5371 & ~n5471 ) ;
  assign n5473 = n1435 & ~n2326 ;
  assign n5474 = n248 & ~n2216 ;
  assign n5475 = n4024 & ~n5474 ;
  assign n5476 = n2620 ^ n2492 ^ 1'b0 ;
  assign n5477 = ~n2495 & n5476 ;
  assign n5478 = n3636 ^ n387 ^ 1'b0 ;
  assign n5479 = n5453 | n5478 ;
  assign n5480 = n1499 ^ n673 ^ 1'b0 ;
  assign n5481 = n516 & n5480 ;
  assign n5482 = n2287 & n5481 ;
  assign n5483 = n5043 ^ x57 ^ 1'b0 ;
  assign n5487 = ~n2142 & n4663 ;
  assign n5485 = n2827 | n4106 ;
  assign n5484 = n1399 | n2632 ;
  assign n5486 = n5485 ^ n5484 ^ 1'b0 ;
  assign n5488 = n5487 ^ n5486 ^ 1'b0 ;
  assign n5489 = n381 & n3910 ;
  assign n5490 = n5489 ^ n1943 ^ 1'b0 ;
  assign n5491 = n2661 | n5490 ;
  assign n5492 = n2339 ^ n1582 ^ 1'b0 ;
  assign n5493 = ( n844 & n977 ) | ( n844 & ~n5492 ) | ( n977 & ~n5492 ) ;
  assign n5494 = n3479 ^ n1824 ^ 1'b0 ;
  assign n5495 = n454 & n5494 ;
  assign n5496 = n5495 ^ x39 ^ 1'b0 ;
  assign n5497 = ~n3766 & n5496 ;
  assign n5498 = n4436 ^ n1489 ^ 1'b0 ;
  assign n5499 = n220 | n5498 ;
  assign n5500 = ~n1185 & n4560 ;
  assign n5501 = n555 & n5500 ;
  assign n5503 = n4020 & ~n4125 ;
  assign n5502 = ~n1101 & n1586 ;
  assign n5504 = n5503 ^ n5502 ^ 1'b0 ;
  assign n5505 = n2184 | n5504 ;
  assign n5506 = n3679 & n5505 ;
  assign n5507 = n5506 ^ n3038 ^ 1'b0 ;
  assign n5508 = ~n4088 & n4625 ;
  assign n5509 = n1634 & n5508 ;
  assign n5510 = n5507 | n5509 ;
  assign n5511 = n5501 & ~n5510 ;
  assign n5512 = n594 ^ n558 ^ 1'b0 ;
  assign n5513 = n1697 & ~n5512 ;
  assign n5514 = n2398 & n5513 ;
  assign n5515 = n5514 ^ n2738 ^ n359 ;
  assign n5516 = n539 & ~n1514 ;
  assign n5517 = ~n840 & n5516 ;
  assign n5518 = n2552 & n5517 ;
  assign n5519 = ~n2839 & n5518 ;
  assign n5520 = n2819 | n5519 ;
  assign n5521 = n2102 | n2531 ;
  assign n5522 = n5521 ^ n4522 ^ 1'b0 ;
  assign n5523 = x25 & n5522 ;
  assign n5524 = ( x29 & ~n5520 ) | ( x29 & n5523 ) | ( ~n5520 & n5523 ) ;
  assign n5525 = n692 & n3345 ;
  assign n5530 = ( n500 & ~n935 ) | ( n500 & n3185 ) | ( ~n935 & n3185 ) ;
  assign n5526 = n2782 ^ n2543 ^ 1'b0 ;
  assign n5527 = n3037 & n5526 ;
  assign n5528 = n2909 & ~n3524 ;
  assign n5529 = ~n5527 & n5528 ;
  assign n5531 = n5530 ^ n5529 ^ 1'b0 ;
  assign n5532 = ~n5525 & n5531 ;
  assign n5533 = n2223 & n5532 ;
  assign n5534 = x83 & ~n762 ;
  assign n5535 = n2777 ^ n1305 ^ 1'b0 ;
  assign n5536 = ( n769 & ~n1599 ) | ( n769 & n4502 ) | ( ~n1599 & n4502 ) ;
  assign n5537 = n1652 & n2907 ;
  assign n5538 = n5536 & n5537 ;
  assign n5539 = ( n3153 & n5535 ) | ( n3153 & n5538 ) | ( n5535 & n5538 ) ;
  assign n5540 = n5534 & ~n5539 ;
  assign n5541 = n5540 ^ n494 ^ 1'b0 ;
  assign n5542 = n5541 ^ n1848 ^ 1'b0 ;
  assign n5543 = ~n2863 & n3139 ;
  assign n5544 = n5543 ^ n325 ^ 1'b0 ;
  assign n5545 = n5544 ^ n563 ^ 1'b0 ;
  assign n5546 = n2980 ^ n1193 ^ 1'b0 ;
  assign n5547 = n5546 ^ n3926 ^ 1'b0 ;
  assign n5548 = n3615 & ~n4880 ;
  assign n5549 = n1648 & ~n3232 ;
  assign n5550 = n2553 ^ n386 ^ 1'b0 ;
  assign n5551 = n1237 & ~n5550 ;
  assign n5552 = ~n4121 & n5551 ;
  assign n5553 = n5552 ^ n3082 ^ n1234 ;
  assign n5554 = n450 & ~n2152 ;
  assign n5555 = n893 ^ n830 ^ 1'b0 ;
  assign n5556 = n5554 & n5555 ;
  assign n5557 = n1519 ^ n135 ^ 1'b0 ;
  assign n5558 = ~n4359 & n5557 ;
  assign n5559 = ~n3489 & n5558 ;
  assign n5560 = n2866 ^ n1842 ^ 1'b0 ;
  assign n5561 = n1171 | n5560 ;
  assign n5562 = n1710 & n5561 ;
  assign n5563 = ( n1387 & ~n2170 ) | ( n1387 & n2214 ) | ( ~n2170 & n2214 ) ;
  assign n5564 = ~n2681 & n5563 ;
  assign n5565 = ~n3058 & n5564 ;
  assign n5566 = ~n616 & n1585 ;
  assign n5567 = ~n403 & n5566 ;
  assign n5568 = n638 | n3429 ;
  assign n5569 = n5568 ^ n1594 ^ 1'b0 ;
  assign n5570 = ~n2973 & n5569 ;
  assign n5571 = n5570 ^ n2005 ^ 1'b0 ;
  assign n5572 = x13 | n4071 ;
  assign n5573 = n508 & ~n1292 ;
  assign n5574 = n2679 | n5573 ;
  assign n5575 = n1509 | n5574 ;
  assign n5576 = n3380 & n5575 ;
  assign n5577 = ~n370 & n5576 ;
  assign n5578 = n276 & n1380 ;
  assign n5579 = n5578 ^ n3747 ^ 1'b0 ;
  assign n5580 = ~n454 & n5579 ;
  assign n5582 = n2726 | n4055 ;
  assign n5583 = n2146 & ~n5582 ;
  assign n5581 = n2837 ^ n2169 ^ 1'b0 ;
  assign n5584 = n5583 ^ n5581 ^ 1'b0 ;
  assign n5585 = n4443 ^ n2001 ^ 1'b0 ;
  assign n5586 = n129 | n5585 ;
  assign n5587 = ( n2204 & n5584 ) | ( n2204 & ~n5586 ) | ( n5584 & ~n5586 ) ;
  assign n5588 = n720 & n2845 ;
  assign n5592 = n811 | n2937 ;
  assign n5593 = n586 & n5592 ;
  assign n5594 = ~n2926 & n5593 ;
  assign n5595 = n5594 ^ n470 ^ 1'b0 ;
  assign n5589 = n1116 & ~n2098 ;
  assign n5590 = ~n1918 & n5589 ;
  assign n5591 = n5590 ^ n2692 ^ 1'b0 ;
  assign n5596 = n5595 ^ n5591 ^ 1'b0 ;
  assign n5597 = n3261 ^ n427 ^ 1'b0 ;
  assign n5602 = ( n134 & n208 ) | ( n134 & n442 ) | ( n208 & n442 ) ;
  assign n5603 = n4662 & n5602 ;
  assign n5598 = n1343 ^ n1077 ^ 1'b0 ;
  assign n5599 = n5598 ^ n5346 ^ 1'b0 ;
  assign n5600 = n4214 & n5520 ;
  assign n5601 = n5599 & n5600 ;
  assign n5604 = n5603 ^ n5601 ^ 1'b0 ;
  assign n5605 = n4131 ^ n2632 ^ 1'b0 ;
  assign n5606 = n1373 & n5605 ;
  assign n5608 = n1313 & n2589 ;
  assign n5609 = x87 & n5608 ;
  assign n5607 = x100 & n1637 ;
  assign n5610 = n5609 ^ n5607 ^ 1'b0 ;
  assign n5611 = n3840 & ~n4826 ;
  assign n5612 = ~n3340 & n4567 ;
  assign n5613 = n4162 ^ n671 ^ 1'b0 ;
  assign n5614 = n4509 | n5613 ;
  assign n5615 = n5614 ^ n3567 ^ 1'b0 ;
  assign n5616 = n2929 | n5615 ;
  assign n5617 = n3005 & n3536 ;
  assign n5618 = n1588 & n5617 ;
  assign n5619 = n4481 | n5618 ;
  assign n5620 = n5619 ^ n4683 ^ 1'b0 ;
  assign n5627 = ~n909 & n1100 ;
  assign n5628 = n167 & n5627 ;
  assign n5629 = n5628 ^ n2199 ^ 1'b0 ;
  assign n5630 = n2893 & n5629 ;
  assign n5621 = x72 | n5530 ;
  assign n5622 = n5621 ^ n1614 ^ 1'b0 ;
  assign n5623 = ~n4620 & n5622 ;
  assign n5624 = ~n785 & n5623 ;
  assign n5625 = ~n946 & n5624 ;
  assign n5626 = n5625 ^ n5168 ^ 1'b0 ;
  assign n5631 = n5630 ^ n5626 ^ n2855 ;
  assign n5632 = n3862 ^ n3061 ^ 1'b0 ;
  assign n5633 = n2766 & ~n2979 ;
  assign n5634 = n1591 | n5633 ;
  assign n5635 = n5634 ^ n2089 ^ 1'b0 ;
  assign n5636 = n1599 | n2115 ;
  assign n5637 = n5636 ^ n1427 ^ 1'b0 ;
  assign n5638 = n3066 & n3503 ;
  assign n5639 = n1629 | n5638 ;
  assign n5640 = n2675 & ~n5639 ;
  assign n5641 = n1198 ^ n279 ^ 1'b0 ;
  assign n5642 = ~n3208 & n5641 ;
  assign n5645 = ~n1603 & n2738 ;
  assign n5643 = n2366 ^ n279 ^ 1'b0 ;
  assign n5644 = x63 & n5643 ;
  assign n5646 = n5645 ^ n5644 ^ 1'b0 ;
  assign n5647 = x27 & n5646 ;
  assign n5648 = n5647 ^ n3673 ^ 1'b0 ;
  assign n5649 = n3807 & ~n5648 ;
  assign n5650 = ~n5642 & n5649 ;
  assign n5651 = n935 & ~n994 ;
  assign n5652 = n5651 ^ n3587 ^ 1'b0 ;
  assign n5653 = n934 & ~n5652 ;
  assign n5654 = n5653 ^ n2104 ^ n1278 ;
  assign n5655 = n1420 & n4270 ;
  assign n5656 = n939 & n3373 ;
  assign n5658 = n327 & ~n2276 ;
  assign n5659 = n5658 ^ n1387 ^ 1'b0 ;
  assign n5657 = n2636 ^ x67 ^ 1'b0 ;
  assign n5660 = n5659 ^ n5657 ^ 1'b0 ;
  assign n5661 = n892 & ~n5660 ;
  assign n5662 = n5661 ^ n3608 ^ n1746 ;
  assign n5663 = n1101 ^ x0 ^ 1'b0 ;
  assign n5664 = n2063 & ~n5663 ;
  assign n5665 = n980 & ~n4420 ;
  assign n5666 = n5665 ^ n190 ^ 1'b0 ;
  assign n5667 = ~n3724 & n5666 ;
  assign n5668 = n5667 ^ x14 ^ 1'b0 ;
  assign n5669 = n433 & n5668 ;
  assign n5670 = n2850 ^ n2067 ^ n1217 ;
  assign n5671 = ( n1109 & n1938 ) | ( n1109 & n3838 ) | ( n1938 & n3838 ) ;
  assign n5672 = n1406 & n5671 ;
  assign n5673 = ~n5670 & n5672 ;
  assign n5674 = n1463 & ~n5673 ;
  assign n5675 = n5674 ^ n5098 ^ 1'b0 ;
  assign n5680 = n1621 | n3323 ;
  assign n5676 = n482 ^ x116 ^ 1'b0 ;
  assign n5677 = n1168 & n5676 ;
  assign n5678 = x32 & ~n3204 ;
  assign n5679 = n5677 & n5678 ;
  assign n5681 = n5680 ^ n5679 ^ 1'b0 ;
  assign n5682 = ( n260 & n673 ) | ( n260 & ~n753 ) | ( n673 & ~n753 ) ;
  assign n5683 = n5682 ^ n2836 ^ 1'b0 ;
  assign n5686 = ( n332 & n854 ) | ( n332 & ~n1021 ) | ( n854 & ~n1021 ) ;
  assign n5687 = ( n314 & n1811 ) | ( n314 & n5686 ) | ( n1811 & n5686 ) ;
  assign n5684 = n1752 & ~n1843 ;
  assign n5685 = n5684 ^ n2045 ^ 1'b0 ;
  assign n5688 = n5687 ^ n5685 ^ 1'b0 ;
  assign n5689 = n5683 & ~n5688 ;
  assign n5690 = n2476 & n5689 ;
  assign n5691 = n5690 ^ n4933 ^ 1'b0 ;
  assign n5692 = x64 & n3584 ;
  assign n5693 = n2164 ^ n1714 ^ n1476 ;
  assign n5694 = n1792 & n5693 ;
  assign n5695 = n2517 & n5694 ;
  assign n5696 = n2843 | n5695 ;
  assign n5697 = n3182 ^ n1189 ^ 1'b0 ;
  assign n5698 = ~n3412 & n5697 ;
  assign n5699 = ~n1472 & n5698 ;
  assign n5700 = n1496 & ~n4895 ;
  assign n5701 = n5551 & n5700 ;
  assign n5702 = n4216 & ~n5701 ;
  assign n5703 = n3861 | n4047 ;
  assign n5704 = n241 & n2525 ;
  assign n5705 = n5704 ^ n1476 ^ 1'b0 ;
  assign n5706 = ( n1072 & n4365 ) | ( n1072 & ~n5705 ) | ( n4365 & ~n5705 ) ;
  assign n5707 = n5706 ^ n2206 ^ 1'b0 ;
  assign n5708 = ~n2636 & n5707 ;
  assign n5709 = n2728 & ~n3930 ;
  assign n5710 = n5709 ^ n1489 ^ 1'b0 ;
  assign n5711 = n4443 & n5710 ;
  assign n5713 = n148 | n2652 ;
  assign n5714 = n3599 | n5713 ;
  assign n5712 = n2414 ^ n857 ^ 1'b0 ;
  assign n5715 = n5714 ^ n5712 ^ n4354 ;
  assign n5716 = n1074 & n4075 ;
  assign n5717 = n5584 & n5716 ;
  assign n5718 = n4625 ^ n2293 ^ 1'b0 ;
  assign n5719 = n4748 | n5718 ;
  assign n5720 = n1033 | n5719 ;
  assign n5721 = n5720 ^ n2266 ^ 1'b0 ;
  assign n5722 = n5213 ^ n196 ^ 1'b0 ;
  assign n5723 = ( n220 & ~n1016 ) | ( n220 & n1851 ) | ( ~n1016 & n1851 ) ;
  assign n5724 = ( n2032 & n5501 ) | ( n2032 & n5723 ) | ( n5501 & n5723 ) ;
  assign n5725 = n1827 & n3773 ;
  assign n5726 = n2070 ^ n490 ^ 1'b0 ;
  assign n5727 = n3743 & n3940 ;
  assign n5728 = ~n1580 & n5727 ;
  assign n5729 = n1841 | n2020 ;
  assign n5730 = n5729 ^ n1231 ^ 1'b0 ;
  assign n5731 = ( n259 & n590 ) | ( n259 & n5730 ) | ( n590 & n5730 ) ;
  assign n5732 = ~n179 & n3931 ;
  assign n5733 = n1013 & n5732 ;
  assign n5734 = ( n555 & n5731 ) | ( n555 & ~n5733 ) | ( n5731 & ~n5733 ) ;
  assign n5735 = n260 | n2482 ;
  assign n5736 = n5735 ^ n416 ^ 1'b0 ;
  assign n5737 = n456 & ~n2591 ;
  assign n5738 = ~n5468 & n5737 ;
  assign n5739 = n1610 & n5738 ;
  assign n5740 = ~n3617 & n3967 ;
  assign n5741 = n5740 ^ n3842 ^ x25 ;
  assign n5742 = n3622 ^ n346 ^ 1'b0 ;
  assign n5754 = n3285 ^ n1125 ^ 1'b0 ;
  assign n5755 = ( n2463 & n4320 ) | ( n2463 & n5754 ) | ( n4320 & n5754 ) ;
  assign n5744 = x91 & n2290 ;
  assign n5745 = ~n323 & n5744 ;
  assign n5743 = n1871 & n2484 ;
  assign n5746 = n5745 ^ n5743 ^ 1'b0 ;
  assign n5748 = ~n1837 & n5592 ;
  assign n5749 = n5748 ^ n150 ^ 1'b0 ;
  assign n5747 = n4432 ^ n2830 ^ 1'b0 ;
  assign n5750 = n5749 ^ n5747 ^ n3805 ;
  assign n5751 = n494 | n5750 ;
  assign n5752 = n3942 | n5751 ;
  assign n5753 = ~n5746 & n5752 ;
  assign n5756 = n5755 ^ n5753 ^ 1'b0 ;
  assign n5757 = x121 & ~n1081 ;
  assign n5758 = n3229 & n5757 ;
  assign n5759 = n5381 & ~n5758 ;
  assign n5760 = ~x29 & n5759 ;
  assign n5761 = ( n408 & ~n1082 ) | ( n408 & n2969 ) | ( ~n1082 & n2969 ) ;
  assign n5762 = n1425 | n4815 ;
  assign n5763 = n2409 | n5762 ;
  assign n5764 = ~n1370 & n3372 ;
  assign n5765 = n2330 & n5764 ;
  assign n5766 = n2901 & n3277 ;
  assign n5767 = n5766 ^ n4639 ^ 1'b0 ;
  assign n5768 = ~n2547 & n5767 ;
  assign n5769 = n3797 ^ n1480 ^ 1'b0 ;
  assign n5770 = n5768 | n5769 ;
  assign n5771 = n3224 ^ n1337 ^ 1'b0 ;
  assign n5772 = ( n750 & n4298 ) | ( n750 & n5771 ) | ( n4298 & n5771 ) ;
  assign n5773 = n2541 ^ n1860 ^ 1'b0 ;
  assign n5774 = n2703 ^ n1885 ^ 1'b0 ;
  assign n5775 = n5774 ^ n4449 ^ 1'b0 ;
  assign n5776 = n2857 & n5775 ;
  assign n5777 = n630 & n654 ;
  assign n5778 = n5777 ^ n4173 ^ 1'b0 ;
  assign n5779 = n5567 ^ n4483 ^ 1'b0 ;
  assign n5780 = n5778 & n5779 ;
  assign n5781 = n3752 ^ n1682 ^ 1'b0 ;
  assign n5782 = n5781 ^ n2409 ^ 1'b0 ;
  assign n5783 = n4911 & n5782 ;
  assign n5784 = n5126 ^ n4995 ^ n2258 ;
  assign n5785 = n248 ^ x24 ^ 1'b0 ;
  assign n5786 = n5785 ^ n1980 ^ 1'b0 ;
  assign n5787 = n2638 & n4367 ;
  assign n5788 = ~n2552 & n5787 ;
  assign n5789 = n3861 | n5788 ;
  assign n5790 = n5786 | n5789 ;
  assign n5791 = n854 ^ n478 ^ 1'b0 ;
  assign n5792 = ( n3576 & n5790 ) | ( n3576 & n5791 ) | ( n5790 & n5791 ) ;
  assign n5793 = n758 & ~n4327 ;
  assign n5794 = ~n3476 & n5793 ;
  assign n5795 = n1064 | n1855 ;
  assign n5796 = n5795 ^ n3048 ^ 1'b0 ;
  assign n5797 = n919 & ~n1819 ;
  assign n5798 = n3689 ^ n1009 ^ 1'b0 ;
  assign n5799 = n5797 & n5798 ;
  assign n5800 = n199 & n5799 ;
  assign n5801 = n1791 & ~n2255 ;
  assign n5802 = n5800 & n5801 ;
  assign n5803 = n4186 ^ n635 ^ 1'b0 ;
  assign n5804 = n3116 | n5803 ;
  assign n5805 = n5804 ^ n799 ^ 1'b0 ;
  assign n5806 = n1996 | n2333 ;
  assign n5807 = ~n2440 & n4276 ;
  assign n5808 = n5807 ^ n1880 ^ 1'b0 ;
  assign n5809 = n5808 ^ n1033 ^ 1'b0 ;
  assign n5810 = n5806 & ~n5809 ;
  assign n5811 = ( ~n245 & n2534 ) | ( ~n245 & n5810 ) | ( n2534 & n5810 ) ;
  assign n5812 = n3127 ^ n2420 ^ 1'b0 ;
  assign n5813 = n4720 | n4948 ;
  assign n5814 = n5813 ^ n3107 ^ 1'b0 ;
  assign n5815 = n435 | n4826 ;
  assign n5816 = n3989 ^ n879 ^ 1'b0 ;
  assign n5817 = n4663 ^ n3485 ^ 1'b0 ;
  assign n5818 = n5817 ^ n1585 ^ n189 ;
  assign n5819 = n3306 & n5818 ;
  assign n5820 = n3292 & n5819 ;
  assign n5821 = n5820 ^ n1721 ^ 1'b0 ;
  assign n5822 = n1762 & n5821 ;
  assign n5823 = n690 | n4204 ;
  assign n5824 = n584 & ~n2544 ;
  assign n5825 = ~n2073 & n5824 ;
  assign n5826 = n5825 ^ n3395 ^ 1'b0 ;
  assign n5827 = ~n4150 & n5293 ;
  assign n5828 = ~n3142 & n5101 ;
  assign n5829 = n4503 & n5828 ;
  assign n5830 = n2388 & ~n4442 ;
  assign n5831 = n3340 & n5830 ;
  assign n5832 = ~n1099 & n3230 ;
  assign n5833 = n755 & n5832 ;
  assign n5838 = n3203 ^ n1630 ^ 1'b0 ;
  assign n5839 = n2429 & ~n5838 ;
  assign n5834 = ~n1131 & n1218 ;
  assign n5835 = n2762 ^ x107 ^ 1'b0 ;
  assign n5836 = n5834 & n5835 ;
  assign n5837 = ~n3757 & n5836 ;
  assign n5840 = n5839 ^ n5837 ^ n5255 ;
  assign n5841 = n5840 ^ n3442 ^ n1950 ;
  assign n5842 = ~n1243 & n5841 ;
  assign n5843 = ~n4648 & n5156 ;
  assign n5844 = n5843 ^ n923 ^ 1'b0 ;
  assign n5845 = n5842 & n5844 ;
  assign n5846 = ~n1002 & n3624 ;
  assign n5847 = n592 & n1111 ;
  assign n5848 = ~n261 & n5847 ;
  assign n5849 = n1945 & ~n5848 ;
  assign n5850 = ~n2593 & n5849 ;
  assign n5851 = n5850 ^ n1698 ^ 1'b0 ;
  assign n5852 = n169 | n5851 ;
  assign n5853 = n2922 | n3758 ;
  assign n5854 = n5852 & ~n5853 ;
  assign n5855 = n5352 ^ n3885 ^ 1'b0 ;
  assign n5856 = n1971 | n5855 ;
  assign n5857 = n5856 ^ n431 ^ 1'b0 ;
  assign n5858 = ~n5833 & n5857 ;
  assign n5859 = n3119 ^ n429 ^ 1'b0 ;
  assign n5860 = n3834 & n5859 ;
  assign n5861 = n1014 & n5860 ;
  assign n5862 = ~n471 & n1858 ;
  assign n5863 = ~n1549 & n5862 ;
  assign n5864 = ~n1457 & n5863 ;
  assign n5865 = n5864 ^ n2506 ^ 1'b0 ;
  assign n5866 = ( n786 & ~n4291 ) | ( n786 & n5865 ) | ( ~n4291 & n5865 ) ;
  assign n5867 = n1234 | n1869 ;
  assign n5868 = n1815 | n5867 ;
  assign n5869 = n548 ^ n510 ^ 1'b0 ;
  assign n5870 = n1175 & ~n5869 ;
  assign n5871 = n5868 & n5870 ;
  assign n5872 = n4713 & n5871 ;
  assign n5873 = n452 | n4552 ;
  assign n5874 = n5873 ^ n4984 ^ 1'b0 ;
  assign n5875 = n4115 ^ n1989 ^ n1716 ;
  assign n5876 = n5875 ^ n2796 ^ n1895 ;
  assign n5877 = n722 & ~n1713 ;
  assign n5878 = n974 & n5877 ;
  assign n5880 = n539 & ~n2115 ;
  assign n5881 = n5880 ^ n3834 ^ 1'b0 ;
  assign n5879 = n994 ^ n513 ^ 1'b0 ;
  assign n5882 = n5881 ^ n5879 ^ n452 ;
  assign n5883 = n826 ^ n407 ^ 1'b0 ;
  assign n5884 = n5883 ^ n2001 ^ 1'b0 ;
  assign n5885 = ~n5882 & n5884 ;
  assign n5886 = ~n5878 & n5885 ;
  assign n5887 = n4916 ^ n3952 ^ 1'b0 ;
  assign n5888 = n3844 ^ n2225 ^ 1'b0 ;
  assign n5889 = n3214 ^ n3015 ^ 1'b0 ;
  assign n5890 = ( n4658 & n5312 ) | ( n4658 & ~n5573 ) | ( n5312 & ~n5573 ) ;
  assign n5891 = n5333 ^ n245 ^ 1'b0 ;
  assign n5892 = n765 ^ n141 ^ 1'b0 ;
  assign n5895 = n5335 ^ n1805 ^ 1'b0 ;
  assign n5893 = n2926 ^ n664 ^ 1'b0 ;
  assign n5894 = ~n3643 & n5893 ;
  assign n5896 = n5895 ^ n5894 ^ 1'b0 ;
  assign n5897 = n2426 ^ n134 ^ 1'b0 ;
  assign n5898 = ( ~n1374 & n4088 ) | ( ~n1374 & n4466 ) | ( n4088 & n4466 ) ;
  assign n5899 = ( n1582 & ~n2634 ) | ( n1582 & n5898 ) | ( ~n2634 & n5898 ) ;
  assign n5900 = n2035 ^ n1945 ^ 1'b0 ;
  assign n5902 = n773 ^ n664 ^ x55 ;
  assign n5901 = n4815 ^ n1168 ^ n903 ;
  assign n5903 = n5902 ^ n5901 ^ 1'b0 ;
  assign n5904 = n4209 & ~n5903 ;
  assign n5905 = n395 & n5904 ;
  assign n5906 = ~n5900 & n5905 ;
  assign n5907 = n1791 & n3286 ;
  assign n5908 = ~n1800 & n5907 ;
  assign n5909 = n2612 | n5837 ;
  assign n5910 = n3639 ^ n1656 ^ 1'b0 ;
  assign n5911 = n5910 ^ n3976 ^ n1679 ;
  assign n5912 = n4104 & ~n5896 ;
  assign n5913 = n5912 ^ n1291 ^ 1'b0 ;
  assign n5914 = n842 & n1179 ;
  assign n5915 = ~n1406 & n5914 ;
  assign n5916 = ~n896 & n1617 ;
  assign n5917 = ~n4593 & n5916 ;
  assign n5918 = n5917 ^ n3900 ^ 1'b0 ;
  assign n5919 = n3845 ^ n3452 ^ 1'b0 ;
  assign n5920 = n2758 & n5919 ;
  assign n5921 = n5534 & n5920 ;
  assign n5922 = n5918 & n5921 ;
  assign n5923 = n923 | n3963 ;
  assign n5924 = n2157 | n5923 ;
  assign n5926 = n2636 ^ n1936 ^ 1'b0 ;
  assign n5927 = n1300 & ~n5850 ;
  assign n5928 = n5926 | n5927 ;
  assign n5925 = ~n842 & n1309 ;
  assign n5929 = n5928 ^ n5925 ^ n4846 ;
  assign n5932 = n731 ^ x117 ^ 1'b0 ;
  assign n5933 = n3354 & ~n5932 ;
  assign n5934 = ~n3015 & n5933 ;
  assign n5935 = n5934 ^ n1472 ^ 1'b0 ;
  assign n5936 = ~n2903 & n5935 ;
  assign n5930 = n3354 | n5487 ;
  assign n5931 = n4780 & n5930 ;
  assign n5937 = n5936 ^ n5931 ^ 1'b0 ;
  assign n5938 = n5937 ^ n4857 ^ n4104 ;
  assign n5939 = n5938 ^ n4955 ^ 1'b0 ;
  assign n5940 = x23 & n5939 ;
  assign n5941 = n1856 ^ n801 ^ 1'b0 ;
  assign n5942 = n5941 ^ n4846 ^ n1246 ;
  assign n5943 = n5942 ^ n5471 ^ 1'b0 ;
  assign n5944 = n1599 & ~n5943 ;
  assign n5945 = n1477 & n2368 ;
  assign n5946 = n835 & ~n3202 ;
  assign n5947 = n960 & ~n4191 ;
  assign n5948 = n2802 ^ n2380 ^ 1'b0 ;
  assign n5949 = n5947 & ~n5948 ;
  assign n5950 = n5949 ^ n1608 ^ 1'b0 ;
  assign n5951 = n3519 ^ n1818 ^ n1713 ;
  assign n5952 = ( n925 & n3997 ) | ( n925 & ~n5951 ) | ( n3997 & ~n5951 ) ;
  assign n5953 = n1781 & n3644 ;
  assign n5954 = n3574 & n5953 ;
  assign n5955 = n5952 & n5954 ;
  assign n5956 = n2558 & n4989 ;
  assign n5957 = ~n918 & n5956 ;
  assign n5958 = n5514 ^ n4850 ^ n3943 ;
  assign n5959 = n5958 ^ n4475 ^ 1'b0 ;
  assign n5960 = n1288 ^ n653 ^ n391 ;
  assign n5961 = ~n642 & n5960 ;
  assign n5962 = n5734 & n5961 ;
  assign n5963 = n5641 & n5941 ;
  assign n5964 = n2490 & n4048 ;
  assign n5966 = n1445 & n3149 ;
  assign n5967 = ~n1867 & n5966 ;
  assign n5968 = n678 | n5967 ;
  assign n5965 = n3188 ^ n487 ^ 1'b0 ;
  assign n5969 = n5968 ^ n5965 ^ 1'b0 ;
  assign n5970 = n2921 | n5969 ;
  assign n5971 = n1260 ^ n173 ^ 1'b0 ;
  assign n5972 = ~n4699 & n5971 ;
  assign n5973 = n2334 | n2715 ;
  assign n5974 = n5973 ^ n1399 ^ 1'b0 ;
  assign n5975 = n668 & n5974 ;
  assign n5976 = n1871 & n5975 ;
  assign n5977 = n5976 ^ n1109 ^ 1'b0 ;
  assign n5978 = ~n1879 & n4187 ;
  assign n5979 = n5978 ^ n3380 ^ 1'b0 ;
  assign n5980 = n5979 ^ n1601 ^ 1'b0 ;
  assign n5982 = n1435 & n1800 ;
  assign n5983 = n5982 ^ n1033 ^ 1'b0 ;
  assign n5981 = ~n3057 & n3776 ;
  assign n5984 = n5983 ^ n5981 ^ 1'b0 ;
  assign n5985 = ~n5980 & n5984 ;
  assign n5986 = n5750 ^ n4246 ^ 1'b0 ;
  assign n5987 = n5534 ^ n1753 ^ 1'b0 ;
  assign n5988 = n2782 | n5987 ;
  assign n5989 = n3240 ^ n3121 ^ n1633 ;
  assign n5990 = ( n650 & ~n3845 ) | ( n650 & n5989 ) | ( ~n3845 & n5989 ) ;
  assign n5991 = n1667 ^ n1611 ^ 1'b0 ;
  assign n5992 = n210 & ~n1875 ;
  assign n5993 = n5992 ^ n620 ^ 1'b0 ;
  assign n5994 = ( n2577 & ~n5991 ) | ( n2577 & n5993 ) | ( ~n5991 & n5993 ) ;
  assign n5995 = n273 | n1627 ;
  assign n5996 = ( ~n773 & n845 ) | ( ~n773 & n3022 ) | ( n845 & n3022 ) ;
  assign n5997 = n5996 ^ n872 ^ 1'b0 ;
  assign n5998 = n5997 ^ n2809 ^ 1'b0 ;
  assign n5999 = n5995 | n5998 ;
  assign n6000 = n5999 ^ n1512 ^ n1067 ;
  assign n6001 = n1127 ^ n335 ^ x89 ;
  assign n6002 = n4207 ^ n1626 ^ 1'b0 ;
  assign n6003 = ( n494 & n2449 ) | ( n494 & n6002 ) | ( n2449 & n6002 ) ;
  assign n6004 = ( ~n763 & n6001 ) | ( ~n763 & n6003 ) | ( n6001 & n6003 ) ;
  assign n6005 = n3788 | n3858 ;
  assign n6006 = n507 & n929 ;
  assign n6007 = n6006 ^ n3011 ^ 1'b0 ;
  assign n6008 = n2765 ^ n2033 ^ n621 ;
  assign n6009 = n5778 & n6008 ;
  assign n6010 = ~n6007 & n6009 ;
  assign n6011 = n1721 & ~n3492 ;
  assign n6012 = n6011 ^ n1791 ^ 1'b0 ;
  assign n6013 = n6012 ^ n2343 ^ 1'b0 ;
  assign n6014 = n3586 ^ n1124 ^ 1'b0 ;
  assign n6015 = n586 & n2293 ;
  assign n6016 = n6015 ^ n1408 ^ 1'b0 ;
  assign n6017 = n2155 & n5395 ;
  assign n6018 = ~n1776 & n6017 ;
  assign n6019 = n3020 & ~n6018 ;
  assign n6020 = n6019 ^ n135 ^ 1'b0 ;
  assign n6021 = n1171 ^ n561 ^ 1'b0 ;
  assign n6022 = n4297 | n6021 ;
  assign n6023 = n2342 ^ n1652 ^ 1'b0 ;
  assign n6025 = n1124 | n1198 ;
  assign n6026 = n2016 | n6025 ;
  assign n6024 = ~n2888 & n3795 ;
  assign n6027 = n6026 ^ n6024 ^ 1'b0 ;
  assign n6028 = n6023 & ~n6027 ;
  assign n6029 = n5885 ^ n2759 ^ 1'b0 ;
  assign n6030 = n1749 & n1917 ;
  assign n6031 = n145 & n3076 ;
  assign n6032 = n3583 | n5895 ;
  assign n6033 = n6031 | n6032 ;
  assign n6034 = n3044 & ~n6033 ;
  assign n6035 = n4805 ^ n3189 ^ 1'b0 ;
  assign n6036 = x20 | n2887 ;
  assign n6037 = n2152 & ~n6036 ;
  assign n6038 = n933 & n6037 ;
  assign n6039 = n6038 ^ n4675 ^ n3361 ;
  assign n6044 = n5546 ^ n3752 ^ 1'b0 ;
  assign n6045 = n4288 & n6044 ;
  assign n6041 = n1418 ^ n1070 ^ 1'b0 ;
  assign n6042 = n215 | n6041 ;
  assign n6043 = n3476 & ~n6042 ;
  assign n6040 = ( ~n1489 & n2438 ) | ( ~n1489 & n4195 ) | ( n2438 & n4195 ) ;
  assign n6046 = n6045 ^ n6043 ^ n6040 ;
  assign n6047 = ( n3353 & n3929 ) | ( n3353 & ~n4006 ) | ( n3929 & ~n4006 ) ;
  assign n6048 = n3966 & ~n4518 ;
  assign n6049 = n3440 ^ n997 ^ n691 ;
  assign n6050 = n6049 ^ n1324 ^ n1323 ;
  assign n6051 = n3175 & ~n6050 ;
  assign n6052 = n3756 & n6051 ;
  assign n6053 = ( n686 & n6048 ) | ( n686 & ~n6052 ) | ( n6048 & ~n6052 ) ;
  assign n6054 = n5150 ^ n1687 ^ 1'b0 ;
  assign n6055 = n3860 & n6054 ;
  assign n6056 = ~n3320 & n5501 ;
  assign n6057 = n3918 ^ n2886 ^ 1'b0 ;
  assign n6058 = n2094 | n6057 ;
  assign n6059 = n5036 ^ n4076 ^ 1'b0 ;
  assign n6060 = n6058 | n6059 ;
  assign n6061 = n1661 & ~n4005 ;
  assign n6062 = n4368 ^ n2130 ^ 1'b0 ;
  assign n6063 = ~n2645 & n6062 ;
  assign n6064 = n1213 & n6063 ;
  assign n6065 = ~n5592 & n6064 ;
  assign n6066 = ( n5205 & n5871 ) | ( n5205 & n6065 ) | ( n5871 & n6065 ) ;
  assign n6067 = n4247 ^ n1791 ^ n196 ;
  assign n6068 = n1549 | n4487 ;
  assign n6069 = n6068 ^ n3537 ^ 1'b0 ;
  assign n6070 = n1585 & n6069 ;
  assign n6074 = n3584 ^ n1420 ^ 1'b0 ;
  assign n6075 = ~n4716 & n6074 ;
  assign n6076 = n6075 ^ n2006 ^ 1'b0 ;
  assign n6071 = n1401 & ~n5595 ;
  assign n6072 = n6071 ^ n2431 ^ 1'b0 ;
  assign n6073 = ( n372 & n1758 ) | ( n372 & n6072 ) | ( n1758 & n6072 ) ;
  assign n6077 = n6076 ^ n6073 ^ 1'b0 ;
  assign n6078 = n6070 & n6077 ;
  assign n6079 = ~n3363 & n3879 ;
  assign n6080 = n4870 | n6079 ;
  assign n6081 = n6080 ^ n1084 ^ 1'b0 ;
  assign n6082 = n509 & ~n1232 ;
  assign n6083 = n1286 & n6082 ;
  assign n6084 = ~n2733 & n4090 ;
  assign n6085 = n943 & n6084 ;
  assign n6086 = n6083 | n6085 ;
  assign n6087 = n5822 | n6086 ;
  assign n6088 = x66 | n2544 ;
  assign n6089 = n1033 | n2954 ;
  assign n6090 = x20 & ~n6089 ;
  assign n6091 = n2207 & ~n6090 ;
  assign n6092 = n6091 ^ n1848 ^ 1'b0 ;
  assign n6093 = n6092 ^ n4833 ^ 1'b0 ;
  assign n6094 = n188 & n3595 ;
  assign n6095 = n319 & n6094 ;
  assign n6096 = ~n1177 & n5330 ;
  assign n6097 = n6096 ^ n2564 ^ 1'b0 ;
  assign n6098 = n6095 | n6097 ;
  assign n6099 = n6098 ^ n760 ^ 1'b0 ;
  assign n6100 = x84 & ~n1634 ;
  assign n6101 = n6100 ^ n3924 ^ 1'b0 ;
  assign n6102 = n1452 & ~n4525 ;
  assign n6103 = n1016 | n6102 ;
  assign n6104 = n6103 ^ n1171 ^ 1'b0 ;
  assign n6105 = n4895 | n6104 ;
  assign n6106 = n2706 & ~n6105 ;
  assign n6107 = n4065 | n4933 ;
  assign n6108 = n1906 ^ n691 ^ 1'b0 ;
  assign n6109 = n1173 & ~n6108 ;
  assign n6110 = n3216 & n6109 ;
  assign n6111 = n6110 ^ n717 ^ 1'b0 ;
  assign n6112 = ~n3329 & n4468 ;
  assign n6113 = x118 & n306 ;
  assign n6114 = n1387 & n6113 ;
  assign n6115 = n6114 ^ n577 ^ 1'b0 ;
  assign n6116 = n135 & ~n6115 ;
  assign n6117 = n1853 & n1914 ;
  assign n6118 = n1305 ^ n899 ^ 1'b0 ;
  assign n6119 = n1238 & ~n6118 ;
  assign n6120 = ( n499 & ~n1586 ) | ( n499 & n3171 ) | ( ~n1586 & n3171 ) ;
  assign n6121 = n3267 ^ n1264 ^ 1'b0 ;
  assign n6122 = ~n6120 & n6121 ;
  assign n6123 = n6122 ^ n3674 ^ 1'b0 ;
  assign n6124 = n6119 & ~n6123 ;
  assign n6125 = n6124 ^ n1720 ^ 1'b0 ;
  assign n6126 = ~n640 & n6125 ;
  assign n6127 = n2256 ^ n1335 ^ 1'b0 ;
  assign n6128 = ~n2453 & n6127 ;
  assign n6129 = ~n273 & n6128 ;
  assign n6130 = n6129 ^ x88 ^ 1'b0 ;
  assign n6131 = n5715 ^ n2701 ^ x88 ;
  assign n6132 = n967 & ~n3429 ;
  assign n6133 = n2160 ^ n1394 ^ 1'b0 ;
  assign n6134 = ~n1749 & n6133 ;
  assign n6135 = n6134 ^ n1803 ^ 1'b0 ;
  assign n6136 = n1703 & n6135 ;
  assign n6137 = n1097 & ~n3887 ;
  assign n6138 = n6137 ^ n1288 ^ 1'b0 ;
  assign n6139 = n5523 & ~n6138 ;
  assign n6140 = n1134 ^ n1036 ^ 1'b0 ;
  assign n6141 = ~n1396 & n6140 ;
  assign n6142 = n3239 | n6141 ;
  assign n6143 = n6139 & ~n6142 ;
  assign n6144 = ~n3344 & n4995 ;
  assign n6145 = n2051 | n3089 ;
  assign n6146 = n4380 & n6145 ;
  assign n6147 = ~n1261 & n1513 ;
  assign n6148 = n6147 ^ n452 ^ 1'b0 ;
  assign n6149 = ( n3781 & n4357 ) | ( n3781 & ~n6148 ) | ( n4357 & ~n6148 ) ;
  assign n6150 = n425 & n6149 ;
  assign n6151 = ~x30 & n6150 ;
  assign n6152 = n4382 ^ n706 ^ 1'b0 ;
  assign n6153 = ~n236 & n6152 ;
  assign n6154 = n6153 ^ n3627 ^ 1'b0 ;
  assign n6155 = n2597 & n6154 ;
  assign n6156 = n1161 & ~n1973 ;
  assign n6157 = n1692 ^ n1630 ^ 1'b0 ;
  assign n6158 = n1877 | n6157 ;
  assign n6159 = n6158 ^ n2987 ^ 1'b0 ;
  assign n6160 = n3608 & ~n6159 ;
  assign n6161 = n6160 ^ n403 ^ 1'b0 ;
  assign n6162 = ( n487 & ~n6156 ) | ( n487 & n6161 ) | ( ~n6156 & n6161 ) ;
  assign n6163 = n5108 ^ n1186 ^ 1'b0 ;
  assign n6164 = ~n4159 & n6163 ;
  assign n6165 = n3607 ^ n1467 ^ 1'b0 ;
  assign n6166 = ~n1008 & n6165 ;
  assign n6167 = n1760 & n3074 ;
  assign n6168 = ~n6166 & n6167 ;
  assign n6170 = n3738 ^ n1306 ^ 1'b0 ;
  assign n6169 = n129 & n3064 ;
  assign n6171 = n6170 ^ n6169 ^ 1'b0 ;
  assign n6172 = ( n503 & n2406 ) | ( n503 & n3017 ) | ( n2406 & n3017 ) ;
  assign n6173 = n3111 ^ n1817 ^ 1'b0 ;
  assign n6174 = x76 & n6173 ;
  assign n6175 = n1251 & n6174 ;
  assign n6176 = n6175 ^ n5970 ^ 1'b0 ;
  assign n6177 = n3051 | n4333 ;
  assign n6178 = n6177 ^ n1730 ^ 1'b0 ;
  assign n6179 = n6178 ^ x61 ^ 1'b0 ;
  assign n6180 = n6179 ^ n1633 ^ 1'b0 ;
  assign n6181 = n3633 & n6180 ;
  assign n6182 = n1171 & n6181 ;
  assign n6189 = ( n1219 & n1291 ) | ( n1219 & n1572 ) | ( n1291 & n1572 ) ;
  assign n6188 = ~n393 & n925 ;
  assign n6190 = n6189 ^ n6188 ^ 1'b0 ;
  assign n6187 = n1186 & n4833 ;
  assign n6183 = n3304 ^ n3043 ^ 1'b0 ;
  assign n6184 = n6183 ^ n892 ^ 1'b0 ;
  assign n6185 = ~n3654 & n6184 ;
  assign n6186 = n6185 ^ n863 ^ 1'b0 ;
  assign n6191 = n6190 ^ n6187 ^ n6186 ;
  assign n6192 = n516 | n5241 ;
  assign n6193 = ~n877 & n6192 ;
  assign n6194 = n2603 & ~n3085 ;
  assign n6195 = n3901 | n6194 ;
  assign n6196 = n1281 & n2509 ;
  assign n6197 = ( n1378 & n6195 ) | ( n1378 & ~n6196 ) | ( n6195 & ~n6196 ) ;
  assign n6198 = n3557 ^ n1670 ^ n1106 ;
  assign n6199 = n494 & n6198 ;
  assign n6200 = n6199 ^ n4044 ^ 1'b0 ;
  assign n6201 = n6200 ^ n6079 ^ n2823 ;
  assign n6202 = n5041 ^ n1611 ^ 1'b0 ;
  assign n6203 = n6201 | n6202 ;
  assign n6204 = n4534 & ~n6203 ;
  assign n6205 = n1434 ^ n939 ^ 1'b0 ;
  assign n6207 = n2608 ^ n2187 ^ 1'b0 ;
  assign n6208 = ~n1222 & n6207 ;
  assign n6209 = ~n779 & n6208 ;
  assign n6210 = n6209 ^ n1887 ^ 1'b0 ;
  assign n6211 = n4475 | n6210 ;
  assign n6206 = n3470 ^ n1079 ^ 1'b0 ;
  assign n6212 = n6211 ^ n6206 ^ 1'b0 ;
  assign n6214 = ( n148 & n1302 ) | ( n148 & ~n1654 ) | ( n1302 & ~n1654 ) ;
  assign n6213 = ~x111 & n451 ;
  assign n6215 = n6214 ^ n6213 ^ 1'b0 ;
  assign n6216 = ~n6157 & n6215 ;
  assign n6217 = n1457 & n6216 ;
  assign n6218 = n4391 ^ n1338 ^ 1'b0 ;
  assign n6219 = n986 & ~n6218 ;
  assign n6220 = n6219 ^ n6187 ^ 1'b0 ;
  assign n6221 = n5225 ^ n2036 ^ 1'b0 ;
  assign n6223 = ( ~n910 & n1208 ) | ( ~n910 & n3249 ) | ( n1208 & n3249 ) ;
  assign n6224 = n439 | n6223 ;
  assign n6225 = n4189 | n6224 ;
  assign n6226 = n6225 ^ n461 ^ 1'b0 ;
  assign n6222 = n343 & ~n1231 ;
  assign n6227 = n6226 ^ n6222 ^ n3369 ;
  assign n6228 = x93 & ~n788 ;
  assign n6229 = n4740 | n6228 ;
  assign n6230 = n2128 & ~n6229 ;
  assign n6231 = n3760 ^ n484 ^ 1'b0 ;
  assign n6232 = n6013 ^ n2143 ^ n1312 ;
  assign n6233 = ( n1081 & n2476 ) | ( n1081 & ~n3814 ) | ( n2476 & ~n3814 ) ;
  assign n6234 = n4453 ^ n299 ^ 1'b0 ;
  assign n6235 = n6233 & ~n6234 ;
  assign n6236 = n3550 ^ n1979 ^ 1'b0 ;
  assign n6237 = x45 & ~n408 ;
  assign n6238 = n5106 & ~n6237 ;
  assign n6239 = n2632 ^ n510 ^ 1'b0 ;
  assign n6240 = n1486 ^ n1380 ^ 1'b0 ;
  assign n6241 = n425 | n6240 ;
  assign n6242 = n923 | n6241 ;
  assign n6243 = n6242 ^ n1734 ^ 1'b0 ;
  assign n6244 = n2886 | n3340 ;
  assign n6245 = n6244 ^ n1436 ^ 1'b0 ;
  assign n6247 = n1375 | n2496 ;
  assign n6246 = n149 | n1924 ;
  assign n6248 = n6247 ^ n6246 ^ 1'b0 ;
  assign n6249 = n6248 ^ n2393 ^ 1'b0 ;
  assign n6250 = n6245 & ~n6249 ;
  assign n6251 = n6250 ^ n2599 ^ 1'b0 ;
  assign n6252 = n630 ^ n527 ^ 1'b0 ;
  assign n6253 = n6252 ^ n2467 ^ n623 ;
  assign n6254 = n6253 ^ n3631 ^ 1'b0 ;
  assign n6255 = n482 & ~n6254 ;
  assign n6256 = x64 & ~n1511 ;
  assign n6257 = ~x20 & n6256 ;
  assign n6258 = n483 & ~n6257 ;
  assign n6259 = n688 & n6258 ;
  assign n6260 = n6259 ^ n1608 ^ 1'b0 ;
  assign n6261 = n4216 | n6260 ;
  assign n6262 = n2903 & ~n4667 ;
  assign n6263 = n223 ^ x58 ^ 1'b0 ;
  assign n6264 = ~n838 & n6263 ;
  assign n6265 = n975 | n6264 ;
  assign n6266 = ~n6262 & n6265 ;
  assign n6267 = n4757 & ~n5948 ;
  assign n6268 = n6267 ^ n650 ^ 1'b0 ;
  assign n6269 = n1220 & ~n3374 ;
  assign n6270 = n5979 ^ n277 ^ 1'b0 ;
  assign n6271 = n2815 & n6270 ;
  assign n6272 = n1553 | n2146 ;
  assign n6273 = n6272 ^ n6119 ^ 1'b0 ;
  assign n6274 = n5797 ^ n4868 ^ 1'b0 ;
  assign n6275 = n1520 & n6274 ;
  assign n6276 = n3111 & n6275 ;
  assign n6277 = n6276 ^ n2236 ^ 1'b0 ;
  assign n6278 = n2279 ^ n1036 ^ n239 ;
  assign n6279 = ( ~n3688 & n4745 ) | ( ~n3688 & n6278 ) | ( n4745 & n6278 ) ;
  assign n6280 = ( n2154 & n3820 ) | ( n2154 & ~n6279 ) | ( n3820 & ~n6279 ) ;
  assign n6281 = n1033 | n5902 ;
  assign n6282 = n6281 ^ n311 ^ 1'b0 ;
  assign n6283 = n3419 | n6282 ;
  assign n6284 = n5043 | n6283 ;
  assign n6285 = n5892 ^ n5415 ^ n5326 ;
  assign n6286 = n1585 & ~n5096 ;
  assign n6287 = n6286 ^ n5097 ^ n4620 ;
  assign n6288 = ( n337 & n379 ) | ( n337 & ~n3590 ) | ( n379 & ~n3590 ) ;
  assign n6289 = n5404 ^ n808 ^ 1'b0 ;
  assign n6290 = n5217 ^ n3842 ^ 1'b0 ;
  assign n6291 = n673 & n889 ;
  assign n6292 = n459 | n6291 ;
  assign n6293 = n6292 ^ n859 ^ 1'b0 ;
  assign n6294 = n925 & ~n6293 ;
  assign n6295 = ~n3910 & n6294 ;
  assign n6296 = ( ~n161 & n683 ) | ( ~n161 & n3334 ) | ( n683 & n3334 ) ;
  assign n6297 = n4637 ^ n3151 ^ 1'b0 ;
  assign n6298 = n5581 & n6297 ;
  assign n6299 = n6298 ^ n3139 ^ 1'b0 ;
  assign n6300 = n2330 ^ n2109 ^ 1'b0 ;
  assign n6301 = ( n309 & n2930 ) | ( n309 & ~n6300 ) | ( n2930 & ~n6300 ) ;
  assign n6302 = n1520 & n6301 ;
  assign n6303 = n5468 ^ n385 ^ 1'b0 ;
  assign n6304 = n4171 ^ n618 ^ 1'b0 ;
  assign n6305 = n6303 & n6304 ;
  assign n6306 = n6302 & n6305 ;
  assign n6307 = n2805 | n4085 ;
  assign n6308 = ( ~n395 & n650 ) | ( ~n395 & n2225 ) | ( n650 & n2225 ) ;
  assign n6309 = n6308 ^ n1762 ^ 1'b0 ;
  assign n6310 = n3418 & ~n6309 ;
  assign n6311 = n1031 | n1667 ;
  assign n6312 = n2221 & ~n6311 ;
  assign n6313 = n3761 & n6312 ;
  assign n6314 = ~n3349 & n6313 ;
  assign n6315 = ( ~n674 & n869 ) | ( ~n674 & n4677 ) | ( n869 & n4677 ) ;
  assign n6316 = n248 & n2873 ;
  assign n6317 = n2588 & n6316 ;
  assign n6318 = n1139 & ~n6317 ;
  assign n6319 = n6318 ^ n3791 ^ 1'b0 ;
  assign n6320 = ( n1570 & n2243 ) | ( n1570 & ~n4931 ) | ( n2243 & ~n4931 ) ;
  assign n6321 = n4353 ^ n1619 ^ 1'b0 ;
  assign n6322 = n2487 & ~n6321 ;
  assign n6323 = n2091 & ~n2569 ;
  assign n6324 = n362 & n4382 ;
  assign n6325 = ~n1673 & n6324 ;
  assign n6326 = n3940 & ~n6325 ;
  assign n6327 = n2461 & n6326 ;
  assign n6328 = n3067 ^ n1153 ^ x3 ;
  assign n6329 = n6328 ^ n3398 ^ 1'b0 ;
  assign n6330 = n920 & n3358 ;
  assign n6331 = ~n2780 & n6330 ;
  assign n6332 = n4485 & n6331 ;
  assign n6333 = n1489 & ~n6332 ;
  assign n6334 = ~n4178 & n6333 ;
  assign n6335 = n199 & n6334 ;
  assign n6336 = n2021 | n6335 ;
  assign n6337 = n4181 ^ x15 ^ 1'b0 ;
  assign n6338 = ( n2692 & n2706 ) | ( n2692 & ~n6337 ) | ( n2706 & ~n6337 ) ;
  assign n6339 = n3617 ^ n3424 ^ 1'b0 ;
  assign n6340 = n6339 ^ n1476 ^ 1'b0 ;
  assign n6341 = n6338 | n6340 ;
  assign n6342 = ~n202 & n1305 ;
  assign n6343 = n6342 ^ n1892 ^ 1'b0 ;
  assign n6344 = ~n1590 & n3358 ;
  assign n6345 = n2782 | n4839 ;
  assign n6346 = n6345 ^ n3653 ^ 1'b0 ;
  assign n6347 = n5001 ^ n4004 ^ 1'b0 ;
  assign n6348 = n742 | n6347 ;
  assign n6349 = n1309 & n3363 ;
  assign n6350 = n6349 ^ n5435 ^ n5002 ;
  assign n6351 = n6350 ^ n4441 ^ n1237 ;
  assign n6359 = n1246 & ~n1684 ;
  assign n6352 = n2107 & n3557 ;
  assign n6353 = n6352 ^ n3885 ^ 1'b0 ;
  assign n6354 = n3413 & ~n6353 ;
  assign n6355 = x94 & n6354 ;
  assign n6356 = n532 & n6355 ;
  assign n6357 = ~n5936 & n6356 ;
  assign n6358 = ( n1629 & n4915 ) | ( n1629 & n6357 ) | ( n4915 & n6357 ) ;
  assign n6360 = n6359 ^ n6358 ^ 1'b0 ;
  assign n6361 = n4183 ^ n733 ^ 1'b0 ;
  assign n6362 = n5076 & ~n6361 ;
  assign n6363 = n336 & n5432 ;
  assign n6364 = n5251 & n6363 ;
  assign n6365 = n132 | n1382 ;
  assign n6366 = n1406 & ~n6365 ;
  assign n6367 = n6366 ^ n331 ^ 1'b0 ;
  assign n6368 = n4750 & n6367 ;
  assign n6369 = n6368 ^ n6164 ^ 1'b0 ;
  assign n6370 = n6297 ^ n403 ^ 1'b0 ;
  assign n6371 = n1275 & ~n6370 ;
  assign n6373 = n3152 ^ n2028 ^ 1'b0 ;
  assign n6374 = n1031 | n6373 ;
  assign n6372 = n1955 ^ n979 ^ n764 ;
  assign n6375 = n6374 ^ n6372 ^ n1479 ;
  assign n6376 = n2106 | n6375 ;
  assign n6377 = n3059 ^ n1512 ^ 1'b0 ;
  assign n6378 = n5001 | n6377 ;
  assign n6379 = ( n1181 & n1306 ) | ( n1181 & ~n5725 ) | ( n1306 & ~n5725 ) ;
  assign n6380 = ( n2137 & ~n3357 ) | ( n2137 & n5772 ) | ( ~n3357 & n5772 ) ;
  assign n6381 = n217 | n6336 ;
  assign n6382 = n4406 ^ n3930 ^ 1'b0 ;
  assign n6383 = ( n1621 & n5858 ) | ( n1621 & n6382 ) | ( n5858 & n6382 ) ;
  assign n6384 = ~n3781 & n3874 ;
  assign n6385 = n3188 & n6384 ;
  assign n6386 = n429 | n4879 ;
  assign n6387 = n683 & ~n3712 ;
  assign n6388 = n6387 ^ n562 ^ 1'b0 ;
  assign n6389 = n6388 ^ n4972 ^ 1'b0 ;
  assign n6390 = n6386 & ~n6389 ;
  assign n6391 = ( n2558 & n3439 ) | ( n2558 & n5546 ) | ( n3439 & n5546 ) ;
  assign n6392 = n698 & n3285 ;
  assign n6393 = n6392 ^ n2558 ^ 1'b0 ;
  assign n6394 = n6393 ^ n4796 ^ n3340 ;
  assign n6396 = n2522 ^ n1070 ^ 1'b0 ;
  assign n6397 = n1776 & n6396 ;
  assign n6395 = n2826 & n5154 ;
  assign n6398 = n6397 ^ n6395 ^ x21 ;
  assign n6399 = ( n767 & n2978 ) | ( n767 & n3468 ) | ( n2978 & n3468 ) ;
  assign n6400 = n6399 ^ n6034 ^ 1'b0 ;
  assign n6401 = ( n730 & ~n1191 ) | ( n730 & n3163 ) | ( ~n1191 & n3163 ) ;
  assign n6402 = n4593 ^ n2666 ^ 1'b0 ;
  assign n6403 = ( x63 & n3583 ) | ( x63 & n6402 ) | ( n3583 & n6402 ) ;
  assign n6405 = n892 & ~n1067 ;
  assign n6406 = n6405 ^ n938 ^ 1'b0 ;
  assign n6404 = n415 & n725 ;
  assign n6407 = n6406 ^ n6404 ^ 1'b0 ;
  assign n6408 = n6403 & ~n6407 ;
  assign n6409 = n146 & ~n2299 ;
  assign n6410 = n6409 ^ n590 ^ 1'b0 ;
  assign n6411 = n146 & n5179 ;
  assign n6412 = ( n1875 & ~n4813 ) | ( n1875 & n6411 ) | ( ~n4813 & n6411 ) ;
  assign n6413 = n4358 & n5922 ;
  assign n6416 = n1519 | n2350 ;
  assign n6417 = n2350 & ~n6416 ;
  assign n6414 = x54 & n1714 ;
  assign n6415 = ~n1758 & n6414 ;
  assign n6418 = n6417 ^ n6415 ^ 1'b0 ;
  assign n6419 = n548 | n6418 ;
  assign n6420 = ~n785 & n1979 ;
  assign n6421 = n3055 ^ n908 ^ 1'b0 ;
  assign n6422 = n3297 & n6421 ;
  assign n6423 = n6422 ^ n3678 ^ 1'b0 ;
  assign n6424 = ~n6420 & n6423 ;
  assign n6425 = n753 | n6063 ;
  assign n6426 = n6425 ^ n483 ^ 1'b0 ;
  assign n6427 = n3728 | n3893 ;
  assign n6428 = n6427 ^ n3485 ^ 1'b0 ;
  assign n6429 = ~n6426 & n6428 ;
  assign n6430 = n6429 ^ n1581 ^ 1'b0 ;
  assign n6431 = n5745 ^ n2861 ^ n480 ;
  assign n6432 = n2429 ^ n1948 ^ 1'b0 ;
  assign n6433 = n3457 & ~n6432 ;
  assign n6434 = n6431 & n6433 ;
  assign n6435 = n3359 & ~n5785 ;
  assign n6436 = n4165 & ~n4874 ;
  assign n6437 = ~n4548 & n5755 ;
  assign n6438 = ~n994 & n6437 ;
  assign n6439 = n3440 ^ n176 ^ 1'b0 ;
  assign n6440 = n5389 ^ n3130 ^ n2293 ;
  assign n6441 = n1479 & n6440 ;
  assign n6442 = n5517 ^ n2793 ^ n638 ;
  assign n6443 = n6442 ^ n2682 ^ 1'b0 ;
  assign n6444 = ~n2627 & n6443 ;
  assign n6445 = n3556 ^ n2069 ^ 1'b0 ;
  assign n6446 = n6444 & n6445 ;
  assign n6452 = n1987 ^ n145 ^ 1'b0 ;
  assign n6449 = n2444 & ~n2583 ;
  assign n6450 = n859 & n6449 ;
  assign n6451 = ( n1949 & n4948 ) | ( n1949 & n6450 ) | ( n4948 & n6450 ) ;
  assign n6447 = n745 | n3710 ;
  assign n6448 = n6447 ^ n4394 ^ 1'b0 ;
  assign n6453 = n6452 ^ n6451 ^ n6448 ;
  assign n6457 = n3292 ^ n3015 ^ n2723 ;
  assign n6458 = n6457 ^ n1382 ^ 1'b0 ;
  assign n6454 = n3602 ^ n1936 ^ 1'b0 ;
  assign n6455 = x69 & n6454 ;
  assign n6456 = n6455 ^ n1498 ^ n955 ;
  assign n6459 = n6458 ^ n6456 ^ n4391 ;
  assign n6460 = ~n1382 & n2260 ;
  assign n6461 = n6460 ^ n706 ^ 1'b0 ;
  assign n6462 = n433 & n1966 ;
  assign n6463 = n521 & n6462 ;
  assign n6464 = x16 | n6463 ;
  assign n6465 = n2149 & n6464 ;
  assign n6466 = n6465 ^ n4757 ^ 1'b0 ;
  assign n6467 = n3708 ^ n1353 ^ 1'b0 ;
  assign n6468 = n4252 & n6467 ;
  assign n6469 = ~n3152 & n5144 ;
  assign n6470 = n6469 ^ n1714 ^ 1'b0 ;
  assign n6471 = ~x19 & n1161 ;
  assign n6472 = n2051 | n6471 ;
  assign n6473 = ( n189 & ~n1347 ) | ( n189 & n6215 ) | ( ~n1347 & n6215 ) ;
  assign n6474 = n1002 ^ x51 ^ 1'b0 ;
  assign n6475 = n4975 & n6474 ;
  assign n6476 = n6475 ^ n4819 ^ 1'b0 ;
  assign n6477 = n3712 ^ n510 ^ 1'b0 ;
  assign n6478 = ~n3617 & n6477 ;
  assign n6479 = n6478 ^ n3465 ^ 1'b0 ;
  assign n6480 = n1489 | n4570 ;
  assign n6481 = n6480 ^ n2896 ^ 1'b0 ;
  assign n6482 = n2331 ^ n2119 ^ 1'b0 ;
  assign n6483 = ( ~n2632 & n4594 ) | ( ~n2632 & n6482 ) | ( n4594 & n6482 ) ;
  assign n6484 = n4149 ^ n2250 ^ 1'b0 ;
  assign n6485 = n1155 | n6484 ;
  assign n6486 = n3567 | n6337 ;
  assign n6487 = n6485 & ~n6486 ;
  assign n6488 = ( x55 & ~n701 ) | ( x55 & n6487 ) | ( ~n701 & n6487 ) ;
  assign n6489 = n6488 ^ n2310 ^ 1'b0 ;
  assign n6490 = n1080 ^ x15 ^ 1'b0 ;
  assign n6491 = n5527 ^ n2221 ^ n1885 ;
  assign n6492 = n2162 & ~n6491 ;
  assign n6493 = n6490 & n6492 ;
  assign n6494 = n4159 ^ n3281 ^ n2147 ;
  assign n6495 = n2406 & ~n4675 ;
  assign n6496 = n6495 ^ n2316 ^ 1'b0 ;
  assign n6497 = n6496 ^ n6195 ^ n1700 ;
  assign n6498 = n6497 ^ x110 ^ x89 ;
  assign n6499 = ~n1525 & n5116 ;
  assign n6500 = n4306 ^ n956 ^ 1'b0 ;
  assign n6501 = n5526 & ~n6500 ;
  assign n6502 = ~n174 & n977 ;
  assign n6503 = n6502 ^ n3103 ^ n972 ;
  assign n6504 = n6382 & ~n6503 ;
  assign n6505 = n3211 ^ n2549 ^ 1'b0 ;
  assign n6506 = n1940 & n6505 ;
  assign n6507 = n3583 | n4106 ;
  assign n6508 = n5078 & ~n6507 ;
  assign n6509 = n6506 & ~n6508 ;
  assign n6511 = n1953 ^ n670 ^ x78 ;
  assign n6510 = n1268 & n1449 ;
  assign n6512 = n6511 ^ n6510 ^ 1'b0 ;
  assign n6513 = n530 & n1776 ;
  assign n6514 = n6512 & n6513 ;
  assign n6515 = n6514 ^ n6479 ^ 1'b0 ;
  assign n6516 = n3310 ^ n1141 ^ 1'b0 ;
  assign n6517 = ~n4927 & n5291 ;
  assign n6518 = n2915 | n5255 ;
  assign n6519 = n6518 ^ n1605 ^ n150 ;
  assign n6520 = ~x37 & x45 ;
  assign n6521 = n2142 & ~n6520 ;
  assign n6522 = ( n644 & n1690 ) | ( n644 & n6521 ) | ( n1690 & n6521 ) ;
  assign n6525 = n612 & ~n2176 ;
  assign n6526 = ~n307 & n6525 ;
  assign n6523 = n676 & ~n1411 ;
  assign n6524 = ~n3270 & n6523 ;
  assign n6527 = n6526 ^ n6524 ^ 1'b0 ;
  assign n6528 = n640 & n6527 ;
  assign n6529 = n5553 | n6528 ;
  assign n6530 = n6529 ^ n5702 ^ n1197 ;
  assign n6531 = n6522 & n6530 ;
  assign n6532 = n6519 & n6531 ;
  assign n6533 = n2231 ^ n899 ^ 1'b0 ;
  assign n6534 = ( n565 & n5750 ) | ( n565 & ~n6533 ) | ( n5750 & ~n6533 ) ;
  assign n6535 = n854 | n6534 ;
  assign n6536 = n6535 ^ n5053 ^ 1'b0 ;
  assign n6537 = n5705 ^ n5281 ^ 1'b0 ;
  assign n6538 = n1251 & n5514 ;
  assign n6539 = n6538 ^ n303 ^ 1'b0 ;
  assign n6540 = n2592 & n6539 ;
  assign n6541 = ~n706 & n6540 ;
  assign n6542 = n6541 ^ n1811 ^ 1'b0 ;
  assign n6543 = ~n2529 & n6542 ;
  assign n6544 = n6543 ^ n681 ^ 1'b0 ;
  assign n6545 = ~n2159 & n6544 ;
  assign n6546 = n3561 & n6122 ;
  assign n6547 = ~n438 & n1570 ;
  assign n6548 = n6546 | n6547 ;
  assign n6549 = x102 & n4362 ;
  assign n6550 = ~n1138 & n3755 ;
  assign n6551 = n681 & n5842 ;
  assign n6552 = n6551 ^ n4613 ^ 1'b0 ;
  assign n6553 = n3110 & ~n3320 ;
  assign n6554 = ~n1023 & n4705 ;
  assign n6555 = n6554 ^ n1486 ^ 1'b0 ;
  assign n6556 = n1033 | n2622 ;
  assign n6557 = n4705 | n6556 ;
  assign n6558 = n6533 ^ n5453 ^ n1792 ;
  assign n6559 = n6558 ^ n1197 ^ 1'b0 ;
  assign n6560 = n6557 & ~n6559 ;
  assign n6564 = ~n734 & n1566 ;
  assign n6565 = x87 & ~n6564 ;
  assign n6566 = n4587 & n6565 ;
  assign n6561 = n2551 & n3637 ;
  assign n6562 = n6561 ^ n2675 ^ 1'b0 ;
  assign n6563 = n4847 | n6562 ;
  assign n6567 = n6566 ^ n6563 ^ n703 ;
  assign n6568 = n497 & n2282 ;
  assign n6569 = ~n5839 & n6568 ;
  assign n6570 = ( n1742 & ~n4931 ) | ( n1742 & n6569 ) | ( ~n4931 & n6569 ) ;
  assign n6571 = n692 & ~n5677 ;
  assign n6572 = n6571 ^ n581 ^ 1'b0 ;
  assign n6573 = n4526 | n6572 ;
  assign n6574 = ~n319 & n2928 ;
  assign n6575 = n6574 ^ n4221 ^ 1'b0 ;
  assign n6576 = ~n2007 & n3422 ;
  assign n6577 = n2737 & ~n3467 ;
  assign n6578 = n6576 & n6577 ;
  assign n6579 = n2756 & ~n6578 ;
  assign n6580 = n2487 ^ n380 ^ 1'b0 ;
  assign n6588 = n2987 ^ n1954 ^ n871 ;
  assign n6589 = x44 & ~n6588 ;
  assign n6590 = n375 & n6589 ;
  assign n6584 = n4550 ^ n2645 ^ n947 ;
  assign n6585 = n2821 | n5144 ;
  assign n6586 = n6584 | n6585 ;
  assign n6581 = n5778 ^ n713 ^ 1'b0 ;
  assign n6582 = ~n1242 & n6581 ;
  assign n6583 = ~n4123 & n6582 ;
  assign n6587 = n6586 ^ n6583 ^ 1'b0 ;
  assign n6591 = n6590 ^ n6587 ^ n4858 ;
  assign n6592 = ~n1743 & n3113 ;
  assign n6593 = ~n3970 & n6592 ;
  assign n6595 = x9 & n691 ;
  assign n6596 = n701 & n6595 ;
  assign n6594 = n1125 & n1154 ;
  assign n6597 = n6596 ^ n6594 ^ 1'b0 ;
  assign n6598 = ~n372 & n6597 ;
  assign n6599 = n6598 ^ n4749 ^ 1'b0 ;
  assign n6600 = n6599 ^ n602 ^ 1'b0 ;
  assign n6601 = x110 | n3529 ;
  assign n6602 = n3369 & ~n6601 ;
  assign n6603 = ( n769 & ~n2842 ) | ( n769 & n6217 ) | ( ~n2842 & n6217 ) ;
  assign n6604 = ( n3904 & n6602 ) | ( n3904 & n6603 ) | ( n6602 & n6603 ) ;
  assign n6605 = n3853 & n6604 ;
  assign n6606 = n764 & ~n1654 ;
  assign n6607 = n6606 ^ n1183 ^ 1'b0 ;
  assign n6608 = ~n1072 & n4354 ;
  assign n6609 = n6607 & n6608 ;
  assign n6610 = ~n3532 & n6609 ;
  assign n6611 = n1067 & ~n6610 ;
  assign n6612 = ~n319 & n2897 ;
  assign n6613 = n2069 & ~n6612 ;
  assign n6614 = ~n1832 & n6613 ;
  assign n6615 = n6614 ^ n859 ^ 1'b0 ;
  assign n6616 = ~n1600 & n6615 ;
  assign n6617 = ( n5316 & n5804 ) | ( n5316 & ~n6616 ) | ( n5804 & ~n6616 ) ;
  assign n6618 = n1169 ^ n483 ^ 1'b0 ;
  assign n6619 = n2926 & ~n6618 ;
  assign n6620 = n248 & n6619 ;
  assign n6621 = n6620 ^ n4445 ^ 1'b0 ;
  assign n6622 = x123 | n1917 ;
  assign n6623 = n3188 | n4874 ;
  assign n6624 = n6623 ^ n5840 ^ n5473 ;
  assign n6631 = ( x41 & ~n404 ) | ( x41 & n1218 ) | ( ~n404 & n1218 ) ;
  assign n6625 = n1607 ^ x60 ^ 1'b0 ;
  assign n6626 = n3362 ^ n202 ^ 1'b0 ;
  assign n6627 = n3138 & n6626 ;
  assign n6628 = n6627 ^ n577 ^ 1'b0 ;
  assign n6629 = n6625 & n6628 ;
  assign n6630 = ~n425 & n6629 ;
  assign n6632 = n6631 ^ n6630 ^ 1'b0 ;
  assign n6633 = n6632 ^ n4704 ^ n454 ;
  assign n6634 = n1072 | n6633 ;
  assign n6635 = n2299 & ~n6590 ;
  assign n6636 = n6635 ^ n2355 ^ 1'b0 ;
  assign n6637 = n1972 & ~n2932 ;
  assign n6638 = n6119 ^ n783 ^ n236 ;
  assign n6639 = ( n6374 & ~n6637 ) | ( n6374 & n6638 ) | ( ~n6637 & n6638 ) ;
  assign n6640 = n5255 ^ n2014 ^ 1'b0 ;
  assign n6641 = n2817 | n6640 ;
  assign n6642 = n1837 | n5594 ;
  assign n6643 = n1599 ^ n819 ^ 1'b0 ;
  assign n6644 = n1583 | n1784 ;
  assign n6645 = n4481 | n6644 ;
  assign n6646 = n6645 ^ n4959 ^ 1'b0 ;
  assign n6647 = n1356 | n1611 ;
  assign n6648 = n5790 & ~n6635 ;
  assign n6649 = n5826 & n6648 ;
  assign n6650 = n4498 & ~n6649 ;
  assign n6651 = n6451 & n6650 ;
  assign n6653 = n850 ^ n764 ^ 1'b0 ;
  assign n6652 = ~n3050 & n4380 ;
  assign n6654 = n6653 ^ n6652 ^ 1'b0 ;
  assign n6655 = ~n4337 & n6654 ;
  assign n6656 = ( n1283 & ~n3057 ) | ( n1283 & n4983 ) | ( ~n3057 & n4983 ) ;
  assign n6657 = n1448 ^ n438 ^ 1'b0 ;
  assign n6658 = n6657 ^ n1150 ^ n764 ;
  assign n6659 = n4283 ^ n2958 ^ 1'b0 ;
  assign n6660 = n6391 & n6659 ;
  assign n6661 = n6635 ^ n3471 ^ n2184 ;
  assign n6662 = n6661 ^ n828 ^ 1'b0 ;
  assign n6663 = n4442 ^ n854 ^ 1'b0 ;
  assign n6664 = n325 & ~n3998 ;
  assign n6665 = n6664 ^ n2151 ^ 1'b0 ;
  assign n6666 = n6337 ^ n731 ^ 1'b0 ;
  assign n6667 = ( n891 & n2103 ) | ( n891 & n6666 ) | ( n2103 & n6666 ) ;
  assign n6668 = ~n6665 & n6667 ;
  assign n6669 = n6668 ^ n6532 ^ 1'b0 ;
  assign n6670 = n5399 ^ n422 ^ 1'b0 ;
  assign n6671 = n6670 ^ n4391 ^ 1'b0 ;
  assign n6672 = n3930 ^ n1899 ^ 1'b0 ;
  assign n6673 = ~n3709 & n6672 ;
  assign n6674 = ~n1791 & n6673 ;
  assign n6675 = n3211 | n5916 ;
  assign n6676 = n6675 ^ n3546 ^ 1'b0 ;
  assign n6677 = n5396 & n6676 ;
  assign n6678 = ~n3265 & n6677 ;
  assign n6679 = n130 & ~n3172 ;
  assign n6680 = n6679 ^ n4879 ^ 1'b0 ;
  assign n6681 = ( n973 & ~n1273 ) | ( n973 & n4968 ) | ( ~n1273 & n4968 ) ;
  assign n6682 = n1746 ^ n764 ^ 1'b0 ;
  assign n6683 = n4451 ^ n687 ^ 1'b0 ;
  assign n6686 = n6602 ^ n4596 ^ 1'b0 ;
  assign n6687 = n6686 ^ n771 ^ 1'b0 ;
  assign n6684 = ( n1594 & ~n2217 ) | ( n1594 & n3070 ) | ( ~n2217 & n3070 ) ;
  assign n6685 = ~n2999 & n6684 ;
  assign n6688 = n6687 ^ n6685 ^ 1'b0 ;
  assign n6689 = n1521 & ~n3292 ;
  assign n6690 = ( n335 & n485 ) | ( n335 & ~n6689 ) | ( n485 & ~n6689 ) ;
  assign n6691 = ( n4543 & ~n6291 ) | ( n4543 & n6690 ) | ( ~n6291 & n6690 ) ;
  assign n6692 = n4131 ^ n2019 ^ n588 ;
  assign n6693 = n2947 & ~n4339 ;
  assign n6694 = n6692 & n6693 ;
  assign n6695 = n2780 ^ n2582 ^ 1'b0 ;
  assign n6696 = ~n1403 & n6695 ;
  assign n6699 = n1693 | n6223 ;
  assign n6700 = n2735 & ~n6699 ;
  assign n6701 = n2005 & n6700 ;
  assign n6697 = ~n2605 & n4400 ;
  assign n6698 = n6697 ^ n2750 ^ 1'b0 ;
  assign n6702 = n6701 ^ n6698 ^ n456 ;
  assign n6703 = n5879 & ~n6170 ;
  assign n6704 = n5797 ^ n2236 ^ 1'b0 ;
  assign n6705 = n6704 ^ n6415 ^ n960 ;
  assign n6706 = n6703 & ~n6705 ;
  assign n6707 = x34 & ~n5133 ;
  assign n6708 = ~n245 & n946 ;
  assign n6709 = n934 & ~n1743 ;
  assign n6710 = ~n2507 & n6709 ;
  assign n6711 = n6710 ^ n1181 ^ 1'b0 ;
  assign n6712 = n6711 ^ n5059 ^ n3304 ;
  assign n6713 = ~n3571 & n6712 ;
  assign n6714 = n3714 & n6713 ;
  assign n6715 = n2566 & ~n5855 ;
  assign n6716 = n6715 ^ n1906 ^ 1'b0 ;
  assign n6717 = ~n498 & n2634 ;
  assign n6718 = n1324 & ~n2118 ;
  assign n6719 = n2634 & n6718 ;
  assign n6720 = n6719 ^ n1766 ^ 1'b0 ;
  assign n6721 = n6717 | n6720 ;
  assign n6722 = ( n576 & n2170 ) | ( n576 & ~n3323 ) | ( n2170 & ~n3323 ) ;
  assign n6723 = n6722 ^ n2892 ^ 1'b0 ;
  assign n6724 = n2046 & ~n6723 ;
  assign n6725 = n3440 & n6724 ;
  assign n6726 = n6725 ^ n5067 ^ 1'b0 ;
  assign n6727 = ~n725 & n5281 ;
  assign n6728 = n6727 ^ n462 ^ 1'b0 ;
  assign n6729 = n6728 ^ n3367 ^ 1'b0 ;
  assign n6733 = n1961 & n2476 ;
  assign n6734 = n2968 & n6733 ;
  assign n6735 = n4752 | n6734 ;
  assign n6730 = n1976 ^ n663 ^ 1'b0 ;
  assign n6731 = n1827 | n6730 ;
  assign n6732 = n5606 & ~n6731 ;
  assign n6736 = n6735 ^ n6732 ^ 1'b0 ;
  assign n6737 = n2825 ^ n1998 ^ 1'b0 ;
  assign n6738 = n2133 | n6737 ;
  assign n6739 = n3542 & ~n6738 ;
  assign n6740 = n1041 | n3014 ;
  assign n6741 = n6740 ^ n3752 ^ 1'b0 ;
  assign n6742 = n6741 ^ n2206 ^ 1'b0 ;
  assign n6743 = ~n496 & n5328 ;
  assign n6744 = n5212 | n6134 ;
  assign n6745 = n3755 | n6744 ;
  assign n6746 = n3351 ^ n373 ^ 1'b0 ;
  assign n6749 = n615 & n4584 ;
  assign n6748 = ( n1094 & n4902 ) | ( n1094 & ~n5391 ) | ( n4902 & ~n5391 ) ;
  assign n6747 = ~n1138 & n1909 ;
  assign n6750 = n6749 ^ n6748 ^ n6747 ;
  assign n6751 = n4346 ^ n2569 ^ n2547 ;
  assign n6752 = n3820 ^ n1655 ^ 1'b0 ;
  assign n6753 = n5327 | n6752 ;
  assign n6754 = n2105 & ~n6753 ;
  assign n6755 = n6754 ^ n3641 ^ 1'b0 ;
  assign n6756 = n2428 | n4593 ;
  assign n6757 = n6756 ^ n4859 ^ 1'b0 ;
  assign n6758 = n3893 | n6757 ;
  assign n6759 = ( n2331 & n2513 ) | ( n2331 & n3436 ) | ( n2513 & n3436 ) ;
  assign n6760 = ~n673 & n1749 ;
  assign n6761 = n6760 ^ n5712 ^ 1'b0 ;
  assign n6762 = n1668 ^ n681 ^ 1'b0 ;
  assign n6763 = n483 & ~n6762 ;
  assign n6764 = ~n3057 & n6763 ;
  assign n6765 = ~n3079 & n6764 ;
  assign n6766 = n6765 ^ n1279 ^ 1'b0 ;
  assign n6767 = n4306 & ~n6766 ;
  assign n6768 = n6706 ^ n1570 ^ 1'b0 ;
  assign n6769 = n3552 ^ n1023 ^ n383 ;
  assign n6770 = ( ~n1134 & n3244 ) | ( ~n1134 & n6769 ) | ( n3244 & n6769 ) ;
  assign n6771 = n6770 ^ n3871 ^ n1150 ;
  assign n6772 = n6687 ^ n6508 ^ 1'b0 ;
  assign n6773 = ~n6771 & n6772 ;
  assign n6776 = ( ~n2682 & n2706 ) | ( ~n2682 & n2831 ) | ( n2706 & n2831 ) ;
  assign n6775 = ~n2262 & n2710 ;
  assign n6777 = n6776 ^ n6775 ^ 1'b0 ;
  assign n6774 = n175 & ~n4494 ;
  assign n6778 = n6777 ^ n6774 ^ 1'b0 ;
  assign n6779 = n4441 ^ n1843 ^ 1'b0 ;
  assign n6780 = n6569 ^ n3323 ^ 1'b0 ;
  assign n6781 = n6779 & n6780 ;
  assign n6782 = n4048 ^ n3653 ^ 1'b0 ;
  assign n6783 = n6782 ^ x20 ^ 1'b0 ;
  assign n6784 = n2795 | n6783 ;
  assign n6785 = n1099 & ~n3476 ;
  assign n6786 = ( n930 & n3429 ) | ( n930 & ~n5043 ) | ( n3429 & ~n5043 ) ;
  assign n6787 = x71 & ~n6786 ;
  assign n6788 = ~n3063 & n3537 ;
  assign n6789 = ~n6787 & n6788 ;
  assign n6790 = ~n840 & n2958 ;
  assign n6791 = ~n2024 & n2339 ;
  assign n6792 = n202 & ~n2045 ;
  assign n6793 = n1106 ^ n231 ^ 1'b0 ;
  assign n6794 = ~n6792 & n6793 ;
  assign n6795 = ( n2415 & ~n6791 ) | ( n2415 & n6794 ) | ( ~n6791 & n6794 ) ;
  assign n6796 = ( n575 & ~n3363 ) | ( n575 & n4048 ) | ( ~n3363 & n4048 ) ;
  assign n6799 = ~n2882 & n3862 ;
  assign n6797 = ( n363 & n1597 ) | ( n363 & ~n6363 ) | ( n1597 & ~n6363 ) ;
  assign n6798 = n6797 ^ n3284 ^ 1'b0 ;
  assign n6800 = n6799 ^ n6798 ^ 1'b0 ;
  assign n6801 = n6796 & n6800 ;
  assign n6802 = ( n2333 & ~n3519 ) | ( n2333 & n4581 ) | ( ~n3519 & n4581 ) ;
  assign n6804 = n479 & ~n2125 ;
  assign n6803 = n642 | n4868 ;
  assign n6805 = n6804 ^ n6803 ^ 1'b0 ;
  assign n6806 = n2951 ^ n2877 ^ 1'b0 ;
  assign n6807 = n4225 ^ n1559 ^ n763 ;
  assign n6808 = n5618 & n6807 ;
  assign n6809 = n6806 & n6808 ;
  assign n6810 = n1106 & ~n3524 ;
  assign n6811 = ~n4323 & n6810 ;
  assign n6812 = n884 & n6411 ;
  assign n6813 = n6198 ^ n670 ^ 1'b0 ;
  assign n6814 = n6813 ^ n1535 ^ 1'b0 ;
  assign n6815 = n5416 | n6814 ;
  assign n6816 = ( n2325 & n3525 ) | ( n2325 & ~n6815 ) | ( n3525 & ~n6815 ) ;
  assign n6817 = n6816 ^ n4311 ^ 1'b0 ;
  assign n6818 = ( n1372 & n2140 ) | ( n1372 & ~n5247 ) | ( n2140 & ~n5247 ) ;
  assign n6819 = n2178 ^ n381 ^ 1'b0 ;
  assign n6820 = n3509 ^ n2260 ^ n1617 ;
  assign n6821 = ~n1385 & n1798 ;
  assign n6822 = n6821 ^ n5900 ^ 1'b0 ;
  assign n6823 = ~n5267 & n6822 ;
  assign n6824 = ( n1498 & n6122 ) | ( n1498 & n6823 ) | ( n6122 & n6823 ) ;
  assign n6825 = ~n6820 & n6824 ;
  assign n6826 = n2970 ^ n1823 ^ n770 ;
  assign n6827 = n6826 ^ n664 ^ 1'b0 ;
  assign n6828 = ~n6046 & n6827 ;
  assign n6832 = n2357 & n4777 ;
  assign n6833 = n6832 ^ n442 ^ 1'b0 ;
  assign n6831 = ~n790 & n1766 ;
  assign n6834 = n6833 ^ n6831 ^ 1'b0 ;
  assign n6829 = ( n730 & n1193 ) | ( n730 & n1805 ) | ( n1193 & n1805 ) ;
  assign n6830 = n6829 ^ n1818 ^ 1'b0 ;
  assign n6835 = n6834 ^ n6830 ^ n3319 ;
  assign n6836 = n2307 & n5528 ;
  assign n6837 = n6836 ^ n3395 ^ 1'b0 ;
  assign n6838 = n6837 ^ n507 ^ 1'b0 ;
  assign n6839 = n1356 | n6838 ;
  assign n6840 = n247 & ~n6839 ;
  assign n6841 = n2744 & n6840 ;
  assign n6842 = n2703 & ~n5013 ;
  assign n6843 = n719 & ~n1171 ;
  assign n6844 = n6843 ^ n627 ^ 1'b0 ;
  assign n6845 = n6844 ^ n3990 ^ 1'b0 ;
  assign n6846 = n2495 ^ n2383 ^ n919 ;
  assign n6847 = n4884 ^ n3217 ^ n2612 ;
  assign n6848 = ~n6846 & n6847 ;
  assign n6849 = n1097 & ~n2276 ;
  assign n6850 = ~n2668 & n6849 ;
  assign n6851 = n407 | n1482 ;
  assign n6852 = n755 & ~n6851 ;
  assign n6853 = n415 & n726 ;
  assign n6854 = n3651 & n6853 ;
  assign n6855 = n5219 & n6854 ;
  assign n6856 = x93 & ~n6855 ;
  assign n6857 = n1041 & ~n3308 ;
  assign n6858 = ~n659 & n6857 ;
  assign n6859 = ( x117 & n2729 ) | ( x117 & ~n3738 ) | ( n2729 & ~n3738 ) ;
  assign n6860 = ( n404 & ~n486 ) | ( n404 & n539 ) | ( ~n486 & n539 ) ;
  assign n6861 = x108 & ~n2802 ;
  assign n6862 = ~n6860 & n6861 ;
  assign n6863 = n6133 ^ n1100 ^ 1'b0 ;
  assign n6864 = n6521 & n6863 ;
  assign n6865 = n663 & n4942 ;
  assign n6866 = ~n6864 & n6865 ;
  assign n6867 = n1742 & ~n3561 ;
  assign n6868 = ( x76 & ~n2546 ) | ( x76 & n6867 ) | ( ~n2546 & n6867 ) ;
  assign n6869 = n3358 & ~n6868 ;
  assign n6870 = ~n6128 & n6869 ;
  assign n6873 = x89 & n1998 ;
  assign n6874 = n3036 & n6873 ;
  assign n6871 = ~n1374 & n3612 ;
  assign n6872 = n6871 ^ n1479 ^ 1'b0 ;
  assign n6875 = n6874 ^ n6872 ^ n3875 ;
  assign n6876 = n4504 ^ n3334 ^ 1'b0 ;
  assign n6877 = n6876 ^ n5839 ^ 1'b0 ;
  assign n6878 = n4420 ^ n471 ^ 1'b0 ;
  assign n6879 = n6878 ^ n450 ^ 1'b0 ;
  assign n6880 = n6877 | n6879 ;
  assign n6881 = n2329 & ~n3172 ;
  assign n6882 = n6881 ^ n1743 ^ 1'b0 ;
  assign n6883 = ~n1705 & n2549 ;
  assign n6884 = n6883 ^ n1135 ^ 1'b0 ;
  assign n6885 = n6884 ^ n3617 ^ 1'b0 ;
  assign n6886 = n744 & ~n4718 ;
  assign n6890 = n1650 & n2800 ;
  assign n6891 = ~n2621 & n6890 ;
  assign n6887 = n521 | n2513 ;
  assign n6888 = n6887 ^ n4875 ^ 1'b0 ;
  assign n6889 = n4812 & n6888 ;
  assign n6892 = n6891 ^ n6889 ^ 1'b0 ;
  assign n6893 = ( n635 & n3095 ) | ( n635 & n6892 ) | ( n3095 & n6892 ) ;
  assign n6894 = n4257 ^ n882 ^ 1'b0 ;
  assign n6895 = ~n1619 & n6894 ;
  assign n6896 = n6895 ^ n2509 ^ 1'b0 ;
  assign n6897 = n3631 | n5240 ;
  assign n6900 = n2226 | n3516 ;
  assign n6898 = n336 & ~n2409 ;
  assign n6899 = n6898 ^ n1885 ^ n452 ;
  assign n6901 = n6900 ^ n6899 ^ n6502 ;
  assign n6908 = n1549 ^ n1192 ^ 1'b0 ;
  assign n6909 = n436 & n725 ;
  assign n6910 = n1181 | n6909 ;
  assign n6911 = n6908 | n6910 ;
  assign n6906 = n3015 ^ n2558 ^ n1959 ;
  assign n6902 = ~n1226 & n2411 ;
  assign n6903 = n6902 ^ n5677 ^ 1'b0 ;
  assign n6904 = n2908 & ~n6903 ;
  assign n6905 = n2007 & n6904 ;
  assign n6907 = n6906 ^ n6905 ^ 1'b0 ;
  assign n6912 = n6911 ^ n6907 ^ n6524 ;
  assign n6913 = n6296 ^ x118 ^ 1'b0 ;
  assign n6914 = n5909 & ~n6913 ;
  assign n6915 = n661 ^ n370 ^ 1'b0 ;
  assign n6916 = ( n487 & n6834 ) | ( n487 & ~n6915 ) | ( n6834 & ~n6915 ) ;
  assign n6917 = n2466 | n3310 ;
  assign n6918 = n6917 ^ n3892 ^ 1'b0 ;
  assign n6919 = n6918 ^ n6297 ^ 1'b0 ;
  assign n6922 = n2767 ^ n742 ^ 1'b0 ;
  assign n6923 = ( n1971 & ~n2789 ) | ( n1971 & n6922 ) | ( ~n2789 & n6922 ) ;
  assign n6920 = n4625 ^ n984 ^ 1'b0 ;
  assign n6921 = n6614 | n6920 ;
  assign n6924 = n6923 ^ n6921 ^ 1'b0 ;
  assign n6925 = n288 | n6924 ;
  assign n6926 = ~n2419 & n4876 ;
  assign n6927 = n5090 | n6114 ;
  assign n6928 = n6927 ^ n5733 ^ 1'b0 ;
  assign n6929 = n5953 ^ n4557 ^ 1'b0 ;
  assign n6930 = n6407 | n6929 ;
  assign n6931 = n478 | n4291 ;
  assign n6936 = x53 | n1308 ;
  assign n6937 = n2693 | n6936 ;
  assign n6938 = n690 & n6937 ;
  assign n6939 = ~n2246 & n6938 ;
  assign n6932 = n1200 | n2323 ;
  assign n6933 = n6932 ^ n4399 ^ 1'b0 ;
  assign n6934 = ~n6844 & n6933 ;
  assign n6935 = n2393 & ~n6934 ;
  assign n6940 = n6939 ^ n6935 ^ 1'b0 ;
  assign n6941 = ~n3946 & n4491 ;
  assign n6942 = n6941 ^ n1212 ^ 1'b0 ;
  assign n6943 = n6940 & ~n6942 ;
  assign n6944 = n4367 ^ n755 ^ 1'b0 ;
  assign n6945 = n4367 & ~n6944 ;
  assign n6946 = n6945 ^ n4716 ^ 1'b0 ;
  assign n6947 = n763 | n6946 ;
  assign n6948 = n6947 ^ n1086 ^ 1'b0 ;
  assign n6949 = n1571 & n5994 ;
  assign n6950 = n6949 ^ n3027 ^ 1'b0 ;
  assign n6951 = n4088 | n6950 ;
  assign n6952 = n3047 & ~n5293 ;
  assign n6953 = ~n3619 & n6952 ;
  assign n6954 = n6953 ^ n6923 ^ 1'b0 ;
  assign n6955 = ~n173 & n5410 ;
  assign n6957 = n5927 ^ n3876 ^ 1'b0 ;
  assign n6958 = x55 & n6957 ;
  assign n6956 = ~n1487 & n2649 ;
  assign n6959 = n6958 ^ n6956 ^ 1'b0 ;
  assign n6960 = n5517 ^ n2660 ^ 1'b0 ;
  assign n6961 = n5968 & ~n6960 ;
  assign n6962 = ~n5583 & n6961 ;
  assign n6963 = n6959 & n6962 ;
  assign n6964 = n6789 & ~n6963 ;
  assign n6965 = x116 & ~n4185 ;
  assign n6966 = n6965 ^ n673 ^ 1'b0 ;
  assign n6967 = n3572 | n6966 ;
  assign n6968 = n4420 | n6967 ;
  assign n6969 = ( n1799 & ~n5400 ) | ( n1799 & n6968 ) | ( ~n5400 & n6968 ) ;
  assign n6974 = n1113 | n4109 ;
  assign n6970 = n1239 & n1995 ;
  assign n6971 = n6318 & n6970 ;
  assign n6972 = n5375 | n6971 ;
  assign n6973 = n6381 | n6972 ;
  assign n6975 = n6974 ^ n6973 ^ 1'b0 ;
  assign n6976 = n1240 | n1501 ;
  assign n6977 = n6976 ^ x0 ^ 1'b0 ;
  assign n6978 = n6977 ^ n3172 ^ 1'b0 ;
  assign n6979 = ( n1467 & n1736 ) | ( n1467 & ~n2295 ) | ( n1736 & ~n2295 ) ;
  assign n6980 = n6979 ^ n6534 ^ n6128 ;
  assign n6981 = n1501 & ~n2969 ;
  assign n6982 = n6031 & ~n6981 ;
  assign n6983 = ( n341 & ~n6980 ) | ( n341 & n6982 ) | ( ~n6980 & n6982 ) ;
  assign n6984 = ~n2864 & n4270 ;
  assign n6985 = n1036 & n6984 ;
  assign n6986 = n6985 ^ n4813 ^ 1'b0 ;
  assign n6987 = n3674 | n6986 ;
  assign n6988 = n1780 | n3492 ;
  assign n6989 = n6609 ^ n858 ^ 1'b0 ;
  assign n6990 = n6408 | n6989 ;
  assign n6992 = n4064 ^ n466 ^ 1'b0 ;
  assign n6993 = n4076 & n6992 ;
  assign n6994 = ~n165 & n6637 ;
  assign n6995 = n6993 & n6994 ;
  assign n6996 = ( n4186 & n4752 ) | ( n4186 & ~n6995 ) | ( n4752 & ~n6995 ) ;
  assign n6991 = ~n821 & n1856 ;
  assign n6997 = n6996 ^ n6991 ^ 1'b0 ;
  assign n6998 = n1903 & ~n6997 ;
  assign n6999 = n6998 ^ n6255 ^ 1'b0 ;
  assign n7000 = x94 & n5283 ;
  assign n7001 = n7000 ^ n3729 ^ n1433 ;
  assign n7002 = n729 & ~n7001 ;
  assign n7003 = n7002 ^ n1697 ^ 1'b0 ;
  assign n7004 = n1496 & ~n2501 ;
  assign n7005 = n7004 ^ n6627 ^ n536 ;
  assign n7006 = n1472 & n7005 ;
  assign n7007 = n6614 & n7006 ;
  assign n7008 = n5485 & ~n7007 ;
  assign n7009 = x38 & n3022 ;
  assign n7010 = n7009 ^ n696 ^ 1'b0 ;
  assign n7012 = n3861 ^ n1374 ^ 1'b0 ;
  assign n7011 = n475 | n2744 ;
  assign n7013 = n7012 ^ n7011 ^ 1'b0 ;
  assign n7014 = n7013 ^ n2538 ^ 1'b0 ;
  assign n7015 = n7010 & n7014 ;
  assign n7016 = n3752 ^ n3612 ^ 1'b0 ;
  assign n7017 = n4765 & n7016 ;
  assign n7018 = n3169 & n7017 ;
  assign n7019 = n1465 | n7018 ;
  assign n7020 = ~n5633 & n7019 ;
  assign n7021 = n7020 ^ n1821 ^ 1'b0 ;
  assign n7022 = n5561 ^ n310 ^ 1'b0 ;
  assign n7023 = ( n6426 & n7021 ) | ( n6426 & n7022 ) | ( n7021 & n7022 ) ;
  assign n7024 = n990 & ~n2575 ;
  assign n7025 = ~n7023 & n7024 ;
  assign n7027 = n480 & ~n2897 ;
  assign n7028 = n1083 | n7027 ;
  assign n7029 = ( n3594 & n3657 ) | ( n3594 & ~n5933 ) | ( n3657 & ~n5933 ) ;
  assign n7030 = n7028 & n7029 ;
  assign n7031 = n7030 ^ x84 ^ 1'b0 ;
  assign n7026 = x118 | n5050 ;
  assign n7032 = n7031 ^ n7026 ^ 1'b0 ;
  assign n7033 = n2525 ^ n1765 ^ 1'b0 ;
  assign n7034 = n3343 & ~n7033 ;
  assign n7035 = n7034 ^ n2467 ^ 1'b0 ;
  assign n7036 = n5876 ^ n3428 ^ 1'b0 ;
  assign n7037 = n7035 & ~n7036 ;
  assign n7038 = n7037 ^ n1122 ^ 1'b0 ;
  assign n7039 = n4734 | n4864 ;
  assign n7040 = n408 | n7039 ;
  assign n7041 = n3922 ^ n1165 ^ n498 ;
  assign n7042 = ( n650 & n2348 ) | ( n650 & ~n7041 ) | ( n2348 & ~n7041 ) ;
  assign n7043 = n3948 & ~n4246 ;
  assign n7044 = n7042 & n7043 ;
  assign n7046 = n668 & n5928 ;
  assign n7045 = n2195 | n2654 ;
  assign n7047 = n7046 ^ n7045 ^ 1'b0 ;
  assign n7054 = n3212 ^ n2719 ^ 1'b0 ;
  assign n7048 = n1295 | n5459 ;
  assign n7050 = n2417 | n3151 ;
  assign n7051 = n2231 | n7050 ;
  assign n7049 = n4917 | n6552 ;
  assign n7052 = n7051 ^ n7049 ^ 1'b0 ;
  assign n7053 = n7048 & n7052 ;
  assign n7055 = n7054 ^ n7053 ^ 1'b0 ;
  assign n7056 = ( n398 & n1809 ) | ( n398 & ~n3554 ) | ( n1809 & ~n3554 ) ;
  assign n7057 = ( n290 & n4720 ) | ( n290 & ~n7056 ) | ( n4720 & ~n7056 ) ;
  assign n7058 = n986 | n5816 ;
  assign n7059 = n3247 & ~n7058 ;
  assign n7060 = n406 & ~n2346 ;
  assign n7061 = ~n3494 & n7060 ;
  assign n7062 = n6675 & n7061 ;
  assign n7063 = n150 & ~n5274 ;
  assign n7064 = ~n2236 & n7063 ;
  assign n7065 = n7064 ^ n3820 ^ 1'b0 ;
  assign n7066 = ~n269 & n2201 ;
  assign n7067 = n7066 ^ n4915 ^ 1'b0 ;
  assign n7068 = n7067 ^ n5754 ^ 1'b0 ;
  assign n7069 = ~n4703 & n4861 ;
  assign n7070 = ~n872 & n3436 ;
  assign n7071 = n7070 ^ n917 ^ 1'b0 ;
  assign n7076 = ~n1370 & n6223 ;
  assign n7072 = n1045 ^ n920 ^ x33 ;
  assign n7073 = n1516 ^ n806 ^ 1'b0 ;
  assign n7074 = n7072 & ~n7073 ;
  assign n7075 = n7074 ^ n3576 ^ 1'b0 ;
  assign n7077 = n7076 ^ n7075 ^ 1'b0 ;
  assign n7078 = n1639 | n7077 ;
  assign n7080 = n1742 & ~n2041 ;
  assign n7079 = n809 & n1010 ;
  assign n7081 = n7080 ^ n7079 ^ x100 ;
  assign n7082 = n1314 & n2866 ;
  assign n7083 = n7082 ^ n938 ^ 1'b0 ;
  assign n7084 = n5222 | n7083 ;
  assign n7085 = n1782 & ~n5040 ;
  assign n7086 = n2886 & ~n7085 ;
  assign n7087 = n236 | n2070 ;
  assign n7088 = n450 & n7087 ;
  assign n7089 = ~n1486 & n1757 ;
  assign n7090 = n2289 ^ n1514 ^ n1103 ;
  assign n7091 = n7090 ^ x109 ^ 1'b0 ;
  assign n7097 = n5745 ^ n1688 ^ 1'b0 ;
  assign n7098 = n7076 & n7097 ;
  assign n7093 = n5933 ^ n1026 ^ x25 ;
  assign n7094 = n7093 ^ n6451 ^ n1652 ;
  assign n7092 = ~n337 & n521 ;
  assign n7095 = n7094 ^ n7092 ^ 1'b0 ;
  assign n7096 = n1652 & n7095 ;
  assign n7099 = n7098 ^ n7096 ^ 1'b0 ;
  assign n7100 = ~n3997 & n6874 ;
  assign n7101 = ( n642 & ~n6687 ) | ( n642 & n7100 ) | ( ~n6687 & n7100 ) ;
  assign n7102 = n2046 & ~n5039 ;
  assign n7103 = n7102 ^ n4318 ^ 1'b0 ;
  assign n7104 = n7103 ^ n3374 ^ 1'b0 ;
  assign n7105 = n5924 ^ n4379 ^ 1'b0 ;
  assign n7106 = n7104 & n7105 ;
  assign n7108 = n2354 ^ n1658 ^ 1'b0 ;
  assign n7109 = ( n1224 & n1766 ) | ( n1224 & ~n7108 ) | ( n1766 & ~n7108 ) ;
  assign n7110 = n5431 | n7109 ;
  assign n7111 = n7110 ^ n3040 ^ 1'b0 ;
  assign n7107 = n3296 ^ n2736 ^ n805 ;
  assign n7112 = n7111 ^ n7107 ^ 1'b0 ;
  assign n7113 = n3488 | n3767 ;
  assign n7114 = ~n5342 & n7113 ;
  assign n7115 = n257 & n603 ;
  assign n7116 = n7115 ^ n2200 ^ 1'b0 ;
  assign n7117 = ~n657 & n7116 ;
  assign n7118 = n3151 & n5357 ;
  assign n7119 = ( n3259 & n7117 ) | ( n3259 & ~n7118 ) | ( n7117 & ~n7118 ) ;
  assign n7120 = ~n1839 & n2746 ;
  assign n7121 = n6821 & ~n7120 ;
  assign n7123 = n2234 ^ n1165 ^ 1'b0 ;
  assign n7122 = n1095 & n1320 ;
  assign n7124 = n7123 ^ n7122 ^ 1'b0 ;
  assign n7125 = n4762 & n7124 ;
  assign n7126 = n7125 ^ n2750 ^ 1'b0 ;
  assign n7127 = ( n1010 & n3419 ) | ( n1010 & n3887 ) | ( n3419 & n3887 ) ;
  assign n7128 = n7127 ^ n681 ^ 1'b0 ;
  assign n7129 = x84 & ~n692 ;
  assign n7130 = n3946 & ~n7129 ;
  assign n7131 = n1674 & ~n3829 ;
  assign n7132 = ~n1854 & n7131 ;
  assign n7133 = n7132 ^ n861 ^ 1'b0 ;
  assign n7134 = n3479 & n5010 ;
  assign n7135 = ~n6310 & n7134 ;
  assign n7136 = ~n1235 & n4156 ;
  assign n7137 = n7136 ^ n6116 ^ 1'b0 ;
  assign n7138 = ~n3705 & n7137 ;
  assign n7141 = n6700 ^ n3674 ^ 1'b0 ;
  assign n7142 = ~n3117 & n7141 ;
  assign n7139 = n5307 ^ n764 ^ 1'b0 ;
  assign n7140 = ~n5278 & n7139 ;
  assign n7143 = n7142 ^ n7140 ^ 1'b0 ;
  assign n7144 = n754 & n2151 ;
  assign n7145 = ~x58 & n7144 ;
  assign n7146 = n1117 & ~n3626 ;
  assign n7147 = n2582 ^ n1989 ^ 1'b0 ;
  assign n7148 = ~n1781 & n2354 ;
  assign n7149 = n7148 ^ n2291 ^ 1'b0 ;
  assign n7150 = n7147 & n7149 ;
  assign n7151 = ~n849 & n3153 ;
  assign n7152 = n661 & n7151 ;
  assign n7153 = ~n7150 & n7152 ;
  assign n7154 = n683 | n2157 ;
  assign n7155 = x114 & ~n1318 ;
  assign n7156 = n7155 ^ n395 ^ 1'b0 ;
  assign n7157 = n3424 & n4777 ;
  assign n7158 = n7156 & n7157 ;
  assign n7159 = n1805 | n3036 ;
  assign n7160 = n7159 ^ n343 ^ 1'b0 ;
  assign n7161 = n1373 & ~n7160 ;
  assign n7162 = n3145 & n7161 ;
  assign n7163 = ( ~n2543 & n4202 ) | ( ~n2543 & n7162 ) | ( n4202 & n7162 ) ;
  assign n7164 = n7163 ^ n899 ^ 1'b0 ;
  assign n7165 = n6602 | n7164 ;
  assign n7166 = ~n7158 & n7165 ;
  assign n7167 = n5050 ^ n4693 ^ 1'b0 ;
  assign n7168 = n3567 ^ n2112 ^ 1'b0 ;
  assign n7169 = n7167 & n7168 ;
  assign n7170 = n5897 ^ n5461 ^ 1'b0 ;
  assign n7171 = n6488 ^ n6190 ^ 1'b0 ;
  assign n7172 = n3026 ^ n2922 ^ 1'b0 ;
  assign n7173 = n1589 & n4406 ;
  assign n7174 = n3694 ^ n368 ^ 1'b0 ;
  assign n7175 = n2791 ^ x110 ^ 1'b0 ;
  assign n7176 = n835 & ~n7175 ;
  assign n7177 = n7176 ^ n3546 ^ n2316 ;
  assign n7178 = n7174 & ~n7177 ;
  assign n7184 = n3633 ^ n2334 ^ 1'b0 ;
  assign n7185 = ~n2696 & n7184 ;
  assign n7180 = x10 & n1151 ;
  assign n7181 = n7180 ^ n5318 ^ 1'b0 ;
  assign n7179 = x47 & ~n4796 ;
  assign n7182 = n7181 ^ n7179 ^ 1'b0 ;
  assign n7183 = n4909 & n7182 ;
  assign n7186 = n7185 ^ n7183 ^ 1'b0 ;
  assign n7187 = n7178 & ~n7186 ;
  assign n7188 = n2137 ^ n555 ^ 1'b0 ;
  assign n7189 = n2729 & n7188 ;
  assign n7190 = n7189 ^ n2507 ^ 1'b0 ;
  assign n7191 = n2818 ^ x3 ^ 1'b0 ;
  assign n7192 = n671 | n7191 ;
  assign n7193 = ~n6790 & n7192 ;
  assign n7194 = n6194 ^ n2021 ^ 1'b0 ;
  assign n7195 = n2393 & ~n7194 ;
  assign n7196 = n1408 | n7195 ;
  assign n7197 = n2147 | n7196 ;
  assign n7198 = n6520 ^ n1741 ^ 1'b0 ;
  assign n7199 = n6114 & n7198 ;
  assign n7200 = n1143 & n7199 ;
  assign n7201 = n3243 & ~n4071 ;
  assign n7202 = n740 | n7201 ;
  assign n7203 = n7200 & ~n7202 ;
  assign n7204 = n256 & n5870 ;
  assign n7207 = n462 ^ n220 ^ 1'b0 ;
  assign n7205 = ~n1072 & n1258 ;
  assign n7206 = n7205 ^ n6782 ^ 1'b0 ;
  assign n7208 = n7207 ^ n7206 ^ 1'b0 ;
  assign n7209 = n2917 | n5387 ;
  assign n7210 = n1796 & ~n7209 ;
  assign n7211 = n4453 | n6758 ;
  assign n7212 = n7211 ^ n4231 ^ 1'b0 ;
  assign n7213 = n1341 & ~n3583 ;
  assign n7214 = n7213 ^ n5247 ^ 1'b0 ;
  assign n7215 = ~n2061 & n7214 ;
  assign n7216 = n6511 ^ x108 ^ 1'b0 ;
  assign n7217 = n651 & n7216 ;
  assign n7218 = n5523 & n7217 ;
  assign n7219 = n4217 ^ n1122 ^ 1'b0 ;
  assign n7220 = ( n2112 & ~n3610 ) | ( n2112 & n7219 ) | ( ~n3610 & n7219 ) ;
  assign n7221 = x118 & ~n6049 ;
  assign n7222 = n1193 & n7221 ;
  assign n7223 = n1057 | n7222 ;
  assign n7224 = n2380 ^ n466 ^ 1'b0 ;
  assign n7225 = n7223 & n7224 ;
  assign n7226 = n2667 & ~n2818 ;
  assign n7227 = n2355 & ~n5742 ;
  assign n7228 = n421 & ~n475 ;
  assign n7229 = ~x71 & n7228 ;
  assign n7230 = n3751 & ~n7229 ;
  assign n7231 = n7230 ^ n290 ^ 1'b0 ;
  assign n7232 = n4241 | n4847 ;
  assign n7233 = ~n7231 & n7232 ;
  assign n7234 = n3655 ^ n348 ^ 1'b0 ;
  assign n7235 = ~n686 & n7234 ;
  assign n7236 = x46 & ~n311 ;
  assign n7237 = n2958 ^ n2827 ^ 1'b0 ;
  assign n7238 = ~n2132 & n7237 ;
  assign n7239 = n4902 ^ n1153 ^ 1'b0 ;
  assign n7240 = ~n1990 & n3861 ;
  assign n7241 = n2334 ^ n539 ^ n461 ;
  assign n7242 = n6532 ^ n4220 ^ 1'b0 ;
  assign n7243 = n4762 ^ n2058 ^ x121 ;
  assign n7244 = n2340 & n6221 ;
  assign n7245 = n7243 & n7244 ;
  assign n7246 = ~n2389 & n2908 ;
  assign n7247 = n7246 ^ n6908 ^ 1'b0 ;
  assign n7248 = n7247 ^ n3488 ^ 1'b0 ;
  assign n7249 = ~n5583 & n7248 ;
  assign n7250 = n6049 ^ n3474 ^ 1'b0 ;
  assign n7251 = n2257 & ~n7250 ;
  assign n7252 = n1260 | n2039 ;
  assign n7253 = n7252 ^ n1021 ^ 1'b0 ;
  assign n7254 = ~n7251 & n7253 ;
  assign n7255 = n1637 ^ n938 ^ 1'b0 ;
  assign n7257 = n2036 ^ n1407 ^ 1'b0 ;
  assign n7258 = n928 | n7257 ;
  assign n7256 = n5084 ^ x59 ^ 1'b0 ;
  assign n7259 = n7258 ^ n7256 ^ 1'b0 ;
  assign n7260 = ~n3687 & n4249 ;
  assign n7261 = x12 & ~n2853 ;
  assign n7262 = ~n3170 & n7261 ;
  assign n7263 = n4817 ^ n1749 ^ 1'b0 ;
  assign n7264 = n652 | n5188 ;
  assign n7265 = n3808 | n7264 ;
  assign n7266 = n3585 & ~n7265 ;
  assign n7267 = n7266 ^ n1000 ^ 1'b0 ;
  assign n7268 = n2081 | n7267 ;
  assign n7269 = n2270 & n6968 ;
  assign n7270 = x125 & n7269 ;
  assign n7271 = n2189 & n7270 ;
  assign n7272 = n2681 & n3474 ;
  assign n7273 = n1695 | n7272 ;
  assign n7274 = n7271 & ~n7273 ;
  assign n7275 = ( x114 & ~n1713 ) | ( x114 & n4902 ) | ( ~n1713 & n4902 ) ;
  assign n7276 = n7275 ^ n5941 ^ 1'b0 ;
  assign n7277 = n5452 & n7276 ;
  assign n7278 = x21 & n7277 ;
  assign n7279 = n7274 & n7278 ;
  assign n7280 = n6787 ^ n3947 ^ 1'b0 ;
  assign n7281 = n1627 & n3434 ;
  assign n7282 = n7087 & n7281 ;
  assign n7283 = ~n2451 & n2824 ;
  assign n7284 = n7282 & n7283 ;
  assign n7285 = n2064 | n7284 ;
  assign n7286 = n7280 & ~n7285 ;
  assign n7287 = n3563 | n4404 ;
  assign n7288 = n2099 & n2930 ;
  assign n7289 = n5116 ^ n4989 ^ 1'b0 ;
  assign n7290 = n5149 ^ n3200 ^ n383 ;
  assign n7291 = n367 & n3058 ;
  assign n7292 = n2064 & n7291 ;
  assign n7293 = n7292 ^ n5444 ^ 1'b0 ;
  assign n7294 = ~n1303 & n7293 ;
  assign n7295 = n2063 ^ n988 ^ 1'b0 ;
  assign n7296 = ~n5632 & n7295 ;
  assign n7297 = n2529 ^ n1855 ^ n236 ;
  assign n7298 = n5935 & n6860 ;
  assign n7299 = n2760 ^ n2544 ^ 1'b0 ;
  assign n7300 = ~n605 & n4695 ;
  assign n7301 = n7300 ^ n4085 ^ 1'b0 ;
  assign n7302 = n7301 ^ n2706 ^ 1'b0 ;
  assign n7303 = n7299 & ~n7302 ;
  assign n7304 = n6791 ^ n1481 ^ 1'b0 ;
  assign n7305 = n6627 ^ n664 ^ 1'b0 ;
  assign n7306 = n7305 ^ n1532 ^ 1'b0 ;
  assign n7307 = n5371 & ~n6746 ;
  assign n7308 = n7307 ^ n1765 ^ 1'b0 ;
  assign n7309 = n1375 | n7191 ;
  assign n7310 = ~n2036 & n2391 ;
  assign n7311 = ~n2649 & n7310 ;
  assign n7312 = n7311 ^ n979 ^ n436 ;
  assign n7313 = ( n6196 & n7035 ) | ( n6196 & ~n7312 ) | ( n7035 & ~n7312 ) ;
  assign n7314 = n1372 & ~n6145 ;
  assign n7315 = n7033 ^ n1981 ^ 1'b0 ;
  assign n7316 = ( n6049 & n7314 ) | ( n6049 & ~n7315 ) | ( n7314 & ~n7315 ) ;
  assign n7317 = n1050 & ~n5093 ;
  assign n7318 = n1452 | n7317 ;
  assign n7319 = n7318 ^ n7114 ^ 1'b0 ;
  assign n7320 = n2252 & n7319 ;
  assign n7321 = n2945 ^ n2850 ^ x47 ;
  assign n7322 = n5249 ^ n1459 ^ 1'b0 ;
  assign n7323 = ~n3470 & n7322 ;
  assign n7324 = n4186 | n7323 ;
  assign n7325 = n3363 ^ n3259 ^ 1'b0 ;
  assign n7326 = ( ~n2334 & n3625 ) | ( ~n2334 & n5492 ) | ( n3625 & n5492 ) ;
  assign n7327 = n4082 & ~n4503 ;
  assign n7328 = n2554 & n7327 ;
  assign n7329 = n4946 | n7328 ;
  assign n7330 = n6687 ^ n5425 ^ n2397 ;
  assign n7331 = ~n1757 & n2676 ;
  assign n7332 = n2720 & n7331 ;
  assign n7333 = n2229 & ~n7332 ;
  assign n7334 = n7332 & n7333 ;
  assign n7335 = n909 | n2428 ;
  assign n7336 = n910 & ~n7335 ;
  assign n7337 = n7336 ^ n2064 ^ 1'b0 ;
  assign n7338 = ( n907 & ~n7334 ) | ( n907 & n7337 ) | ( ~n7334 & n7337 ) ;
  assign n7339 = n2823 & ~n3208 ;
  assign n7340 = n3243 & ~n3966 ;
  assign n7341 = ( n551 & n616 ) | ( n551 & ~n1490 ) | ( n616 & ~n1490 ) ;
  assign n7348 = n1799 & ~n6771 ;
  assign n7349 = n7348 ^ n2527 ^ 1'b0 ;
  assign n7350 = n1861 & ~n7349 ;
  assign n7346 = n1399 ^ n590 ^ 1'b0 ;
  assign n7344 = n2451 & n4537 ;
  assign n7342 = ~x81 & n5900 ;
  assign n7343 = n3574 & n7342 ;
  assign n7345 = n7344 ^ n7343 ^ 1'b0 ;
  assign n7347 = n7346 ^ n7345 ^ 1'b0 ;
  assign n7351 = n7350 ^ n7347 ^ n2706 ;
  assign n7352 = n4023 & ~n4933 ;
  assign n7353 = n376 & n5758 ;
  assign n7354 = n2041 & ~n4159 ;
  assign n7355 = n3525 & n7354 ;
  assign n7356 = n5941 & ~n7355 ;
  assign n7357 = n7353 & n7356 ;
  assign n7358 = n406 & n7093 ;
  assign n7362 = ~n1860 & n3583 ;
  assign n7359 = n2694 & n2959 ;
  assign n7360 = n3766 | n7359 ;
  assign n7361 = n1445 | n7360 ;
  assign n7363 = n7362 ^ n7361 ^ 1'b0 ;
  assign n7364 = n6287 & n7363 ;
  assign n7365 = n7358 & n7364 ;
  assign n7366 = n3080 & ~n5971 ;
  assign n7367 = n7366 ^ n3055 ^ 1'b0 ;
  assign n7368 = n4270 ^ n3775 ^ n463 ;
  assign n7369 = ~n6058 & n7368 ;
  assign n7370 = n7369 ^ n1476 ^ 1'b0 ;
  assign n7371 = n7370 ^ n4952 ^ 1'b0 ;
  assign n7372 = ~n3447 & n7371 ;
  assign n7373 = n725 & ~n1610 ;
  assign n7374 = ~n370 & n7373 ;
  assign n7375 = n1416 ^ n730 ^ 1'b0 ;
  assign n7376 = n850 | n7375 ;
  assign n7377 = n7376 ^ n4777 ^ 1'b0 ;
  assign n7378 = n1436 ^ n1335 ^ 1'b0 ;
  assign n7379 = n7377 & n7378 ;
  assign n7380 = n7379 ^ n4868 ^ n2246 ;
  assign n7381 = x3 & n4782 ;
  assign n7382 = n1014 & n7381 ;
  assign n7383 = n2859 & n6694 ;
  assign n7384 = n840 & n2256 ;
  assign n7385 = n1771 ^ n1594 ^ 1'b0 ;
  assign n7386 = n5986 & ~n7385 ;
  assign n7387 = n794 | n5466 ;
  assign n7388 = n2754 & ~n7387 ;
  assign n7389 = n7388 ^ n6607 ^ x51 ;
  assign n7390 = n6087 ^ n2329 ^ 1'b0 ;
  assign n7391 = n6109 ^ n3082 ^ 1'b0 ;
  assign n7392 = n6807 & n7391 ;
  assign n7393 = n4025 & n7392 ;
  assign n7395 = n4184 ^ n3253 ^ 1'b0 ;
  assign n7396 = n431 & n2186 ;
  assign n7397 = n7396 ^ n5503 ^ 1'b0 ;
  assign n7398 = n7395 | n7397 ;
  assign n7394 = n808 | n4791 ;
  assign n7399 = n7398 ^ n7394 ^ 1'b0 ;
  assign n7400 = n2354 & ~n4898 ;
  assign n7401 = ~n569 & n858 ;
  assign n7402 = n7401 ^ n4340 ^ 1'b0 ;
  assign n7403 = n5113 & ~n7402 ;
  assign n7404 = n3783 & n5598 ;
  assign n7405 = ~n3783 & n7404 ;
  assign n7406 = n6862 | n7405 ;
  assign n7407 = n7403 & ~n7406 ;
  assign n7408 = n3070 ^ n1966 ^ n1765 ;
  assign n7409 = n5255 ^ n2304 ^ 1'b0 ;
  assign n7410 = n7408 | n7409 ;
  assign n7411 = n7410 ^ n748 ^ 1'b0 ;
  assign n7412 = n1450 & n7411 ;
  assign n7413 = n7412 ^ n4919 ^ 1'b0 ;
  assign n7414 = n694 | n798 ;
  assign n7415 = n3857 & ~n7414 ;
  assign n7416 = n7415 ^ n895 ^ 1'b0 ;
  assign n7417 = n7416 ^ n1539 ^ 1'b0 ;
  assign n7418 = ~n3794 & n7417 ;
  assign n7420 = n821 & ~n4012 ;
  assign n7419 = n283 & ~n3187 ;
  assign n7421 = n7420 ^ n7419 ^ 1'b0 ;
  assign n7422 = n1607 | n5463 ;
  assign n7423 = ~n984 & n4572 ;
  assign n7424 = n2608 & n7423 ;
  assign n7425 = n3868 ^ n2051 ^ n1711 ;
  assign n7426 = n3562 ^ n138 ^ 1'b0 ;
  assign n7427 = ~n7425 & n7426 ;
  assign n7428 = ~n2577 & n7427 ;
  assign n7429 = ( ~n385 & n3354 ) | ( ~n385 & n3710 ) | ( n3354 & n3710 ) ;
  assign n7430 = n4749 | n7429 ;
  assign n7431 = n2783 | n6742 ;
  assign n7432 = n7430 & ~n7431 ;
  assign n7434 = n2283 ^ n869 ^ 1'b0 ;
  assign n7435 = n2642 | n7434 ;
  assign n7436 = n7435 ^ n2581 ^ 1'b0 ;
  assign n7433 = n5013 | n6308 ;
  assign n7437 = n7436 ^ n7433 ^ 1'b0 ;
  assign n7438 = ~n3316 & n7437 ;
  assign n7439 = n4347 ^ n2873 ^ n485 ;
  assign n7440 = ( x69 & ~n1352 ) | ( x69 & n1596 ) | ( ~n1352 & n1596 ) ;
  assign n7441 = n7440 ^ n2233 ^ 1'b0 ;
  assign n7442 = n7439 & ~n7441 ;
  assign n7443 = ~n2694 & n3583 ;
  assign n7444 = n4972 & n7443 ;
  assign n7445 = n2304 ^ n431 ^ x126 ;
  assign n7446 = x38 & n7445 ;
  assign n7447 = n7444 & ~n7446 ;
  assign n7448 = n7447 ^ n6815 ^ 1'b0 ;
  assign n7449 = ~n4085 & n4462 ;
  assign n7450 = n5514 ^ n967 ^ 1'b0 ;
  assign n7451 = n7403 & ~n7450 ;
  assign n7452 = n2811 ^ n717 ^ 1'b0 ;
  assign n7453 = n7452 ^ n1880 ^ 1'b0 ;
  assign n7454 = n3117 ^ n1205 ^ 1'b0 ;
  assign n7455 = ( x2 & n331 ) | ( x2 & n7454 ) | ( n331 & n7454 ) ;
  assign n7456 = n2839 & ~n3332 ;
  assign n7457 = ~n1938 & n7456 ;
  assign n7458 = ( x18 & ~x92 ) | ( x18 & n2760 ) | ( ~x92 & n2760 ) ;
  assign n7459 = n5536 ^ n570 ^ 1'b0 ;
  assign n7460 = n7458 & n7459 ;
  assign n7462 = n918 | n2346 ;
  assign n7461 = n1610 & ~n3857 ;
  assign n7463 = n7462 ^ n7461 ^ n454 ;
  assign n7464 = n3596 | n4061 ;
  assign n7465 = n5059 | n7464 ;
  assign n7466 = n2055 & ~n2341 ;
  assign n7467 = n7466 ^ n3699 ^ 1'b0 ;
  assign n7468 = n191 & n2729 ;
  assign n7469 = n7468 ^ n615 ^ 1'b0 ;
  assign n7470 = n3662 & ~n4655 ;
  assign n7471 = ~n1962 & n7470 ;
  assign n7472 = n3619 ^ n367 ^ 1'b0 ;
  assign n7473 = n7472 ^ n1914 ^ n1471 ;
  assign n7474 = n1374 | n7473 ;
  assign n7475 = n3057 & ~n7474 ;
  assign n7476 = ( ~n7469 & n7471 ) | ( ~n7469 & n7475 ) | ( n7471 & n7475 ) ;
  assign n7477 = n2485 & n7476 ;
  assign n7478 = ~n7467 & n7477 ;
  assign n7479 = ( ~n467 & n5523 ) | ( ~n467 & n6397 ) | ( n5523 & n6397 ) ;
  assign n7480 = n2384 & ~n2632 ;
  assign n7481 = n7480 ^ n4042 ^ n3857 ;
  assign n7482 = ~n1935 & n7481 ;
  assign n7484 = n3340 ^ n1443 ^ 1'b0 ;
  assign n7483 = n1450 & n5361 ;
  assign n7485 = n7484 ^ n7483 ^ 1'b0 ;
  assign n7486 = n849 | n3688 ;
  assign n7487 = n7486 ^ n2016 ^ 1'b0 ;
  assign n7488 = n1839 & n7487 ;
  assign n7489 = ~n3033 & n4385 ;
  assign n7490 = ( n1578 & n5338 ) | ( n1578 & ~n5848 ) | ( n5338 & ~n5848 ) ;
  assign n7491 = ( n5166 & ~n7489 ) | ( n5166 & n7490 ) | ( ~n7489 & n7490 ) ;
  assign n7492 = n2197 ^ n408 ^ 1'b0 ;
  assign n7493 = n1794 & n7492 ;
  assign n7494 = ~n2706 & n7493 ;
  assign n7495 = n7494 ^ n1802 ^ 1'b0 ;
  assign n7496 = n7495 ^ n2321 ^ 1'b0 ;
  assign n7501 = n2529 ^ n372 ^ 1'b0 ;
  assign n7497 = n1379 ^ x91 ^ 1'b0 ;
  assign n7498 = n2299 | n5875 ;
  assign n7499 = n7498 ^ n5347 ^ 1'b0 ;
  assign n7500 = n7497 & ~n7499 ;
  assign n7502 = n7501 ^ n7500 ^ 1'b0 ;
  assign n7503 = n6523 ^ n1123 ^ n625 ;
  assign n7504 = n7503 ^ n2085 ^ 1'b0 ;
  assign n7505 = ~n3618 & n7504 ;
  assign n7506 = ~n370 & n7505 ;
  assign n7507 = n283 & ~n7506 ;
  assign n7508 = n6018 & n7507 ;
  assign n7509 = ~n1424 & n7508 ;
  assign n7510 = n6264 ^ n4343 ^ 1'b0 ;
  assign n7511 = ~n7509 & n7510 ;
  assign n7513 = n4211 ^ n3345 ^ n2433 ;
  assign n7512 = x57 & ~n4373 ;
  assign n7514 = n7513 ^ n7512 ^ 1'b0 ;
  assign n7515 = ~n1029 & n1966 ;
  assign n7516 = n7515 ^ n3044 ^ 1'b0 ;
  assign n7517 = n6248 ^ n1171 ^ 1'b0 ;
  assign n7518 = n3727 & n7517 ;
  assign n7519 = n1046 & ~n1366 ;
  assign n7520 = n899 & n7519 ;
  assign n7521 = n2380 & ~n7520 ;
  assign n7522 = ( x118 & n4398 ) | ( x118 & ~n7521 ) | ( n4398 & ~n7521 ) ;
  assign n7523 = ( ~n3770 & n7033 ) | ( ~n3770 & n7522 ) | ( n7033 & n7522 ) ;
  assign n7524 = ( n5999 & n7518 ) | ( n5999 & n7523 ) | ( n7518 & n7523 ) ;
  assign n7525 = n5812 ^ n2969 ^ n1291 ;
  assign n7526 = n1837 | n5551 ;
  assign n7527 = n7027 ^ n5630 ^ 1'b0 ;
  assign n7532 = n2467 | n3163 ;
  assign n7533 = n3138 | n7532 ;
  assign n7528 = n1528 ^ n1514 ^ 1'b0 ;
  assign n7529 = n3712 & ~n7528 ;
  assign n7530 = n7529 ^ n236 ^ 1'b0 ;
  assign n7531 = n6399 & n7530 ;
  assign n7534 = n7533 ^ n7531 ^ 1'b0 ;
  assign n7535 = n4777 & ~n7534 ;
  assign n7536 = n7535 ^ n3315 ^ 1'b0 ;
  assign n7537 = ~n1033 & n1134 ;
  assign n7538 = n186 & n7537 ;
  assign n7539 = n3679 | n7538 ;
  assign n7540 = n259 | n1013 ;
  assign n7541 = n1013 & ~n7540 ;
  assign n7542 = n279 & n1961 ;
  assign n7543 = ~n1961 & n7542 ;
  assign n7544 = n7541 & ~n7543 ;
  assign n7545 = ( ~n2958 & n6497 ) | ( ~n2958 & n7544 ) | ( n6497 & n7544 ) ;
  assign n7546 = n593 & n2574 ;
  assign n7547 = n190 | n7546 ;
  assign n7548 = n362 & n1732 ;
  assign n7549 = ~x79 & n7548 ;
  assign n7550 = x76 & n7549 ;
  assign n7551 = n4975 & n7550 ;
  assign n7552 = n5250 & n7551 ;
  assign n7553 = n7552 ^ n4071 ^ 1'b0 ;
  assign n7554 = n4123 | n5459 ;
  assign n7555 = n7506 & ~n7554 ;
  assign n7556 = n3277 & n7555 ;
  assign n7557 = ~n7553 & n7556 ;
  assign n7558 = ~n509 & n962 ;
  assign n7559 = ( ~n549 & n1637 ) | ( ~n549 & n7558 ) | ( n1637 & n7558 ) ;
  assign n7560 = n6770 ^ x2 ^ 1'b0 ;
  assign n7561 = ( n1175 & n1450 ) | ( n1175 & n5188 ) | ( n1450 & n5188 ) ;
  assign n7562 = n7561 ^ n3384 ^ 1'b0 ;
  assign n7563 = n3630 & ~n3694 ;
  assign n7564 = n7563 ^ n4806 ^ 1'b0 ;
  assign n7565 = ( ~n1213 & n2840 ) | ( ~n1213 & n5813 ) | ( n2840 & n5813 ) ;
  assign n7566 = n7565 ^ n770 ^ 1'b0 ;
  assign n7567 = ( n4913 & n7564 ) | ( n4913 & n7566 ) | ( n7564 & n7566 ) ;
  assign n7568 = n1462 | n3878 ;
  assign n7569 = n7568 ^ n3111 ^ 1'b0 ;
  assign n7570 = n4883 & ~n7569 ;
  assign n7571 = n3788 ^ n802 ^ 1'b0 ;
  assign n7572 = n6287 & ~n7571 ;
  assign n7573 = n7572 ^ n2489 ^ 1'b0 ;
  assign n7574 = n7528 ^ n4110 ^ 1'b0 ;
  assign n7575 = n5687 | n7574 ;
  assign n7576 = n7575 ^ n6959 ^ 1'b0 ;
  assign n7577 = ~n2673 & n3559 ;
  assign n7578 = ( n2170 & n3179 ) | ( n2170 & ~n4860 ) | ( n3179 & ~n4860 ) ;
  assign n7579 = ~n571 & n7578 ;
  assign n7580 = ( n399 & n7577 ) | ( n399 & n7579 ) | ( n7577 & n7579 ) ;
  assign n7581 = n7528 ^ n7129 ^ n2868 ;
  assign n7582 = n7581 ^ n5592 ^ n5331 ;
  assign n7583 = n7582 ^ n510 ^ 1'b0 ;
  assign n7584 = n1033 ^ n403 ^ 1'b0 ;
  assign n7585 = n7584 ^ n4286 ^ 1'b0 ;
  assign n7586 = ~n6797 & n7585 ;
  assign n7587 = n7586 ^ n6685 ^ 1'b0 ;
  assign n7588 = n643 ^ x103 ^ 1'b0 ;
  assign n7589 = n3339 ^ n2102 ^ 1'b0 ;
  assign n7590 = n7589 ^ n725 ^ 1'b0 ;
  assign n7591 = n7588 & n7590 ;
  assign n7592 = n1407 ^ n1203 ^ 1'b0 ;
  assign n7593 = n3156 & ~n7592 ;
  assign n7594 = ~n7591 & n7593 ;
  assign n7595 = n6991 ^ n2292 ^ 1'b0 ;
  assign n7596 = n3079 & ~n4150 ;
  assign n7597 = ~n2570 & n7596 ;
  assign n7598 = n7362 | n7597 ;
  assign n7599 = n7598 ^ n227 ^ 1'b0 ;
  assign n7600 = ~n369 & n1876 ;
  assign n7601 = n366 & n7600 ;
  assign n7602 = n483 & ~n616 ;
  assign n7603 = n7601 | n7602 ;
  assign n7604 = n7599 & ~n7603 ;
  assign n7605 = n2199 | n2376 ;
  assign n7606 = n4828 | n7605 ;
  assign n7607 = n243 & n4765 ;
  assign n7608 = n7606 | n7607 ;
  assign n7609 = n280 & ~n1175 ;
  assign n7612 = ~n369 & n7123 ;
  assign n7613 = ~n2663 & n7612 ;
  assign n7610 = n6488 & n6647 ;
  assign n7611 = n5258 & ~n7610 ;
  assign n7614 = n7613 ^ n7611 ^ 1'b0 ;
  assign n7615 = n3182 & ~n4337 ;
  assign n7616 = n2325 & n7615 ;
  assign n7617 = n1961 & n5675 ;
  assign n7618 = ~n703 & n7617 ;
  assign n7619 = n1958 ^ n490 ^ 1'b0 ;
  assign n7620 = ( n5141 & n5165 ) | ( n5141 & ~n6304 ) | ( n5165 & ~n6304 ) ;
  assign n7621 = n1868 ^ n185 ^ 1'b0 ;
  assign n7622 = n7620 & ~n7621 ;
  assign n7623 = n3414 | n5256 ;
  assign n7624 = n2164 | n7370 ;
  assign n7625 = n1236 | n7624 ;
  assign n7626 = ( n1088 & ~n3055 ) | ( n1088 & n7200 ) | ( ~n3055 & n7200 ) ;
  assign n7627 = n680 | n3759 ;
  assign n7628 = n7626 & n7627 ;
  assign n7629 = ~n7005 & n7628 ;
  assign n7630 = n2490 | n7629 ;
  assign n7631 = n7038 ^ n4279 ^ n383 ;
  assign n7632 = ( n149 & ~n179 ) | ( n149 & n1003 ) | ( ~n179 & n1003 ) ;
  assign n7633 = n4469 & n7632 ;
  assign n7634 = n3989 ^ n1970 ^ 1'b0 ;
  assign n7635 = n7633 | n7634 ;
  assign n7636 = ~x16 & n5223 ;
  assign n7637 = n7636 ^ n3217 ^ 1'b0 ;
  assign n7638 = n7637 ^ n863 ^ 1'b0 ;
  assign n7639 = ( n1630 & n2780 ) | ( n1630 & ~n4585 ) | ( n2780 & ~n4585 ) ;
  assign n7640 = n1258 | n7639 ;
  assign n7641 = n6691 | n7640 ;
  assign n7644 = n2180 ^ n1519 ^ 1'b0 ;
  assign n7645 = n2209 & ~n7644 ;
  assign n7646 = n7645 ^ n2622 ^ 1'b0 ;
  assign n7647 = n7646 ^ n4247 ^ n3453 ;
  assign n7642 = n1906 & n6102 ;
  assign n7643 = n2637 | n7642 ;
  assign n7648 = n7647 ^ n7643 ^ 1'b0 ;
  assign n7649 = n7312 ^ n1957 ^ n1208 ;
  assign n7652 = ( n2837 & n3906 ) | ( n2837 & n4038 ) | ( n3906 & n4038 ) ;
  assign n7653 = n2229 ^ n182 ^ 1'b0 ;
  assign n7654 = ~n3916 & n7653 ;
  assign n7655 = n5078 | n7654 ;
  assign n7656 = n1879 & ~n7655 ;
  assign n7657 = n6571 & n7656 ;
  assign n7658 = n7652 & ~n7657 ;
  assign n7650 = n4006 ^ n904 ^ 1'b0 ;
  assign n7651 = ( n193 & n6271 ) | ( n193 & ~n7650 ) | ( n6271 & ~n7650 ) ;
  assign n7659 = n7658 ^ n7651 ^ 1'b0 ;
  assign n7660 = x15 & n7659 ;
  assign n7661 = n6829 ^ n1655 ^ 1'b0 ;
  assign n7662 = n4194 | n7661 ;
  assign n7663 = ~n1656 & n7662 ;
  assign n7664 = ~n350 & n7663 ;
  assign n7665 = ~n3307 & n7664 ;
  assign n7666 = n3961 | n7665 ;
  assign n7667 = n7251 ^ n2768 ^ 1'b0 ;
  assign n7668 = n1784 & ~n1827 ;
  assign n7669 = n7444 ^ n4667 ^ 1'b0 ;
  assign n7670 = n842 & ~n7669 ;
  assign n7671 = ~n7581 & n7670 ;
  assign n7672 = ~n7668 & n7671 ;
  assign n7673 = n5326 & n5923 ;
  assign n7678 = ~n707 & n6895 ;
  assign n7679 = n7678 ^ n3367 ^ 1'b0 ;
  assign n7680 = n346 | n7679 ;
  assign n7681 = n1236 & n7680 ;
  assign n7674 = n4272 & ~n7504 ;
  assign n7675 = n2717 ^ n1644 ^ 1'b0 ;
  assign n7676 = n7674 & ~n7675 ;
  assign n7677 = n4844 & n7676 ;
  assign n7682 = n7681 ^ n7677 ^ 1'b0 ;
  assign n7683 = n6530 ^ n6196 ^ n5326 ;
  assign n7684 = n6497 ^ n3041 ^ 1'b0 ;
  assign n7685 = n4479 & n7684 ;
  assign n7686 = n2622 | n2671 ;
  assign n7687 = n1572 | n7686 ;
  assign n7688 = n5029 ^ n3838 ^ 1'b0 ;
  assign n7689 = n7688 ^ n5265 ^ 1'b0 ;
  assign n7690 = n2751 | n3869 ;
  assign n7691 = n7690 ^ n1297 ^ 1'b0 ;
  assign n7692 = n7165 | n7691 ;
  assign n7693 = n6261 ^ n323 ^ 1'b0 ;
  assign n7694 = n7693 ^ n3267 ^ 1'b0 ;
  assign n7695 = n3595 | n7694 ;
  assign n7696 = n1237 & ~n3958 ;
  assign n7697 = n7696 ^ n793 ^ 1'b0 ;
  assign n7698 = ( ~n2746 & n6707 ) | ( ~n2746 & n7697 ) | ( n6707 & n7697 ) ;
  assign n7699 = n750 | n5264 ;
  assign n7700 = n7699 ^ n7007 ^ 1'b0 ;
  assign n7701 = n362 | n1784 ;
  assign n7702 = n6176 & n7701 ;
  assign n7703 = n5423 & n7702 ;
  assign n7704 = n1072 ^ x120 ^ 1'b0 ;
  assign n7705 = n1008 | n7704 ;
  assign n7706 = n5369 & ~n7705 ;
  assign n7707 = n7706 ^ n4404 ^ 1'b0 ;
  assign n7708 = n7229 ^ n2169 ^ 1'b0 ;
  assign n7709 = ~n821 & n7708 ;
  assign n7710 = ~n1031 & n7709 ;
  assign n7711 = ~n2649 & n7710 ;
  assign n7712 = n7707 | n7711 ;
  assign n7713 = n7712 ^ n3528 ^ 1'b0 ;
  assign n7714 = n5567 ^ n1971 ^ n1109 ;
  assign n7715 = ( ~n692 & n6631 ) | ( ~n692 & n7714 ) | ( n6631 & n7714 ) ;
  assign n7716 = ( n1385 & ~n2090 ) | ( n1385 & n2420 ) | ( ~n2090 & n2420 ) ;
  assign n7717 = ( n977 & n2340 ) | ( n977 & ~n2900 ) | ( n2340 & ~n2900 ) ;
  assign n7718 = n4773 ^ n3556 ^ n957 ;
  assign n7719 = ~n3602 & n7718 ;
  assign n7720 = ( n7716 & n7717 ) | ( n7716 & n7719 ) | ( n7717 & n7719 ) ;
  assign n7721 = ( n738 & n2194 ) | ( n738 & ~n2699 ) | ( n2194 & ~n2699 ) ;
  assign n7722 = n1501 & ~n4462 ;
  assign n7723 = n7722 ^ n3237 ^ 1'b0 ;
  assign n7724 = n4674 ^ n3766 ^ n3401 ;
  assign n7725 = n3515 ^ n979 ^ 1'b0 ;
  assign n7726 = ~n5881 & n7725 ;
  assign n7727 = n3610 ^ n1912 ^ 1'b0 ;
  assign n7728 = n7727 ^ n5784 ^ 1'b0 ;
  assign n7729 = n7726 & n7728 ;
  assign n7730 = n1159 & n3569 ;
  assign n7731 = n7730 ^ n4306 ^ 1'b0 ;
  assign n7732 = n7124 ^ n1935 ^ 1'b0 ;
  assign n7733 = ~n4369 & n7732 ;
  assign n7734 = ~n7731 & n7733 ;
  assign n7735 = n7734 ^ n614 ^ 1'b0 ;
  assign n7736 = ( ~n161 & n3728 ) | ( ~n161 & n7528 ) | ( n3728 & n7528 ) ;
  assign n7737 = n7736 ^ n2354 ^ n1513 ;
  assign n7738 = n5608 ^ n1839 ^ 1'b0 ;
  assign n7739 = n4499 & n7738 ;
  assign n7740 = ( n1611 & n1626 ) | ( n1611 & ~n5517 ) | ( n1626 & ~n5517 ) ;
  assign n7741 = n1656 | n2831 ;
  assign n7742 = n7741 ^ n4650 ^ 1'b0 ;
  assign n7743 = n1977 & n7396 ;
  assign n7744 = n7743 ^ n7391 ^ n1097 ;
  assign n7745 = ~n6499 & n7744 ;
  assign n7746 = n7742 & n7745 ;
  assign n7747 = n2658 ^ n923 ^ 1'b0 ;
  assign n7748 = n2307 & n7747 ;
  assign n7749 = n2476 & n3252 ;
  assign n7750 = n409 & n7749 ;
  assign n7751 = n6840 & ~n7750 ;
  assign n7752 = n7751 ^ n2350 ^ 1'b0 ;
  assign n7753 = n2444 ^ n1673 ^ 1'b0 ;
  assign n7754 = n2154 & n7753 ;
  assign n7755 = ~n6662 & n7754 ;
  assign n7756 = n7755 ^ n4916 ^ 1'b0 ;
  assign n7757 = n2101 | n3574 ;
  assign n7758 = n2547 & n5913 ;
  assign n7759 = ( n4263 & n6247 ) | ( n4263 & ~n7758 ) | ( n6247 & ~n7758 ) ;
  assign n7760 = n1864 & n4623 ;
  assign n7761 = n7760 ^ n2074 ^ 1'b0 ;
  assign n7762 = n4850 ^ n2926 ^ n2053 ;
  assign n7763 = ~n331 & n7762 ;
  assign n7764 = ( n1742 & n2020 ) | ( n1742 & ~n7763 ) | ( n2020 & ~n7763 ) ;
  assign n7765 = n6036 | n7764 ;
  assign n7766 = n4610 | n7765 ;
  assign n7767 = n612 | n4821 ;
  assign n7768 = n2621 | n7767 ;
  assign n7769 = ( n2026 & n5166 ) | ( n2026 & n7768 ) | ( n5166 & n7768 ) ;
  assign n7770 = n7766 & n7769 ;
  assign n7771 = n7761 & n7770 ;
  assign n7772 = n2538 ^ n1669 ^ 1'b0 ;
  assign n7773 = ~n3028 & n7772 ;
  assign n7774 = ~n2462 & n6156 ;
  assign n7775 = n4835 ^ n4006 ^ 1'b0 ;
  assign n7776 = n6632 | n7775 ;
  assign n7777 = n2256 & ~n4701 ;
  assign n7778 = ~n6911 & n7777 ;
  assign n7779 = ~n5293 & n5785 ;
  assign n7780 = n7778 & n7779 ;
  assign n7781 = n5330 ^ n3879 ^ 1'b0 ;
  assign n7782 = n256 & ~n293 ;
  assign n7783 = n5813 & ~n7782 ;
  assign n7784 = n5416 & n7783 ;
  assign n7785 = ( ~n469 & n7781 ) | ( ~n469 & n7784 ) | ( n7781 & n7784 ) ;
  assign n7788 = n3422 & ~n4472 ;
  assign n7789 = n7788 ^ n4084 ^ 1'b0 ;
  assign n7786 = n1423 ^ n398 ^ 1'b0 ;
  assign n7787 = x16 | n7786 ;
  assign n7790 = n7789 ^ n7787 ^ n3298 ;
  assign n7791 = n7571 ^ n3216 ^ n1679 ;
  assign n7792 = ( ~n3518 & n3540 ) | ( ~n3518 & n4241 ) | ( n3540 & n4241 ) ;
  assign n7793 = n6143 ^ n3788 ^ n2222 ;
  assign n7794 = n7793 ^ n256 ^ 1'b0 ;
  assign n7796 = n325 & ~n3247 ;
  assign n7795 = n5541 ^ n1915 ^ 1'b0 ;
  assign n7797 = n7796 ^ n7795 ^ n1449 ;
  assign n7798 = ~n627 & n4222 ;
  assign n7799 = ( ~n135 & n2277 ) | ( ~n135 & n6353 ) | ( n2277 & n6353 ) ;
  assign n7800 = n7799 ^ n4511 ^ 1'b0 ;
  assign n7801 = n2206 & ~n5788 ;
  assign n7802 = n6877 | n7801 ;
  assign n7803 = ~n4032 & n5591 ;
  assign n7804 = n4204 ^ n876 ^ 1'b0 ;
  assign n7805 = n909 | n2024 ;
  assign n7806 = n7805 ^ n7253 ^ 1'b0 ;
  assign n7807 = n7806 ^ x92 ^ 1'b0 ;
  assign n7808 = n7804 & n7807 ;
  assign n7809 = ~n6168 & n7808 ;
  assign n7810 = n7809 ^ n2667 ^ 1'b0 ;
  assign n7811 = n7810 ^ n6954 ^ 1'b0 ;
  assign n7812 = ~n5316 & n7811 ;
  assign n7813 = n3158 ^ n2663 ^ 1'b0 ;
  assign n7814 = n3396 & n3433 ;
  assign n7815 = n7814 ^ n2187 ^ 1'b0 ;
  assign n7816 = n6683 | n7815 ;
  assign n7819 = n5440 ^ n3608 ^ n3185 ;
  assign n7817 = x70 | n1157 ;
  assign n7818 = n306 | n7817 ;
  assign n7820 = n7819 ^ n7818 ^ n1450 ;
  assign n7822 = n306 | n5113 ;
  assign n7823 = n7822 ^ n3143 ^ 1'b0 ;
  assign n7824 = n7823 ^ n2945 ^ 1'b0 ;
  assign n7821 = ~n664 & n3480 ;
  assign n7825 = n7824 ^ n7821 ^ 1'b0 ;
  assign n7826 = ~n4297 & n5941 ;
  assign n7827 = n7826 ^ n3021 ^ 1'b0 ;
  assign n7828 = ~n7769 & n7827 ;
  assign n7829 = n7079 ^ n4253 ^ 1'b0 ;
  assign n7830 = ~n1880 & n5621 ;
  assign n7831 = n7830 ^ n3679 ^ 1'b0 ;
  assign n7832 = n4452 & ~n5734 ;
  assign n7833 = ~n2592 & n7832 ;
  assign n7834 = ( ~n6526 & n7831 ) | ( ~n6526 & n7833 ) | ( n7831 & n7833 ) ;
  assign n7835 = ( n651 & n7829 ) | ( n651 & n7834 ) | ( n7829 & n7834 ) ;
  assign n7836 = ~n2750 & n3244 ;
  assign n7837 = ( n3675 & ~n7019 ) | ( n3675 & n7836 ) | ( ~n7019 & n7836 ) ;
  assign n7838 = n4570 ^ n3625 ^ 1'b0 ;
  assign n7839 = n2209 & n7838 ;
  assign n7840 = ( n1907 & ~n3775 ) | ( n1907 & n6563 ) | ( ~n3775 & n6563 ) ;
  assign n7841 = n6395 ^ n5495 ^ n3089 ;
  assign n7842 = x74 | n518 ;
  assign n7843 = ~n4291 & n7842 ;
  assign n7844 = n2903 & n7843 ;
  assign n7845 = n3876 ^ n1418 ^ n539 ;
  assign n7846 = n7845 ^ n1162 ^ 1'b0 ;
  assign n7847 = n7844 | n7846 ;
  assign n7848 = ~n959 & n7847 ;
  assign n7849 = n134 & ~n650 ;
  assign n7850 = ~n739 & n7849 ;
  assign n7855 = n1244 & n3342 ;
  assign n7851 = n4985 & ~n5074 ;
  assign n7852 = n5784 & ~n7851 ;
  assign n7853 = n4185 & n7852 ;
  assign n7854 = n3387 | n7853 ;
  assign n7856 = n7855 ^ n7854 ^ 1'b0 ;
  assign n7857 = n7850 & ~n7856 ;
  assign n7858 = n4811 ^ n1234 ^ 1'b0 ;
  assign n7859 = n2658 ^ n1403 ^ 1'b0 ;
  assign n7860 = n726 & n778 ;
  assign n7861 = n7860 ^ n524 ^ 1'b0 ;
  assign n7862 = n1089 | n2426 ;
  assign n7863 = ( n174 & n3670 ) | ( n174 & n7862 ) | ( n3670 & n7862 ) ;
  assign n7864 = ( n3113 & n3916 ) | ( n3113 & n7863 ) | ( n3916 & n7863 ) ;
  assign n7865 = n7032 ^ n4550 ^ n3961 ;
  assign n7866 = n4675 ^ n3515 ^ 1'b0 ;
  assign n7867 = n6218 & n7866 ;
  assign n7868 = n4786 & n6133 ;
  assign n7869 = ~n3464 & n3485 ;
  assign n7870 = n7182 ^ n6514 ^ 1'b0 ;
  assign n7871 = n7869 | n7870 ;
  assign n7872 = ~n1430 & n1736 ;
  assign n7873 = n4165 & ~n4245 ;
  assign n7874 = n2880 & n4232 ;
  assign n7875 = n719 & ~n872 ;
  assign n7876 = ~n2180 & n7875 ;
  assign n7877 = n3025 & ~n7876 ;
  assign n7878 = ( n5392 & n7874 ) | ( n5392 & n7877 ) | ( n7874 & n7877 ) ;
  assign n7879 = n1326 | n1835 ;
  assign n7880 = n2804 & n7879 ;
  assign n7881 = n746 & n1197 ;
  assign n7882 = n7880 | n7881 ;
  assign n7883 = n5852 ^ n4962 ^ n4123 ;
  assign n7884 = n7883 ^ n2647 ^ 1'b0 ;
  assign n7885 = n3593 | n7884 ;
  assign n7886 = n1471 & n3468 ;
  assign n7887 = n7886 ^ n2291 ^ 1'b0 ;
  assign n7888 = ~n912 & n7887 ;
  assign n7889 = n597 & n1265 ;
  assign n7890 = n7889 ^ n1109 ^ 1'b0 ;
  assign n7891 = n7890 ^ n4408 ^ 1'b0 ;
  assign n7892 = ~n2851 & n5774 ;
  assign n7893 = n3402 & n7892 ;
  assign n7894 = ( ~n2401 & n3189 ) | ( ~n2401 & n4127 ) | ( n3189 & n4127 ) ;
  assign n7895 = ~n7893 & n7894 ;
  assign n7896 = n7895 ^ n4716 ^ 1'b0 ;
  assign n7897 = n341 & ~n2438 ;
  assign n7904 = n1639 | n6337 ;
  assign n7901 = n5307 ^ n2105 ^ 1'b0 ;
  assign n7902 = ~n1605 & n7901 ;
  assign n7903 = n3691 & n7902 ;
  assign n7905 = n7904 ^ n7903 ^ 1'b0 ;
  assign n7906 = n1407 & ~n6625 ;
  assign n7907 = n2268 & ~n7906 ;
  assign n7908 = ~n7905 & n7907 ;
  assign n7898 = n4775 ^ n3958 ^ 1'b0 ;
  assign n7899 = n359 | n7898 ;
  assign n7900 = n7899 ^ n3535 ^ 1'b0 ;
  assign n7909 = n7908 ^ n7900 ^ 1'b0 ;
  assign n7910 = ~n740 & n3068 ;
  assign n7911 = n7910 ^ x104 ^ 1'b0 ;
  assign n7912 = n1534 & ~n6687 ;
  assign n7913 = n7328 & n7912 ;
  assign n7918 = n3857 ^ n982 ^ n532 ;
  assign n7919 = n7789 & n7918 ;
  assign n7920 = n7919 ^ n4379 ^ 1'b0 ;
  assign n7921 = n7920 ^ n6283 ^ 1'b0 ;
  assign n7914 = n3472 ^ n507 ^ 1'b0 ;
  assign n7915 = n2697 & n7914 ;
  assign n7916 = ( n421 & n4191 ) | ( n421 & n7915 ) | ( n4191 & n7915 ) ;
  assign n7917 = n2456 & n7916 ;
  assign n7922 = n7921 ^ n7917 ^ 1'b0 ;
  assign n7923 = x58 & ~n5882 ;
  assign n7924 = n2999 & n7923 ;
  assign n7925 = n7924 ^ n398 ^ 1'b0 ;
  assign n7926 = ~n4285 & n5611 ;
  assign n7927 = ~n7925 & n7926 ;
  assign n7929 = n3872 ^ n758 ^ 1'b0 ;
  assign n7930 = n159 | n7929 ;
  assign n7928 = n1655 | n5687 ;
  assign n7931 = n7930 ^ n7928 ^ n642 ;
  assign n7932 = n3114 & n4325 ;
  assign n7933 = n7931 & n7932 ;
  assign n7934 = ( n3827 & n4932 ) | ( n3827 & ~n6018 ) | ( n4932 & ~n6018 ) ;
  assign n7935 = n571 & ~n4783 ;
  assign n7939 = ~n395 & n711 ;
  assign n7940 = n5076 & ~n7939 ;
  assign n7941 = n7940 ^ n6259 ^ 1'b0 ;
  assign n7936 = ~n1436 & n5183 ;
  assign n7937 = n6122 & ~n7936 ;
  assign n7938 = ~n994 & n7937 ;
  assign n7942 = n7941 ^ n7938 ^ 1'b0 ;
  assign n7943 = n1175 & ~n7942 ;
  assign n7944 = ~n1644 & n6319 ;
  assign n7945 = ~n2014 & n2592 ;
  assign n7946 = n7945 ^ n4919 ^ n4817 ;
  assign n7947 = ~n4641 & n7113 ;
  assign n7948 = n4400 ^ n1440 ^ 1'b0 ;
  assign n7949 = n6374 | n7948 ;
  assign n7950 = n5523 & ~n7949 ;
  assign n7951 = n7950 ^ n7569 ^ 1'b0 ;
  assign n7952 = n3450 & ~n5092 ;
  assign n7953 = n3906 & n7952 ;
  assign n7954 = n7953 ^ n4022 ^ n3528 ;
  assign n7955 = n6829 ^ n1283 ^ 1'b0 ;
  assign n7956 = n1191 | n7955 ;
  assign n7957 = n7956 ^ n2839 ^ 1'b0 ;
  assign n7958 = ~n1600 & n2490 ;
  assign n7959 = x12 | n4739 ;
  assign n7960 = ~n1120 & n1342 ;
  assign n7961 = n4364 | n7960 ;
  assign n7962 = n7959 | n7961 ;
  assign n7963 = x38 | n6578 ;
  assign n7964 = n5944 ^ n5714 ^ 1'b0 ;
  assign n7966 = n1339 | n3000 ;
  assign n7967 = n7966 ^ n4826 ^ 1'b0 ;
  assign n7965 = x124 & n2500 ;
  assign n7968 = n7967 ^ n7965 ^ 1'b0 ;
  assign n7969 = n7083 ^ n4912 ^ 1'b0 ;
  assign n7970 = ( n3755 & n5338 ) | ( n3755 & n5871 ) | ( n5338 & n5871 ) ;
  assign n7971 = n1405 & ~n3036 ;
  assign n7972 = n7970 & ~n7971 ;
  assign n7973 = n5580 & n7972 ;
  assign n7974 = n2632 ^ n350 ^ 1'b0 ;
  assign n7975 = ~n3607 & n6523 ;
  assign n7976 = n7975 ^ n1829 ^ 1'b0 ;
  assign n7977 = n4202 ^ n671 ^ 1'b0 ;
  assign n7978 = n1002 | n7977 ;
  assign n7979 = n5878 ^ n1601 ^ 1'b0 ;
  assign n7980 = n7979 ^ n2744 ^ 1'b0 ;
  assign n7981 = n7978 & n7980 ;
  assign n7982 = n7976 & n7981 ;
  assign n7983 = ( ~n6692 & n7974 ) | ( ~n6692 & n7982 ) | ( n7974 & n7982 ) ;
  assign n7984 = x3 | n1608 ;
  assign n7985 = n4526 | n7984 ;
  assign n7986 = n2403 & ~n7985 ;
  assign n7987 = n605 & n3999 ;
  assign n7988 = n1940 ^ x14 ^ 1'b0 ;
  assign n7989 = ( ~n2119 & n4247 ) | ( ~n2119 & n7988 ) | ( n4247 & n7988 ) ;
  assign n7990 = n5353 ^ n4907 ^ x79 ;
  assign n7991 = n3986 | n6002 ;
  assign n7992 = ~n161 & n1953 ;
  assign n7993 = n3033 ^ n2184 ^ 1'b0 ;
  assign n7994 = ~n493 & n567 ;
  assign n7995 = ( ~n3457 & n6934 ) | ( ~n3457 & n7994 ) | ( n6934 & n7994 ) ;
  assign n7996 = n2365 ^ n696 ^ 1'b0 ;
  assign n7997 = n886 & ~n7996 ;
  assign n7998 = n2966 & n7997 ;
  assign n7999 = n7998 ^ n508 ^ 1'b0 ;
  assign n8000 = ~n6665 & n7999 ;
  assign n8001 = n8000 ^ n5037 ^ 1'b0 ;
  assign n8002 = n3931 ^ n3396 ^ 1'b0 ;
  assign n8003 = n8002 ^ x3 ^ 1'b0 ;
  assign n8004 = n2859 & n8003 ;
  assign n8005 = x58 | n1987 ;
  assign n8006 = n3643 & ~n6341 ;
  assign n8007 = n5432 & ~n7251 ;
  assign n8008 = n8006 | n8007 ;
  assign n8009 = ~n738 & n2164 ;
  assign n8010 = n2928 & n3216 ;
  assign n8011 = n2882 & n8010 ;
  assign n8012 = n1962 & ~n3290 ;
  assign n8013 = n8011 & n8012 ;
  assign n8014 = n2092 | n8013 ;
  assign n8015 = n3006 | n8014 ;
  assign n8019 = n2791 ^ n2703 ^ 1'b0 ;
  assign n8020 = n2711 & n8019 ;
  assign n8016 = n947 & ~n1155 ;
  assign n8017 = n8016 ^ n177 ^ 1'b0 ;
  assign n8018 = ~n3203 & n8017 ;
  assign n8021 = n8020 ^ n8018 ^ 1'b0 ;
  assign n8022 = n702 & n769 ;
  assign n8023 = n615 | n8022 ;
  assign n8024 = n8023 ^ n4189 ^ 1'b0 ;
  assign n8025 = n3931 ^ n875 ^ 1'b0 ;
  assign n8026 = n575 & n8025 ;
  assign n8027 = ~n3340 & n8026 ;
  assign n8028 = ~n8024 & n8027 ;
  assign n8029 = n8021 & ~n8028 ;
  assign n8030 = n2836 & ~n3814 ;
  assign n8034 = n7546 ^ n4627 ^ 1'b0 ;
  assign n8035 = ~n363 & n8034 ;
  assign n8031 = n1027 | n3053 ;
  assign n8032 = n8031 ^ n856 ^ 1'b0 ;
  assign n8033 = n6176 & ~n8032 ;
  assign n8036 = n8035 ^ n8033 ^ 1'b0 ;
  assign n8037 = n8036 ^ n1500 ^ 1'b0 ;
  assign n8038 = n4188 & n8037 ;
  assign n8039 = n6823 ^ n1652 ^ 1'b0 ;
  assign n8040 = ~n2933 & n8039 ;
  assign n8041 = ~n2988 & n7887 ;
  assign n8042 = n1360 & n8041 ;
  assign n8043 = n1561 & ~n8042 ;
  assign n8044 = n8043 ^ n1505 ^ 1'b0 ;
  assign n8045 = n6686 ^ n4358 ^ 1'b0 ;
  assign n8046 = n8044 & n8045 ;
  assign n8047 = n1952 ^ n1860 ^ 1'b0 ;
  assign n8048 = ~n4070 & n8047 ;
  assign n8049 = n8048 ^ n2166 ^ 1'b0 ;
  assign n8053 = n4365 ^ n3169 ^ 1'b0 ;
  assign n8050 = x42 & n1291 ;
  assign n8051 = ~n581 & n777 ;
  assign n8052 = ~n8050 & n8051 ;
  assign n8054 = n8053 ^ n8052 ^ n7452 ;
  assign n8055 = ( n745 & ~n8049 ) | ( n745 & n8054 ) | ( ~n8049 & n8054 ) ;
  assign n8056 = n4985 | n6148 ;
  assign n8057 = n299 & n5480 ;
  assign n8058 = n8057 ^ n5818 ^ 1'b0 ;
  assign n8059 = ( x55 & ~n1540 ) | ( x55 & n8058 ) | ( ~n1540 & n8058 ) ;
  assign n8060 = n1677 ^ n742 ^ 1'b0 ;
  assign n8061 = ~n8059 & n8060 ;
  assign n8062 = n2826 ^ n1930 ^ 1'b0 ;
  assign n8063 = n1476 & ~n7223 ;
  assign n8064 = n5397 ^ n3729 ^ 1'b0 ;
  assign n8066 = n134 & ~n3741 ;
  assign n8067 = n8066 ^ n6524 ^ 1'b0 ;
  assign n8068 = n5013 | n5024 ;
  assign n8069 = n8067 & n8068 ;
  assign n8065 = n3064 | n4222 ;
  assign n8070 = n8069 ^ n8065 ^ 1'b0 ;
  assign n8071 = ~n8064 & n8070 ;
  assign n8075 = n3291 ^ n2690 ^ 1'b0 ;
  assign n8072 = n5959 & ~n7408 ;
  assign n8073 = ~n812 & n8072 ;
  assign n8074 = n8073 ^ n3950 ^ n2747 ;
  assign n8076 = n8075 ^ n8074 ^ 1'b0 ;
  assign n8077 = n2414 | n8076 ;
  assign n8078 = n7085 | n8077 ;
  assign n8079 = ~n2371 & n5407 ;
  assign n8081 = n4537 ^ n4062 ^ n3967 ;
  assign n8080 = ( n346 & ~n1251 ) | ( n346 & n1920 ) | ( ~n1251 & n1920 ) ;
  assign n8082 = n8081 ^ n8080 ^ n7887 ;
  assign n8083 = n1568 & n6232 ;
  assign n8084 = n1607 & n1809 ;
  assign n8085 = n8084 ^ n4964 ^ 1'b0 ;
  assign n8086 = n2805 & ~n8085 ;
  assign n8087 = n6067 ^ n1316 ^ 1'b0 ;
  assign n8088 = x51 | n342 ;
  assign n8089 = n590 & ~n8088 ;
  assign n8090 = n3289 | n8089 ;
  assign n8091 = n5608 & n8090 ;
  assign n8092 = ~n486 & n4827 ;
  assign n8093 = n2973 & n8092 ;
  assign n8094 = n247 | n4845 ;
  assign n8095 = n142 | n1784 ;
  assign n8096 = n8095 ^ n1784 ^ 1'b0 ;
  assign n8097 = n8096 ^ n4968 ^ n1771 ;
  assign n8098 = n185 & n1239 ;
  assign n8099 = n1991 & n8098 ;
  assign n8100 = n8099 ^ n5520 ^ n3684 ;
  assign n8101 = n5561 ^ n4457 ^ 1'b0 ;
  assign n8102 = ~n6534 & n8101 ;
  assign n8103 = ( ~n1475 & n3411 ) | ( ~n1475 & n8102 ) | ( n3411 & n8102 ) ;
  assign n8105 = n1892 ^ n538 ^ 1'b0 ;
  assign n8106 = n3221 & n8105 ;
  assign n8104 = n7632 ^ n3847 ^ n1135 ;
  assign n8107 = n8106 ^ n8104 ^ 1'b0 ;
  assign n8108 = ( n3265 & n3812 ) | ( n3265 & ~n5648 ) | ( n3812 & ~n5648 ) ;
  assign n8109 = ~n1576 & n8108 ;
  assign n8110 = n8109 ^ n7956 ^ 1'b0 ;
  assign n8111 = n1779 & ~n4648 ;
  assign n8112 = n4966 & n8111 ;
  assign n8113 = ( n509 & n8110 ) | ( n509 & n8112 ) | ( n8110 & n8112 ) ;
  assign n8114 = n393 & ~n521 ;
  assign n8115 = x21 & n4150 ;
  assign n8116 = ~n1637 & n7493 ;
  assign n8117 = n5415 ^ n2517 ^ 1'b0 ;
  assign n8118 = ~n1743 & n8117 ;
  assign n8119 = ~n536 & n1263 ;
  assign n8120 = n8119 ^ n4627 ^ 1'b0 ;
  assign n8121 = n3838 & ~n7260 ;
  assign n8122 = n2924 ^ n2051 ^ 1'b0 ;
  assign n8123 = ( ~n4570 & n5699 ) | ( ~n4570 & n8122 ) | ( n5699 & n8122 ) ;
  assign n8124 = ~n2051 & n5147 ;
  assign n8125 = n4705 ^ n1264 ^ 1'b0 ;
  assign n8126 = n8124 & n8125 ;
  assign n8127 = ( n651 & n4339 ) | ( n651 & ~n6131 ) | ( n4339 & ~n6131 ) ;
  assign n8128 = n7616 ^ n5936 ^ n905 ;
  assign n8129 = n4833 ^ n3433 ^ n2695 ;
  assign n8130 = ( n1927 & ~n5074 ) | ( n1927 & n8129 ) | ( ~n5074 & n8129 ) ;
  assign n8131 = n5516 ^ n485 ^ 1'b0 ;
  assign n8132 = n8130 & ~n8131 ;
  assign n8133 = n6671 ^ n706 ^ 1'b0 ;
  assign n8134 = n8132 & n8133 ;
  assign n8135 = n5602 ^ n3785 ^ 1'b0 ;
  assign n8136 = n5101 ^ n2189 ^ 1'b0 ;
  assign n8137 = n5839 ^ n3737 ^ 1'b0 ;
  assign n8138 = n6138 ^ n5425 ^ n288 ;
  assign n8139 = n8138 ^ n544 ^ 1'b0 ;
  assign n8140 = ~n5002 & n8139 ;
  assign n8141 = n7674 ^ n4402 ^ 1'b0 ;
  assign n8143 = n4946 ^ n4669 ^ n4147 ;
  assign n8142 = n3524 ^ n342 ^ 1'b0 ;
  assign n8144 = n8143 ^ n8142 ^ n4479 ;
  assign n8145 = n8144 ^ n1374 ^ 1'b0 ;
  assign n8146 = n7911 ^ n3587 ^ 1'b0 ;
  assign n8147 = ( n1992 & n2051 ) | ( n1992 & ~n6420 ) | ( n2051 & ~n6420 ) ;
  assign n8148 = n3492 ^ n2190 ^ n1895 ;
  assign n8149 = n8148 ^ n683 ^ 1'b0 ;
  assign n8150 = n638 | n8149 ;
  assign n8151 = n8150 ^ n3472 ^ 1'b0 ;
  assign n8152 = n1041 | n8151 ;
  assign n8153 = n612 & ~n8152 ;
  assign n8154 = ~n3565 & n8153 ;
  assign n8155 = n1134 & ~n6432 ;
  assign n8156 = n8155 ^ n4745 ^ 1'b0 ;
  assign n8157 = ( n1470 & n3887 ) | ( n1470 & n4209 ) | ( n3887 & n4209 ) ;
  assign n8158 = n1272 | n8157 ;
  assign n8159 = n8158 ^ n4853 ^ 1'b0 ;
  assign n8160 = n3746 & n8159 ;
  assign n8161 = n8156 & n8160 ;
  assign n8162 = n6848 & n8161 ;
  assign n8163 = ~n4037 & n4768 ;
  assign n8164 = n8163 ^ n3596 ^ x13 ;
  assign n8165 = n8164 ^ n1940 ^ 1'b0 ;
  assign n8166 = n3691 & ~n4942 ;
  assign n8167 = n4714 ^ n3437 ^ 1'b0 ;
  assign n8168 = n2589 & n6251 ;
  assign n8169 = ~n4330 & n8168 ;
  assign n8170 = n3583 & ~n8169 ;
  assign n8171 = n5353 & ~n5573 ;
  assign n8172 = n3076 & n7347 ;
  assign n8179 = n1624 & ~n1927 ;
  assign n8177 = n2074 ^ n905 ^ 1'b0 ;
  assign n8173 = ~x95 & x103 ;
  assign n8174 = n8173 ^ n2172 ^ 1'b0 ;
  assign n8175 = n309 & ~n8174 ;
  assign n8176 = ~n2791 & n8175 ;
  assign n8178 = n8177 ^ n8176 ^ 1'b0 ;
  assign n8180 = n8179 ^ n8178 ^ 1'b0 ;
  assign n8181 = n2366 ^ n1512 ^ n1462 ;
  assign n8182 = n3627 | n8181 ;
  assign n8183 = ~n2736 & n7869 ;
  assign n8184 = n1193 | n1973 ;
  assign n8185 = n558 & ~n8184 ;
  assign n8186 = n7415 | n8185 ;
  assign n8187 = n7222 & ~n8186 ;
  assign n8188 = x55 & ~n8187 ;
  assign n8189 = n8188 ^ n4071 ^ 1'b0 ;
  assign n8192 = n7749 ^ n367 ^ 1'b0 ;
  assign n8190 = n806 & n7905 ;
  assign n8191 = n8190 ^ n6255 ^ n4487 ;
  assign n8193 = n8192 ^ n8191 ^ 1'b0 ;
  assign n8194 = n1944 & n7854 ;
  assign n8195 = n8194 ^ n5458 ^ 1'b0 ;
  assign n8196 = n4109 & ~n4393 ;
  assign n8197 = ~n819 & n8196 ;
  assign n8198 = n5079 ^ n404 ^ 1'b0 ;
  assign n8199 = n6821 | n8198 ;
  assign n8200 = ~n217 & n4199 ;
  assign n8201 = n3545 | n6610 ;
  assign n8202 = n2198 | n8201 ;
  assign n8203 = n4963 & n8202 ;
  assign n8204 = n6512 & n8203 ;
  assign n8205 = n3901 ^ n2096 ^ 1'b0 ;
  assign n8206 = x9 & ~n8205 ;
  assign n8207 = ~n2295 & n5778 ;
  assign n8208 = n1494 & ~n8207 ;
  assign n8209 = ~n1234 & n2596 ;
  assign n8210 = n8209 ^ n4631 ^ 1'b0 ;
  assign n8211 = n4498 & ~n6374 ;
  assign n8212 = n8211 ^ n1746 ^ 1'b0 ;
  assign n8213 = n8212 ^ n5890 ^ 1'b0 ;
  assign n8214 = ~n3310 & n3701 ;
  assign n8215 = n337 & n1017 ;
  assign n8216 = n8215 ^ n867 ^ 1'b0 ;
  assign n8217 = n8216 ^ n2932 ^ n2775 ;
  assign n8218 = ~n1654 & n8217 ;
  assign n8219 = n8218 ^ n6570 ^ 1'b0 ;
  assign n8220 = ~n6382 & n8219 ;
  assign n8221 = n4634 ^ n1330 ^ 1'b0 ;
  assign n8222 = n7918 & ~n8221 ;
  assign n8223 = ( n457 & n2534 ) | ( n457 & n6402 ) | ( n2534 & n6402 ) ;
  assign n8224 = x64 ^ x14 ^ 1'b0 ;
  assign n8225 = n1626 & n8224 ;
  assign n8226 = n8225 ^ n4410 ^ 1'b0 ;
  assign n8227 = ( ~n5435 & n8223 ) | ( ~n5435 & n8226 ) | ( n8223 & n8226 ) ;
  assign n8228 = n8166 ^ n494 ^ 1'b0 ;
  assign n8229 = n2208 & n8228 ;
  assign n8230 = n3058 ^ n2590 ^ n912 ;
  assign n8231 = n748 & n8230 ;
  assign n8232 = ( n134 & ~n3795 ) | ( n134 & n8231 ) | ( ~n3795 & n8231 ) ;
  assign n8233 = n1946 ^ n648 ^ 1'b0 ;
  assign n8234 = n374 & ~n393 ;
  assign n8235 = ~n374 & n8234 ;
  assign n8236 = n1547 | n3124 ;
  assign n8237 = n3124 & ~n8236 ;
  assign n8238 = n2964 | n8237 ;
  assign n8239 = n2964 & ~n8238 ;
  assign n8240 = n2062 | n8239 ;
  assign n8241 = n2062 & ~n8240 ;
  assign n8242 = n1422 & ~n8241 ;
  assign n8243 = n8235 & n8242 ;
  assign n8244 = n8243 ^ n2189 ^ 1'b0 ;
  assign n8245 = ~n8233 & n8244 ;
  assign n8246 = n1392 | n4110 ;
  assign n8247 = n8246 ^ n2903 ^ 1'b0 ;
  assign n8248 = ~n2673 & n8247 ;
  assign n8249 = n2024 | n5967 ;
  assign n8250 = n3723 | n8249 ;
  assign n8251 = n301 | n2122 ;
  assign n8252 = n8251 ^ n1547 ^ 1'b0 ;
  assign n8253 = n1506 | n3542 ;
  assign n8254 = n8253 ^ n7181 ^ n2201 ;
  assign n8255 = n1506 & n8254 ;
  assign n8256 = n8255 ^ n4725 ^ 1'b0 ;
  assign n8259 = n4898 ^ n2271 ^ n954 ;
  assign n8257 = n4636 ^ n3879 ^ n466 ;
  assign n8258 = n8257 ^ n3521 ^ 1'b0 ;
  assign n8260 = n8259 ^ n8258 ^ n5840 ;
  assign n8261 = ( ~n1085 & n1953 ) | ( ~n1085 & n2315 ) | ( n1953 & n2315 ) ;
  assign n8262 = n8261 ^ n3073 ^ 1'b0 ;
  assign n8263 = n3861 & n5857 ;
  assign n8264 = n8263 ^ n7430 ^ 1'b0 ;
  assign n8265 = x8 & n667 ;
  assign n8266 = n4054 ^ n615 ^ 1'b0 ;
  assign n8267 = n8265 & n8266 ;
  assign n8268 = n8267 ^ n7048 ^ 1'b0 ;
  assign n8269 = n5069 | n8268 ;
  assign n8270 = n2203 & n5034 ;
  assign n8271 = ~n2444 & n8270 ;
  assign n8272 = n8271 ^ n2322 ^ 1'b0 ;
  assign n8273 = n2546 ^ n1571 ^ n1450 ;
  assign n8274 = ~n2780 & n5248 ;
  assign n8275 = n8273 & n8274 ;
  assign n8276 = n7317 ^ n1248 ^ 1'b0 ;
  assign n8277 = n1242 & n8276 ;
  assign n8278 = n374 & ~n4111 ;
  assign n8279 = n1123 ^ n639 ^ 1'b0 ;
  assign n8280 = n8279 ^ n1217 ^ 1'b0 ;
  assign n8281 = n3865 | n8280 ;
  assign n8282 = n8281 ^ n892 ^ 1'b0 ;
  assign n8283 = n4948 ^ n657 ^ 1'b0 ;
  assign n8284 = n665 | n8283 ;
  assign n8285 = n8284 ^ n193 ^ 1'b0 ;
  assign n8286 = ~n7819 & n8285 ;
  assign n8287 = n3999 ^ x126 ^ 1'b0 ;
  assign n8288 = n8287 ^ n5382 ^ n3355 ;
  assign n8289 = n482 & ~n7653 ;
  assign n8290 = n4531 ^ n2342 ^ 1'b0 ;
  assign n8291 = ~n8289 & n8290 ;
  assign n8292 = n1671 & n8291 ;
  assign n8293 = n8292 ^ n7651 ^ 1'b0 ;
  assign n8295 = n2167 ^ n881 ^ 1'b0 ;
  assign n8294 = ( n4359 & n4732 ) | ( n4359 & ~n6888 ) | ( n4732 & ~n6888 ) ;
  assign n8296 = n8295 ^ n8294 ^ n7605 ;
  assign n8300 = n4091 ^ n283 ^ 1'b0 ;
  assign n8301 = n8300 ^ n3315 ^ n2456 ;
  assign n8298 = n6654 ^ n5761 ^ 1'b0 ;
  assign n8297 = n4400 & n6386 ;
  assign n8299 = n8298 ^ n8297 ^ 1'b0 ;
  assign n8302 = n8301 ^ n8299 ^ 1'b0 ;
  assign n8303 = ~n1658 & n4346 ;
  assign n8304 = n6882 ^ n5262 ^ 1'b0 ;
  assign n8305 = n6201 | n8304 ;
  assign n8306 = n4946 ^ n2605 ^ 1'b0 ;
  assign n8307 = n2760 & ~n4247 ;
  assign n8308 = n456 & n8307 ;
  assign n8309 = n992 & ~n6104 ;
  assign n8310 = n920 & n8309 ;
  assign n8311 = n2296 | n8310 ;
  assign n8312 = n3836 | n8311 ;
  assign n8313 = n5600 | n8312 ;
  assign n8314 = n8313 ^ n442 ^ 1'b0 ;
  assign n8315 = n8308 | n8314 ;
  assign n8316 = n2272 ^ n470 ^ 1'b0 ;
  assign n8317 = n2113 | n8316 ;
  assign n8318 = ~n206 & n5608 ;
  assign n8319 = n8318 ^ n2930 ^ 1'b0 ;
  assign n8320 = ( n2186 & n3103 ) | ( n2186 & n8319 ) | ( n3103 & n8319 ) ;
  assign n8321 = n8317 & n8320 ;
  assign n8322 = ~n7925 & n8321 ;
  assign n8323 = n3791 & n6093 ;
  assign n8324 = n8323 ^ n5490 ^ 1'b0 ;
  assign n8325 = n1711 ^ n1283 ^ 1'b0 ;
  assign n8326 = n6464 & n8325 ;
  assign n8327 = n2167 & n5356 ;
  assign n8328 = n8327 ^ n2634 ^ 1'b0 ;
  assign n8329 = n1985 & n6908 ;
  assign n8330 = n7408 ^ n7111 ^ n368 ;
  assign n8331 = n1775 | n7205 ;
  assign n8332 = ( n7504 & n8330 ) | ( n7504 & ~n8331 ) | ( n8330 & ~n8331 ) ;
  assign n8333 = ~n5915 & n7550 ;
  assign n8334 = ~n1998 & n8333 ;
  assign n8335 = n1585 ^ x54 ^ 1'b0 ;
  assign n8336 = ~n1420 & n8335 ;
  assign n8337 = n922 | n8336 ;
  assign n8338 = n8337 ^ n3169 ^ 1'b0 ;
  assign n8339 = n8338 ^ n4765 ^ 1'b0 ;
  assign n8340 = ~n8334 & n8339 ;
  assign n8341 = n2345 ^ n821 ^ n452 ;
  assign n8342 = n8341 ^ n5573 ^ n750 ;
  assign n8343 = n3958 ^ n3752 ^ x11 ;
  assign n8344 = ( x48 & n828 ) | ( x48 & ~n8343 ) | ( n828 & ~n8343 ) ;
  assign n8345 = n2266 & ~n5551 ;
  assign n8346 = n1481 & ~n5278 ;
  assign n8347 = n5705 & n8346 ;
  assign n8348 = n3276 & ~n8347 ;
  assign n8349 = n8348 ^ n1689 ^ 1'b0 ;
  assign n8350 = n5378 ^ n3882 ^ 1'b0 ;
  assign n8351 = n4456 & n8350 ;
  assign n8352 = n961 | n1634 ;
  assign n8353 = n7210 & ~n8352 ;
  assign n8354 = n2787 | n8353 ;
  assign n8355 = n3033 | n6455 ;
  assign n8356 = n8355 ^ n320 ^ 1'b0 ;
  assign n8357 = n2750 ^ n2670 ^ 1'b0 ;
  assign n8358 = n8357 ^ n2472 ^ 1'b0 ;
  assign n8359 = ~n2627 & n6936 ;
  assign n8360 = n8359 ^ n3614 ^ 1'b0 ;
  assign n8361 = n746 & n2756 ;
  assign n8362 = n3929 & n8361 ;
  assign n8363 = n606 & n8362 ;
  assign n8364 = n8360 & ~n8363 ;
  assign n8365 = n8358 & n8364 ;
  assign n8366 = n2806 | n8365 ;
  assign n8367 = n1915 & ~n2527 ;
  assign n8368 = n8140 ^ n2087 ^ 1'b0 ;
  assign n8369 = ( n1207 & n2796 ) | ( n1207 & n3619 ) | ( n2796 & n3619 ) ;
  assign n8371 = n837 ^ n248 ^ 1'b0 ;
  assign n8370 = n3113 | n4701 ;
  assign n8372 = n8371 ^ n8370 ^ 1'b0 ;
  assign n8373 = n5523 & n8372 ;
  assign n8374 = n8373 ^ n5061 ^ 1'b0 ;
  assign n8375 = n3590 ^ n1062 ^ 1'b0 ;
  assign n8376 = ~n1634 & n8375 ;
  assign n8377 = n535 | n8376 ;
  assign n8378 = n8377 ^ n3694 ^ n3034 ;
  assign n8379 = n3657 & ~n8378 ;
  assign n8380 = ~n3727 & n8379 ;
  assign n8381 = n4042 ^ n1471 ^ 1'b0 ;
  assign n8382 = n6353 ^ n544 ^ 1'b0 ;
  assign n8383 = n7549 ^ n4000 ^ 1'b0 ;
  assign n8384 = ~n2863 & n8383 ;
  assign n8385 = n1907 & n2326 ;
  assign n8386 = n5168 ^ n4751 ^ 1'b0 ;
  assign n8387 = n6586 & ~n8386 ;
  assign n8389 = n1405 & n4104 ;
  assign n8390 = n3437 ^ n280 ^ 1'b0 ;
  assign n8391 = n4703 & n8390 ;
  assign n8392 = ~n8389 & n8391 ;
  assign n8388 = ~n3015 & n4869 ;
  assign n8393 = n8392 ^ n8388 ^ 1'b0 ;
  assign n8394 = ~n443 & n1291 ;
  assign n8395 = n8394 ^ n5092 ^ 1'b0 ;
  assign n8396 = n3158 | n3698 ;
  assign n8397 = n8396 ^ x110 ^ 1'b0 ;
  assign n8398 = n3265 & n8397 ;
  assign n8399 = ~n8395 & n8398 ;
  assign n8400 = n2209 & ~n3089 ;
  assign n8401 = n1954 & n8400 ;
  assign n8402 = x27 & ~n7348 ;
  assign n8403 = n8401 & n8402 ;
  assign n8404 = n8403 ^ n3872 ^ 1'b0 ;
  assign n8405 = n1511 & n1708 ;
  assign n8406 = ~n2841 & n6070 ;
  assign n8407 = ~n8405 & n8406 ;
  assign n8408 = n7581 & n8407 ;
  assign n8409 = n8408 ^ n4216 ^ 1'b0 ;
  assign n8410 = n5336 & ~n8409 ;
  assign n8411 = ~n2165 & n2721 ;
  assign n8412 = n8411 ^ n1224 ^ 1'b0 ;
  assign n8413 = n8412 ^ n2485 ^ 1'b0 ;
  assign n8414 = n8278 & n8413 ;
  assign n8415 = ~n8410 & n8414 ;
  assign n8419 = n3312 ^ n3026 ^ 1'b0 ;
  assign n8416 = n2602 ^ n1368 ^ 1'b0 ;
  assign n8417 = ~n2508 & n8416 ;
  assign n8418 = n2018 & n8417 ;
  assign n8420 = n8419 ^ n8418 ^ 1'b0 ;
  assign n8421 = n6026 & n8420 ;
  assign n8422 = n3256 & n8421 ;
  assign n8423 = n2747 & ~n8422 ;
  assign n8424 = n8423 ^ n7796 ^ 1'b0 ;
  assign n8425 = ~n1008 & n1465 ;
  assign n8426 = n8425 ^ n5783 ^ n509 ;
  assign n8427 = n2003 ^ n1314 ^ 1'b0 ;
  assign n8428 = n8427 ^ n2824 ^ x126 ;
  assign n8429 = n8081 ^ n3221 ^ 1'b0 ;
  assign n8431 = ( n319 & n2238 ) | ( n319 & n3358 ) | ( n2238 & n3358 ) ;
  assign n8430 = n1761 | n2765 ;
  assign n8432 = n8431 ^ n8430 ^ 1'b0 ;
  assign n8433 = ~n969 & n8432 ;
  assign n8434 = n8433 ^ n1610 ^ 1'b0 ;
  assign n8435 = ~n4468 & n6047 ;
  assign n8436 = n8435 ^ n7217 ^ 1'b0 ;
  assign n8437 = n2028 | n8058 ;
  assign n8438 = ~n2812 & n8437 ;
  assign n8439 = n7944 | n8438 ;
  assign n8440 = n8439 ^ n1061 ^ 1'b0 ;
  assign n8441 = n8440 ^ n2151 ^ n285 ;
  assign n8442 = ~n1111 & n1434 ;
  assign n8443 = n8442 ^ n399 ^ 1'b0 ;
  assign n8446 = n6631 & n6821 ;
  assign n8447 = n8446 ^ n1720 ^ 1'b0 ;
  assign n8444 = n2645 & n7558 ;
  assign n8445 = n5027 & ~n8444 ;
  assign n8448 = n8447 ^ n8445 ^ 1'b0 ;
  assign n8449 = n8443 & n8448 ;
  assign n8450 = n683 & n6657 ;
  assign n8451 = n4180 | n8450 ;
  assign n8452 = n2221 | n8451 ;
  assign n8453 = n6934 ^ n2450 ^ 1'b0 ;
  assign n8454 = n3950 ^ n996 ^ 1'b0 ;
  assign n8457 = n865 | n6265 ;
  assign n8458 = n8457 ^ n3467 ^ 1'b0 ;
  assign n8455 = n7589 ^ x54 ^ 1'b0 ;
  assign n8456 = ~n2349 & n8455 ;
  assign n8459 = n8458 ^ n8456 ^ 1'b0 ;
  assign n8460 = n1687 & ~n3053 ;
  assign n8461 = n8460 ^ n3775 ^ 1'b0 ;
  assign n8462 = n4489 & ~n6187 ;
  assign n8463 = n8355 ^ n1703 ^ 1'b0 ;
  assign n8464 = n350 | n8463 ;
  assign n8465 = n1226 | n4734 ;
  assign n8466 = n8465 ^ n2038 ^ 1'b0 ;
  assign n8467 = n5785 & n8466 ;
  assign n8468 = ~n2675 & n3230 ;
  assign n8469 = n8468 ^ n1940 ^ 1'b0 ;
  assign n8470 = n7432 ^ n5783 ^ n461 ;
  assign n8471 = n8341 ^ n3297 ^ 1'b0 ;
  assign n8472 = n7242 ^ n2451 ^ 1'b0 ;
  assign n8473 = ~n4161 & n8472 ;
  assign n8474 = ~n2793 & n5126 ;
  assign n8475 = ~n7764 & n8474 ;
  assign n8476 = ~n8473 & n8475 ;
  assign n8477 = ~n2594 & n5603 ;
  assign n8478 = n8477 ^ n175 ^ 1'b0 ;
  assign n8479 = n1062 & n2165 ;
  assign n8480 = ~n6357 & n8479 ;
  assign n8481 = n5204 ^ n4165 ^ 1'b0 ;
  assign n8482 = n5492 ^ n4221 ^ 1'b0 ;
  assign n8483 = n4490 & n8482 ;
  assign n8484 = n8481 & n8483 ;
  assign n8485 = n6010 ^ n4471 ^ 1'b0 ;
  assign n8486 = n3906 | n8485 ;
  assign n8487 = n1795 | n2839 ;
  assign n8488 = ~n2670 & n8487 ;
  assign n8489 = n5475 ^ n5342 ^ 1'b0 ;
  assign n8490 = ~n8488 & n8489 ;
  assign n8491 = n1086 ^ n445 ^ 1'b0 ;
  assign n8492 = n8491 ^ n1205 ^ 1'b0 ;
  assign n8493 = n8492 ^ n6385 ^ n3943 ;
  assign n8494 = n1670 & n7528 ;
  assign n8495 = n8494 ^ n1482 ^ 1'b0 ;
  assign n8496 = ~n4979 & n8495 ;
  assign n8498 = n574 & ~n8150 ;
  assign n8497 = n5435 ^ n1408 ^ 1'b0 ;
  assign n8499 = n8498 ^ n8497 ^ 1'b0 ;
  assign n8500 = n2800 & ~n6597 ;
  assign n8501 = n1794 & n5059 ;
  assign n8502 = n5248 ^ n396 ^ 1'b0 ;
  assign n8503 = ( n729 & n8501 ) | ( n729 & ~n8502 ) | ( n8501 & ~n8502 ) ;
  assign n8504 = n1885 & n4449 ;
  assign n8505 = n3562 & ~n8502 ;
  assign n8506 = n978 | n6537 ;
  assign n8507 = n8506 ^ n6847 ^ 1'b0 ;
  assign n8508 = n593 & ~n7061 ;
  assign n8509 = n8508 ^ n2403 ^ 1'b0 ;
  assign n8510 = ~n4293 & n8509 ;
  assign n8511 = n909 ^ n277 ^ 1'b0 ;
  assign n8512 = n910 & n8511 ;
  assign n8513 = n1411 | n8512 ;
  assign n8514 = n8513 ^ n7358 ^ 1'b0 ;
  assign n8515 = n6663 | n8258 ;
  assign n8516 = n8415 ^ n1601 ^ 1'b0 ;
  assign n8518 = n6218 ^ n5473 ^ 1'b0 ;
  assign n8519 = ~n508 & n8518 ;
  assign n8517 = n2304 | n5724 ;
  assign n8520 = n8519 ^ n8517 ^ 1'b0 ;
  assign n8521 = n2951 & ~n8500 ;
  assign n8522 = ~n8520 & n8521 ;
  assign n8523 = n3021 ^ n2249 ^ 1'b0 ;
  assign n8524 = n4543 ^ n804 ^ 1'b0 ;
  assign n8525 = n8523 | n8524 ;
  assign n8526 = ~n5014 & n8525 ;
  assign n8527 = n8319 ^ n2178 ^ 1'b0 ;
  assign n8528 = ~n2350 & n8527 ;
  assign n8529 = n6631 ^ n1772 ^ 1'b0 ;
  assign n8530 = n2560 | n8529 ;
  assign n8531 = n944 | n8530 ;
  assign n8532 = n8531 ^ n6786 ^ n2106 ;
  assign n8533 = n8528 & n8532 ;
  assign n8534 = n8533 ^ n8017 ^ 1'b0 ;
  assign n8541 = n5018 ^ n593 ^ 1'b0 ;
  assign n8542 = n3792 & ~n8541 ;
  assign n8543 = n5310 & n8542 ;
  assign n8535 = n1425 | n2726 ;
  assign n8536 = n8535 ^ n2642 ^ 1'b0 ;
  assign n8537 = ~n5125 & n8536 ;
  assign n8538 = ( n190 & n1776 ) | ( n190 & n8537 ) | ( n1776 & n8537 ) ;
  assign n8539 = ~n1876 & n8538 ;
  assign n8540 = n1724 & n8539 ;
  assign n8544 = n8543 ^ n8540 ^ 1'b0 ;
  assign n8545 = n897 ^ n574 ^ 1'b0 ;
  assign n8546 = ( x32 & n5391 ) | ( x32 & n7057 ) | ( n5391 & n7057 ) ;
  assign n8547 = n2857 | n8546 ;
  assign n8548 = ( ~n5606 & n8545 ) | ( ~n5606 & n8547 ) | ( n8545 & n8547 ) ;
  assign n8549 = n3148 ^ n1486 ^ 1'b0 ;
  assign n8550 = ( n4376 & n5516 ) | ( n4376 & ~n8549 ) | ( n5516 & ~n8549 ) ;
  assign n8552 = n2501 ^ n424 ^ 1'b0 ;
  assign n8551 = ~n1081 & n7726 ;
  assign n8553 = n8552 ^ n8551 ^ 1'b0 ;
  assign n8554 = n461 & n6165 ;
  assign n8555 = n8554 ^ n654 ^ 1'b0 ;
  assign n8556 = ( n1974 & ~n4803 ) | ( n1974 & n8555 ) | ( ~n4803 & n8555 ) ;
  assign n8557 = n488 & ~n3584 ;
  assign n8558 = n8557 ^ n5947 ^ 1'b0 ;
  assign n8559 = n8317 ^ n5312 ^ 1'b0 ;
  assign n8560 = n6991 ^ n1907 ^ 1'b0 ;
  assign n8561 = n5783 ^ n1461 ^ 1'b0 ;
  assign n8562 = n7422 ^ n1726 ^ 1'b0 ;
  assign n8563 = n8562 ^ n3662 ^ 1'b0 ;
  assign n8565 = ~n2972 & n3844 ;
  assign n8564 = ~n3933 & n6582 ;
  assign n8566 = n8565 ^ n8564 ^ 1'b0 ;
  assign n8567 = n5810 ^ n174 ^ x13 ;
  assign n8568 = n8567 ^ n8289 ^ n182 ;
  assign n8569 = n4330 ^ n3647 ^ 1'b0 ;
  assign n8570 = n571 & n8569 ;
  assign n8571 = ~n651 & n1362 ;
  assign n8572 = ~n523 & n8571 ;
  assign n8573 = n3717 & n8572 ;
  assign n8574 = n6968 ^ x21 ^ 1'b0 ;
  assign n8575 = n1380 & n3497 ;
  assign n8576 = n625 & n8575 ;
  assign n8577 = n8576 ^ n1603 ^ 1'b0 ;
  assign n8578 = n4195 ^ n665 ^ 1'b0 ;
  assign n8579 = ~n2829 & n8578 ;
  assign n8580 = n4382 & n4640 ;
  assign n8581 = n8580 ^ n4662 ^ 1'b0 ;
  assign n8582 = ~n3419 & n5207 ;
  assign n8583 = n5249 | n8582 ;
  assign n8584 = n8583 ^ n2335 ^ 1'b0 ;
  assign n8585 = n1288 | n3742 ;
  assign n8586 = n8585 ^ n1251 ^ 1'b0 ;
  assign n8587 = n8586 ^ n3853 ^ n970 ;
  assign n8588 = n2280 & ~n8587 ;
  assign n8589 = n750 | n8588 ;
  assign n8590 = n8584 & ~n8589 ;
  assign n8591 = n1808 | n5397 ;
  assign n8592 = n2594 | n8591 ;
  assign n8593 = n500 | n6639 ;
  assign n8594 = n3091 | n8593 ;
  assign n8595 = n1722 ^ n625 ^ 1'b0 ;
  assign n8596 = n8594 & ~n8595 ;
  assign n8597 = n1820 & n5117 ;
  assign n8598 = n4575 ^ n852 ^ 1'b0 ;
  assign n8599 = ~n3812 & n3927 ;
  assign n8600 = n8599 ^ n215 ^ 1'b0 ;
  assign n8601 = ~n6874 & n7021 ;
  assign n8602 = n8601 ^ n6070 ^ 1'b0 ;
  assign n8603 = n3576 ^ n1944 ^ 1'b0 ;
  assign n8604 = n5395 & ~n8603 ;
  assign n8605 = n8604 ^ n532 ^ 1'b0 ;
  assign n8606 = n3399 & n3960 ;
  assign n8607 = n8605 & ~n8606 ;
  assign n8608 = ~n7192 & n8607 ;
  assign n8609 = n2886 | n8608 ;
  assign n8610 = ( n3074 & n5814 ) | ( n3074 & n8609 ) | ( n5814 & n8609 ) ;
  assign n8611 = n6570 & n8610 ;
  assign n8612 = n1406 & n7005 ;
  assign n8613 = n8612 ^ n4368 ^ 1'b0 ;
  assign n8614 = n288 | n4456 ;
  assign n8615 = n8614 ^ n8089 ^ 1'b0 ;
  assign n8618 = n2090 | n2833 ;
  assign n8616 = n1945 ^ n1449 ^ 1'b0 ;
  assign n8617 = n7481 & n8616 ;
  assign n8619 = n8618 ^ n8617 ^ n5382 ;
  assign n8620 = ( ~n398 & n2602 ) | ( ~n398 & n8619 ) | ( n2602 & n8619 ) ;
  assign n8621 = ( n1844 & n3830 ) | ( n1844 & ~n8620 ) | ( n3830 & ~n8620 ) ;
  assign n8622 = n5834 ^ n3113 ^ 1'b0 ;
  assign n8623 = ~n3439 & n8622 ;
  assign n8624 = n8623 ^ n505 ^ n288 ;
  assign n8625 = n1702 | n8624 ;
  assign n8626 = n8625 ^ n8512 ^ 1'b0 ;
  assign n8627 = n391 | n7222 ;
  assign n8628 = n8627 ^ n5113 ^ 1'b0 ;
  assign n8629 = n2027 | n8628 ;
  assign n8630 = n3793 | n8629 ;
  assign n8631 = n5879 ^ n1086 ^ 1'b0 ;
  assign n8632 = n2800 & ~n8631 ;
  assign n8633 = n5742 & n8632 ;
  assign n8634 = n8633 ^ n8365 ^ 1'b0 ;
  assign n8635 = n1364 & n8395 ;
  assign n8636 = n8635 ^ n2790 ^ 1'b0 ;
  assign n8637 = n7890 ^ n3189 ^ n1473 ;
  assign n8638 = ~n5067 & n8637 ;
  assign n8639 = ~n474 & n2226 ;
  assign n8640 = n8639 ^ n992 ^ 1'b0 ;
  assign n8641 = n8640 ^ n7271 ^ 1'b0 ;
  assign n8642 = n1077 & n2149 ;
  assign n8643 = ~n2065 & n8642 ;
  assign n8644 = n1442 & ~n8643 ;
  assign n8645 = n8644 ^ x51 ^ 1'b0 ;
  assign n8646 = n8641 | n8645 ;
  assign n8647 = n4446 | n8646 ;
  assign n8648 = n7420 | n7635 ;
  assign n8649 = n8647 | n8648 ;
  assign n8650 = n8181 ^ n1815 ^ 1'b0 ;
  assign n8651 = n1861 & ~n6891 ;
  assign n8652 = n8650 & n8651 ;
  assign n8653 = n319 & n7557 ;
  assign n8654 = n7945 ^ n7863 ^ n2364 ;
  assign n8655 = ( n4380 & n7968 ) | ( n4380 & n8654 ) | ( n7968 & n8654 ) ;
  assign n8656 = n7345 ^ n1791 ^ 1'b0 ;
  assign n8657 = n8152 | n8656 ;
  assign n8658 = n7647 ^ n3641 ^ 1'b0 ;
  assign n8659 = ~n7867 & n8658 ;
  assign n8660 = n6041 ^ n5504 ^ n3041 ;
  assign n8661 = n6028 ^ n2350 ^ n929 ;
  assign n8662 = n7879 ^ n4259 ^ 1'b0 ;
  assign n8663 = ~n8661 & n8662 ;
  assign n8664 = n1553 & ~n4407 ;
  assign n8665 = ( ~n169 & n1892 ) | ( ~n169 & n5614 ) | ( n1892 & n5614 ) ;
  assign n8666 = n7916 ^ n7323 ^ 1'b0 ;
  assign n8667 = n803 & n3434 ;
  assign n8668 = n8667 ^ x40 ^ 1'b0 ;
  assign n8669 = n1806 & n8668 ;
  assign n8670 = n2354 & ~n8029 ;
  assign n8671 = n8670 ^ n7701 ^ 1'b0 ;
  assign n8672 = ~x110 & n1222 ;
  assign n8673 = n8672 ^ n2547 ^ 1'b0 ;
  assign n8674 = n8673 ^ n8377 ^ 1'b0 ;
  assign n8676 = n664 & n1742 ;
  assign n8675 = n4054 | n4833 ;
  assign n8677 = n8676 ^ n8675 ^ 1'b0 ;
  assign n8678 = n8677 ^ n7370 ^ 1'b0 ;
  assign n8679 = n7999 ^ n477 ^ 1'b0 ;
  assign n8680 = n5767 & n8679 ;
  assign n8681 = n8680 ^ n4989 ^ 1'b0 ;
  assign n8682 = n6134 | n8681 ;
  assign n8683 = n6310 ^ n6265 ^ n371 ;
  assign n8684 = x2 & ~n8683 ;
  assign n8689 = n1197 & ~n3815 ;
  assign n8690 = ~n5012 & n8689 ;
  assign n8685 = n5281 ^ n3127 ^ n1670 ;
  assign n8686 = n3104 ^ n998 ^ 1'b0 ;
  assign n8687 = n5740 | n8686 ;
  assign n8688 = n8685 | n8687 ;
  assign n8691 = n8690 ^ n8688 ^ 1'b0 ;
  assign n8692 = n2435 & n8691 ;
  assign n8693 = ~n2414 & n8372 ;
  assign n8694 = n8693 ^ n5901 ^ 1'b0 ;
  assign n8695 = n3151 ^ n2219 ^ n576 ;
  assign n8696 = ~n1399 & n8695 ;
  assign n8697 = n859 & n8696 ;
  assign n8698 = n8697 ^ n2914 ^ 1'b0 ;
  assign n8699 = n8694 | n8698 ;
  assign n8700 = n5613 | n8699 ;
  assign n8701 = n4751 ^ n4011 ^ 1'b0 ;
  assign n8702 = n175 & n1374 ;
  assign n8703 = ~n8701 & n8702 ;
  assign n8704 = n1150 ^ n901 ^ 1'b0 ;
  assign n8705 = n567 & n8704 ;
  assign n8706 = n6337 ^ n3870 ^ n2636 ;
  assign n8707 = n8706 ^ x63 ^ 1'b0 ;
  assign n8709 = n202 & ~n928 ;
  assign n8710 = n2656 | n8709 ;
  assign n8711 = n8710 ^ n2932 ^ 1'b0 ;
  assign n8708 = n1716 | n7056 ;
  assign n8712 = n8711 ^ n8708 ^ 1'b0 ;
  assign n8713 = n5857 ^ n1421 ^ 1'b0 ;
  assign n8714 = n2923 | n8713 ;
  assign n8715 = n8714 ^ n5925 ^ 1'b0 ;
  assign n8716 = n3856 ^ n842 ^ 1'b0 ;
  assign n8717 = n4827 ^ n1927 ^ 1'b0 ;
  assign n8718 = n2379 ^ n1829 ^ 1'b0 ;
  assign n8719 = x106 & n3516 ;
  assign n8720 = n8719 ^ n5667 ^ 1'b0 ;
  assign n8721 = n8720 ^ n4927 ^ 1'b0 ;
  assign n8722 = ( n935 & n1013 ) | ( n935 & ~n8721 ) | ( n1013 & ~n8721 ) ;
  assign n8723 = n8145 ^ n2912 ^ 1'b0 ;
  assign n8724 = n2673 | n3705 ;
  assign n8725 = n8724 ^ n4017 ^ 1'b0 ;
  assign n8726 = n1829 ^ n1025 ^ 1'b0 ;
  assign n8727 = n756 | n8726 ;
  assign n8728 = n2870 & ~n4474 ;
  assign n8729 = n8727 & n8728 ;
  assign n8730 = n3831 | n7245 ;
  assign n8731 = n6658 ^ n5972 ^ 1'b0 ;
  assign n8732 = n4584 | n8731 ;
  assign n8733 = n6734 ^ n398 ^ 1'b0 ;
  assign n8734 = n1567 | n5092 ;
  assign n8735 = ( n1496 & n1501 ) | ( n1496 & n2034 ) | ( n1501 & n2034 ) ;
  assign n8736 = n297 & n8735 ;
  assign n8737 = n6588 & n8736 ;
  assign n8738 = n1473 & n7528 ;
  assign n8739 = n8737 | n8738 ;
  assign n8740 = n7904 | n8739 ;
  assign n8741 = n3249 | n5105 ;
  assign n8742 = n8741 ^ n4199 ^ 1'b0 ;
  assign n8743 = n7893 ^ n442 ^ 1'b0 ;
  assign n8744 = n5546 ^ n683 ^ 1'b0 ;
  assign n8745 = ~n978 & n8744 ;
  assign n8746 = n4755 ^ n621 ^ 1'b0 ;
  assign n8747 = n8745 & ~n8746 ;
  assign n8748 = n6250 ^ n1869 ^ n1481 ;
  assign n8749 = ~n7888 & n8748 ;
  assign n8750 = n1711 ^ x69 ^ 1'b0 ;
  assign n8751 = n935 & ~n8750 ;
  assign n8752 = n8751 ^ n3379 ^ n2658 ;
  assign n8753 = ~n5765 & n8752 ;
  assign n8755 = n691 & ~n3140 ;
  assign n8754 = n1265 & n5326 ;
  assign n8756 = n8755 ^ n8754 ^ 1'b0 ;
  assign n8757 = n2459 | n3906 ;
  assign n8758 = n7990 | n8757 ;
  assign n8759 = ( n1062 & n3372 ) | ( n1062 & ~n5785 ) | ( n3372 & ~n5785 ) ;
  assign n8760 = n8759 ^ n6363 ^ 1'b0 ;
  assign n8761 = n535 | n8760 ;
  assign n8762 = n2694 | n8761 ;
  assign n8763 = n1231 | n8762 ;
  assign n8764 = n8763 ^ n5316 ^ 1'b0 ;
  assign n8765 = n4596 ^ n1597 ^ n1436 ;
  assign n8766 = ( ~n569 & n2020 ) | ( ~n569 & n2529 ) | ( n2020 & n2529 ) ;
  assign n8767 = n8765 & n8766 ;
  assign n8768 = ( n357 & ~n3871 ) | ( n357 & n8767 ) | ( ~n3871 & n8767 ) ;
  assign n8769 = n8768 ^ n3532 ^ 1'b0 ;
  assign n8770 = n7672 | n8769 ;
  assign n8771 = n8770 ^ n8096 ^ 1'b0 ;
  assign n8772 = n8145 ^ n654 ^ 1'b0 ;
  assign n8773 = n8771 | n8772 ;
  assign n8774 = n2442 | n5057 ;
  assign n8775 = n8774 ^ n8479 ^ n6829 ;
  assign n8776 = n1224 ^ n487 ^ 1'b0 ;
  assign n8777 = n8776 ^ n7421 ^ n5985 ;
  assign n8778 = n3089 ^ n1607 ^ 1'b0 ;
  assign n8779 = n7328 | n8778 ;
  assign n8783 = n5745 ^ n1494 ^ n1471 ;
  assign n8784 = n1714 & ~n8783 ;
  assign n8785 = n8784 ^ n4806 ^ 1'b0 ;
  assign n8786 = n8785 ^ n3901 ^ 1'b0 ;
  assign n8780 = n984 ^ n849 ^ n473 ;
  assign n8781 = ~n8548 & n8780 ;
  assign n8782 = n5963 & n8781 ;
  assign n8787 = n8786 ^ n8782 ^ n4801 ;
  assign n8790 = n2473 | n5110 ;
  assign n8791 = n8790 ^ n623 ^ 1'b0 ;
  assign n8792 = n1906 | n8791 ;
  assign n8788 = n674 | n8358 ;
  assign n8789 = n4224 | n8788 ;
  assign n8793 = n8792 ^ n8789 ^ 1'b0 ;
  assign n8794 = n8793 ^ n5503 ^ n2897 ;
  assign n8795 = n2648 & n2847 ;
  assign n8796 = n2694 & n8795 ;
  assign n8797 = ~n2858 & n8796 ;
  assign n8798 = n8797 ^ n3003 ^ 1'b0 ;
  assign n8799 = n6807 ^ n644 ^ 1'b0 ;
  assign n8800 = n1312 ^ n722 ^ 1'b0 ;
  assign n8801 = ~n8799 & n8800 ;
  assign n8802 = n8223 ^ n6226 ^ 1'b0 ;
  assign n8803 = n1248 & ~n8802 ;
  assign n8804 = ( n3567 & n3793 ) | ( n3567 & ~n4127 ) | ( n3793 & ~n4127 ) ;
  assign n8805 = n8804 ^ n5817 ^ n726 ;
  assign n8806 = n8805 ^ n4087 ^ 1'b0 ;
  assign n8807 = n188 & n8806 ;
  assign n8808 = n483 & n2886 ;
  assign n8809 = n8808 ^ n2145 ^ 1'b0 ;
  assign n8810 = n6663 | n7262 ;
  assign n8811 = n4084 | n8810 ;
  assign n8812 = n6493 ^ n1106 ^ 1'b0 ;
  assign n8813 = ~n8084 & n8812 ;
  assign n8814 = n1113 & n1388 ;
  assign n8815 = n8814 ^ n1708 ^ 1'b0 ;
  assign n8816 = n2526 | n8815 ;
  assign n8817 = ( n799 & n8562 ) | ( n799 & n8816 ) | ( n8562 & n8816 ) ;
  assign n8818 = ( ~n607 & n2965 ) | ( ~n607 & n5848 ) | ( n2965 & n5848 ) ;
  assign n8819 = ~n3666 & n8818 ;
  assign n8820 = ~n3636 & n8819 ;
  assign n8821 = n5964 | n7888 ;
  assign n8825 = n2160 | n2996 ;
  assign n8826 = n6165 | n8825 ;
  assign n8823 = n2218 ^ n2036 ^ 1'b0 ;
  assign n8822 = n5633 | n7312 ;
  assign n8824 = n8823 ^ n8822 ^ 1'b0 ;
  assign n8827 = n8826 ^ n8824 ^ 1'b0 ;
  assign n8828 = n8267 & n8827 ;
  assign n8829 = n1863 & ~n6381 ;
  assign n8830 = ( ~n5488 & n6117 ) | ( ~n5488 & n8829 ) | ( n6117 & n8829 ) ;
  assign n8831 = n7874 & n8830 ;
  assign n8839 = n3954 | n4584 ;
  assign n8840 = n8265 | n8839 ;
  assign n8832 = n2362 ^ n1779 ^ n617 ;
  assign n8833 = n949 | n8832 ;
  assign n8836 = n415 & ~n7321 ;
  assign n8834 = n1162 & ~n3519 ;
  assign n8835 = n8834 ^ n7957 ^ n5516 ;
  assign n8837 = n8836 ^ n8835 ^ 1'b0 ;
  assign n8838 = n8833 & n8837 ;
  assign n8841 = n8840 ^ n8838 ^ 1'b0 ;
  assign n8842 = n3200 ^ n305 ^ 1'b0 ;
  assign n8843 = n4532 ^ n2045 ^ 1'b0 ;
  assign n8844 = n5786 & n8843 ;
  assign n8845 = n7622 & ~n8844 ;
  assign n8846 = n1077 & ~n1963 ;
  assign n8847 = n8846 ^ n7169 ^ 1'b0 ;
  assign n8848 = n8767 ^ n4075 ^ n2909 ;
  assign n8849 = ( ~n1014 & n2692 ) | ( ~n1014 & n8848 ) | ( n2692 & n8848 ) ;
  assign n8850 = n3339 ^ n1006 ^ 1'b0 ;
  assign n8851 = ~n8120 & n8850 ;
  assign n8852 = n1054 & n8851 ;
  assign n8853 = n6208 ^ n1485 ^ 1'b0 ;
  assign n8854 = n1846 & n8853 ;
  assign n8855 = ~n7714 & n8854 ;
  assign n8856 = n8855 ^ n8055 ^ 1'b0 ;
  assign n8857 = n7018 & n8856 ;
  assign n8858 = n1140 & n4859 ;
  assign n8859 = n8858 ^ n2609 ^ 1'b0 ;
  assign n8860 = n2151 ^ x72 ^ 1'b0 ;
  assign n8861 = n849 & ~n8860 ;
  assign n8862 = n8861 ^ n6602 ^ 1'b0 ;
  assign n8863 = n5114 & ~n8862 ;
  assign n8864 = n8863 ^ n196 ^ 1'b0 ;
  assign n8865 = n3396 | n8864 ;
  assign n8866 = n8859 | n8865 ;
  assign n8867 = n8866 ^ n4502 ^ 1'b0 ;
  assign n8868 = n7566 ^ n377 ^ 1'b0 ;
  assign n8869 = n5806 & ~n8868 ;
  assign n8872 = n5326 ^ n1111 ^ 1'b0 ;
  assign n8870 = n2687 & ~n6053 ;
  assign n8871 = ~n3953 & n8870 ;
  assign n8873 = n8872 ^ n8871 ^ 1'b0 ;
  assign n8874 = n5641 ^ n1772 ^ 1'b0 ;
  assign n8875 = ( n1505 & n5395 ) | ( n1505 & n5637 ) | ( n5395 & n5637 ) ;
  assign n8876 = n8875 ^ n6959 ^ 1'b0 ;
  assign n8877 = n6421 | n8876 ;
  assign n8878 = n8877 ^ n7304 ^ 1'b0 ;
  assign n8879 = ( n254 & n5407 ) | ( n254 & n7048 ) | ( n5407 & n7048 ) ;
  assign n8880 = ( n5466 & n7785 ) | ( n5466 & ~n8879 ) | ( n7785 & ~n8879 ) ;
  assign n8882 = n6102 ^ n906 ^ 1'b0 ;
  assign n8883 = n8882 ^ n4911 ^ n3933 ;
  assign n8881 = ~n5897 & n6164 ;
  assign n8884 = n8883 ^ n8881 ^ 1'b0 ;
  assign n8885 = n4548 | n7613 ;
  assign n8886 = n8885 ^ n7108 ^ 1'b0 ;
  assign n8887 = n1842 | n2348 ;
  assign n8888 = n3571 ^ n1086 ^ 1'b0 ;
  assign n8889 = ~n8818 & n8888 ;
  assign n8890 = n8887 & n8889 ;
  assign n8891 = n3117 | n4297 ;
  assign n8892 = n6157 & ~n8891 ;
  assign n8893 = n8892 ^ n5915 ^ 1'b0 ;
  assign n8894 = n6926 & n8893 ;
  assign n8895 = ( ~n1741 & n5250 ) | ( ~n1741 & n7305 ) | ( n5250 & n7305 ) ;
  assign n8896 = n8895 ^ n7638 ^ 1'b0 ;
  assign n8899 = n3391 | n5692 ;
  assign n8897 = n5118 | n5123 ;
  assign n8898 = n1250 | n8897 ;
  assign n8900 = n8899 ^ n8898 ^ n5219 ;
  assign n8901 = n8885 | n8900 ;
  assign n8902 = n8901 ^ n6288 ^ 1'b0 ;
  assign n8908 = n3710 | n5960 ;
  assign n8903 = ( n275 & n1338 ) | ( n275 & n5659 ) | ( n1338 & n5659 ) ;
  assign n8904 = n2049 & ~n8903 ;
  assign n8905 = n786 & n8904 ;
  assign n8906 = n3758 ^ n2803 ^ 1'b0 ;
  assign n8907 = ~n8905 & n8906 ;
  assign n8909 = n8908 ^ n8907 ^ 1'b0 ;
  assign n8910 = n2521 ^ n1679 ^ 1'b0 ;
  assign n8911 = n5391 | n8910 ;
  assign n8912 = ~n4806 & n8911 ;
  assign n8913 = n1976 & n8912 ;
  assign n8914 = n3232 ^ n135 ^ 1'b0 ;
  assign n8915 = n8914 ^ n1013 ^ 1'b0 ;
  assign n8919 = n2833 ^ n1730 ^ n151 ;
  assign n8916 = n854 | n7352 ;
  assign n8917 = n8916 ^ n4292 ^ 1'b0 ;
  assign n8918 = ~n3694 & n8917 ;
  assign n8920 = n8919 ^ n8918 ^ 1'b0 ;
  assign n8921 = ~n3347 & n8920 ;
  assign n8922 = ~n8915 & n8921 ;
  assign n8923 = n4165 & n6564 ;
  assign n8924 = n1505 ^ n250 ^ 1'b0 ;
  assign n8925 = n8923 & n8924 ;
  assign n8926 = n5083 ^ n909 ^ 1'b0 ;
  assign n8927 = n8925 & ~n8926 ;
  assign n8928 = n8927 ^ n196 ^ 1'b0 ;
  assign n8929 = n6257 ^ n1791 ^ n419 ;
  assign n8930 = ~n2509 & n8929 ;
  assign n8931 = n8930 ^ n2692 ^ 1'b0 ;
  assign n8932 = n7691 ^ n2063 ^ 1'b0 ;
  assign n8933 = n8931 & n8932 ;
  assign n8934 = n8933 ^ n8856 ^ x13 ;
  assign n8935 = n8303 | n8934 ;
  assign n8936 = n8935 ^ n2727 ^ 1'b0 ;
  assign n8937 = n7177 ^ n3265 ^ 1'b0 ;
  assign n8938 = x115 & ~n1286 ;
  assign n8939 = n2675 | n8938 ;
  assign n8940 = n569 & n8939 ;
  assign n8941 = n3587 & ~n3878 ;
  assign n8942 = ~n1791 & n8941 ;
  assign n8943 = n5815 | n8942 ;
  assign n8944 = n8170 & ~n8943 ;
  assign n8945 = ~n1991 & n3630 ;
  assign n8946 = x107 | n149 ;
  assign n8947 = ~n1601 & n5574 ;
  assign n8948 = n8947 ^ n1238 ^ 1'b0 ;
  assign n8949 = n8948 ^ n7450 ^ 1'b0 ;
  assign n8950 = n7915 & n8766 ;
  assign n8951 = n8949 & ~n8950 ;
  assign n8952 = ~n8946 & n8951 ;
  assign n8953 = n7368 ^ n1012 ^ 1'b0 ;
  assign n8954 = n6982 & n8953 ;
  assign n8955 = ~n5840 & n8954 ;
  assign n8956 = n4180 ^ n3219 ^ 1'b0 ;
  assign n8957 = n8956 ^ n4662 ^ 1'b0 ;
  assign n8958 = n5742 ^ n5446 ^ 1'b0 ;
  assign n8959 = n5850 ^ n1652 ^ n1384 ;
  assign n8960 = n1876 & n3353 ;
  assign n8961 = n4348 ^ n748 ^ 1'b0 ;
  assign n8962 = n8259 & ~n8961 ;
  assign n8963 = n8960 & ~n8962 ;
  assign n8964 = n1998 & n5175 ;
  assign n8965 = n8964 ^ n6550 ^ 1'b0 ;
  assign n8966 = n7625 | n8965 ;
  assign n8967 = ( n196 & ~n8867 ) | ( n196 & n8966 ) | ( ~n8867 & n8966 ) ;
  assign n8968 = ~n5517 & n5791 ;
  assign n8969 = n8968 ^ n3633 ^ 1'b0 ;
  assign n8970 = n6478 ^ n3243 ^ 1'b0 ;
  assign n8971 = ~n8500 & n8970 ;
  assign n8972 = n3342 ^ n1440 ^ 1'b0 ;
  assign n8974 = ~n548 & n1621 ;
  assign n8977 = n2175 ^ n361 ^ 1'b0 ;
  assign n8975 = n4169 ^ n3830 ^ 1'b0 ;
  assign n8976 = n5683 & ~n8975 ;
  assign n8978 = n8977 ^ n8976 ^ n7806 ;
  assign n8979 = ( n431 & n8974 ) | ( n431 & n8978 ) | ( n8974 & n8978 ) ;
  assign n8973 = ~n3576 & n8765 ;
  assign n8980 = n8979 ^ n8973 ^ 1'b0 ;
  assign n8986 = n1222 & ~n2451 ;
  assign n8987 = ~n1222 & n8986 ;
  assign n8988 = n8987 ^ n4419 ^ 1'b0 ;
  assign n8981 = n3217 & ~n4259 ;
  assign n8982 = n1534 ^ n1410 ^ n166 ;
  assign n8983 = n8982 ^ n466 ^ 1'b0 ;
  assign n8984 = n8981 | n8983 ;
  assign n8985 = n6759 | n8984 ;
  assign n8989 = n8988 ^ n8985 ^ 1'b0 ;
  assign n8990 = n521 | n1634 ;
  assign n8991 = n8990 ^ n832 ^ 1'b0 ;
  assign n8992 = n2859 & n8991 ;
  assign n8993 = n8992 ^ n2206 ^ n1591 ;
  assign n8994 = n1788 ^ n1443 ^ 1'b0 ;
  assign n8995 = n4684 ^ n439 ^ 1'b0 ;
  assign n8996 = n8994 & n8995 ;
  assign n8997 = n8996 ^ n5394 ^ 1'b0 ;
  assign n8998 = n775 | n8997 ;
  assign n8999 = ~n4358 & n4454 ;
  assign n9002 = n1084 | n6829 ;
  assign n9000 = n7484 & ~n8628 ;
  assign n9001 = n3739 & n9000 ;
  assign n9003 = n9002 ^ n9001 ^ 1'b0 ;
  assign n9004 = n196 | n6654 ;
  assign n9005 = n9004 ^ n2692 ^ 1'b0 ;
  assign n9006 = n496 ^ x116 ^ 1'b0 ;
  assign n9007 = n2246 & ~n9006 ;
  assign n9008 = n9007 ^ n2040 ^ 1'b0 ;
  assign n9009 = n9008 ^ n6563 ^ n1664 ;
  assign n9010 = n1420 & ~n9009 ;
  assign n9011 = n3849 ^ n1045 ^ 1'b0 ;
  assign n9012 = ~n918 & n1861 ;
  assign n9013 = n3876 & ~n9012 ;
  assign n9014 = n9011 | n9013 ;
  assign n9015 = n9010 & ~n9014 ;
  assign n9016 = n408 & ~n849 ;
  assign n9017 = ~n8341 & n9016 ;
  assign n9018 = n9017 ^ n369 ^ 1'b0 ;
  assign n9019 = n703 & ~n9018 ;
  assign n9020 = n1613 & n9019 ;
  assign n9021 = n4757 | n9020 ;
  assign n9022 = n9021 ^ n7666 ^ 1'b0 ;
  assign n9023 = n5361 ^ n5231 ^ 1'b0 ;
  assign n9024 = n2019 & n9023 ;
  assign n9025 = n1948 | n2089 ;
  assign n9026 = n9025 ^ n3586 ^ 1'b0 ;
  assign n9027 = n9026 ^ n4136 ^ 1'b0 ;
  assign n9028 = ~n1637 & n2623 ;
  assign n9029 = n2140 & n9028 ;
  assign n9030 = ( n4963 & n9027 ) | ( n4963 & ~n9029 ) | ( n9027 & ~n9029 ) ;
  assign n9031 = n7791 ^ n738 ^ 1'b0 ;
  assign n9032 = n9030 & ~n9031 ;
  assign n9033 = n9032 ^ n8878 ^ 1'b0 ;
  assign n9034 = n4125 & n7004 ;
  assign n9035 = n6633 & n9034 ;
  assign n9045 = n681 ^ n512 ^ 1'b0 ;
  assign n9038 = n4522 ^ n1997 ^ 1'b0 ;
  assign n9039 = n8531 | n9038 ;
  assign n9036 = n4026 | n6705 ;
  assign n9037 = n3313 | n9036 ;
  assign n9040 = n9039 ^ n9037 ^ 1'b0 ;
  assign n9041 = n3831 & ~n9040 ;
  assign n9042 = n9041 ^ n2742 ^ 1'b0 ;
  assign n9043 = n245 & n9042 ;
  assign n9044 = n6668 & n9043 ;
  assign n9046 = n9045 ^ n9044 ^ 1'b0 ;
  assign n9047 = n1106 | n9046 ;
  assign n9048 = n4594 & ~n9047 ;
  assign n9049 = ~n3026 & n3931 ;
  assign n9050 = n9049 ^ n3981 ^ 1'b0 ;
  assign n9051 = ~n3724 & n9050 ;
  assign n9052 = ~n2193 & n9051 ;
  assign n9053 = n8657 | n9052 ;
  assign n9054 = n8621 | n9053 ;
  assign n9055 = n4859 ^ n2715 ^ x56 ;
  assign n9056 = ( x14 & n3697 ) | ( x14 & ~n5737 ) | ( n3697 & ~n5737 ) ;
  assign n9057 = n9056 ^ n3224 ^ 1'b0 ;
  assign n9058 = n3153 & ~n6770 ;
  assign n9059 = n4467 & n9058 ;
  assign n9060 = ( x30 & ~n9057 ) | ( x30 & n9059 ) | ( ~n9057 & n9059 ) ;
  assign n9061 = n9060 ^ n3678 ^ 1'b0 ;
  assign n9062 = n6299 & ~n8076 ;
  assign n9063 = ( n744 & n1490 ) | ( n744 & ~n5911 ) | ( n1490 & ~n5911 ) ;
  assign n9064 = ~n876 & n9063 ;
  assign n9065 = ~n984 & n5017 ;
  assign n9066 = n9065 ^ n6711 ^ 1'b0 ;
  assign n9069 = ~x89 & n748 ;
  assign n9067 = n7160 ^ n2214 ^ 1'b0 ;
  assign n9068 = n6168 & n9067 ;
  assign n9070 = n9069 ^ n9068 ^ 1'b0 ;
  assign n9071 = n1903 & n9070 ;
  assign n9074 = ~n1580 & n3985 ;
  assign n9072 = ~n956 & n6195 ;
  assign n9073 = n8413 & n9072 ;
  assign n9075 = n9074 ^ n9073 ^ 1'b0 ;
  assign n9076 = n1314 & ~n6590 ;
  assign n9077 = n9076 ^ n3794 ^ 1'b0 ;
  assign n9078 = n5968 ^ n2562 ^ n1843 ;
  assign n9079 = n9078 ^ n7416 ^ 1'b0 ;
  assign n9080 = n4771 ^ n373 ^ 1'b0 ;
  assign n9081 = n5137 & n9080 ;
  assign n9082 = n7921 & n9081 ;
  assign n9083 = n9082 ^ n3838 ^ 1'b0 ;
  assign n9084 = n7089 ^ n1422 ^ 1'b0 ;
  assign n9085 = n9084 ^ n4725 ^ 1'b0 ;
  assign n9086 = ( n2173 & ~n3979 ) | ( n2173 & n5790 ) | ( ~n3979 & n5790 ) ;
  assign n9087 = n9086 ^ n6166 ^ 1'b0 ;
  assign n9088 = n9085 & ~n9087 ;
  assign n9089 = ~n1138 & n3414 ;
  assign n9090 = n1540 & n9089 ;
  assign n9091 = ~n1489 & n1990 ;
  assign n9092 = n9091 ^ n1963 ^ 1'b0 ;
  assign n9093 = n1909 & ~n9092 ;
  assign n9094 = ~n8501 & n9093 ;
  assign n9095 = n3628 | n9094 ;
  assign n9096 = n9090 & ~n9095 ;
  assign n9097 = x26 & n908 ;
  assign n9098 = ~x26 & n9097 ;
  assign n9099 = n242 & n1746 ;
  assign n9100 = ~n242 & n9099 ;
  assign n9101 = n536 | n9100 ;
  assign n9102 = n9100 & ~n9101 ;
  assign n9103 = x73 & ~n1197 ;
  assign n9104 = ~x73 & n9103 ;
  assign n9105 = n9102 & ~n9104 ;
  assign n9106 = x89 & ~n237 ;
  assign n9107 = ~x89 & n9106 ;
  assign n9108 = n419 & ~n9107 ;
  assign n9109 = n9107 & n9108 ;
  assign n9110 = n1795 ^ n1295 ^ 1'b0 ;
  assign n9111 = n9109 | n9110 ;
  assign n9112 = ( ~n9098 & n9105 ) | ( ~n9098 & n9111 ) | ( n9105 & n9111 ) ;
  assign n9113 = n917 | n1690 ;
  assign n9114 = n917 & ~n9113 ;
  assign n9115 = x3 & ~n9114 ;
  assign n9119 = x62 & x71 ;
  assign n9120 = ~x71 & n9119 ;
  assign n9121 = n533 | n9120 ;
  assign n9122 = n9120 & ~n9121 ;
  assign n9116 = ~n295 & n1905 ;
  assign n9117 = n295 & n9116 ;
  assign n9118 = n642 | n9117 ;
  assign n9123 = n9122 ^ n9118 ^ 1'b0 ;
  assign n9124 = n9115 & ~n9123 ;
  assign n9125 = n9112 & n9124 ;
  assign n9126 = n736 | n3369 ;
  assign n9127 = n3369 & ~n9126 ;
  assign n9128 = n5487 | n9127 ;
  assign n9129 = n9125 & ~n9128 ;
  assign n9130 = n7761 ^ n2057 ^ n208 ;
  assign n9131 = n8227 ^ n5116 ^ 1'b0 ;
  assign n9134 = n3354 ^ n1718 ^ 1'b0 ;
  assign n9132 = n1961 ^ n150 ^ 1'b0 ;
  assign n9133 = n146 & n9132 ;
  assign n9135 = n9134 ^ n9133 ^ 1'b0 ;
  assign n9136 = n1062 & n1330 ;
  assign n9137 = n965 & n9136 ;
  assign n9138 = n2453 & ~n9137 ;
  assign n9139 = n2384 & n4761 ;
  assign n9140 = n9139 ^ n2011 ^ 1'b0 ;
  assign n9142 = n3107 & n3791 ;
  assign n9141 = x15 & ~n7709 ;
  assign n9143 = n9142 ^ n9141 ^ 1'b0 ;
  assign n9144 = ( n143 & n2142 ) | ( n143 & n3643 ) | ( n2142 & n3643 ) ;
  assign n9145 = n259 | n9144 ;
  assign n9146 = n7142 ^ n2770 ^ 1'b0 ;
  assign n9147 = n9145 | n9146 ;
  assign n9148 = n9147 ^ n3886 ^ 1'b0 ;
  assign n9149 = n3516 | n9148 ;
  assign n9150 = n9149 ^ n7129 ^ 1'b0 ;
  assign n9151 = n6689 | n8154 ;
  assign n9152 = n8920 | n9151 ;
  assign n9153 = n1165 & ~n6018 ;
  assign n9154 = n9153 ^ n7178 ^ 1'b0 ;
  assign n9155 = n1669 & ~n9154 ;
  assign n9156 = n2579 & n9155 ;
  assign n9160 = n3038 & ~n4141 ;
  assign n9161 = n1498 & n9160 ;
  assign n9162 = n4921 & ~n9161 ;
  assign n9157 = n6206 ^ n3578 ^ 1'b0 ;
  assign n9158 = n2035 & ~n9157 ;
  assign n9159 = ( ~n4748 & n6023 ) | ( ~n4748 & n9158 ) | ( n6023 & n9158 ) ;
  assign n9163 = n9162 ^ n9159 ^ 1'b0 ;
  assign n9164 = ( n225 & ~n2112 ) | ( n225 & n3742 ) | ( ~n2112 & n3742 ) ;
  assign n9165 = n7195 & ~n9164 ;
  assign n9166 = ~n6769 & n9165 ;
  assign n9167 = n8903 ^ n4441 ^ n4076 ;
  assign n9168 = n4337 | n8157 ;
  assign n9169 = n3717 | n9168 ;
  assign n9170 = n9169 ^ n324 ^ 1'b0 ;
  assign n9171 = n9167 & n9170 ;
  assign n9172 = n4710 | n9171 ;
  assign n9176 = ~n4120 & n6114 ;
  assign n9173 = n1559 & ~n2549 ;
  assign n9174 = n4131 & n9173 ;
  assign n9175 = n9174 ^ n3927 ^ n2021 ;
  assign n9177 = n9176 ^ n9175 ^ 1'b0 ;
  assign n9178 = n716 & ~n2234 ;
  assign n9179 = n9178 ^ n3235 ^ x78 ;
  assign n9180 = n6140 ^ n5945 ^ 1'b0 ;
  assign n9181 = n4207 ^ n1243 ^ 1'b0 ;
  assign n9182 = n706 & ~n775 ;
  assign n9183 = ( n9180 & ~n9181 ) | ( n9180 & n9182 ) | ( ~n9181 & n9182 ) ;
  assign n9184 = n3903 & n9183 ;
  assign n9185 = n150 & ~n9184 ;
  assign n9186 = n5957 & n9185 ;
  assign n9187 = n7328 ^ n2007 ^ 1'b0 ;
  assign n9191 = n2649 & n2737 ;
  assign n9192 = n9191 ^ n3739 ^ 1'b0 ;
  assign n9188 = x31 & ~n4362 ;
  assign n9189 = ~n5139 & n9188 ;
  assign n9190 = n5651 | n9189 ;
  assign n9193 = n9192 ^ n9190 ^ 1'b0 ;
  assign n9194 = n5165 ^ n2802 ^ x103 ;
  assign n9195 = n6350 ^ n3308 ^ 1'b0 ;
  assign n9196 = ~n2386 & n9195 ;
  assign n9197 = n4998 ^ n1894 ^ 1'b0 ;
  assign n9198 = ~n3365 & n3434 ;
  assign n9199 = ( n2912 & n6135 ) | ( n2912 & ~n9198 ) | ( n6135 & ~n9198 ) ;
  assign n9200 = n6998 & n9199 ;
  assign n9201 = n9200 ^ n618 ^ 1'b0 ;
  assign n9202 = n6846 ^ n1860 ^ 1'b0 ;
  assign n9203 = n484 & ~n9202 ;
  assign n9204 = n9203 ^ n493 ^ 1'b0 ;
  assign n9205 = n1970 | n9204 ;
  assign n9206 = n9205 ^ n1057 ^ 1'b0 ;
  assign n9207 = n5036 | n6079 ;
  assign n9208 = n221 & ~n9207 ;
  assign n9209 = n6102 ^ n4429 ^ n4088 ;
  assign n9210 = n9209 ^ n5505 ^ 1'b0 ;
  assign n9211 = n9210 ^ n2354 ^ 1'b0 ;
  assign n9212 = n2741 & ~n7376 ;
  assign n9213 = ~n4002 & n9212 ;
  assign n9214 = ~n7561 & n9213 ;
  assign n9215 = n9214 ^ n305 ^ 1'b0 ;
  assign n9216 = ( ~n2928 & n3918 ) | ( ~n2928 & n8013 ) | ( n3918 & n8013 ) ;
  assign n9217 = n9216 ^ n380 ^ 1'b0 ;
  assign n9218 = ~n7305 & n9217 ;
  assign n9219 = n529 | n8289 ;
  assign n9220 = n9219 ^ n3441 ^ 1'b0 ;
  assign n9221 = ~n612 & n1953 ;
  assign n9222 = n9221 ^ n143 ^ 1'b0 ;
  assign n9223 = n7176 ^ n4385 ^ n2979 ;
  assign n9224 = n9223 ^ n2485 ^ 1'b0 ;
  assign n9225 = ~n8582 & n9224 ;
  assign n9226 = n9222 & n9225 ;
  assign n9227 = ~n4765 & n5053 ;
  assign n9228 = n856 & ~n1578 ;
  assign n9229 = ~n1553 & n5318 ;
  assign n9230 = n4876 ^ n194 ^ 1'b0 ;
  assign n9231 = ~n3710 & n9230 ;
  assign n9232 = x72 & n6131 ;
  assign n9233 = n9232 ^ n6087 ^ 1'b0 ;
  assign n9234 = n9233 ^ n7737 ^ 1'b0 ;
  assign n9235 = n7812 & ~n9234 ;
  assign n9236 = ~n9231 & n9235 ;
  assign n9237 = n1286 ^ n442 ^ 1'b0 ;
  assign n9238 = ( n1008 & ~n1202 ) | ( n1008 & n5633 ) | ( ~n1202 & n5633 ) ;
  assign n9239 = ( n939 & ~n6867 ) | ( n939 & n9238 ) | ( ~n6867 & n9238 ) ;
  assign n9240 = n1097 & ~n9239 ;
  assign n9241 = n3025 | n3734 ;
  assign n9242 = ~n2223 & n5179 ;
  assign n9243 = n2780 & n9242 ;
  assign n9244 = n9243 ^ n672 ^ 1'b0 ;
  assign n9245 = n9241 & ~n9244 ;
  assign n9246 = n5701 ^ n817 ^ 1'b0 ;
  assign n9247 = n148 | n9246 ;
  assign n9248 = n7521 ^ n4503 ^ 1'b0 ;
  assign n9249 = ~n9247 & n9248 ;
  assign n9250 = n7967 ^ x90 ^ 1'b0 ;
  assign n9251 = n245 & n9250 ;
  assign n9252 = ~n6514 & n9251 ;
  assign n9253 = n9252 ^ n852 ^ 1'b0 ;
  assign n9254 = n1459 | n8541 ;
  assign n9255 = n8156 | n9254 ;
  assign n9256 = n9255 ^ n6421 ^ 1'b0 ;
  assign n9257 = n6571 & ~n9256 ;
  assign n9258 = n5171 & ~n6402 ;
  assign n9259 = n3978 ^ n2996 ^ 1'b0 ;
  assign n9260 = n5051 | n9259 ;
  assign n9261 = n3666 & n8104 ;
  assign n9262 = n9261 ^ n319 ^ 1'b0 ;
  assign n9263 = n6402 ^ n2755 ^ 1'b0 ;
  assign n9264 = n1794 & ~n2721 ;
  assign n9265 = ~n3482 & n9264 ;
  assign n9266 = n5211 | n9265 ;
  assign n9267 = n3379 | n9266 ;
  assign n9268 = ~n1992 & n5213 ;
  assign n9269 = n4449 ^ n1895 ^ 1'b0 ;
  assign n9270 = ~n9268 & n9269 ;
  assign n9271 = n2568 & ~n9270 ;
  assign n9272 = n6830 ^ n6157 ^ 1'b0 ;
  assign n9273 = ~n265 & n9272 ;
  assign n9274 = n9273 ^ n3868 ^ 1'b0 ;
  assign n9275 = n992 & ~n3794 ;
  assign n9276 = n2668 & ~n9275 ;
  assign n9277 = n9276 ^ n801 ^ 1'b0 ;
  assign n9278 = x94 & n9277 ;
  assign n9279 = n6813 & n9278 ;
  assign n9280 = ~n1100 & n9279 ;
  assign n9281 = n5314 ^ n508 ^ 1'b0 ;
  assign n9282 = n7178 | n9281 ;
  assign n9283 = n2861 & n7869 ;
  assign n9284 = n9282 | n9283 ;
  assign n9285 = n3403 ^ n2254 ^ n579 ;
  assign n9286 = n9285 ^ n2809 ^ 1'b0 ;
  assign n9287 = n256 & n9286 ;
  assign n9288 = ~n6238 & n7812 ;
  assign n9289 = n6040 & n9288 ;
  assign n9290 = n3480 & ~n9289 ;
  assign n9291 = n9290 ^ n4865 ^ 1'b0 ;
  assign n9292 = n786 & n5006 ;
  assign n9293 = n2479 | n8567 ;
  assign n9294 = n9292 | n9293 ;
  assign n9295 = ~n439 & n9294 ;
  assign n9296 = n6716 & n9295 ;
  assign n9297 = x119 & ~n7161 ;
  assign n9298 = ~n2266 & n9297 ;
  assign n9299 = n9298 ^ n2940 ^ 1'b0 ;
  assign n9300 = n179 & ~n5261 ;
  assign n9301 = ~n1601 & n2455 ;
  assign n9302 = n9301 ^ n2654 ^ 1'b0 ;
  assign n9303 = n2404 & ~n9302 ;
  assign n9304 = n2959 | n5169 ;
  assign n9305 = ( n234 & ~n9303 ) | ( n234 & n9304 ) | ( ~n9303 & n9304 ) ;
  assign n9306 = n4597 ^ x80 ^ 1'b0 ;
  assign n9307 = n8124 & n9306 ;
  assign n9308 = n9307 ^ n4121 ^ 1'b0 ;
  assign n9309 = n5339 ^ n2815 ^ 1'b0 ;
  assign n9310 = n5456 & n9309 ;
  assign n9311 = x25 & n5356 ;
  assign n9312 = ~n9310 & n9311 ;
  assign n9313 = n4802 ^ n1197 ^ 1'b0 ;
  assign n9314 = n7866 & ~n9313 ;
  assign n9315 = n1943 & ~n8705 ;
  assign n9316 = n4186 ^ n3335 ^ 1'b0 ;
  assign n9317 = n5952 | n9316 ;
  assign n9318 = ( n4740 & n5185 ) | ( n4740 & n6642 ) | ( n5185 & n6642 ) ;
  assign n9319 = n1501 & ~n1872 ;
  assign n9320 = n9319 ^ n2023 ^ 1'b0 ;
  assign n9321 = n3016 & ~n9320 ;
  assign n9322 = n9321 ^ n4091 ^ n2256 ;
  assign n9323 = n4589 | n5767 ;
  assign n9324 = n8011 ^ n2048 ^ 1'b0 ;
  assign n9325 = ( n969 & n9323 ) | ( n969 & ~n9324 ) | ( n9323 & ~n9324 ) ;
  assign n9326 = ( n1571 & n1989 ) | ( n1571 & ~n3276 ) | ( n1989 & ~n3276 ) ;
  assign n9327 = x97 | n9326 ;
  assign n9328 = n4227 | n9327 ;
  assign n9329 = n5848 ^ n3213 ^ 1'b0 ;
  assign n9330 = ~n4612 & n9329 ;
  assign n9331 = n9330 ^ n1700 ^ 1'b0 ;
  assign n9332 = ~n9328 & n9331 ;
  assign n9333 = n9332 ^ n398 ^ 1'b0 ;
  assign n9334 = x60 & n9333 ;
  assign n9335 = n7479 | n9334 ;
  assign n9336 = n3003 & ~n8480 ;
  assign n9337 = n9336 ^ n2980 ^ 1'b0 ;
  assign n9343 = ( n480 & ~n1594 ) | ( n480 & n5677 ) | ( ~n1594 & n5677 ) ;
  assign n9338 = n1619 | n1982 ;
  assign n9339 = n2329 | n9338 ;
  assign n9340 = n9339 ^ n1687 ^ 1'b0 ;
  assign n9341 = n3999 & ~n9340 ;
  assign n9342 = n9341 ^ n892 ^ 1'b0 ;
  assign n9344 = n9343 ^ n9342 ^ n3608 ;
  assign n9345 = n8340 ^ n191 ^ 1'b0 ;
  assign n9346 = ~n7707 & n9345 ;
  assign n9347 = n2231 & ~n2275 ;
  assign n9348 = n9347 ^ n210 ^ 1'b0 ;
  assign n9349 = n9348 ^ n4422 ^ n1935 ;
  assign n9350 = n2437 ^ n982 ^ 1'b0 ;
  assign n9351 = n4298 | n9350 ;
  assign n9352 = n9349 & ~n9351 ;
  assign n9356 = n8737 ^ n586 ^ 1'b0 ;
  assign n9353 = n3191 ^ n2479 ^ 1'b0 ;
  assign n9354 = n565 & n9353 ;
  assign n9355 = n8681 & n9354 ;
  assign n9357 = n9356 ^ n9355 ^ 1'b0 ;
  assign n9358 = n1418 | n8720 ;
  assign n9359 = n1418 & ~n9358 ;
  assign n9360 = n937 | n9359 ;
  assign n9361 = n1403 | n9360 ;
  assign n9362 = n9361 ^ n1440 ^ 1'b0 ;
  assign n9363 = n833 & ~n4475 ;
  assign n9364 = n8905 ^ n1935 ^ n374 ;
  assign n9365 = n5837 & ~n9364 ;
  assign n9366 = n2255 & n9365 ;
  assign n9367 = n9366 ^ x15 ^ 1'b0 ;
  assign n9368 = n452 | n9367 ;
  assign n9370 = n2595 ^ x23 ^ 1'b0 ;
  assign n9369 = n2151 & n8887 ;
  assign n9371 = n9370 ^ n9369 ^ n235 ;
  assign n9372 = ~n256 & n1364 ;
  assign n9373 = n9372 ^ n1841 ^ 1'b0 ;
  assign n9374 = n2152 & n9373 ;
  assign n9375 = n9374 ^ x8 ^ 1'b0 ;
  assign n9376 = ~n2323 & n3440 ;
  assign n9377 = n3189 & ~n8156 ;
  assign n9378 = n9376 & n9377 ;
  assign n9379 = n3893 & n9378 ;
  assign n9380 = n167 | n2801 ;
  assign n9381 = n9380 ^ n8487 ^ 1'b0 ;
  assign n9382 = ~n8565 & n9381 ;
  assign n9383 = n9382 ^ n3608 ^ 1'b0 ;
  assign n9384 = n2642 | n9383 ;
  assign n9385 = n3340 | n3406 ;
  assign n9386 = n6162 & ~n9349 ;
  assign n9387 = ~n2331 & n9386 ;
  assign n9388 = n1880 | n4071 ;
  assign n9389 = n4231 & ~n9388 ;
  assign n9390 = n9389 ^ n6782 ^ 1'b0 ;
  assign n9391 = n9204 ^ n4380 ^ x57 ;
  assign n9392 = ~n6738 & n9391 ;
  assign n9393 = ~n8613 & n9392 ;
  assign n9394 = n7563 ^ n5014 ^ 1'b0 ;
  assign n9395 = n516 & ~n9394 ;
  assign n9397 = n2675 | n4362 ;
  assign n9398 = n5396 | n9397 ;
  assign n9396 = n3860 & n5712 ;
  assign n9399 = n9398 ^ n9396 ^ n373 ;
  assign n9400 = n7688 ^ n4407 ^ 1'b0 ;
  assign n9401 = n2755 & n9400 ;
  assign n9402 = n9401 ^ n2106 ^ 1'b0 ;
  assign n9403 = n9402 ^ n493 ^ 1'b0 ;
  assign n9404 = n5034 ^ n3250 ^ 1'b0 ;
  assign n9405 = ( n935 & n9403 ) | ( n935 & n9404 ) | ( n9403 & n9404 ) ;
  assign n9406 = n3744 & n4601 ;
  assign n9407 = n5017 & n9406 ;
  assign n9408 = n7342 & n9133 ;
  assign n9409 = n2793 & n9408 ;
  assign n9410 = n5989 & ~n9409 ;
  assign n9411 = n5088 & n9410 ;
  assign n9412 = ( n288 & n840 ) | ( n288 & n2780 ) | ( n840 & n2780 ) ;
  assign n9413 = ( n891 & n1311 ) | ( n891 & ~n9412 ) | ( n1311 & ~n9412 ) ;
  assign n9414 = n9413 ^ n4776 ^ 1'b0 ;
  assign n9415 = n6986 & n9414 ;
  assign n9416 = n4497 ^ n1314 ^ 1'b0 ;
  assign n9417 = ~n1994 & n9416 ;
  assign n9418 = n1771 ^ n503 ^ 1'b0 ;
  assign n9419 = n9418 ^ n2981 ^ 1'b0 ;
  assign n9420 = n9417 & n9419 ;
  assign n9421 = ~n1619 & n8424 ;
  assign n9422 = ~n5216 & n9421 ;
  assign n9423 = n8999 ^ n5046 ^ 1'b0 ;
  assign n9424 = n4102 | n9423 ;
  assign n9425 = ~n654 & n3975 ;
  assign n9426 = ( x118 & n1125 ) | ( x118 & ~n9425 ) | ( n1125 & ~n9425 ) ;
  assign n9427 = n2509 | n9426 ;
  assign n9428 = n5511 & n7666 ;
  assign n9429 = n7731 | n8598 ;
  assign n9430 = n4778 | n9429 ;
  assign n9431 = n2102 | n8372 ;
  assign n9432 = ~n355 & n6771 ;
  assign n9433 = n2036 | n9432 ;
  assign n9434 = n9433 ^ n4186 ^ 1'b0 ;
  assign n9435 = ~n3525 & n8124 ;
  assign n9436 = n5006 ^ n1347 ^ 1'b0 ;
  assign n9437 = n4879 | n9436 ;
  assign n9438 = n9437 ^ n8024 ^ 1'b0 ;
  assign n9439 = n9438 ^ n5262 ^ 1'b0 ;
  assign n9440 = x37 & ~n9439 ;
  assign n9441 = ( ~n6950 & n9435 ) | ( ~n6950 & n9440 ) | ( n9435 & n9440 ) ;
  assign n9442 = n8509 ^ n6524 ^ n1115 ;
  assign n9443 = n3296 | n9442 ;
  assign n9444 = n6970 & ~n9443 ;
  assign n9445 = n1757 | n3875 ;
  assign n9446 = n9445 ^ n5373 ^ 1'b0 ;
  assign n9447 = n1619 ^ n188 ^ 1'b0 ;
  assign n9448 = n9446 | n9447 ;
  assign n9449 = n3256 & n4107 ;
  assign n9459 = n3698 ^ n935 ^ 1'b0 ;
  assign n9456 = n4209 ^ x97 ^ 1'b0 ;
  assign n9457 = n9456 ^ n4502 ^ n1295 ;
  assign n9450 = n2212 & ~n2720 ;
  assign n9451 = n9450 ^ n1628 ^ n781 ;
  assign n9452 = n9451 ^ n7571 ^ 1'b0 ;
  assign n9453 = n4131 | n9452 ;
  assign n9454 = n9453 ^ n2432 ^ 1'b0 ;
  assign n9455 = n3191 | n9454 ;
  assign n9458 = n9457 ^ n9455 ^ 1'b0 ;
  assign n9460 = n9459 ^ n9458 ^ 1'b0 ;
  assign n9461 = ( n383 & n681 ) | ( n383 & ~n4006 ) | ( n681 & ~n4006 ) ;
  assign n9462 = n461 & ~n3618 ;
  assign n9463 = ~n9461 & n9462 ;
  assign n9464 = ( ~n777 & n1643 ) | ( ~n777 & n7716 ) | ( n1643 & n7716 ) ;
  assign n9465 = ~n571 & n858 ;
  assign n9466 = n9464 & n9465 ;
  assign n9467 = ( n1362 & ~n9141 ) | ( n1362 & n9466 ) | ( ~n9141 & n9466 ) ;
  assign n9468 = n316 & n1905 ;
  assign n9469 = n3345 | n9468 ;
  assign n9470 = n9469 ^ n5323 ^ 1'b0 ;
  assign n9471 = n7786 ^ n3110 ^ 1'b0 ;
  assign n9472 = ( n708 & n9470 ) | ( n708 & n9471 ) | ( n9470 & n9471 ) ;
  assign n9473 = n2103 & n2667 ;
  assign n9474 = ~n1684 & n9473 ;
  assign n9475 = ( n1559 & n6145 ) | ( n1559 & ~n9474 ) | ( n6145 & ~n9474 ) ;
  assign n9477 = ~n7521 & n7984 ;
  assign n9476 = n6008 ^ n5556 ^ 1'b0 ;
  assign n9478 = n9477 ^ n9476 ^ n1765 ;
  assign n9480 = n1432 & ~n3933 ;
  assign n9481 = ~n6709 & n9480 ;
  assign n9482 = n9481 ^ n245 ^ 1'b0 ;
  assign n9479 = n4651 & n5060 ;
  assign n9483 = n9482 ^ n9479 ^ 1'b0 ;
  assign n9485 = n2022 ^ n231 ^ 1'b0 ;
  assign n9484 = ( n4404 & ~n5654 ) | ( n4404 & n8218 ) | ( ~n5654 & n8218 ) ;
  assign n9486 = n9485 ^ n9484 ^ n355 ;
  assign n9487 = n6319 & n9486 ;
  assign n9488 = n3217 ^ n1200 ^ 1'b0 ;
  assign n9489 = n1565 & n9488 ;
  assign n9490 = n8653 & n9489 ;
  assign n9491 = ~n5990 & n9490 ;
  assign n9492 = n9273 & n9334 ;
  assign n9493 = n236 & n597 ;
  assign n9494 = n7513 ^ n4253 ^ 1'b0 ;
  assign n9495 = n4844 & ~n9494 ;
  assign n9496 = n8639 ^ n1427 ^ 1'b0 ;
  assign n9497 = n9496 ^ n6435 ^ 1'b0 ;
  assign n9498 = n674 & ~n4931 ;
  assign n9499 = n9498 ^ n4426 ^ 1'b0 ;
  assign n9500 = ~n1610 & n2623 ;
  assign n9501 = n9500 ^ n8143 ^ 1'b0 ;
  assign n9502 = n210 | n852 ;
  assign n9503 = n3641 | n6968 ;
  assign n9504 = n2590 & n7379 ;
  assign n9505 = ~n2933 & n9504 ;
  assign n9506 = n5106 ^ n529 ^ 1'b0 ;
  assign n9507 = ~n6893 & n9506 ;
  assign n9508 = n1380 & ~n8859 ;
  assign n9509 = ~n9507 & n9508 ;
  assign n9511 = ~n3350 & n5326 ;
  assign n9512 = n4503 | n9511 ;
  assign n9513 = n2312 | n9512 ;
  assign n9510 = ~n5957 & n8342 ;
  assign n9514 = n9513 ^ n9510 ^ 1'b0 ;
  assign n9515 = n6068 ^ n1364 ^ 1'b0 ;
  assign n9516 = n2940 & n9515 ;
  assign n9517 = ~n174 & n9200 ;
  assign n9518 = ~n4732 & n9517 ;
  assign n9519 = n373 | n3810 ;
  assign n9520 = ( n1526 & n6651 ) | ( n1526 & n9519 ) | ( n6651 & n9519 ) ;
  assign n9521 = ( n3245 & n5212 ) | ( n3245 & n6369 ) | ( n5212 & n6369 ) ;
  assign n9522 = n4027 ^ n496 ^ 1'b0 ;
  assign n9523 = n671 & n3556 ;
  assign n9524 = n9523 ^ n2062 ^ 1'b0 ;
  assign n9525 = n9524 ^ n2978 ^ 1'b0 ;
  assign n9526 = n7219 & ~n9525 ;
  assign n9527 = ~n4004 & n9526 ;
  assign n9528 = n9527 ^ n7927 ^ n4156 ;
  assign n9529 = ( n6483 & n9522 ) | ( n6483 & n9528 ) | ( n9522 & n9528 ) ;
  assign n9530 = n9478 ^ n2291 ^ 1'b0 ;
  assign n9531 = n3525 | n3688 ;
  assign n9532 = n3208 & ~n9531 ;
  assign n9533 = n4232 & ~n9532 ;
  assign n9534 = n9381 & n9533 ;
  assign n9535 = n1600 | n8412 ;
  assign n9536 = n4075 ^ n2805 ^ n1440 ;
  assign n9537 = ~n3735 & n4762 ;
  assign n9538 = n9537 ^ n1948 ^ 1'b0 ;
  assign n9539 = n1339 & ~n3814 ;
  assign n9540 = n9539 ^ n623 ^ 1'b0 ;
  assign n9541 = ~n422 & n9540 ;
  assign n9542 = n3896 ^ n707 ^ 1'b0 ;
  assign n9543 = n5993 ^ n2737 ^ 1'b0 ;
  assign n9544 = ~n3567 & n9543 ;
  assign n9545 = n1079 & n4362 ;
  assign n9546 = n767 & ~n9545 ;
  assign n9547 = ~n1829 & n7314 ;
  assign n9548 = n3244 & n9547 ;
  assign n9549 = n9548 ^ n2608 ^ 1'b0 ;
  assign n9550 = n4449 ^ n1589 ^ 1'b0 ;
  assign n9551 = ~n8169 & n9550 ;
  assign n9552 = ~n1753 & n5300 ;
  assign n9553 = ~n342 & n835 ;
  assign n9554 = n9553 ^ n150 ^ 1'b0 ;
  assign n9555 = n9554 ^ n7921 ^ 1'b0 ;
  assign n9556 = n8040 ^ n5396 ^ 1'b0 ;
  assign n9557 = n9390 | n9556 ;
  assign n9558 = n1195 ^ n673 ^ x119 ;
  assign n9559 = ( n3195 & n5509 ) | ( n3195 & ~n9558 ) | ( n5509 & ~n9558 ) ;
  assign n9560 = n9559 ^ n6023 ^ 1'b0 ;
  assign n9561 = n6856 ^ n891 ^ 1'b0 ;
  assign n9562 = n6808 & ~n9561 ;
  assign n9563 = n9562 ^ n1946 ^ 1'b0 ;
  assign n9564 = ~n7646 & n9563 ;
  assign n9565 = n3365 ^ n1903 ^ n1134 ;
  assign n9566 = n1390 & ~n6392 ;
  assign n9567 = n6878 ^ n579 ^ 1'b0 ;
  assign n9568 = n5771 ^ n2328 ^ 1'b0 ;
  assign n9569 = n3954 | n9568 ;
  assign n9570 = n5034 ^ n3918 ^ 1'b0 ;
  assign n9571 = ~n876 & n8424 ;
  assign n9572 = ~n8450 & n9571 ;
  assign n9573 = n5039 | n8278 ;
  assign n9574 = n7754 ^ n848 ^ 1'b0 ;
  assign n9575 = n9574 ^ n2770 ^ n1053 ;
  assign n9576 = n9575 ^ n3662 ^ 1'b0 ;
  assign n9577 = n4812 | n9576 ;
  assign n9578 = ~n673 & n9577 ;
  assign n9579 = n1309 | n4639 ;
  assign n9580 = n210 | n9579 ;
  assign n9581 = ~n5545 & n9580 ;
  assign n9582 = ~n9578 & n9581 ;
  assign n9583 = n742 ^ n713 ^ 1'b0 ;
  assign n9584 = n3617 | n9583 ;
  assign n9585 = n9584 ^ n6678 ^ 1'b0 ;
  assign n9586 = ~n4584 & n9585 ;
  assign n9587 = n8603 ^ x116 ^ 1'b0 ;
  assign n9588 = n521 | n8121 ;
  assign n9589 = n9587 | n9588 ;
  assign n9590 = x88 & n3480 ;
  assign n9591 = n9590 ^ n3561 ^ 1'b0 ;
  assign n9592 = ~n5415 & n9591 ;
  assign n9594 = n3706 & n6124 ;
  assign n9593 = n3861 & ~n4282 ;
  assign n9595 = n9594 ^ n9593 ^ n6647 ;
  assign n9596 = n1677 ^ n778 ^ n413 ;
  assign n9597 = n9596 ^ n3452 ^ 1'b0 ;
  assign n9598 = n6895 & ~n9597 ;
  assign n9599 = n4534 ^ n3955 ^ 1'b0 ;
  assign n9600 = n387 & n3684 ;
  assign n9601 = ~n9599 & n9600 ;
  assign n9602 = n9601 ^ n8692 ^ 1'b0 ;
  assign n9603 = n7284 & n9602 ;
  assign n9604 = n254 & ~n1094 ;
  assign n9605 = n7581 ^ n5741 ^ n5016 ;
  assign n9606 = n2186 & ~n9605 ;
  assign n9607 = ( ~x31 & n1432 ) | ( ~x31 & n3284 ) | ( n1432 & n3284 ) ;
  assign n9608 = n9402 | n9607 ;
  assign n9609 = n7953 ^ n4270 ^ 1'b0 ;
  assign n9610 = x74 & ~n9609 ;
  assign n9611 = n9610 ^ n3835 ^ n2053 ;
  assign n9612 = n6496 ^ n1356 ^ 1'b0 ;
  assign n9613 = n3666 ^ x97 ^ 1'b0 ;
  assign n9614 = n3994 & n8519 ;
  assign n9615 = n9052 & n9614 ;
  assign n9616 = ( ~n2283 & n5461 ) | ( ~n2283 & n6633 ) | ( n5461 & n6633 ) ;
  assign n9617 = ( n4532 & n5926 ) | ( n4532 & ~n7953 ) | ( n5926 & ~n7953 ) ;
  assign n9618 = n5548 ^ n2419 ^ 1'b0 ;
  assign n9619 = n9617 & n9618 ;
  assign n9620 = n1309 | n2549 ;
  assign n9621 = n3937 & ~n9620 ;
  assign n9622 = n5881 | n9621 ;
  assign n9623 = n9622 ^ n4303 ^ 1'b0 ;
  assign n9624 = n3755 & n5056 ;
  assign n9625 = n433 & ~n5834 ;
  assign n9626 = n2649 & n6473 ;
  assign n9627 = n9626 ^ n8390 ^ 1'b0 ;
  assign n9628 = ~n9625 & n9627 ;
  assign n9629 = n3684 ^ n2155 ^ 1'b0 ;
  assign n9630 = ~n2482 & n9629 ;
  assign n9631 = n9630 ^ n612 ^ 1'b0 ;
  assign n9632 = n8206 & n9631 ;
  assign n9633 = n5361 ^ n424 ^ 1'b0 ;
  assign n9634 = n9632 & n9633 ;
  assign n9635 = n2777 ^ n833 ^ n447 ;
  assign n9637 = n614 & n1463 ;
  assign n9638 = n4067 & n9637 ;
  assign n9639 = n4115 & n7200 ;
  assign n9640 = n5591 & n9639 ;
  assign n9641 = n9638 & n9640 ;
  assign n9636 = ( n1026 & ~n1578 ) | ( n1026 & n6273 ) | ( ~n1578 & n6273 ) ;
  assign n9642 = n9641 ^ n9636 ^ n4932 ;
  assign n9647 = n2313 | n8598 ;
  assign n9643 = ~n850 & n3304 ;
  assign n9644 = ~x3 & n9643 ;
  assign n9645 = ~n7801 & n9644 ;
  assign n9646 = n5947 & ~n9645 ;
  assign n9648 = n9647 ^ n9646 ^ 1'b0 ;
  assign n9649 = n2622 & ~n9645 ;
  assign n9650 = n9649 ^ n142 ^ 1'b0 ;
  assign n9651 = n9484 | n9650 ;
  assign n9656 = n2212 ^ n2109 ^ 1'b0 ;
  assign n9652 = n9007 ^ n1848 ^ 1'b0 ;
  assign n9653 = n1418 | n9652 ;
  assign n9654 = n2423 | n9653 ;
  assign n9655 = n6350 & ~n9654 ;
  assign n9657 = n9656 ^ n9655 ^ n4972 ;
  assign n9658 = n9657 ^ n6170 ^ n576 ;
  assign n9659 = ~n1030 & n5862 ;
  assign n9660 = ~n3070 & n9659 ;
  assign n9661 = ~n1766 & n9660 ;
  assign n9662 = n1703 & ~n9592 ;
  assign n9663 = ( ~n3036 & n5723 ) | ( ~n3036 & n6547 ) | ( n5723 & n6547 ) ;
  assign n9664 = n9663 ^ n9522 ^ 1'b0 ;
  assign n9665 = ~n6295 & n7481 ;
  assign n9666 = n9664 & n9665 ;
  assign n9667 = ( ~x47 & n1708 ) | ( ~x47 & n3547 ) | ( n1708 & n3547 ) ;
  assign n9668 = n9520 | n9667 ;
  assign n9669 = n5866 | n9668 ;
  assign n9670 = n1843 & n7905 ;
  assign n9671 = ~n2964 & n4597 ;
  assign n9672 = n7555 & n9671 ;
  assign n9673 = n9672 ^ n3906 ^ 1'b0 ;
  assign n9674 = n3223 & n9673 ;
  assign n9675 = n9670 & n9674 ;
  assign n9676 = n9675 ^ n3656 ^ 1'b0 ;
  assign n9677 = n8929 ^ n1918 ^ n306 ;
  assign n9678 = n9677 ^ n2647 ^ 1'b0 ;
  assign n9679 = ~n1970 & n9678 ;
  assign n9680 = n2710 ^ n363 ^ 1'b0 ;
  assign n9681 = n4052 & ~n9680 ;
  assign n9682 = n4305 ^ n2236 ^ 1'b0 ;
  assign n9683 = n2437 | n3247 ;
  assign n9684 = n9683 ^ n1339 ^ 1'b0 ;
  assign n9685 = ~n1668 & n9684 ;
  assign n9686 = ~n1333 & n9685 ;
  assign n9687 = ( n373 & n2912 ) | ( n373 & n9686 ) | ( n2912 & n9686 ) ;
  assign n9688 = n7243 ^ n3482 ^ 1'b0 ;
  assign n9689 = n9687 | n9688 ;
  assign n9690 = n1679 & ~n9689 ;
  assign n9691 = ~n5076 & n9690 ;
  assign n9692 = n5181 & n7201 ;
  assign n9693 = ~n442 & n890 ;
  assign n9694 = n1135 & n1321 ;
  assign n9695 = n8502 | n9694 ;
  assign n9696 = n9695 ^ n7872 ^ 1'b0 ;
  assign n9697 = n899 & n3065 ;
  assign n9698 = n4183 & n9697 ;
  assign n9699 = n9698 ^ n7595 ^ 1'b0 ;
  assign n9700 = n8548 | n9699 ;
  assign n9701 = n4639 | n8882 ;
  assign n9702 = n9701 ^ n6933 ^ 1'b0 ;
  assign n9703 = ( ~n3857 & n4293 ) | ( ~n3857 & n9702 ) | ( n4293 & n9702 ) ;
  assign n9704 = n9703 ^ n6569 ^ 1'b0 ;
  assign n9705 = n1527 & n7019 ;
  assign n9706 = n9705 ^ n7008 ^ 1'b0 ;
  assign n9707 = n176 & ~n8471 ;
  assign n9708 = n7160 ^ n3220 ^ n3151 ;
  assign n9709 = n9708 ^ n6515 ^ n2289 ;
  assign n9710 = n9709 ^ n1106 ^ 1'b0 ;
  assign n9711 = n6434 ^ n2970 ^ n2579 ;
  assign n9712 = n7978 & ~n8641 ;
  assign n9713 = ~n1445 & n9712 ;
  assign n9714 = n3934 | n8887 ;
  assign n9715 = ~n3484 & n7154 ;
  assign n9719 = n290 & ~n3626 ;
  assign n9716 = n4380 ^ n1462 ^ 1'b0 ;
  assign n9717 = n4419 & n9716 ;
  assign n9718 = n1652 & n9717 ;
  assign n9720 = n9719 ^ n9718 ^ 1'b0 ;
  assign n9721 = n5657 ^ n3446 ^ 1'b0 ;
  assign n9722 = n4123 | n9721 ;
  assign n9723 = n7784 ^ n5981 ^ 1'b0 ;
  assign n9724 = n9722 | n9723 ;
  assign n9725 = n5263 & ~n6408 ;
  assign n9726 = n9724 & n9725 ;
  assign n9727 = x69 & ~n9726 ;
  assign n9728 = n159 & n9727 ;
  assign n9729 = n1762 | n4087 ;
  assign n9730 = ( n2532 & ~n5734 ) | ( n2532 & n9729 ) | ( ~n5734 & n9729 ) ;
  assign n9731 = n2216 | n5431 ;
  assign n9732 = n324 | n8860 ;
  assign n9733 = n1511 & ~n9732 ;
  assign n9734 = n3672 ^ n606 ^ 1'b0 ;
  assign n9735 = ~n9733 & n9734 ;
  assign n9736 = ~n1171 & n2756 ;
  assign n9737 = n8455 ^ n8419 ^ n764 ;
  assign n9738 = n4548 & ~n4668 ;
  assign n9739 = ( n4313 & ~n9737 ) | ( n4313 & n9738 ) | ( ~n9737 & n9738 ) ;
  assign n9740 = n2012 & n3732 ;
  assign n9741 = n9740 ^ n5796 ^ 1'b0 ;
  assign n9743 = ( n161 & n595 ) | ( n161 & ~n5281 ) | ( n595 & ~n5281 ) ;
  assign n9742 = ~n1258 & n4625 ;
  assign n9744 = n9743 ^ n9742 ^ 1'b0 ;
  assign n9745 = n1990 | n3568 ;
  assign n9746 = n2275 & ~n9745 ;
  assign n9747 = ~n9141 & n9746 ;
  assign n9748 = ~n2912 & n9747 ;
  assign n9749 = n2579 | n4810 ;
  assign n9750 = n778 & n6979 ;
  assign n9751 = n1410 & n9750 ;
  assign n9752 = n9751 ^ n4543 ^ 1'b0 ;
  assign n9753 = x1 & n299 ;
  assign n9754 = n9753 ^ n5786 ^ 1'b0 ;
  assign n9755 = n9754 ^ n6846 ^ 1'b0 ;
  assign n9756 = n6876 | n9755 ;
  assign n9757 = n1423 | n4439 ;
  assign n9758 = n9757 ^ n4667 ^ 1'b0 ;
  assign n9759 = ( ~n8559 & n9756 ) | ( ~n8559 & n9758 ) | ( n9756 & n9758 ) ;
  assign n9760 = n879 | n5863 ;
  assign n9761 = n1599 | n3137 ;
  assign n9762 = n9760 & n9761 ;
  assign n9763 = n9762 ^ n4460 ^ 1'b0 ;
  assign n9764 = n5476 ^ n3134 ^ 1'b0 ;
  assign n9765 = n5194 ^ n3480 ^ 1'b0 ;
  assign n9770 = n2214 ^ n668 ^ 1'b0 ;
  assign n9771 = n1123 & n9770 ;
  assign n9772 = n1972 & n9771 ;
  assign n9773 = ~n7462 & n9772 ;
  assign n9769 = n1452 & n2310 ;
  assign n9774 = n9773 ^ n9769 ^ 1'b0 ;
  assign n9766 = ( n1413 & n3705 ) | ( n1413 & n5132 ) | ( n3705 & n5132 ) ;
  assign n9767 = n842 & ~n9766 ;
  assign n9768 = n9767 ^ n2638 ^ 1'b0 ;
  assign n9775 = n9774 ^ n9768 ^ n744 ;
  assign n9776 = n7146 ^ n5981 ^ 1'b0 ;
  assign n9777 = n2850 ^ n1080 ^ 1'b0 ;
  assign n9778 = ( n1765 & n5351 ) | ( n1765 & n7192 ) | ( n5351 & n7192 ) ;
  assign n9779 = ( n1552 & ~n9777 ) | ( n1552 & n9778 ) | ( ~n9777 & n9778 ) ;
  assign n9780 = n1352 & n7296 ;
  assign n9781 = n9780 ^ n3849 ^ 1'b0 ;
  assign n9782 = ~n9013 & n9524 ;
  assign n9783 = n7325 & n9782 ;
  assign n9784 = n9656 ^ n2841 ^ 1'b0 ;
  assign n9785 = ~n6526 & n9784 ;
  assign n9786 = ~n1421 & n7161 ;
  assign n9787 = n1286 | n9786 ;
  assign n9788 = n9787 ^ n1692 ^ 1'b0 ;
  assign n9789 = n4000 ^ n570 ^ 1'b0 ;
  assign n9790 = n2634 | n9789 ;
  assign n9791 = n9790 ^ n3011 ^ n135 ;
  assign n9792 = n750 & ~n3828 ;
  assign n9793 = ~n1533 & n9792 ;
  assign n9794 = n3176 ^ n1438 ^ 1'b0 ;
  assign n9795 = ~n4954 & n9794 ;
  assign n9796 = n9795 ^ n8110 ^ 1'b0 ;
  assign n9797 = n1630 & n8553 ;
  assign n9798 = ~n333 & n9702 ;
  assign n9799 = n9798 ^ n3153 ^ 1'b0 ;
  assign n9800 = ~n2447 & n9799 ;
  assign n9801 = ~n1384 & n9800 ;
  assign n9802 = n1384 & n9801 ;
  assign n9803 = ~n3149 & n5870 ;
  assign n9804 = n1582 | n4631 ;
  assign n9805 = n9803 & ~n9804 ;
  assign n9806 = n388 & ~n2447 ;
  assign n9807 = n6941 & n9806 ;
  assign n9808 = n6212 ^ n1306 ^ 1'b0 ;
  assign n9809 = n1023 | n9808 ;
  assign n9810 = n4653 ^ n1263 ^ 1'b0 ;
  assign n9811 = n2437 | n9810 ;
  assign n9812 = n9811 ^ n9088 ^ 1'b0 ;
  assign n9813 = n8576 | n9812 ;
  assign n9814 = n2289 & n8619 ;
  assign n9815 = n8523 ^ n1943 ^ 1'b0 ;
  assign n9816 = ~n5063 & n9815 ;
  assign n9817 = n9816 ^ n4725 ^ n1463 ;
  assign n9818 = n9467 ^ n8512 ^ n5945 ;
  assign n9819 = n5406 ^ n582 ^ 1'b0 ;
  assign n9820 = n3431 | n9819 ;
  assign n9821 = n9820 ^ n3295 ^ 1'b0 ;
  assign n9822 = n1841 ^ x5 ^ 1'b0 ;
  assign n9823 = ~n702 & n9822 ;
  assign n9824 = n9823 ^ n7094 ^ 1'b0 ;
  assign n9825 = n3929 & ~n9824 ;
  assign n9826 = ~n9821 & n9825 ;
  assign n9827 = n9826 ^ n9014 ^ 1'b0 ;
  assign n9828 = ~n2375 & n6162 ;
  assign n9829 = ~n3513 & n9828 ;
  assign n9830 = ~x57 & n9418 ;
  assign n9831 = n7608 ^ n3901 ^ 1'b0 ;
  assign n9832 = n9830 | n9831 ;
  assign n9833 = n3895 & ~n9832 ;
  assign n9834 = n9829 & n9833 ;
  assign n9835 = n2959 & n8229 ;
  assign n9836 = ~n2017 & n9835 ;
  assign n9837 = n3646 | n4327 ;
  assign n9838 = n1945 | n9837 ;
  assign n9839 = n1106 | n6784 ;
  assign n9840 = n6557 ^ n1559 ^ 1'b0 ;
  assign n9841 = n9840 ^ n4145 ^ n3067 ;
  assign n9842 = n9841 ^ n2495 ^ 1'b0 ;
  assign n9843 = ~n9839 & n9842 ;
  assign n9844 = x42 & n261 ;
  assign n9845 = ~x42 & n9844 ;
  assign n9846 = ~n2687 & n9845 ;
  assign n9847 = n1162 & n9846 ;
  assign n9848 = n1002 | n3308 ;
  assign n9849 = n3308 & ~n9848 ;
  assign n9850 = n9849 ^ n1025 ^ 1'b0 ;
  assign n9851 = n9847 | n9850 ;
  assign n9852 = n4118 & ~n9851 ;
  assign n9853 = n9852 ^ n3476 ^ 1'b0 ;
  assign n9854 = x62 & ~n3964 ;
  assign n9855 = n4108 ^ n1450 ^ 1'b0 ;
  assign n9856 = n4323 & ~n9855 ;
  assign n9857 = n2852 & ~n9856 ;
  assign n9858 = ( n9853 & n9854 ) | ( n9853 & n9857 ) | ( n9854 & n9857 ) ;
  assign n9859 = n2847 & ~n5682 ;
  assign n9860 = n5516 ^ n1085 ^ n671 ;
  assign n9861 = n9860 ^ n6787 ^ 1'b0 ;
  assign n9862 = n4670 & n9861 ;
  assign n9863 = n237 & ~n1003 ;
  assign n9864 = n9863 ^ n2132 ^ 1'b0 ;
  assign n9865 = n9862 & n9864 ;
  assign n9866 = n2112 ^ n925 ^ n471 ;
  assign n9867 = n9866 ^ n8249 ^ n1802 ;
  assign n9868 = n633 ^ n569 ^ 1'b0 ;
  assign n9869 = n2266 | n8200 ;
  assign n9870 = n9868 & ~n9869 ;
  assign n9872 = n3602 ^ n2829 ^ n828 ;
  assign n9871 = n196 | n8879 ;
  assign n9873 = n9872 ^ n9871 ^ 1'b0 ;
  assign n9879 = n1406 & n4295 ;
  assign n9880 = n9879 ^ n939 ^ 1'b0 ;
  assign n9874 = ( n739 & ~n1578 ) | ( n739 & n3678 ) | ( ~n1578 & n3678 ) ;
  assign n9875 = n1943 & n9874 ;
  assign n9876 = n1496 ^ n846 ^ 1'b0 ;
  assign n9877 = ~n9875 & n9876 ;
  assign n9878 = ~n293 & n9877 ;
  assign n9881 = n9880 ^ n9878 ^ 1'b0 ;
  assign n9882 = n4637 ^ n2552 ^ n1656 ;
  assign n9883 = ( n6225 & n8552 ) | ( n6225 & n9882 ) | ( n8552 & n9882 ) ;
  assign n9884 = n6257 ^ n2423 ^ 1'b0 ;
  assign n9885 = ~n5229 & n9884 ;
  assign n9886 = n8541 ^ n202 ^ 1'b0 ;
  assign n9887 = n3862 & n9886 ;
  assign n9888 = ~n5850 & n9887 ;
  assign n9889 = n234 & ~n7518 ;
  assign n9890 = n3753 & ~n9889 ;
  assign n9891 = n9555 ^ n6763 ^ n4996 ;
  assign n9892 = ( n210 & n9890 ) | ( n210 & n9891 ) | ( n9890 & n9891 ) ;
  assign n9893 = ~n786 & n3325 ;
  assign n9894 = n9893 ^ n8541 ^ 1'b0 ;
  assign n9895 = n1775 & n9894 ;
  assign n9896 = n9895 ^ n990 ^ 1'b0 ;
  assign n9897 = n3815 & n4048 ;
  assign n9898 = n7019 & ~n8962 ;
  assign n9899 = n5785 ^ n2673 ^ 1'b0 ;
  assign n9900 = n819 & ~n9899 ;
  assign n9901 = ~n3055 & n9900 ;
  assign n9902 = n1140 & n4405 ;
  assign n9903 = n202 & n4169 ;
  assign n9904 = n179 | n2990 ;
  assign n9905 = n7654 ^ n6801 ^ 1'b0 ;
  assign n9906 = n9904 | n9905 ;
  assign n9907 = ~n1746 & n7674 ;
  assign n9908 = n565 & n9907 ;
  assign n9909 = n7344 ^ x124 ^ 1'b0 ;
  assign n9910 = n2266 | n9909 ;
  assign n9911 = n9908 & n9910 ;
  assign n9912 = ~n9908 & n9911 ;
  assign n9913 = n9884 ^ n4811 ^ 1'b0 ;
  assign n9914 = n9913 ^ n8512 ^ n7974 ;
  assign n9915 = n411 | n5520 ;
  assign n9916 = x88 & ~n3666 ;
  assign n9917 = ~n4748 & n9916 ;
  assign n9918 = ~n969 & n9917 ;
  assign n9920 = n3626 | n6209 ;
  assign n9921 = n316 & ~n9920 ;
  assign n9919 = ( n1203 & ~n2408 ) | ( n1203 & n3482 ) | ( ~n2408 & n3482 ) ;
  assign n9922 = n9921 ^ n9919 ^ n9334 ;
  assign n9923 = n383 | n1855 ;
  assign n9924 = n8552 ^ n5827 ^ 1'b0 ;
  assign n9925 = n3179 & ~n9924 ;
  assign n9933 = x124 & n2253 ;
  assign n9931 = n1906 | n6844 ;
  assign n9932 = n3561 & n9931 ;
  assign n9934 = n9933 ^ n9932 ^ n3317 ;
  assign n9926 = n2826 & ~n5621 ;
  assign n9927 = n9926 ^ n1086 ^ 1'b0 ;
  assign n9928 = n1457 | n7844 ;
  assign n9929 = n9928 ^ n6015 ^ 1'b0 ;
  assign n9930 = ~n9927 & n9929 ;
  assign n9935 = n9934 ^ n9930 ^ 1'b0 ;
  assign n9936 = ( ~n7481 & n9925 ) | ( ~n7481 & n9935 ) | ( n9925 & n9935 ) ;
  assign n9937 = n9923 & ~n9936 ;
  assign n9938 = n2600 & ~n4208 ;
  assign n9939 = ~n1405 & n1940 ;
  assign n9940 = n3176 | n9939 ;
  assign n9941 = n9940 ^ n756 ^ 1'b0 ;
  assign n9942 = n9938 & n9941 ;
  assign n9943 = n4285 ^ n3371 ^ 1'b0 ;
  assign n9944 = n3265 & ~n5519 ;
  assign n9945 = ( n2934 & n3093 ) | ( n2934 & ~n9944 ) | ( n3093 & ~n9944 ) ;
  assign n9946 = n1627 & n9945 ;
  assign n9947 = n5091 & ~n6953 ;
  assign n9948 = n9947 ^ n8873 ^ n5365 ;
  assign n9950 = n3861 ^ n2461 ^ 1'b0 ;
  assign n9951 = ~n3547 & n9950 ;
  assign n9952 = n9951 ^ n4749 ^ 1'b0 ;
  assign n9953 = n299 & ~n9952 ;
  assign n9949 = n6689 ^ n2821 ^ 1'b0 ;
  assign n9954 = n9953 ^ n9949 ^ 1'b0 ;
  assign n9955 = n4842 ^ n2526 ^ 1'b0 ;
  assign n9956 = n4363 | n9955 ;
  assign n9957 = n9956 ^ n8144 ^ n4662 ;
  assign n9958 = n5901 & ~n9957 ;
  assign n9959 = n4921 ^ n2365 ^ 1'b0 ;
  assign n9960 = n3187 | n9959 ;
  assign n9961 = n5999 | n9960 ;
  assign n9962 = n9961 ^ n5380 ^ 1'b0 ;
  assign n9963 = ~n2291 & n4712 ;
  assign n9964 = n9963 ^ n3723 ^ 1'b0 ;
  assign n9965 = n2866 ^ n964 ^ 1'b0 ;
  assign n9966 = n9964 & n9965 ;
  assign n9967 = ~n7231 & n9966 ;
  assign n9968 = n9962 & n9967 ;
  assign n9969 = n4553 & ~n5420 ;
  assign n9970 = ~n1855 & n7668 ;
  assign n9971 = n9970 ^ n4863 ^ 1'b0 ;
  assign n9972 = ( n1795 & n3487 ) | ( n1795 & n9971 ) | ( n3487 & n9971 ) ;
  assign n9973 = ~n1226 & n9972 ;
  assign n9974 = n9973 ^ n2463 ^ 1'b0 ;
  assign n9978 = ~n3705 & n5834 ;
  assign n9979 = n2888 & n9978 ;
  assign n9980 = n3083 ^ n1832 ^ 1'b0 ;
  assign n9981 = ~n9979 & n9980 ;
  assign n9976 = n2368 ^ n1713 ^ 1'b0 ;
  assign n9977 = n8084 | n9976 ;
  assign n9975 = n9352 ^ n1459 ^ 1'b0 ;
  assign n9982 = n9981 ^ n9977 ^ n9975 ;
  assign n9983 = ( ~n193 & n513 ) | ( ~n193 & n7395 ) | ( n513 & n7395 ) ;
  assign n9984 = n7642 ^ n2306 ^ 1'b0 ;
  assign n9985 = n4366 | n9984 ;
  assign n9986 = n9985 ^ n7372 ^ n375 ;
  assign n9987 = n9952 ^ n2871 ^ n2498 ;
  assign n9988 = n7317 & n9987 ;
  assign n9989 = ~n4281 & n9988 ;
  assign n9990 = n636 & n8085 ;
  assign n9991 = ~n9989 & n9990 ;
  assign n9992 = n5739 | n8372 ;
  assign n9993 = n1265 & ~n8330 ;
  assign n9994 = n2656 | n4552 ;
  assign n9995 = n9993 | n9994 ;
  assign n9996 = n5352 ^ n379 ^ 1'b0 ;
  assign n9997 = n4796 | n9996 ;
  assign n9998 = n683 & ~n6339 ;
  assign n9999 = n9998 ^ n6183 ^ 1'b0 ;
  assign n10000 = ~n9997 & n9999 ;
  assign n10001 = ~n6122 & n10000 ;
  assign n10002 = n10001 ^ n9577 ^ n5948 ;
  assign n10003 = ~n835 & n1499 ;
  assign n10004 = n9376 ^ n1806 ^ 1'b0 ;
  assign n10005 = ~n8256 & n10004 ;
  assign n10006 = n4308 ^ n3558 ^ 1'b0 ;
  assign n10007 = n6701 ^ n221 ^ 1'b0 ;
  assign n10008 = n5063 | n10007 ;
  assign n10009 = n1368 | n10008 ;
  assign n10010 = n5577 & ~n10009 ;
  assign n10011 = n10010 ^ n5581 ^ 1'b0 ;
  assign n10012 = n9178 ^ n7170 ^ 1'b0 ;
  assign n10013 = n2608 | n10012 ;
  assign n10014 = n875 & ~n7445 ;
  assign n10015 = n3396 & n10014 ;
  assign n10016 = n3275 ^ n750 ^ 1'b0 ;
  assign n10019 = n2590 ^ n2299 ^ 1'b0 ;
  assign n10017 = n1791 & n4498 ;
  assign n10018 = ~n5248 & n10017 ;
  assign n10020 = n10019 ^ n10018 ^ 1'b0 ;
  assign n10021 = n2527 & n7956 ;
  assign n10022 = n6707 & n10021 ;
  assign n10023 = n7550 | n8816 ;
  assign n10026 = n3896 & n4300 ;
  assign n10027 = n1987 | n3307 ;
  assign n10028 = n10026 & ~n10027 ;
  assign n10029 = n10028 ^ n4033 ^ 1'b0 ;
  assign n10025 = n3003 & n3523 ;
  assign n10030 = n10029 ^ n10025 ^ 1'b0 ;
  assign n10031 = n10030 ^ n340 ^ 1'b0 ;
  assign n10032 = ~n5815 & n10031 ;
  assign n10024 = n4225 & ~n6421 ;
  assign n10033 = n10032 ^ n10024 ^ 1'b0 ;
  assign n10034 = n770 | n2540 ;
  assign n10035 = ~n2738 & n4131 ;
  assign n10036 = n7012 & ~n10035 ;
  assign n10037 = n5552 & n9543 ;
  assign n10038 = ~n345 & n10037 ;
  assign n10039 = n7099 | n10038 ;
  assign n10040 = ~n338 & n7025 ;
  assign n10042 = n643 & ~n1258 ;
  assign n10043 = n10042 ^ n4500 ^ 1'b0 ;
  assign n10044 = n4895 | n10043 ;
  assign n10045 = n7114 & ~n10044 ;
  assign n10041 = n5702 ^ n2647 ^ 1'b0 ;
  assign n10046 = n10045 ^ n10041 ^ n424 ;
  assign n10047 = n7656 & ~n7774 ;
  assign n10048 = ~x6 & n10047 ;
  assign n10049 = n5275 | n10048 ;
  assign n10050 = x13 | n10049 ;
  assign n10051 = n9917 ^ n3760 ^ 1'b0 ;
  assign n10052 = n5850 | n10051 ;
  assign n10053 = n8862 | n10052 ;
  assign n10054 = n10053 ^ n3228 ^ 1'b0 ;
  assign n10055 = n1356 & ~n10054 ;
  assign n10056 = n903 & n3783 ;
  assign n10057 = n3901 & n10056 ;
  assign n10058 = n3825 | n10057 ;
  assign n10059 = n10058 ^ n3128 ^ 1'b0 ;
  assign n10060 = n350 & ~n1971 ;
  assign n10061 = n1139 | n10060 ;
  assign n10062 = n3675 | n10061 ;
  assign n10063 = n3868 | n9941 ;
  assign n10064 = n4562 | n10063 ;
  assign n10065 = n1842 ^ n668 ^ 1'b0 ;
  assign n10066 = n740 | n10065 ;
  assign n10067 = n10066 ^ n884 ^ n141 ;
  assign n10068 = n1905 & ~n5266 ;
  assign n10069 = ( n1592 & n8163 ) | ( n1592 & n10068 ) | ( n8163 & n10068 ) ;
  assign n10070 = n1671 & ~n3148 ;
  assign n10071 = ~x4 & n10070 ;
  assign n10072 = n257 & n10071 ;
  assign n10073 = ( n1123 & ~n7083 ) | ( n1123 & n8343 ) | ( ~n7083 & n8343 ) ;
  assign n10074 = n8085 & n10073 ;
  assign n10075 = n5990 & ~n8919 ;
  assign n10076 = n1039 & n10075 ;
  assign n10077 = ( n2981 & n3786 ) | ( n2981 & ~n5074 ) | ( n3786 & ~n5074 ) ;
  assign n10078 = ~n5376 & n6977 ;
  assign n10079 = n1205 & ~n2341 ;
  assign n10080 = n10079 ^ n6501 ^ 1'b0 ;
  assign n10081 = n2175 | n4044 ;
  assign n10082 = n10081 ^ n2622 ^ 1'b0 ;
  assign n10085 = n130 & ~n6900 ;
  assign n10083 = n6145 ^ n5626 ^ 1'b0 ;
  assign n10084 = n7084 & n10083 ;
  assign n10086 = n10085 ^ n10084 ^ 1'b0 ;
  assign n10087 = n9484 | n10086 ;
  assign n10088 = n8200 ^ n3870 ^ 1'b0 ;
  assign n10089 = n6000 & n8177 ;
  assign n10090 = n8140 ^ x16 ^ 1'b0 ;
  assign n10091 = n7217 & n10090 ;
  assign n10092 = ( n1843 & n10089 ) | ( n1843 & n10091 ) | ( n10089 & n10091 ) ;
  assign n10093 = ~n2167 & n3245 ;
  assign n10094 = n10093 ^ n3476 ^ 1'b0 ;
  assign n10095 = n10094 ^ n5296 ^ 1'b0 ;
  assign n10096 = ( n694 & n848 ) | ( n694 & n8253 ) | ( n848 & n8253 ) ;
  assign n10097 = n10095 & ~n10096 ;
  assign n10098 = ~n5586 & n5806 ;
  assign n10099 = ~n4912 & n10098 ;
  assign n10100 = ( n2581 & n10097 ) | ( n2581 & ~n10099 ) | ( n10097 & ~n10099 ) ;
  assign n10101 = n2886 ^ n2229 ^ 1'b0 ;
  assign n10103 = n1826 ^ n612 ^ 1'b0 ;
  assign n10104 = x11 & ~n10103 ;
  assign n10105 = n10104 ^ n353 ^ 1'b0 ;
  assign n10106 = n1619 | n10105 ;
  assign n10102 = n8196 & ~n8327 ;
  assign n10107 = n10106 ^ n10102 ^ 1'b0 ;
  assign n10108 = n10107 ^ n1150 ^ 1'b0 ;
  assign n10109 = n4642 ^ n391 ^ 1'b0 ;
  assign n10110 = n202 & ~n10109 ;
  assign n10111 = n1764 ^ n1687 ^ n1147 ;
  assign n10112 = n10111 ^ n2634 ^ 1'b0 ;
  assign n10113 = ~n4788 & n10112 ;
  assign n10114 = n636 & ~n10113 ;
  assign n10115 = n1521 | n1654 ;
  assign n10116 = n1654 & ~n10115 ;
  assign n10117 = n1193 | n10116 ;
  assign n10118 = n1193 & ~n10117 ;
  assign n10119 = n6787 | n10118 ;
  assign n10120 = n6787 & ~n10119 ;
  assign n10121 = ~n1033 & n3593 ;
  assign n10122 = n8773 ^ n3434 ^ 1'b0 ;
  assign n10123 = n10121 & ~n10122 ;
  assign n10124 = ~n4858 & n7023 ;
  assign n10125 = n10124 ^ n8960 ^ 1'b0 ;
  assign n10126 = n4487 ^ n4285 ^ 1'b0 ;
  assign n10127 = n10126 ^ n3840 ^ 1'b0 ;
  assign n10128 = n4768 & n9064 ;
  assign n10129 = ~n3990 & n10128 ;
  assign n10130 = n4250 | n9694 ;
  assign n10131 = n10130 ^ n2426 ^ 1'b0 ;
  assign n10132 = n8351 ^ n3385 ^ 1'b0 ;
  assign n10133 = n3719 ^ n3557 ^ 1'b0 ;
  assign n10134 = n1220 & n10133 ;
  assign n10135 = n3738 & n10134 ;
  assign n10136 = n9927 & n10135 ;
  assign n10137 = ( n896 & ~n6117 ) | ( n896 & n10136 ) | ( ~n6117 & n10136 ) ;
  assign n10138 = ( n4785 & n5402 ) | ( n4785 & n7784 ) | ( n5402 & n7784 ) ;
  assign n10139 = n6046 & ~n10138 ;
  assign n10140 = n3536 ^ n920 ^ 1'b0 ;
  assign n10141 = n8210 ^ n4313 ^ 1'b0 ;
  assign n10142 = n10140 & ~n10141 ;
  assign n10143 = n7906 | n9273 ;
  assign n10144 = ~n4106 & n5678 ;
  assign n10145 = ~n10143 & n10144 ;
  assign n10146 = n5661 ^ n1418 ^ 1'b0 ;
  assign n10147 = n129 & ~n10146 ;
  assign n10148 = ~n6386 & n10147 ;
  assign n10149 = n1757 | n9096 ;
  assign n10150 = n10149 ^ n1686 ^ 1'b0 ;
  assign n10151 = n10150 ^ n259 ^ 1'b0 ;
  assign n10152 = n309 & ~n10151 ;
  assign n10153 = n2461 & n2571 ;
  assign n10154 = n10153 ^ n4653 ^ x30 ;
  assign n10155 = n1575 & ~n2317 ;
  assign n10156 = ~x16 & n10155 ;
  assign n10157 = n10156 ^ n2386 ^ 1'b0 ;
  assign n10158 = n863 & n10157 ;
  assign n10159 = n579 | n9149 ;
  assign n10160 = n5123 & ~n10159 ;
  assign n10161 = ( ~n5084 & n5841 ) | ( ~n5084 & n10160 ) | ( n5841 & n10160 ) ;
  assign n10162 = ( ~n1053 & n10158 ) | ( ~n1053 & n10161 ) | ( n10158 & n10161 ) ;
  assign n10163 = ~n6132 & n7972 ;
  assign n10164 = n1288 & n10163 ;
  assign n10165 = n3977 & n6041 ;
  assign n10166 = n10165 ^ n8086 ^ 1'b0 ;
  assign n10167 = n6738 & ~n7086 ;
  assign n10168 = n10167 ^ n6847 ^ n4923 ;
  assign n10169 = n6527 ^ n1085 ^ 1'b0 ;
  assign n10170 = n8279 | n10169 ;
  assign n10171 = n10170 ^ n9216 ^ 1'b0 ;
  assign n10172 = n7637 & n10171 ;
  assign n10173 = n3441 ^ n530 ^ 1'b0 ;
  assign n10174 = n167 | n1196 ;
  assign n10175 = n10173 & ~n10174 ;
  assign n10176 = n10175 ^ n6223 ^ 1'b0 ;
  assign n10177 = n6896 ^ n6657 ^ 1'b0 ;
  assign n10178 = n3759 & n10177 ;
  assign n10179 = n9710 ^ n6532 ^ 1'b0 ;
  assign n10180 = ~n606 & n8674 ;
  assign n10181 = n1794 & n8443 ;
  assign n10182 = ~n4870 & n5353 ;
  assign n10183 = n10181 & n10182 ;
  assign n10184 = n10183 ^ x110 ^ 1'b0 ;
  assign n10185 = ( ~n1079 & n2208 ) | ( ~n1079 & n7123 ) | ( n2208 & n7123 ) ;
  assign n10186 = n3915 ^ n2833 ^ 1'b0 ;
  assign n10187 = ~n2104 & n10186 ;
  assign n10188 = ~n8938 & n10187 ;
  assign n10189 = n3202 ^ n3067 ^ 1'b0 ;
  assign n10190 = n6786 & n10189 ;
  assign n10191 = ~n10188 & n10190 ;
  assign n10192 = ~n10185 & n10191 ;
  assign n10193 = ~n1286 & n3753 ;
  assign n10194 = n10193 ^ n852 ^ 1'b0 ;
  assign n10195 = ~n3433 & n4479 ;
  assign n10196 = n10194 | n10195 ;
  assign n10197 = n2560 | n6308 ;
  assign n10198 = n3471 | n10197 ;
  assign n10199 = n10198 ^ n3448 ^ n1687 ;
  assign n10200 = n777 & n2354 ;
  assign n10201 = n10200 ^ n1785 ^ 1'b0 ;
  assign n10202 = n8121 | n10201 ;
  assign n10203 = n10202 ^ n4658 ^ 1'b0 ;
  assign n10204 = n4565 & n10203 ;
  assign n10205 = ( n3418 & n4011 ) | ( n3418 & n4402 ) | ( n4011 & n4402 ) ;
  assign n10206 = n1924 & ~n7231 ;
  assign n10208 = n6972 & n9072 ;
  assign n10207 = n5433 & n8504 ;
  assign n10209 = n10208 ^ n10207 ^ 1'b0 ;
  assign n10210 = n1459 | n4587 ;
  assign n10211 = n240 | n10210 ;
  assign n10212 = n9639 | n10211 ;
  assign n10213 = n6306 ^ n2621 ^ 1'b0 ;
  assign n10214 = n651 | n10213 ;
  assign n10215 = n3001 & ~n4285 ;
  assign n10216 = n7222 ^ n6050 ^ n3794 ;
  assign n10217 = ( n1256 & n7553 ) | ( n1256 & ~n10216 ) | ( n7553 & ~n10216 ) ;
  assign n10218 = n4574 & ~n9975 ;
  assign n10219 = n4667 & n4749 ;
  assign n10220 = n1581 & ~n10219 ;
  assign n10221 = n10220 ^ n4578 ^ 1'b0 ;
  assign n10222 = n10221 ^ n3265 ^ 1'b0 ;
  assign n10223 = x106 & ~n10222 ;
  assign n10224 = n3474 ^ n182 ^ 1'b0 ;
  assign n10225 = n10224 ^ n7672 ^ 1'b0 ;
  assign n10226 = ( x2 & n431 ) | ( x2 & n2888 ) | ( n431 & n2888 ) ;
  assign n10229 = n1991 ^ n1532 ^ 1'b0 ;
  assign n10227 = n9294 ^ x116 ^ 1'b0 ;
  assign n10228 = n1821 & n10227 ;
  assign n10230 = n10229 ^ n10228 ^ 1'b0 ;
  assign n10231 = n10226 & ~n10230 ;
  assign n10232 = n132 & ~n2138 ;
  assign n10233 = n1094 ^ x3 ^ 1'b0 ;
  assign n10234 = n10233 ^ n8639 ^ 1'b0 ;
  assign n10235 = n5213 ^ n4681 ^ 1'b0 ;
  assign n10236 = n9422 | n10235 ;
  assign n10237 = ~n2642 & n9029 ;
  assign n10238 = n10237 ^ n7914 ^ 1'b0 ;
  assign n10239 = n7974 | n10238 ;
  assign n10240 = n564 & n5717 ;
  assign n10241 = n4668 ^ n3326 ^ 1'b0 ;
  assign n10242 = ( n2631 & n5431 ) | ( n2631 & n10241 ) | ( n5431 & n10241 ) ;
  assign n10243 = n5326 ^ n3264 ^ 1'b0 ;
  assign n10244 = n950 & n10243 ;
  assign n10245 = n10244 ^ n6708 ^ n835 ;
  assign n10246 = n2450 ^ n299 ^ 1'b0 ;
  assign n10247 = n2052 & n4705 ;
  assign n10248 = ~n6243 & n10247 ;
  assign n10249 = n10248 ^ n3299 ^ 1'b0 ;
  assign n10250 = n10246 & n10249 ;
  assign n10251 = n5693 ^ n762 ^ 1'b0 ;
  assign n10252 = n7530 & n10251 ;
  assign n10253 = n10252 ^ n471 ^ 1'b0 ;
  assign n10254 = n5796 ^ n3994 ^ n1505 ;
  assign n10255 = n10254 ^ n6521 ^ 1'b0 ;
  assign n10256 = n1048 & ~n2962 ;
  assign n10257 = ( ~n3991 & n4745 ) | ( ~n3991 & n10256 ) | ( n4745 & n10256 ) ;
  assign n10258 = n508 ^ n407 ^ 1'b0 ;
  assign n10259 = ~n1033 & n10258 ;
  assign n10260 = n10259 ^ n9904 ^ 1'b0 ;
  assign n10261 = ~n10257 & n10260 ;
  assign n10262 = n312 | n5519 ;
  assign n10263 = n10262 ^ n6139 ^ n1267 ;
  assign n10264 = n2409 ^ n145 ^ 1'b0 ;
  assign n10265 = n1736 & n10264 ;
  assign n10266 = n2760 & ~n5736 ;
  assign n10267 = ( n9719 & n10265 ) | ( n9719 & n10266 ) | ( n10265 & n10266 ) ;
  assign n10268 = n9352 ^ n2441 ^ 1'b0 ;
  assign n10269 = n3153 ^ n234 ^ 1'b0 ;
  assign n10270 = n6959 | n10269 ;
  assign n10271 = ( n959 & ~n1329 ) | ( n959 & n9632 ) | ( ~n1329 & n9632 ) ;
  assign n10272 = n3578 ^ n499 ^ 1'b0 ;
  assign n10273 = n10272 ^ n10188 ^ n1371 ;
  assign n10274 = n1526 | n10273 ;
  assign n10275 = n10274 ^ n6849 ^ 1'b0 ;
  assign n10276 = n2672 ^ n1479 ^ 1'b0 ;
  assign n10277 = n892 & ~n10276 ;
  assign n10278 = n1626 & n4770 ;
  assign n10279 = ~n10277 & n10278 ;
  assign n10280 = n2152 & n5515 ;
  assign n10281 = n10279 & n10280 ;
  assign n10282 = n5697 | n10281 ;
  assign n10283 = ~n4462 & n6020 ;
  assign n10284 = n10282 | n10283 ;
  assign n10285 = n10284 ^ n3148 ^ 1'b0 ;
  assign n10286 = n4580 | n10285 ;
  assign n10287 = n8059 ^ n5796 ^ 1'b0 ;
  assign n10288 = n10246 & ~n10287 ;
  assign n10289 = n10288 ^ n1029 ^ 1'b0 ;
  assign n10292 = n1760 & n2476 ;
  assign n10293 = n10292 ^ n1309 ^ 1'b0 ;
  assign n10290 = n1884 & ~n3057 ;
  assign n10291 = n3206 & n10290 ;
  assign n10294 = n10293 ^ n10291 ^ 1'b0 ;
  assign n10295 = n615 & ~n4298 ;
  assign n10296 = ( n3424 & n6094 ) | ( n3424 & n10295 ) | ( n6094 & n10295 ) ;
  assign n10297 = n10296 ^ n10019 ^ n5993 ;
  assign n10299 = n5659 | n9141 ;
  assign n10300 = n10299 ^ n3986 ^ 1'b0 ;
  assign n10298 = n7916 ^ n3053 ^ n1095 ;
  assign n10301 = n10300 ^ n10298 ^ 1'b0 ;
  assign n10305 = ( n1435 & n3476 ) | ( n1435 & ~n3658 ) | ( n3476 & ~n3658 ) ;
  assign n10304 = n6308 | n8676 ;
  assign n10306 = n10305 ^ n10304 ^ 1'b0 ;
  assign n10303 = n194 & ~n5437 ;
  assign n10307 = n10306 ^ n10303 ^ 1'b0 ;
  assign n10302 = n8573 & n9702 ;
  assign n10308 = n10307 ^ n10302 ^ 1'b0 ;
  assign n10309 = n6162 & n10170 ;
  assign n10310 = n3461 | n6217 ;
  assign n10311 = n4500 | n10310 ;
  assign n10312 = n1139 ^ n1113 ^ n856 ;
  assign n10313 = n10312 ^ n5211 ^ 1'b0 ;
  assign n10314 = ~n1248 & n3497 ;
  assign n10315 = n1038 & n10314 ;
  assign n10316 = n2710 & ~n10315 ;
  assign n10317 = n10316 ^ n6891 ^ 1'b0 ;
  assign n10318 = n375 | n403 ;
  assign n10319 = ~n6855 & n10318 ;
  assign n10320 = ~n10317 & n10319 ;
  assign n10321 = n805 & n8915 ;
  assign n10322 = n3401 | n8559 ;
  assign n10323 = n4082 | n10322 ;
  assign n10324 = n1594 & n2249 ;
  assign n10325 = n8106 | n10324 ;
  assign n10326 = n6135 ^ n2393 ^ 1'b0 ;
  assign n10327 = ~n5211 & n8966 ;
  assign n10328 = ~n1250 & n4032 ;
  assign n10329 = n4268 & n10328 ;
  assign n10330 = n10329 ^ n4691 ^ 1'b0 ;
  assign n10331 = ~n8774 & n9321 ;
  assign n10332 = ~n1374 & n1664 ;
  assign n10333 = n1981 & n10332 ;
  assign n10334 = n7388 ^ n5461 ^ 1'b0 ;
  assign n10335 = n10333 & ~n10334 ;
  assign n10336 = ( n4565 & n10331 ) | ( n4565 & ~n10335 ) | ( n10331 & ~n10335 ) ;
  assign n10337 = n10229 ^ n3468 ^ 1'b0 ;
  assign n10339 = n1938 & n2019 ;
  assign n10340 = n10339 ^ n9323 ^ n7723 ;
  assign n10338 = n2809 & ~n6435 ;
  assign n10341 = n10340 ^ n10338 ^ 1'b0 ;
  assign n10342 = n678 & n1679 ;
  assign n10343 = n2376 & n10342 ;
  assign n10344 = n3330 & ~n3342 ;
  assign n10345 = n6052 & n10344 ;
  assign n10346 = n1798 & ~n3998 ;
  assign n10347 = n10345 & n10346 ;
  assign n10348 = ( ~n2693 & n2878 ) | ( ~n2693 & n8512 ) | ( n2878 & n8512 ) ;
  assign n10349 = n10348 ^ n9283 ^ 1'b0 ;
  assign n10350 = ~n10347 & n10349 ;
  assign n10351 = n4983 | n5417 ;
  assign n10352 = n10351 ^ n6868 ^ 1'b0 ;
  assign n10353 = n4428 & ~n5702 ;
  assign n10354 = n1010 & n2823 ;
  assign n10355 = n2333 & n10354 ;
  assign n10356 = n5040 ^ n2642 ^ 1'b0 ;
  assign n10357 = ( ~n2152 & n10355 ) | ( ~n2152 & n10356 ) | ( n10355 & n10356 ) ;
  assign n10358 = n10353 | n10357 ;
  assign n10359 = n3435 & ~n10358 ;
  assign n10360 = n10359 ^ n7352 ^ 1'b0 ;
  assign n10361 = n8586 | n10360 ;
  assign n10362 = n2596 ^ n1565 ^ 1'b0 ;
  assign n10363 = n3755 | n10362 ;
  assign n10364 = n3213 & n9323 ;
  assign n10365 = ~n10363 & n10364 ;
  assign n10366 = n10365 ^ n138 ^ 1'b0 ;
  assign n10369 = n3064 ^ n194 ^ 1'b0 ;
  assign n10370 = n7004 & ~n10369 ;
  assign n10367 = n1928 | n3814 ;
  assign n10368 = n8481 & ~n10367 ;
  assign n10371 = n10370 ^ n10368 ^ 1'b0 ;
  assign n10372 = n4219 | n10371 ;
  assign n10373 = n2321 & n8287 ;
  assign n10374 = ( n1425 & ~n2503 ) | ( n1425 & n3315 ) | ( ~n2503 & n3315 ) ;
  assign n10375 = n10374 ^ n6539 ^ n3383 ;
  assign n10376 = ( n5255 & ~n7388 ) | ( n5255 & n10375 ) | ( ~n7388 & n10375 ) ;
  assign n10377 = n6149 ^ n4239 ^ 1'b0 ;
  assign n10378 = n3107 & ~n10377 ;
  assign n10379 = n8643 & ~n10378 ;
  assign n10380 = n901 & ~n6269 ;
  assign n10381 = n9963 & n10380 ;
  assign n10382 = n6558 & n8733 ;
  assign n10383 = n10381 & n10382 ;
  assign n10384 = n6170 ^ n778 ^ 1'b0 ;
  assign n10385 = n5963 | n10384 ;
  assign n10386 = n2711 & ~n3448 ;
  assign n10387 = ~n1828 & n10386 ;
  assign n10388 = ( n462 & ~n4720 ) | ( n462 & n10387 ) | ( ~n4720 & n10387 ) ;
  assign n10389 = n8584 ^ n5448 ^ 1'b0 ;
  assign n10390 = ~n7345 & n9694 ;
  assign n10391 = n1324 & ~n8516 ;
  assign n10392 = n6312 & n10391 ;
  assign n10393 = n8563 ^ n6815 ^ 1'b0 ;
  assign n10394 = n9069 ^ n1944 ^ 1'b0 ;
  assign n10395 = n683 ^ n652 ^ 1'b0 ;
  assign n10396 = n10395 ^ n1286 ^ 1'b0 ;
  assign n10397 = n5223 & ~n10396 ;
  assign n10398 = n987 & ~n5156 ;
  assign n10399 = n10398 ^ n4535 ^ 1'b0 ;
  assign n10400 = n10397 | n10399 ;
  assign n10401 = n3108 & ~n6310 ;
  assign n10402 = ( n840 & n1034 ) | ( n840 & n6339 ) | ( n1034 & n6339 ) ;
  assign n10403 = n2166 & ~n8863 ;
  assign n10404 = n10403 ^ n9489 ^ 1'b0 ;
  assign n10412 = n512 | n4509 ;
  assign n10405 = n1380 & ~n5641 ;
  assign n10406 = n5641 & n10405 ;
  assign n10407 = ~n2064 & n10406 ;
  assign n10408 = n3240 & n3243 ;
  assign n10409 = ~n3240 & n10408 ;
  assign n10410 = n4759 | n10409 ;
  assign n10411 = n10407 & ~n10410 ;
  assign n10413 = n10412 ^ n10411 ^ 1'b0 ;
  assign n10414 = ( n1286 & n2994 ) | ( n1286 & ~n5927 ) | ( n2994 & ~n5927 ) ;
  assign n10415 = n2109 ^ n846 ^ 1'b0 ;
  assign n10416 = ~n1366 & n5773 ;
  assign n10417 = n7569 ^ n6811 ^ 1'b0 ;
  assign n10418 = n1775 & n10417 ;
  assign n10419 = n3389 & n10418 ;
  assign n10420 = ~n616 & n9907 ;
  assign n10421 = n5878 ^ n5758 ^ 1'b0 ;
  assign n10422 = n370 & ~n2801 ;
  assign n10423 = ~n326 & n10422 ;
  assign n10424 = n10423 ^ n3415 ^ 1'b0 ;
  assign n10425 = n1374 | n6049 ;
  assign n10426 = n10425 ^ n303 ^ 1'b0 ;
  assign n10427 = n416 & ~n10426 ;
  assign n10428 = n10427 ^ n977 ^ 1'b0 ;
  assign n10429 = n10428 ^ n9489 ^ 1'b0 ;
  assign n10430 = ~n10424 & n10429 ;
  assign n10431 = n10430 ^ n3413 ^ 1'b0 ;
  assign n10432 = ~n7547 & n10431 ;
  assign n10433 = n7275 ^ n7269 ^ 1'b0 ;
  assign n10434 = ~n4845 & n10433 ;
  assign n10435 = n1765 & ~n10434 ;
  assign n10436 = n6849 & ~n8055 ;
  assign n10439 = n8948 ^ n4221 ^ 1'b0 ;
  assign n10437 = n2606 | n5031 ;
  assign n10438 = n10437 ^ n4509 ^ 1'b0 ;
  assign n10440 = n10439 ^ n10438 ^ 1'b0 ;
  assign n10441 = n3396 | n5132 ;
  assign n10442 = n10441 ^ n3608 ^ 1'b0 ;
  assign n10443 = n10442 ^ n4637 ^ 1'b0 ;
  assign n10444 = ~n6005 & n10443 ;
  assign n10448 = n3802 ^ n425 ^ 1'b0 ;
  assign n10445 = n1796 ^ n612 ^ 1'b0 ;
  assign n10446 = ( n8389 & ~n10134 ) | ( n8389 & n10445 ) | ( ~n10134 & n10445 ) ;
  assign n10447 = ~n5459 & n10446 ;
  assign n10449 = n10448 ^ n10447 ^ 1'b0 ;
  assign n10450 = ~n5077 & n9067 ;
  assign n10451 = n10450 ^ n2248 ^ 1'b0 ;
  assign n10452 = ( n712 & n1608 ) | ( n712 & ~n5662 ) | ( n1608 & ~n5662 ) ;
  assign n10453 = n10452 ^ n6922 ^ n4303 ;
  assign n10454 = n264 & n4029 ;
  assign n10455 = n10454 ^ n7451 ^ n6353 ;
  assign n10456 = n4853 ^ n2608 ^ 1'b0 ;
  assign n10457 = n672 & n10456 ;
  assign n10458 = n4456 & n10457 ;
  assign n10459 = ( n6958 & n9797 ) | ( n6958 & n10458 ) | ( n9797 & n10458 ) ;
  assign n10460 = n7116 ^ n3649 ^ n1586 ;
  assign n10461 = n10460 ^ n2187 ^ 1'b0 ;
  assign n10462 = n9156 ^ n6012 ^ 1'b0 ;
  assign n10463 = n10461 | n10462 ;
  assign n10464 = n7204 & ~n8086 ;
  assign n10465 = n8823 ^ n5129 ^ 1'b0 ;
  assign n10466 = n488 & ~n10465 ;
  assign n10467 = n10466 ^ n7573 ^ 1'b0 ;
  assign n10468 = n9528 ^ n8818 ^ 1'b0 ;
  assign n10469 = n3794 | n7829 ;
  assign n10470 = ~n997 & n10469 ;
  assign n10471 = n9446 ^ n5554 ^ 1'b0 ;
  assign n10472 = n9133 ^ n5437 ^ x3 ;
  assign n10473 = ~n10471 & n10472 ;
  assign n10474 = n6241 ^ n1130 ^ 1'b0 ;
  assign n10475 = n10473 | n10474 ;
  assign n10476 = n1633 ^ n1286 ^ 1'b0 ;
  assign n10477 = n10476 ^ n6633 ^ 1'b0 ;
  assign n10478 = n9754 ^ n5061 ^ 1'b0 ;
  assign n10479 = n10477 | n10478 ;
  assign n10480 = n5096 ^ n1212 ^ 1'b0 ;
  assign n10481 = n1123 & n10480 ;
  assign n10482 = n10481 ^ n775 ^ n265 ;
  assign n10483 = n1875 & n10482 ;
  assign n10484 = n7506 ^ n2322 ^ 1'b0 ;
  assign n10485 = n10484 ^ n5517 ^ 1'b0 ;
  assign n10486 = n6701 & ~n10485 ;
  assign n10487 = n2318 | n6578 ;
  assign n10488 = n2419 ^ n1136 ^ 1'b0 ;
  assign n10489 = n6884 ^ n3367 ^ 1'b0 ;
  assign n10490 = n9011 & n10489 ;
  assign n10491 = n8437 ^ n4758 ^ 1'b0 ;
  assign n10492 = n4081 & n10491 ;
  assign n10493 = n9074 & n10492 ;
  assign n10494 = ( n1680 & ~n2853 ) | ( n1680 & n3297 ) | ( ~n2853 & n3297 ) ;
  assign n10495 = n1694 & ~n10494 ;
  assign n10496 = ~n4238 & n10495 ;
  assign n10497 = ~n8006 & n10496 ;
  assign n10498 = n3755 ^ n2038 ^ n1629 ;
  assign n10499 = n557 & ~n10498 ;
  assign n10500 = ( n2560 & ~n8922 ) | ( n2560 & n10499 ) | ( ~n8922 & n10499 ) ;
  assign n10501 = n10500 ^ n9131 ^ 1'b0 ;
  assign n10502 = n1714 & ~n10281 ;
  assign n10503 = n1040 & n7796 ;
  assign n10504 = n970 & n10503 ;
  assign n10505 = ( n7727 & n9039 ) | ( n7727 & ~n10504 ) | ( n9039 & ~n10504 ) ;
  assign n10506 = n10505 ^ n5785 ^ 1'b0 ;
  assign n10507 = n2500 & ~n6159 ;
  assign n10508 = ~x2 & n4460 ;
  assign n10509 = n1172 & n1892 ;
  assign n10510 = ~n3339 & n6126 ;
  assign n10511 = n10510 ^ n2906 ^ 1'b0 ;
  assign n10512 = n10018 ^ n4903 ^ 1'b0 ;
  assign n10513 = ~n8818 & n10512 ;
  assign n10514 = n7113 & n7882 ;
  assign n10515 = ~n10513 & n10514 ;
  assign n10516 = ~n1448 & n2041 ;
  assign n10517 = ~n5933 & n10516 ;
  assign n10518 = n9413 & ~n10517 ;
  assign n10519 = n10518 ^ n6870 ^ 1'b0 ;
  assign n10520 = n2019 & ~n9396 ;
  assign n10521 = n10520 ^ n8681 ^ 1'b0 ;
  assign n10522 = n5327 ^ n3014 ^ 1'b0 ;
  assign n10523 = n10522 ^ n909 ^ 1'b0 ;
  assign n10524 = x18 & ~n6821 ;
  assign n10525 = n4211 ^ n871 ^ 1'b0 ;
  assign n10526 = n4209 ^ n1654 ^ 1'b0 ;
  assign n10527 = ~n1517 & n1803 ;
  assign n10528 = n10526 & n10527 ;
  assign n10529 = n10525 | n10528 ;
  assign n10530 = n10529 ^ n8707 ^ 1'b0 ;
  assign n10531 = n10530 ^ n463 ^ 1'b0 ;
  assign n10532 = n1927 & n4942 ;
  assign n10533 = ~n3349 & n10532 ;
  assign n10534 = x121 & ~n3563 ;
  assign n10535 = n10534 ^ n10188 ^ 1'b0 ;
  assign n10536 = n5256 ^ n615 ^ 1'b0 ;
  assign n10537 = n6141 | n10536 ;
  assign n10538 = n6327 ^ n4333 ^ 1'b0 ;
  assign n10539 = n750 & ~n7251 ;
  assign n10540 = n10539 ^ n7440 ^ 1'b0 ;
  assign n10541 = n3277 & n8190 ;
  assign n10542 = ~n5783 & n10541 ;
  assign n10543 = n6145 | n10542 ;
  assign n10544 = x101 | n10543 ;
  assign n10545 = n196 | n7186 ;
  assign n10546 = n6579 | n10545 ;
  assign n10547 = x74 | n5719 ;
  assign n10548 = n5742 & n10547 ;
  assign n10549 = ~n10434 & n10548 ;
  assign n10550 = n508 & ~n10549 ;
  assign n10551 = ( n3200 & n3316 ) | ( n3200 & n10550 ) | ( n3316 & n10550 ) ;
  assign n10552 = n581 | n7046 ;
  assign n10553 = n10552 ^ n3284 ^ 1'b0 ;
  assign n10554 = n4355 & ~n9939 ;
  assign n10555 = n3310 | n10554 ;
  assign n10556 = n5989 & ~n7908 ;
  assign n10557 = n6031 & n10556 ;
  assign n10558 = n10557 ^ n6223 ^ 1'b0 ;
  assign n10559 = n2102 & ~n8405 ;
  assign n10560 = n10559 ^ n10095 ^ 1'b0 ;
  assign n10561 = n4366 ^ n4146 ^ 1'b0 ;
  assign n10562 = n3324 & n5289 ;
  assign n10563 = n10561 & n10562 ;
  assign n10564 = n10563 ^ n8729 ^ 1'b0 ;
  assign n10565 = n2315 ^ n1745 ^ 1'b0 ;
  assign n10566 = n10440 ^ x66 ^ 1'b0 ;
  assign n10567 = ( n1390 & n2291 ) | ( n1390 & n3176 ) | ( n2291 & n3176 ) ;
  assign n10568 = n10567 ^ x28 ^ 1'b0 ;
  assign n10569 = n5034 & n10568 ;
  assign n10570 = n8717 ^ n2930 ^ 1'b0 ;
  assign n10571 = n10569 & ~n10570 ;
  assign n10572 = n6713 ^ n6259 ^ 1'b0 ;
  assign n10573 = n10572 ^ n7461 ^ 1'b0 ;
  assign n10574 = n10571 & ~n10573 ;
  assign n10575 = n7930 ^ n3828 ^ 1'b0 ;
  assign n10576 = ~n3492 & n10575 ;
  assign n10577 = n10576 ^ n9915 ^ 1'b0 ;
  assign n10578 = n886 & n7037 ;
  assign n10579 = n10578 ^ n3929 ^ 1'b0 ;
  assign n10580 = n3026 | n5573 ;
  assign n10581 = n10580 ^ n1465 ^ 1'b0 ;
  assign n10582 = ( n7079 & ~n8967 ) | ( n7079 & n10581 ) | ( ~n8967 & n10581 ) ;
  assign n10583 = n6151 ^ n1521 ^ 1'b0 ;
  assign n10584 = n2279 & ~n10583 ;
  assign n10585 = n3984 & ~n6563 ;
  assign n10586 = ~n6166 & n10585 ;
  assign n10587 = n3272 | n4014 ;
  assign n10588 = n1688 & ~n10587 ;
  assign n10589 = n548 | n10588 ;
  assign n10590 = n10586 & ~n10589 ;
  assign n10591 = n620 & n6264 ;
  assign n10592 = n10591 ^ n4285 ^ 1'b0 ;
  assign n10593 = ~n9898 & n10229 ;
  assign n10594 = n7528 ^ n5749 ^ n1074 ;
  assign n10595 = n2221 | n10594 ;
  assign n10596 = n4347 & ~n7087 ;
  assign n10597 = n10596 ^ n2193 ^ 1'b0 ;
  assign n10598 = n10597 ^ n2677 ^ n818 ;
  assign n10599 = n10598 ^ n7662 ^ 1'b0 ;
  assign n10600 = n2893 & n10599 ;
  assign n10601 = n376 & n2055 ;
  assign n10602 = n10601 ^ n5535 ^ 1'b0 ;
  assign n10603 = n2259 ^ n586 ^ 1'b0 ;
  assign n10604 = n445 | n10603 ;
  assign n10605 = n10604 ^ n2928 ^ 1'b0 ;
  assign n10608 = n1458 ^ n279 ^ 1'b0 ;
  assign n10609 = ~n202 & n10608 ;
  assign n10606 = ( ~n443 & n2098 ) | ( ~n443 & n2998 ) | ( n2098 & n2998 ) ;
  assign n10607 = ~n6214 & n10606 ;
  assign n10610 = n10609 ^ n10607 ^ 1'b0 ;
  assign n10611 = ( ~n5561 & n8573 ) | ( ~n5561 & n10610 ) | ( n8573 & n10610 ) ;
  assign n10612 = n4996 & n8846 ;
  assign n10613 = ( n1422 & n2341 ) | ( n1422 & n10612 ) | ( n2341 & n10612 ) ;
  assign n10614 = n10613 ^ n129 ^ 1'b0 ;
  assign n10615 = n1655 & n10614 ;
  assign n10616 = ( ~n1445 & n1664 ) | ( ~n1445 & n3918 ) | ( n1664 & n3918 ) ;
  assign n10617 = n7391 & n10616 ;
  assign n10618 = n10617 ^ n5808 ^ 1'b0 ;
  assign n10619 = n1669 & n2376 ;
  assign n10620 = ~n2132 & n10619 ;
  assign n10621 = ~n8570 & n10620 ;
  assign n10622 = n6120 ^ n3325 ^ 1'b0 ;
  assign n10623 = n1998 & ~n4358 ;
  assign n10624 = n7402 & ~n9569 ;
  assign n10625 = n379 & n3510 ;
  assign n10626 = n10625 ^ n6675 ^ n2727 ;
  assign n10627 = n10626 ^ n3557 ^ 1'b0 ;
  assign n10628 = n2579 & ~n10306 ;
  assign n10629 = n8863 ^ n1614 ^ 1'b0 ;
  assign n10630 = n6327 | n8584 ;
  assign n10631 = ~n10629 & n10630 ;
  assign n10634 = n1842 & ~n7436 ;
  assign n10635 = n10634 ^ n4368 ^ 1'b0 ;
  assign n10636 = n1652 & n10635 ;
  assign n10637 = n10636 ^ n6157 ^ n5993 ;
  assign n10632 = x110 & ~n3557 ;
  assign n10633 = n5740 & n10632 ;
  assign n10638 = n10637 ^ n10633 ^ n1329 ;
  assign n10639 = n2665 & n6807 ;
  assign n10640 = n10639 ^ n4560 ^ 1'b0 ;
  assign n10641 = n1550 & n10126 ;
  assign n10642 = n10640 & n10641 ;
  assign n10643 = n9904 ^ n6550 ^ n2514 ;
  assign n10644 = n5519 & ~n6199 ;
  assign n10645 = n490 & n2125 ;
  assign n10646 = n680 | n1477 ;
  assign n10647 = n10646 ^ n1101 ^ 1'b0 ;
  assign n10648 = n10647 ^ n1390 ^ 1'b0 ;
  assign n10649 = n906 & ~n10648 ;
  assign n10650 = n7229 | n10649 ;
  assign n10651 = n1001 & ~n6821 ;
  assign n10652 = ( n3055 & ~n3182 ) | ( n3055 & n10651 ) | ( ~n3182 & n10651 ) ;
  assign n10653 = ~n8028 & n10652 ;
  assign n10654 = n8584 ^ n4716 ^ 1'b0 ;
  assign n10655 = n10126 ^ n2819 ^ 1'b0 ;
  assign n10656 = n10654 & n10655 ;
  assign n10657 = n10127 & n10656 ;
  assign n10658 = n4316 ^ n1064 ^ 1'b0 ;
  assign n10659 = n6361 ^ n4545 ^ 1'b0 ;
  assign n10660 = ~n3628 & n10659 ;
  assign n10664 = n5389 ^ n3011 ^ 1'b0 ;
  assign n10665 = n4605 | n10664 ;
  assign n10661 = ~n370 & n5885 ;
  assign n10662 = n396 & n10661 ;
  assign n10663 = ~n5414 & n10662 ;
  assign n10666 = n10665 ^ n10663 ^ 1'b0 ;
  assign n10667 = n3705 | n4219 ;
  assign n10668 = n2500 | n10667 ;
  assign n10669 = n7514 ^ n3776 ^ 1'b0 ;
  assign n10670 = n10668 | n10669 ;
  assign n10671 = ~n5613 & n10542 ;
  assign n10672 = n10671 ^ n10208 ^ n7924 ;
  assign n10673 = n5208 ^ n1698 ^ 1'b0 ;
  assign n10674 = n2665 ^ n1069 ^ 1'b0 ;
  assign n10675 = n2455 & ~n10674 ;
  assign n10676 = n2540 & n10675 ;
  assign n10677 = n3001 & n10676 ;
  assign n10678 = n10673 | n10677 ;
  assign n10679 = n10678 ^ n9760 ^ 1'b0 ;
  assign n10680 = ( n798 & ~n7720 ) | ( n798 & n9287 ) | ( ~n7720 & n9287 ) ;
  assign n10681 = ( n6834 & n8233 ) | ( n6834 & n10680 ) | ( n8233 & n10680 ) ;
  assign n10682 = n8269 ^ n5648 ^ 1'b0 ;
  assign n10683 = ~n686 & n2033 ;
  assign n10684 = n10683 ^ n8709 ^ 1'b0 ;
  assign n10685 = n2980 ^ n891 ^ 1'b0 ;
  assign n10686 = n10684 & ~n10685 ;
  assign n10687 = ~n3618 & n10686 ;
  assign n10688 = n10682 & n10687 ;
  assign n10689 = n3214 & n8148 ;
  assign n10690 = n2328 | n7061 ;
  assign n10691 = n5265 | n10690 ;
  assign n10692 = n7108 ^ x96 ^ 1'b0 ;
  assign n10693 = n10692 ^ n3776 ^ 1'b0 ;
  assign n10694 = n5562 | n10693 ;
  assign n10695 = n10694 ^ n10071 ^ 1'b0 ;
  assign n10696 = ~n763 & n7887 ;
  assign n10697 = n1374 & n10696 ;
  assign n10698 = n10697 ^ n7599 ^ n683 ;
  assign n10699 = n8711 ^ n7930 ^ n3767 ;
  assign n10700 = n10699 ^ n7893 ^ 1'b0 ;
  assign n10701 = n10260 ^ x110 ^ 1'b0 ;
  assign n10702 = n10701 ^ n2038 ^ n1159 ;
  assign n10703 = n6308 ^ n1637 ^ 1'b0 ;
  assign n10704 = n4029 & n6452 ;
  assign n10705 = n10704 ^ n9085 ^ n2199 ;
  assign n10709 = ( ~n1192 & n1983 ) | ( ~n1192 & n2850 ) | ( n1983 & n2850 ) ;
  assign n10706 = n2373 & ~n5169 ;
  assign n10707 = n3444 & n10706 ;
  assign n10708 = n7469 | n10707 ;
  assign n10710 = n10709 ^ n10708 ^ 1'b0 ;
  assign n10711 = n10710 ^ n9751 ^ n7235 ;
  assign n10712 = n1996 & ~n10711 ;
  assign n10713 = n8496 ^ n3989 ^ 1'b0 ;
  assign n10714 = n7238 & n10713 ;
  assign n10715 = ~n2780 & n8938 ;
  assign n10716 = n10715 ^ n4867 ^ 1'b0 ;
  assign n10717 = n5098 ^ n5036 ^ n1747 ;
  assign n10718 = n10716 & ~n10717 ;
  assign n10719 = x126 & ~n1892 ;
  assign n10720 = n5024 ^ n2076 ^ 1'b0 ;
  assign n10721 = ( n7091 & n10719 ) | ( n7091 & ~n10720 ) | ( n10719 & ~n10720 ) ;
  assign n10722 = ( n2297 & n3080 ) | ( n2297 & n3838 ) | ( n3080 & n3838 ) ;
  assign n10723 = ~n7502 & n8934 ;
  assign n10724 = n10723 ^ n5493 ^ 1'b0 ;
  assign n10726 = ~n2529 & n6068 ;
  assign n10727 = n2435 & n10726 ;
  assign n10728 = n10727 ^ n5036 ^ 1'b0 ;
  assign n10729 = ~n6991 & n10728 ;
  assign n10725 = ~n1610 & n8004 ;
  assign n10730 = n10729 ^ n10725 ^ 1'b0 ;
  assign n10731 = n3999 ^ n2851 ^ 1'b0 ;
  assign n10734 = n4509 | n5366 ;
  assign n10735 = n10734 ^ n4851 ^ 1'b0 ;
  assign n10732 = ~n2736 & n10625 ;
  assign n10733 = ~n8206 & n10732 ;
  assign n10736 = n10735 ^ n10733 ^ n3999 ;
  assign n10737 = n4472 & n8419 ;
  assign n10738 = n557 | n10476 ;
  assign n10739 = n10738 ^ n3599 ^ 1'b0 ;
  assign n10740 = ~n5036 & n10739 ;
  assign n10741 = n1853 & n4828 ;
  assign n10742 = n4911 ^ n1113 ^ 1'b0 ;
  assign n10743 = n1722 & n8862 ;
  assign n10744 = n10742 & n10743 ;
  assign n10745 = n10744 ^ n2749 ^ 1'b0 ;
  assign n10746 = n10741 & n10745 ;
  assign n10750 = n2973 ^ x12 ^ 1'b0 ;
  assign n10751 = n10750 ^ n4273 ^ 1'b0 ;
  assign n10752 = n10751 ^ n5632 ^ 1'b0 ;
  assign n10753 = n6533 & n10752 ;
  assign n10747 = n640 | n1582 ;
  assign n10748 = x98 & ~n10747 ;
  assign n10749 = ( n1703 & n8222 ) | ( n1703 & ~n10748 ) | ( n8222 & ~n10748 ) ;
  assign n10754 = n10753 ^ n10749 ^ 1'b0 ;
  assign n10755 = ~n3307 & n10689 ;
  assign n10756 = n10755 ^ n6791 ^ 1'b0 ;
  assign n10757 = n3560 & ~n10251 ;
  assign n10758 = n1171 | n6318 ;
  assign n10759 = n5103 ^ n424 ^ 1'b0 ;
  assign n10760 = n10758 & n10759 ;
  assign n10761 = ( n4957 & n10703 ) | ( n4957 & n10760 ) | ( n10703 & n10760 ) ;
  assign n10762 = n3016 | n5003 ;
  assign n10763 = ~n8512 & n10762 ;
  assign n10764 = ~n6026 & n8361 ;
  assign n10765 = n4778 & n10764 ;
  assign n10766 = ~n5471 & n10765 ;
  assign n10767 = n433 | n4379 ;
  assign n10768 = n2817 & n10767 ;
  assign n10772 = n1411 & n1996 ;
  assign n10769 = n5927 ^ n3059 ^ 1'b0 ;
  assign n10770 = n10769 ^ n5446 ^ n5369 ;
  assign n10771 = n7051 & ~n10770 ;
  assign n10773 = n10772 ^ n10771 ^ n2710 ;
  assign n10775 = n1034 & ~n3872 ;
  assign n10776 = n10775 ^ n8190 ^ n5745 ;
  assign n10774 = n5530 ^ n1837 ^ 1'b0 ;
  assign n10777 = n10776 ^ n10774 ^ 1'b0 ;
  assign n10778 = n10773 & n10777 ;
  assign n10779 = ~n10768 & n10778 ;
  assign n10780 = n3351 | n4819 ;
  assign n10783 = n1428 | n6049 ;
  assign n10781 = n1613 & ~n7099 ;
  assign n10782 = n7784 | n10781 ;
  assign n10784 = n10783 ^ n10782 ^ 1'b0 ;
  assign n10785 = n2490 | n2597 ;
  assign n10786 = ( n2202 & ~n4468 ) | ( n2202 & n10785 ) | ( ~n4468 & n10785 ) ;
  assign n10787 = n10786 ^ n2125 ^ 1'b0 ;
  assign n10788 = n3773 & n10787 ;
  assign n10789 = ~n935 & n2503 ;
  assign n10790 = ( ~n366 & n6083 ) | ( ~n366 & n9381 ) | ( n6083 & n9381 ) ;
  assign n10791 = ~n3304 & n4962 ;
  assign n10792 = ~n10790 & n10791 ;
  assign n10793 = n10792 ^ n7269 ^ 1'b0 ;
  assign n10794 = ( n4291 & ~n7955 ) | ( n4291 & n8437 ) | ( ~n7955 & n8437 ) ;
  assign n10795 = n10071 ^ n6104 ^ 1'b0 ;
  assign n10796 = ~n10794 & n10795 ;
  assign n10797 = n3193 ^ n2622 ^ 1'b0 ;
  assign n10798 = ~n8282 & n10797 ;
  assign n10799 = n7538 & n10798 ;
  assign n10800 = n4347 ^ n984 ^ 1'b0 ;
  assign n10801 = n10800 ^ n5464 ^ 1'b0 ;
  assign n10802 = n4147 & ~n10801 ;
  assign n10803 = n10802 ^ n10028 ^ 1'b0 ;
  assign n10804 = n840 & n10803 ;
  assign n10805 = n707 & ~n1578 ;
  assign n10806 = n10805 ^ n8177 ^ n1127 ;
  assign n10808 = ~n1689 & n2546 ;
  assign n10807 = n2364 & ~n4999 ;
  assign n10809 = n10808 ^ n10807 ^ 1'b0 ;
  assign n10810 = n10809 ^ n8835 ^ n562 ;
  assign n10811 = n1821 & ~n2966 ;
  assign n10812 = n10811 ^ n653 ^ n206 ;
  assign n10813 = x10 & n1476 ;
  assign n10814 = n10813 ^ n6728 ^ 1'b0 ;
  assign n10815 = ( n5412 & n10125 ) | ( n5412 & ~n10814 ) | ( n10125 & ~n10814 ) ;
  assign n10816 = n3631 ^ n1962 ^ 1'b0 ;
  assign n10817 = ~n2964 & n10816 ;
  assign n10818 = n10817 ^ n10188 ^ 1'b0 ;
  assign n10819 = n645 | n10818 ;
  assign n10820 = n10819 ^ n2625 ^ 1'b0 ;
  assign n10821 = n2878 ^ n2817 ^ 1'b0 ;
  assign n10822 = n4602 & ~n9515 ;
  assign n10823 = n2180 ^ x84 ^ 1'b0 ;
  assign n10824 = n4331 | n6088 ;
  assign n10825 = n4330 | n10824 ;
  assign n10829 = n2443 & n3285 ;
  assign n10828 = n3961 & n9440 ;
  assign n10830 = n10829 ^ n10828 ^ 1'b0 ;
  assign n10826 = n3031 | n6408 ;
  assign n10827 = n5155 & ~n10826 ;
  assign n10831 = n10830 ^ n10827 ^ 1'b0 ;
  assign n10832 = n4805 & ~n8530 ;
  assign n10839 = n2701 | n4113 ;
  assign n10840 = n10839 ^ n4672 ^ 1'b0 ;
  assign n10841 = n10840 ^ n4243 ^ n4030 ;
  assign n10833 = ~n4471 & n6597 ;
  assign n10834 = x9 | n10833 ;
  assign n10835 = n6148 ^ n3554 ^ 1'b0 ;
  assign n10836 = n7169 & ~n10835 ;
  assign n10837 = n1654 & n10836 ;
  assign n10838 = ( n1155 & n10834 ) | ( n1155 & n10837 ) | ( n10834 & n10837 ) ;
  assign n10842 = n10841 ^ n10838 ^ 1'b0 ;
  assign n10843 = n7198 ^ n5784 ^ n5783 ;
  assign n10844 = n840 & ~n10843 ;
  assign n10845 = ~n5152 & n10844 ;
  assign n10849 = n6164 & n6543 ;
  assign n10850 = n10849 ^ n7214 ^ 1'b0 ;
  assign n10846 = n4448 ^ n703 ^ 1'b0 ;
  assign n10847 = n5863 & n10846 ;
  assign n10848 = ~n7816 & n10847 ;
  assign n10851 = n10850 ^ n10848 ^ 1'b0 ;
  assign n10852 = n7986 ^ n1338 ^ 1'b0 ;
  assign n10853 = n8028 | n10852 ;
  assign n10854 = ( n614 & n8113 ) | ( n614 & n10853 ) | ( n8113 & n10853 ) ;
  assign n10855 = n2238 & ~n2905 ;
  assign n10856 = n2591 | n4650 ;
  assign n10859 = n2073 | n2111 ;
  assign n10860 = n627 & ~n10859 ;
  assign n10861 = n10860 ^ n2806 ^ 1'b0 ;
  assign n10862 = n935 & ~n10861 ;
  assign n10857 = n2484 ^ n256 ^ 1'b0 ;
  assign n10858 = ~n9758 & n10857 ;
  assign n10863 = n10862 ^ n10858 ^ n2337 ;
  assign n10864 = n2901 ^ n2081 ^ 1'b0 ;
  assign n10865 = n10863 | n10864 ;
  assign n10866 = n4685 & ~n7290 ;
  assign n10867 = ~n2496 & n10866 ;
  assign n10868 = n6165 ^ n4503 ^ 1'b0 ;
  assign n10869 = ( ~n3654 & n10422 ) | ( ~n3654 & n10868 ) | ( n10422 & n10868 ) ;
  assign n10870 = n2428 ^ n1842 ^ 1'b0 ;
  assign n10871 = ~n3686 & n8738 ;
  assign n10873 = n2900 ^ n1479 ^ 1'b0 ;
  assign n10872 = n6974 ^ n2725 ^ 1'b0 ;
  assign n10874 = n10873 ^ n10872 ^ 1'b0 ;
  assign n10875 = n2087 ^ n323 ^ 1'b0 ;
  assign n10876 = n510 & n10875 ;
  assign n10877 = n10876 ^ n1307 ^ 1'b0 ;
  assign n10878 = n7113 ^ n6311 ^ 1'b0 ;
  assign n10881 = ~n1044 & n2414 ;
  assign n10882 = n1800 & ~n2063 ;
  assign n10883 = n10881 & n10882 ;
  assign n10879 = n8052 ^ n3705 ^ 1'b0 ;
  assign n10880 = ~n5699 & n10879 ;
  assign n10884 = n10883 ^ n10880 ^ 1'b0 ;
  assign n10885 = n1818 ^ n1730 ^ 1'b0 ;
  assign n10886 = n8256 ^ n4380 ^ n436 ;
  assign n10887 = n10885 & n10886 ;
  assign n10888 = ~n10884 & n10887 ;
  assign n10889 = ( n167 & n10878 ) | ( n167 & ~n10888 ) | ( n10878 & ~n10888 ) ;
  assign n10890 = ~n771 & n1382 ;
  assign n10891 = ~n7478 & n10890 ;
  assign n10892 = n5030 ^ n4428 ^ 1'b0 ;
  assign n10893 = n9787 & ~n10892 ;
  assign n10894 = ~n4131 & n6031 ;
  assign n10895 = ~n1815 & n10894 ;
  assign n10896 = n10895 ^ n4951 ^ 1'b0 ;
  assign n10897 = ( n5452 & n5514 ) | ( n5452 & n6239 ) | ( n5514 & n6239 ) ;
  assign n10898 = n9228 ^ n4727 ^ n2574 ;
  assign n10899 = n5567 & ~n6435 ;
  assign n10900 = n10899 ^ n299 ^ 1'b0 ;
  assign n10901 = ~n3299 & n3435 ;
  assign n10902 = n10630 | n10901 ;
  assign n10903 = n1540 & ~n10902 ;
  assign n10904 = n325 & n6174 ;
  assign n10905 = n5882 & n10904 ;
  assign n10906 = n3950 ^ n597 ^ 1'b0 ;
  assign n10907 = ( n9217 & n10905 ) | ( n9217 & n10906 ) | ( n10905 & n10906 ) ;
  assign n10908 = n2819 ^ n1918 ^ n1470 ;
  assign n10909 = n3197 & n8293 ;
  assign n10910 = n3324 & n10909 ;
  assign n10911 = n4639 | n10910 ;
  assign n10912 = n10911 ^ n7780 ^ 1'b0 ;
  assign n10920 = n1578 ^ n331 ^ 1'b0 ;
  assign n10921 = n635 | n10920 ;
  assign n10922 = n10921 ^ n7372 ^ 1'b0 ;
  assign n10915 = n6325 ^ n4760 ^ 1'b0 ;
  assign n10916 = n3893 | n10915 ;
  assign n10917 = ~n2639 & n3355 ;
  assign n10918 = n10916 & n10917 ;
  assign n10913 = n7639 ^ n799 ^ 1'b0 ;
  assign n10914 = ~n3872 & n10913 ;
  assign n10919 = n10918 ^ n10914 ^ 1'b0 ;
  assign n10923 = n10922 ^ n10919 ^ 1'b0 ;
  assign n10924 = ~n808 & n2912 ;
  assign n10925 = n10126 & ~n10200 ;
  assign n10926 = n4869 & ~n8422 ;
  assign n10927 = n2287 & n10926 ;
  assign n10928 = n6886 | n9516 ;
  assign n10929 = n10927 & ~n10928 ;
  assign n10930 = ( n2968 & ~n7085 ) | ( n2968 & n10929 ) | ( ~n7085 & n10929 ) ;
  assign n10931 = n254 & n10351 ;
  assign n10932 = n7955 & ~n10200 ;
  assign n10933 = ( ~n5116 & n10499 ) | ( ~n5116 & n10932 ) | ( n10499 & n10932 ) ;
  assign n10934 = n8608 & ~n9567 ;
  assign n10935 = n1981 & n4651 ;
  assign n10936 = n10935 ^ n8996 ^ 1'b0 ;
  assign n10937 = ~n1185 & n10936 ;
  assign n10938 = n10937 ^ n5149 ^ x99 ;
  assign n10939 = n4723 & n6923 ;
  assign n10940 = n1710 ^ n342 ^ 1'b0 ;
  assign n10941 = n10939 & n10940 ;
  assign n10942 = n10941 ^ n6498 ^ 1'b0 ;
  assign n10943 = n1950 & ~n10942 ;
  assign n10944 = n1765 & n10265 ;
  assign n10945 = n3224 ^ n869 ^ 1'b0 ;
  assign n10946 = n4443 | n10945 ;
  assign n10947 = n4665 & n6481 ;
  assign n10948 = n3966 & ~n4686 ;
  assign n10949 = n2864 | n10881 ;
  assign n10950 = n3743 | n10949 ;
  assign n10951 = n10950 ^ n5324 ^ n5039 ;
  assign n10952 = n3340 ^ x49 ^ 1'b0 ;
  assign n10953 = n10951 & ~n10952 ;
  assign n10954 = n6763 ^ n1074 ^ 1'b0 ;
  assign n10955 = ( n1218 & n5266 ) | ( n1218 & ~n10954 ) | ( n5266 & ~n10954 ) ;
  assign n10956 = n804 & ~n10955 ;
  assign n10957 = n10956 ^ n5223 ^ 1'b0 ;
  assign n10958 = n569 | n5223 ;
  assign n10959 = n10958 ^ x69 ^ 1'b0 ;
  assign n10962 = n1714 & n2775 ;
  assign n10963 = ( ~n2472 & n3353 ) | ( ~n2472 & n10962 ) | ( n3353 & n10962 ) ;
  assign n10960 = n4076 & ~n4298 ;
  assign n10961 = n10960 ^ n3958 ^ 1'b0 ;
  assign n10964 = n10963 ^ n10961 ^ 1'b0 ;
  assign n10966 = n1630 & ~n2850 ;
  assign n10967 = n10966 ^ n2482 ^ 1'b0 ;
  assign n10965 = ~n3979 & n9657 ;
  assign n10968 = n10967 ^ n10965 ^ 1'b0 ;
  assign n10969 = n10636 ^ n7616 ^ n7606 ;
  assign n10970 = n2906 ^ n2096 ^ 1'b0 ;
  assign n10971 = ( x41 & n802 ) | ( x41 & ~n10970 ) | ( n802 & ~n10970 ) ;
  assign n10972 = ( ~x57 & n4288 ) | ( ~x57 & n9872 ) | ( n4288 & n9872 ) ;
  assign n10973 = n5048 & ~n10972 ;
  assign n10974 = n6387 & n10973 ;
  assign n10975 = ~n2892 & n5409 ;
  assign n10976 = ~n2469 & n8340 ;
  assign n10977 = n10975 & n10976 ;
  assign n10984 = n2419 | n9872 ;
  assign n10985 = n5979 & ~n10984 ;
  assign n10978 = n4946 ^ n3815 ^ 1'b0 ;
  assign n10979 = n7191 ^ n5306 ^ 1'b0 ;
  assign n10980 = n10978 & n10979 ;
  assign n10981 = ( n4850 & n5487 ) | ( n4850 & n10980 ) | ( n5487 & n10980 ) ;
  assign n10982 = ( ~n1936 & n7972 ) | ( ~n1936 & n10981 ) | ( n7972 & n10981 ) ;
  assign n10983 = n3313 & ~n10982 ;
  assign n10986 = n10985 ^ n10983 ^ 1'b0 ;
  assign n10987 = n10986 ^ n10165 ^ 1'b0 ;
  assign n10988 = ~n10977 & n10987 ;
  assign n10989 = ( n4757 & ~n5415 ) | ( n4757 & n5603 ) | ( ~n5415 & n5603 ) ;
  assign n10990 = n7340 & n10989 ;
  assign n10991 = n678 & n10990 ;
  assign n10992 = n10991 ^ n433 ^ 1'b0 ;
  assign n10993 = n10992 ^ n3766 ^ 1'b0 ;
  assign n10994 = n9093 ^ n5923 ^ 1'b0 ;
  assign n10995 = n6749 & ~n9605 ;
  assign n10996 = n630 & ~n904 ;
  assign n10997 = ( n654 & n1860 ) | ( n654 & n10996 ) | ( n1860 & n10996 ) ;
  assign n10998 = n5016 & ~n10997 ;
  assign n10999 = n10998 ^ n3242 ^ 1'b0 ;
  assign n11000 = n6820 ^ n1839 ^ 1'b0 ;
  assign n11001 = n8505 & ~n10277 ;
  assign n11002 = ~n8175 & n10246 ;
  assign n11003 = n11002 ^ n4180 ^ 1'b0 ;
  assign n11005 = n4776 & ~n6687 ;
  assign n11006 = n11005 ^ n6049 ^ 1'b0 ;
  assign n11004 = n775 & n8503 ;
  assign n11007 = n11006 ^ n11004 ^ 1'b0 ;
  assign n11008 = n10198 ^ n2846 ^ 1'b0 ;
  assign n11009 = n11008 ^ n5875 ^ 1'b0 ;
  assign n11010 = n7230 & n11009 ;
  assign n11011 = n11010 ^ n1609 ^ 1'b0 ;
  assign n11012 = n11007 & n11011 ;
  assign n11013 = n9065 ^ n2325 ^ 1'b0 ;
  assign n11014 = n7219 & ~n11013 ;
  assign n11016 = ~n6308 & n8336 ;
  assign n11017 = n11016 ^ n3367 ^ 1'b0 ;
  assign n11018 = x13 & ~n11017 ;
  assign n11019 = n11018 ^ n6497 ^ 1'b0 ;
  assign n11015 = n1019 & ~n9204 ;
  assign n11020 = n11019 ^ n11015 ^ 1'b0 ;
  assign n11021 = n11020 ^ n5321 ^ n1380 ;
  assign n11022 = n9947 ^ n3441 ^ 1'b0 ;
  assign n11023 = n3768 ^ n892 ^ 1'b0 ;
  assign n11024 = ~n405 & n11023 ;
  assign n11025 = n11024 ^ n7874 ^ 1'b0 ;
  assign n11026 = n11025 ^ n6840 ^ n4133 ;
  assign n11027 = ~n3247 & n11026 ;
  assign n11028 = ~n3972 & n11027 ;
  assign n11029 = n9468 ^ n4079 ^ 1'b0 ;
  assign n11030 = n10439 ^ n5585 ^ 1'b0 ;
  assign n11031 = n7473 | n11030 ;
  assign n11032 = ~n433 & n2667 ;
  assign n11033 = n7226 ^ n7173 ^ n3403 ;
  assign n11034 = n4672 ^ n1610 ^ 1'b0 ;
  assign n11035 = n5126 | n10863 ;
  assign n11036 = n736 | n5459 ;
  assign n11037 = n5300 | n8749 ;
  assign n11038 = ( n3585 & ~n9754 ) | ( n3585 & n9776 ) | ( ~n9754 & n9776 ) ;
  assign n11039 = n9163 ^ n450 ^ 1'b0 ;
  assign n11040 = n4094 | n11039 ;
  assign n11043 = ~n718 & n1265 ;
  assign n11041 = n1079 | n7220 ;
  assign n11042 = n4916 & ~n11041 ;
  assign n11044 = n11043 ^ n11042 ^ n2333 ;
  assign n11045 = n3297 ^ n2438 ^ 1'b0 ;
  assign n11046 = n4264 & n11045 ;
  assign n11047 = ~n11044 & n11046 ;
  assign n11048 = n11047 ^ n6520 ^ 1'b0 ;
  assign n11049 = n4672 ^ n1583 ^ 1'b0 ;
  assign n11050 = n11048 & n11049 ;
  assign n11051 = n8102 ^ n563 ^ 1'b0 ;
  assign n11057 = n4847 ^ n4518 ^ 1'b0 ;
  assign n11053 = n8541 ^ n1811 ^ 1'b0 ;
  assign n11054 = n11053 ^ n2433 ^ 1'b0 ;
  assign n11055 = ~n4129 & n11054 ;
  assign n11056 = ~n1835 & n11055 ;
  assign n11058 = n11057 ^ n11056 ^ 1'b0 ;
  assign n11052 = n2933 & ~n3304 ;
  assign n11059 = n11058 ^ n11052 ^ 1'b0 ;
  assign n11060 = n5671 ^ n485 ^ 1'b0 ;
  assign n11061 = n3415 & ~n11060 ;
  assign n11062 = ( n4777 & n10525 ) | ( n4777 & n11061 ) | ( n10525 & n11061 ) ;
  assign n11063 = n387 & n11062 ;
  assign n11064 = ~n1208 & n11063 ;
  assign n11066 = n6296 ^ n4456 ^ 1'b0 ;
  assign n11067 = n1413 | n11066 ;
  assign n11068 = ~n7816 & n11067 ;
  assign n11069 = ~n3895 & n11068 ;
  assign n11065 = ~n3870 & n6936 ;
  assign n11070 = n11069 ^ n11065 ^ 1'b0 ;
  assign n11071 = n3608 ^ n2866 ^ 1'b0 ;
  assign n11072 = n11071 ^ n2104 ^ 1'b0 ;
  assign n11073 = n279 & ~n11072 ;
  assign n11075 = n1265 & ~n8254 ;
  assign n11074 = n4981 ^ n1482 ^ 1'b0 ;
  assign n11076 = n11075 ^ n11074 ^ n7814 ;
  assign n11077 = n493 & n7787 ;
  assign n11078 = ~n3899 & n11077 ;
  assign n11079 = n6311 ^ n1218 ^ n509 ;
  assign n11080 = ( n2203 & ~n5244 ) | ( n2203 & n9934 ) | ( ~n5244 & n9934 ) ;
  assign n11081 = n11079 & n11080 ;
  assign n11082 = n6496 ^ n1930 ^ x2 ;
  assign n11083 = n1207 | n5238 ;
  assign n11084 = n8378 & ~n11083 ;
  assign n11085 = n4195 ^ n1586 ^ 1'b0 ;
  assign n11086 = n10018 | n11085 ;
  assign n11087 = n11086 ^ n2164 ^ 1'b0 ;
  assign n11088 = ~n973 & n4752 ;
  assign n11089 = n8397 & n11088 ;
  assign n11090 = ~n1623 & n11089 ;
  assign n11091 = n5389 ^ n2104 ^ n362 ;
  assign n11095 = n6425 ^ n3479 ^ 1'b0 ;
  assign n11096 = ( n1941 & ~n8455 ) | ( n1941 & n11095 ) | ( ~n8455 & n11095 ) ;
  assign n11092 = n4308 | n8380 ;
  assign n11093 = n9612 | n11092 ;
  assign n11094 = n9502 | n11093 ;
  assign n11097 = n11096 ^ n11094 ^ 1'b0 ;
  assign n11098 = ( n6872 & n6969 ) | ( n6872 & n8681 ) | ( n6969 & n8681 ) ;
  assign n11099 = n3417 & n8223 ;
  assign n11100 = n11099 ^ n2450 ^ 1'b0 ;
  assign n11101 = n3519 ^ n1888 ^ n202 ;
  assign n11102 = n1209 ^ n386 ^ 1'b0 ;
  assign n11103 = ~x82 & n11102 ;
  assign n11104 = ( ~n11100 & n11101 ) | ( ~n11100 & n11103 ) | ( n11101 & n11103 ) ;
  assign n11105 = n2522 | n4564 ;
  assign n11106 = ~n7062 & n11105 ;
  assign n11107 = n11106 ^ n2706 ^ 1'b0 ;
  assign n11108 = ~n2751 & n7951 ;
  assign n11109 = n6756 & n11108 ;
  assign n11110 = n11109 ^ n9375 ^ 1'b0 ;
  assign n11111 = n410 & n2266 ;
  assign n11112 = n11111 ^ n11109 ^ n4407 ;
  assign n11115 = n997 & n2947 ;
  assign n11116 = n5883 & n11115 ;
  assign n11113 = n7092 ^ n6360 ^ 1'b0 ;
  assign n11114 = n7726 & n11113 ;
  assign n11117 = n11116 ^ n11114 ^ 1'b0 ;
  assign n11118 = n10651 | n11117 ;
  assign n11120 = ( n4797 & n5511 ) | ( n4797 & n5667 ) | ( n5511 & n5667 ) ;
  assign n11121 = n5790 & n7401 ;
  assign n11122 = ~n11120 & n11121 ;
  assign n11119 = ~n2329 & n6892 ;
  assign n11123 = n11122 ^ n11119 ^ 1'b0 ;
  assign n11124 = n11123 ^ n3157 ^ 1'b0 ;
  assign n11125 = n4382 & ~n11124 ;
  assign n11126 = n11125 ^ n4068 ^ 1'b0 ;
  assign n11128 = n7119 ^ n271 ^ 1'b0 ;
  assign n11127 = n1123 & ~n1990 ;
  assign n11129 = n11128 ^ n11127 ^ 1'b0 ;
  assign n11130 = n3395 ^ n3105 ^ n2302 ;
  assign n11131 = ( ~n1155 & n6226 ) | ( ~n1155 & n11130 ) | ( n6226 & n11130 ) ;
  assign n11132 = n7197 ^ n5517 ^ n773 ;
  assign n11147 = ~n447 & n5591 ;
  assign n11148 = ~n1356 & n2290 ;
  assign n11149 = ( n5898 & n11147 ) | ( n5898 & n11148 ) | ( n11147 & n11148 ) ;
  assign n11150 = n8466 & ~n11149 ;
  assign n11151 = ~n8466 & n11150 ;
  assign n11133 = n202 | n425 ;
  assign n11134 = n202 & ~n11133 ;
  assign n11135 = n320 | n11134 ;
  assign n11136 = n11134 & ~n11135 ;
  assign n11137 = x39 & x70 ;
  assign n11138 = ~x39 & n11137 ;
  assign n11139 = x56 & n845 ;
  assign n11140 = n11138 & n11139 ;
  assign n11141 = n805 & n1627 ;
  assign n11142 = n11140 & n11141 ;
  assign n11143 = n3589 | n11142 ;
  assign n11144 = n11142 & ~n11143 ;
  assign n11145 = n11136 | n11144 ;
  assign n11146 = n11145 ^ n914 ^ 1'b0 ;
  assign n11152 = n11151 ^ n11146 ^ n4846 ;
  assign n11153 = n7242 ^ n7085 ^ 1'b0 ;
  assign n11154 = n561 & n2048 ;
  assign n11155 = ~n4844 & n11154 ;
  assign n11157 = n138 & ~n7444 ;
  assign n11158 = n11157 ^ n4704 ^ 1'b0 ;
  assign n11159 = n431 & n11158 ;
  assign n11156 = n3169 | n10368 ;
  assign n11160 = n11159 ^ n11156 ^ 1'b0 ;
  assign n11161 = n9162 ^ n8996 ^ 1'b0 ;
  assign n11162 = n5191 & n11161 ;
  assign n11163 = n6375 ^ n672 ^ 1'b0 ;
  assign n11164 = n678 & n2549 ;
  assign n11165 = n4854 & n11164 ;
  assign n11166 = n11165 ^ n283 ^ 1'b0 ;
  assign n11167 = n11163 | n11166 ;
  assign n11168 = ~n2194 & n7687 ;
  assign n11169 = n7927 ^ x88 ^ 1'b0 ;
  assign n11170 = n1869 | n11169 ;
  assign n11171 = n1000 & ~n7774 ;
  assign n11172 = n3930 & n11171 ;
  assign n11176 = n2877 & ~n2978 ;
  assign n11174 = n3055 ^ n1844 ^ 1'b0 ;
  assign n11175 = ( n5178 & ~n6557 ) | ( n5178 & n11174 ) | ( ~n6557 & n11174 ) ;
  assign n11173 = ( n2290 & ~n3240 ) | ( n2290 & n4023 ) | ( ~n3240 & n4023 ) ;
  assign n11177 = n11176 ^ n11175 ^ n11173 ;
  assign n11178 = n1219 & ~n1382 ;
  assign n11179 = n11178 ^ n2677 ^ n1945 ;
  assign n11180 = n4714 ^ n2926 ^ 1'b0 ;
  assign n11181 = n349 | n11180 ;
  assign n11182 = n11179 & ~n11181 ;
  assign n11183 = n739 ^ n134 ^ 1'b0 ;
  assign n11184 = ~n148 & n11183 ;
  assign n11186 = n726 & n10625 ;
  assign n11187 = n11186 ^ n1378 ^ 1'b0 ;
  assign n11185 = n9952 ^ n6647 ^ n422 ;
  assign n11188 = n11187 ^ n11185 ^ 1'b0 ;
  assign n11189 = n11184 & ~n11188 ;
  assign n11190 = n4363 ^ n4047 ^ 1'b0 ;
  assign n11191 = n11190 ^ n2679 ^ n327 ;
  assign n11192 = ( n3200 & n8887 ) | ( n3200 & ~n11191 ) | ( n8887 & ~n11191 ) ;
  assign n11193 = n7294 & ~n9472 ;
  assign n11199 = ( ~x121 & n398 ) | ( ~x121 & n7904 ) | ( n398 & n7904 ) ;
  assign n11196 = n5053 & ~n6168 ;
  assign n11197 = n3193 ^ n1782 ^ 1'b0 ;
  assign n11198 = n11196 & n11197 ;
  assign n11194 = n389 & n4043 ;
  assign n11195 = ~n5024 & n11194 ;
  assign n11200 = n11199 ^ n11198 ^ n11195 ;
  assign n11205 = n8257 ^ n6451 ^ 1'b0 ;
  assign n11202 = n403 & ~n2864 ;
  assign n11203 = n11202 ^ n1882 ^ 1'b0 ;
  assign n11201 = n988 | n11061 ;
  assign n11204 = n11203 ^ n11201 ^ 1'b0 ;
  assign n11206 = n11205 ^ n11204 ^ n3717 ;
  assign n11207 = ( ~n9559 & n10190 ) | ( ~n9559 & n11206 ) | ( n10190 & n11206 ) ;
  assign n11208 = ~n11200 & n11207 ;
  assign n11209 = ( n888 & n1500 ) | ( n888 & n5468 ) | ( n1500 & n5468 ) ;
  assign n11210 = ( ~n771 & n9960 ) | ( ~n771 & n11209 ) | ( n9960 & n11209 ) ;
  assign n11213 = n5128 ^ n4597 ^ 1'b0 ;
  assign n11214 = n4059 & ~n11213 ;
  assign n11211 = n912 & n2207 ;
  assign n11212 = ~n8225 & n11211 ;
  assign n11215 = n11214 ^ n11212 ^ 1'b0 ;
  assign n11216 = n4275 ^ n3187 ^ 1'b0 ;
  assign n11217 = n7514 & ~n11216 ;
  assign n11218 = ~n3828 & n11217 ;
  assign n11219 = n3856 & n11218 ;
  assign n11220 = n1959 & n6915 ;
  assign n11221 = n11219 & n11220 ;
  assign n11222 = n9756 | n10439 ;
  assign n11223 = n7027 | n10372 ;
  assign n11224 = n7597 | n9894 ;
  assign n11225 = ( n2368 & ~n6018 ) | ( n2368 & n8709 ) | ( ~n6018 & n8709 ) ;
  assign n11226 = n9617 & n11225 ;
  assign n11227 = n8537 ^ n3040 ^ n2030 ;
  assign n11228 = n2091 & n8971 ;
  assign n11229 = n11227 & n11228 ;
  assign n11232 = n1085 & ~n7161 ;
  assign n11233 = n8903 & n11232 ;
  assign n11234 = ~n5761 & n11233 ;
  assign n11230 = ~n7452 & n10136 ;
  assign n11231 = n10318 & ~n11230 ;
  assign n11235 = n11234 ^ n11231 ^ 1'b0 ;
  assign n11236 = x103 & n7647 ;
  assign n11237 = n3529 | n4605 ;
  assign n11238 = n10035 & ~n11237 ;
  assign n11239 = n9259 ^ n869 ^ 1'b0 ;
  assign n11240 = n1671 & n4133 ;
  assign n11241 = n11240 ^ n4294 ^ 1'b0 ;
  assign n11242 = n5600 & ~n11241 ;
  assign n11243 = n2527 ^ n1177 ^ x50 ;
  assign n11244 = n411 ^ n229 ^ 1'b0 ;
  assign n11245 = ~n823 & n11244 ;
  assign n11246 = n1846 ^ n595 ^ 1'b0 ;
  assign n11247 = n11245 & n11246 ;
  assign n11248 = n11247 ^ n7083 ^ n3143 ;
  assign n11249 = n6796 & n11248 ;
  assign n11250 = ~n11243 & n11249 ;
  assign n11251 = n2199 | n3535 ;
  assign n11252 = ~n2845 & n5608 ;
  assign n11253 = n11252 ^ n1664 ^ 1'b0 ;
  assign n11254 = n1503 | n6905 ;
  assign n11255 = n2652 & ~n7309 ;
  assign n11256 = n4907 & ~n8991 ;
  assign n11257 = n5160 & ~n9592 ;
  assign n11258 = ~n5693 & n11257 ;
  assign n11259 = ( n1106 & n1996 ) | ( n1106 & ~n2868 ) | ( n1996 & ~n2868 ) ;
  assign n11260 = n10052 & n11259 ;
  assign n11261 = n2333 ^ x103 ^ 1'b0 ;
  assign n11262 = n4335 & n11261 ;
  assign n11263 = n5076 ^ n1162 ^ 1'b0 ;
  assign n11264 = n1730 & ~n11263 ;
  assign n11265 = n11264 ^ n5144 ^ 1'b0 ;
  assign n11266 = n490 ^ n242 ^ 1'b0 ;
  assign n11267 = n6931 ^ n2607 ^ 1'b0 ;
  assign n11268 = n11266 & ~n11267 ;
  assign n11273 = n6002 ^ n5256 ^ n5213 ;
  assign n11272 = n2637 ^ n681 ^ 1'b0 ;
  assign n11274 = n11273 ^ n11272 ^ n4375 ;
  assign n11275 = n11274 ^ n3340 ^ 1'b0 ;
  assign n11269 = n6672 ^ n2812 ^ 1'b0 ;
  assign n11270 = n6579 & n11269 ;
  assign n11271 = n6081 & ~n11270 ;
  assign n11276 = n11275 ^ n11271 ^ 1'b0 ;
  assign n11277 = n7536 ^ n7422 ^ 1'b0 ;
  assign n11278 = n2299 & n4495 ;
  assign n11279 = n9944 & n11071 ;
  assign n11280 = ( n1811 & n1894 ) | ( n1811 & ~n2694 ) | ( n1894 & ~n2694 ) ;
  assign n11281 = n1853 | n11280 ;
  assign n11282 = ( n1309 & n10308 ) | ( n1309 & n11281 ) | ( n10308 & n11281 ) ;
  assign n11283 = ( n5121 & n6566 ) | ( n5121 & n7601 ) | ( n6566 & n7601 ) ;
  assign n11284 = n7118 & n7594 ;
  assign n11286 = n10967 ^ n4429 ^ 1'b0 ;
  assign n11285 = n5708 & ~n6607 ;
  assign n11287 = n11286 ^ n11285 ^ 1'b0 ;
  assign n11288 = n2551 & ~n11203 ;
  assign n11289 = ~n3328 & n11288 ;
  assign n11290 = ~n11287 & n11289 ;
  assign n11291 = n3687 & ~n4879 ;
  assign n11292 = n6223 ^ n3701 ^ 1'b0 ;
  assign n11293 = n11292 ^ n4306 ^ x122 ;
  assign n11294 = n8466 ^ n5277 ^ 1'b0 ;
  assign n11295 = ( n8501 & ~n10650 ) | ( n8501 & n11294 ) | ( ~n10650 & n11294 ) ;
  assign n11296 = n3770 ^ n1989 ^ 1'b0 ;
  assign n11297 = ~n8899 & n11296 ;
  assign n11298 = n1892 & ~n3938 ;
  assign n11299 = n5790 | n11298 ;
  assign n11300 = n614 & ~n1624 ;
  assign n11301 = n623 | n11300 ;
  assign n11302 = n11301 ^ n9934 ^ 1'b0 ;
  assign n11303 = n1275 | n7960 ;
  assign n11304 = n1150 & ~n7003 ;
  assign n11305 = ( ~n1166 & n2937 ) | ( ~n1166 & n11304 ) | ( n2937 & n11304 ) ;
  assign n11307 = ~n657 & n1435 ;
  assign n11308 = n11307 ^ n1798 ^ 1'b0 ;
  assign n11306 = n6202 ^ n1034 ^ 1'b0 ;
  assign n11309 = n11308 ^ n11306 ^ 1'b0 ;
  assign n11311 = n1197 ^ n217 ^ 1'b0 ;
  assign n11310 = n7514 ^ n1796 ^ 1'b0 ;
  assign n11312 = n11311 ^ n11310 ^ n9470 ;
  assign n11313 = n8652 ^ n5359 ^ 1'b0 ;
  assign n11314 = n11312 | n11313 ;
  assign n11315 = n4374 ^ x110 ^ 1'b0 ;
  assign n11316 = n7199 & n11315 ;
  assign n11317 = ~n3175 & n11316 ;
  assign n11318 = n11317 ^ n2285 ^ 1'b0 ;
  assign n11319 = n3938 ^ n1680 ^ 1'b0 ;
  assign n11320 = n910 | n11319 ;
  assign n11321 = n6797 | n11320 ;
  assign n11322 = n11321 ^ n4895 ^ 1'b0 ;
  assign n11323 = n8859 ^ n6286 ^ 1'b0 ;
  assign n11324 = n451 & n11323 ;
  assign n11325 = n11324 ^ n725 ^ 1'b0 ;
  assign n11326 = ~n1308 & n11325 ;
  assign n11327 = n2625 | n5888 ;
  assign n11328 = ( n6240 & n9294 ) | ( n6240 & n11327 ) | ( n9294 & n11327 ) ;
  assign n11329 = ( n408 & n1044 ) | ( n408 & ~n11328 ) | ( n1044 & ~n11328 ) ;
  assign n11330 = n11329 ^ n8343 ^ n1860 ;
  assign n11331 = n2200 & ~n9189 ;
  assign n11332 = ( n720 & n11330 ) | ( n720 & n11331 ) | ( n11330 & n11331 ) ;
  assign n11333 = n10096 & ~n10681 ;
  assign n11334 = n1300 & n11333 ;
  assign n11335 = ( ~n2033 & n4708 ) | ( ~n2033 & n7723 ) | ( n4708 & n7723 ) ;
  assign n11336 = n6073 | n11335 ;
  assign n11342 = n1940 ^ n129 ^ 1'b0 ;
  assign n11343 = ~n1433 & n11342 ;
  assign n11344 = n11343 ^ n1485 ^ n1042 ;
  assign n11337 = n3369 ^ x127 ^ 1'b0 ;
  assign n11338 = n4912 & ~n11337 ;
  assign n11339 = ( n3599 & ~n5563 ) | ( n3599 & n7142 ) | ( ~n5563 & n7142 ) ;
  assign n11340 = ~n1281 & n11339 ;
  assign n11341 = n11338 & n11340 ;
  assign n11345 = n11344 ^ n11341 ^ n5887 ;
  assign n11346 = ( ~n975 & n3085 ) | ( ~n975 & n7683 ) | ( n3085 & n7683 ) ;
  assign n11347 = n3455 | n6563 ;
  assign n11348 = n5291 & ~n11347 ;
  assign n11349 = n177 | n11348 ;
  assign n11350 = n4861 | n11349 ;
  assign n11351 = n10500 ^ n920 ^ 1'b0 ;
  assign n11352 = n6671 ^ n1639 ^ 1'b0 ;
  assign n11353 = n7865 & n11352 ;
  assign n11354 = n11351 | n11353 ;
  assign n11355 = n5357 ^ n3359 ^ 1'b0 ;
  assign n11356 = n1034 & n11355 ;
  assign n11357 = n5567 | n7855 ;
  assign n11358 = n11356 & ~n11357 ;
  assign n11359 = n5927 | n7665 ;
  assign n11360 = n309 | n11359 ;
  assign n11361 = n1271 | n10229 ;
  assign n11362 = n11361 ^ n2696 ^ 1'b0 ;
  assign n11363 = ( n1567 & n6701 ) | ( n1567 & ~n11362 ) | ( n6701 & ~n11362 ) ;
  assign n11364 = n9144 ^ n1141 ^ 1'b0 ;
  assign n11365 = ( n130 & n11061 ) | ( n130 & ~n11364 ) | ( n11061 & ~n11364 ) ;
  assign n11366 = ~n221 & n750 ;
  assign n11369 = n4439 ^ n723 ^ 1'b0 ;
  assign n11370 = ~n1597 & n11369 ;
  assign n11367 = ~n4632 & n4898 ;
  assign n11368 = n11367 ^ n994 ^ 1'b0 ;
  assign n11371 = n11370 ^ n11368 ^ 1'b0 ;
  assign n11372 = n11366 & ~n11371 ;
  assign n11373 = ~n1150 & n10125 ;
  assign n11374 = n11373 ^ n4407 ^ 1'b0 ;
  assign n11375 = n403 & n9418 ;
  assign n11376 = n11375 ^ n1943 ^ 1'b0 ;
  assign n11377 = n673 & ~n11376 ;
  assign n11378 = ~n408 & n11377 ;
  assign n11379 = ( n1425 & n4110 ) | ( n1425 & ~n11378 ) | ( n4110 & ~n11378 ) ;
  assign n11380 = ~n8488 & n11379 ;
  assign n11381 = n2422 & ~n4870 ;
  assign n11382 = n11381 ^ n1724 ^ 1'b0 ;
  assign n11383 = n548 | n4159 ;
  assign n11384 = n2020 ^ n1311 ^ 1'b0 ;
  assign n11385 = ( ~n1590 & n4698 ) | ( ~n1590 & n11384 ) | ( n4698 & n11384 ) ;
  assign n11386 = n2492 ^ n389 ^ 1'b0 ;
  assign n11396 = n388 & n8639 ;
  assign n11391 = n5116 ^ n729 ^ 1'b0 ;
  assign n11392 = n229 | n11391 ;
  assign n11393 = n11392 ^ n1010 ^ 1'b0 ;
  assign n11394 = ( n1309 & n7534 ) | ( n1309 & n11393 ) | ( n7534 & n11393 ) ;
  assign n11387 = n1575 & ~n2348 ;
  assign n11388 = ~n5820 & n11387 ;
  assign n11389 = ~n1630 & n11388 ;
  assign n11390 = n8488 | n11389 ;
  assign n11395 = n11394 ^ n11390 ^ 1'b0 ;
  assign n11397 = n11396 ^ n11395 ^ n3022 ;
  assign n11398 = ( n3657 & n4457 ) | ( n3657 & n6145 ) | ( n4457 & n6145 ) ;
  assign n11399 = ( n342 & ~n3036 ) | ( n342 & n5598 ) | ( ~n3036 & n5598 ) ;
  assign n11400 = n2703 & ~n11399 ;
  assign n11401 = n11400 ^ n8181 ^ 1'b0 ;
  assign n11402 = n3584 ^ n2892 ^ 1'b0 ;
  assign n11403 = n6940 & ~n11402 ;
  assign n11404 = n5189 & ~n11403 ;
  assign n11405 = ( n3315 & ~n4652 ) | ( n3315 & n11404 ) | ( ~n4652 & n11404 ) ;
  assign n11406 = ~n1980 & n5551 ;
  assign n11407 = ( n3075 & n4185 ) | ( n3075 & ~n11406 ) | ( n4185 & ~n11406 ) ;
  assign n11408 = n11407 ^ n4487 ^ n824 ;
  assign n11409 = n11408 ^ n7130 ^ 1'b0 ;
  assign n11410 = n10016 & ~n11409 ;
  assign n11411 = n2256 & n2465 ;
  assign n11412 = n11411 ^ n5212 ^ 1'b0 ;
  assign n11422 = n2705 ^ n1917 ^ 1'b0 ;
  assign n11423 = ~n9364 & n11422 ;
  assign n11420 = n1292 & ~n1782 ;
  assign n11421 = n11420 ^ n2826 ^ 1'b0 ;
  assign n11416 = n8994 ^ n7218 ^ 1'b0 ;
  assign n11417 = n9662 & n11416 ;
  assign n11418 = n11417 ^ n5316 ^ 1'b0 ;
  assign n11413 = n2510 ^ n1782 ^ 1'b0 ;
  assign n11414 = n4127 & ~n11413 ;
  assign n11415 = ~n8955 & n11414 ;
  assign n11419 = n11418 ^ n11415 ^ 1'b0 ;
  assign n11424 = n11423 ^ n11421 ^ n11419 ;
  assign n11425 = n7559 & ~n10449 ;
  assign n11426 = n6442 | n6792 ;
  assign n11427 = n3596 & ~n11426 ;
  assign n11428 = n11427 ^ n10418 ^ 1'b0 ;
  assign n11429 = n1739 & n8122 ;
  assign n11430 = n7718 | n11429 ;
  assign n11431 = n1564 & n11430 ;
  assign n11432 = n11431 ^ n8214 ^ n3211 ;
  assign n11433 = n11432 ^ n8377 ^ 1'b0 ;
  assign n11434 = ~n9913 & n11433 ;
  assign n11435 = n7229 ^ n7025 ^ 1'b0 ;
  assign n11436 = n11435 ^ n2859 ^ n247 ;
  assign n11437 = n1265 | n5145 ;
  assign n11438 = n1530 | n11437 ;
  assign n11440 = n10099 ^ n6717 ^ 1'b0 ;
  assign n11439 = n1191 & n9984 ;
  assign n11441 = n11440 ^ n11439 ^ 1'b0 ;
  assign n11442 = n4749 & ~n10261 ;
  assign n11443 = n11442 ^ n4439 ^ 1'b0 ;
  assign n11444 = ~n1666 & n1867 ;
  assign n11445 = n11444 ^ n11327 ^ 1'b0 ;
  assign n11446 = n2487 & n4058 ;
  assign n11447 = n11446 ^ n1181 ^ 1'b0 ;
  assign n11448 = n7685 | n11447 ;
  assign n11449 = n7615 ^ n2057 ^ 1'b0 ;
  assign n11450 = n11449 ^ n177 ^ 1'b0 ;
  assign n11451 = ~n5539 & n7726 ;
  assign n11452 = ~n1775 & n11451 ;
  assign n11453 = ( n254 & ~n1751 ) | ( n254 & n2985 ) | ( ~n1751 & n2985 ) ;
  assign n11454 = ~n1809 & n8175 ;
  assign n11455 = ( n10041 & ~n11453 ) | ( n10041 & n11454 ) | ( ~n11453 & n11454 ) ;
  assign n11459 = n517 & n2199 ;
  assign n11460 = n11459 ^ n5863 ^ n4813 ;
  assign n11457 = n2953 | n4202 ;
  assign n11456 = n623 | n9131 ;
  assign n11458 = n11457 ^ n11456 ^ 1'b0 ;
  assign n11461 = n11460 ^ n11458 ^ n4035 ;
  assign n11462 = n1692 | n6503 ;
  assign n11463 = n11462 ^ n2719 ^ 1'b0 ;
  assign n11464 = n11463 ^ n10111 ^ n8669 ;
  assign n11467 = ( n1686 & ~n4752 ) | ( n1686 & n8007 ) | ( ~n4752 & n8007 ) ;
  assign n11465 = n1292 ^ n551 ^ 1'b0 ;
  assign n11466 = n6448 & ~n11465 ;
  assign n11468 = n11467 ^ n11466 ^ n9030 ;
  assign n11469 = n4181 ^ n3414 ^ 1'b0 ;
  assign n11470 = n11469 ^ n4895 ^ 1'b0 ;
  assign n11471 = n1125 & ~n11470 ;
  assign n11474 = n5857 ^ n1123 ^ 1'b0 ;
  assign n11475 = n386 & ~n11474 ;
  assign n11473 = ~n3757 & n5620 ;
  assign n11476 = n11475 ^ n11473 ^ 1'b0 ;
  assign n11472 = n1762 & ~n5746 ;
  assign n11477 = n11476 ^ n11472 ^ 1'b0 ;
  assign n11478 = n11471 & n11477 ;
  assign n11479 = ~n11468 & n11478 ;
  assign n11480 = n8765 & ~n10100 ;
  assign n11481 = n11479 & n11480 ;
  assign n11482 = n6703 ^ n2772 ^ 1'b0 ;
  assign n11483 = n8191 ^ n4204 ^ n324 ;
  assign n11484 = n3173 & n11483 ;
  assign n11485 = n11482 & n11484 ;
  assign n11486 = n6712 & n10356 ;
  assign n11487 = n7882 & n8222 ;
  assign n11488 = n11486 & n11487 ;
  assign n11489 = n2447 & n2926 ;
  assign n11490 = n3047 & n3660 ;
  assign n11491 = ( n2465 & n7438 ) | ( n2465 & ~n11490 ) | ( n7438 & ~n11490 ) ;
  assign n11492 = n11274 ^ n7001 ^ 1'b0 ;
  assign n11493 = n4362 & ~n5316 ;
  assign n11494 = n8428 | n11493 ;
  assign n11495 = n1244 | n11494 ;
  assign n11496 = n671 & n738 ;
  assign n11497 = n11496 ^ n1387 ^ 1'b0 ;
  assign n11498 = ~n3492 & n10482 ;
  assign n11499 = n11102 & n11498 ;
  assign n11500 = n11499 ^ n4651 ^ 1'b0 ;
  assign n11501 = ~n811 & n3185 ;
  assign n11505 = n3656 ^ n1564 ^ 1'b0 ;
  assign n11502 = n5953 & n9402 ;
  assign n11503 = n11502 ^ n3304 ^ 1'b0 ;
  assign n11504 = ~n346 & n11503 ;
  assign n11506 = n11505 ^ n11504 ^ 1'b0 ;
  assign n11507 = n3350 ^ n2448 ^ 1'b0 ;
  assign n11508 = n1416 & ~n11507 ;
  assign n11509 = n11508 ^ n1101 ^ 1'b0 ;
  assign n11510 = n3708 & ~n4455 ;
  assign n11511 = n11510 ^ n630 ^ 1'b0 ;
  assign n11512 = n6687 ^ n5968 ^ 1'b0 ;
  assign n11513 = n11391 | n11512 ;
  assign n11514 = ~n6073 & n11513 ;
  assign n11515 = n2119 | n4325 ;
  assign n11516 = n6717 ^ n4110 ^ n2831 ;
  assign n11517 = n11516 ^ n1829 ^ n1059 ;
  assign n11518 = ( n1168 & n1526 ) | ( n1168 & ~n1535 ) | ( n1526 & ~n1535 ) ;
  assign n11519 = n2118 & n11518 ;
  assign n11520 = n5535 & n11519 ;
  assign n11521 = n7385 & n11520 ;
  assign n11522 = n9333 ^ n1475 ^ 1'b0 ;
  assign n11524 = n9787 ^ n5298 ^ n2312 ;
  assign n11523 = n6616 & ~n7971 ;
  assign n11525 = n11524 ^ n11523 ^ 1'b0 ;
  assign n11526 = n9863 & ~n10827 ;
  assign n11527 = n3821 & n8300 ;
  assign n11528 = n11527 ^ n9496 ^ 1'b0 ;
  assign n11529 = n11528 ^ n9593 ^ 1'b0 ;
  assign n11530 = n5247 ^ n4468 ^ n1040 ;
  assign n11531 = n4261 ^ n1706 ^ 1'b0 ;
  assign n11532 = n4064 & n11531 ;
  assign n11533 = ( n7171 & n11530 ) | ( n7171 & n11532 ) | ( n11530 & n11532 ) ;
  assign n11534 = n1003 | n8214 ;
  assign n11535 = n11534 ^ n188 ^ 1'b0 ;
  assign n11536 = n3728 & ~n11535 ;
  assign n11538 = n9908 & ~n10733 ;
  assign n11539 = n11538 ^ n5450 ^ 1'b0 ;
  assign n11537 = ~n2020 & n10738 ;
  assign n11540 = n11539 ^ n11537 ^ 1'b0 ;
  assign n11541 = n6753 | n11084 ;
  assign n11542 = n11540 & ~n11541 ;
  assign n11543 = n10809 & ~n11058 ;
  assign n11544 = ~n9540 & n11543 ;
  assign n11545 = n2510 & ~n11544 ;
  assign n11546 = ~n9435 & n11545 ;
  assign n11547 = n4750 ^ n1452 ^ n1266 ;
  assign n11548 = n11547 ^ n1425 ^ 1'b0 ;
  assign n11554 = n189 | n3130 ;
  assign n11550 = n7189 ^ n2147 ^ 1'b0 ;
  assign n11551 = n3644 & ~n11550 ;
  assign n11552 = n9243 & n11551 ;
  assign n11553 = n11552 ^ n6777 ^ 1'b0 ;
  assign n11549 = ( n1286 & ~n4078 ) | ( n1286 & n5778 ) | ( ~n4078 & n5778 ) ;
  assign n11555 = n11554 ^ n11553 ^ n11549 ;
  assign n11556 = ~n967 & n11122 ;
  assign n11557 = n3440 ^ n3287 ^ n681 ;
  assign n11558 = n11557 ^ n8914 ^ 1'b0 ;
  assign n11559 = n11556 & n11558 ;
  assign n11560 = ~n4648 & n11559 ;
  assign n11561 = n11560 ^ n809 ^ 1'b0 ;
  assign n11562 = n630 & n8834 ;
  assign n11563 = ~n6050 & n11562 ;
  assign n11564 = ( ~n5680 & n9830 ) | ( ~n5680 & n11563 ) | ( n9830 & n11563 ) ;
  assign n11565 = n5207 | n7503 ;
  assign n11566 = n3036 | n3933 ;
  assign n11567 = n11566 ^ n3199 ^ 1'b0 ;
  assign n11568 = n4946 & ~n11567 ;
  assign n11569 = ~n9988 & n11568 ;
  assign n11570 = n11287 & n11569 ;
  assign n11571 = n7890 & n9063 ;
  assign n11572 = ~n964 & n11571 ;
  assign n11573 = n6311 & n9908 ;
  assign n11574 = ~n2622 & n11573 ;
  assign n11575 = n2690 | n10127 ;
  assign n11576 = ( n5717 & ~n11574 ) | ( n5717 & n11575 ) | ( ~n11574 & n11575 ) ;
  assign n11578 = ~n1207 & n8637 ;
  assign n11579 = n11578 ^ n1949 ^ 1'b0 ;
  assign n11577 = n1048 | n9507 ;
  assign n11580 = n11579 ^ n11577 ^ 1'b0 ;
  assign n11581 = n9771 & ~n11580 ;
  assign n11582 = n11581 ^ n7093 ^ x76 ;
  assign n11583 = n2260 & n7462 ;
  assign n11584 = n11583 ^ x118 ^ 1'b0 ;
  assign n11585 = n11584 ^ n2073 ^ 1'b0 ;
  assign n11586 = ( x69 & ~x103 ) | ( x69 & n2652 ) | ( ~x103 & n2652 ) ;
  assign n11587 = ~n729 & n2366 ;
  assign n11588 = n6106 ^ n5691 ^ 1'b0 ;
  assign n11589 = n11587 & n11588 ;
  assign n11590 = n9193 & n11589 ;
  assign n11591 = n11586 & n11590 ;
  assign n11592 = ( ~n5218 & n5303 ) | ( ~n5218 & n7355 ) | ( n5303 & n7355 ) ;
  assign n11593 = n3253 & ~n11021 ;
  assign n11594 = n11592 & n11593 ;
  assign n11595 = n3652 | n7673 ;
  assign n11596 = n5114 ^ n1762 ^ 1'b0 ;
  assign n11597 = n6201 & ~n11596 ;
  assign n11598 = n11597 ^ n149 ^ 1'b0 ;
  assign n11599 = ~n4124 & n11598 ;
  assign n11600 = n234 | n11599 ;
  assign n11601 = n2671 ^ n581 ^ 1'b0 ;
  assign n11602 = n1414 & ~n11601 ;
  assign n11603 = n5352 ^ n621 ^ 1'b0 ;
  assign n11604 = ~n1420 & n11603 ;
  assign n11605 = n11604 ^ n8282 ^ n869 ;
  assign n11606 = n10039 ^ n6053 ^ x13 ;
  assign n11607 = n8953 ^ n7235 ^ n5057 ;
  assign n11608 = n3673 & ~n11607 ;
  assign n11609 = n11608 ^ n2471 ^ 1'b0 ;
  assign n11610 = n4023 ^ n1095 ^ 1'b0 ;
  assign n11611 = ~n2702 & n11610 ;
  assign n11612 = n11611 ^ n10923 ^ n6092 ;
  assign n11613 = n508 | n8150 ;
  assign n11614 = n11613 ^ n1594 ^ 1'b0 ;
  assign n11615 = n617 | n10707 ;
  assign n11616 = n11615 ^ n11235 ^ 1'b0 ;
  assign n11617 = ~n11614 & n11616 ;
  assign n11618 = n5926 ^ n1059 ^ 1'b0 ;
  assign n11619 = ~n2864 & n11618 ;
  assign n11620 = n11619 ^ n5918 ^ 1'b0 ;
  assign n11621 = ~n4903 & n11620 ;
  assign n11622 = n8422 & n11621 ;
  assign n11623 = n4717 ^ n3340 ^ 1'b0 ;
  assign n11624 = n11622 | n11623 ;
  assign n11625 = n1286 | n3557 ;
  assign n11626 = n4014 ^ x13 ^ 1'b0 ;
  assign n11627 = n11625 & ~n11626 ;
  assign n11628 = n4246 & n11627 ;
  assign n11629 = n11628 ^ n1912 ^ n1560 ;
  assign n11630 = n872 & n5938 ;
  assign n11631 = n4479 & n11630 ;
  assign n11632 = n11631 ^ n10961 ^ 1'b0 ;
  assign n11633 = n7546 ^ n1385 ^ n1171 ;
  assign n11634 = n10031 | n11633 ;
  assign n11635 = n11632 & ~n11634 ;
  assign n11636 = n5734 | n9371 ;
  assign n11637 = n2746 | n9830 ;
  assign n11639 = ( ~n1458 & n1920 ) | ( ~n1458 & n2871 ) | ( n1920 & n2871 ) ;
  assign n11638 = n799 & ~n2489 ;
  assign n11640 = n11639 ^ n11638 ^ 1'b0 ;
  assign n11641 = n11637 | n11640 ;
  assign n11642 = n5149 ^ n3025 ^ 1'b0 ;
  assign n11643 = ~n8597 & n11642 ;
  assign n11644 = ( n1743 & n9180 ) | ( n1743 & ~n10939 ) | ( n9180 & ~n10939 ) ;
  assign n11645 = n2540 & n3236 ;
  assign n11646 = n11645 ^ n5556 ^ 1'b0 ;
  assign n11647 = n8745 & ~n11646 ;
  assign n11648 = n245 & n11647 ;
  assign n11649 = n11648 ^ n1397 ^ 1'b0 ;
  assign n11650 = n9369 | n10026 ;
  assign n11651 = n212 | n11650 ;
  assign n11652 = n6786 & ~n9426 ;
  assign n11653 = n6141 & n11652 ;
  assign n11654 = n5199 | n11653 ;
  assign n11655 = n5349 & ~n11654 ;
  assign n11656 = n359 & ~n3531 ;
  assign n11657 = n826 & ~n11312 ;
  assign n11658 = n11656 & n11657 ;
  assign n11659 = x62 & x117 ;
  assign n11662 = n6047 ^ n4297 ^ n3587 ;
  assign n11660 = ~n148 & n812 ;
  assign n11661 = n7719 & ~n11660 ;
  assign n11663 = n11662 ^ n11661 ^ 1'b0 ;
  assign n11664 = n619 & ~n2236 ;
  assign n11665 = ~n7136 & n11664 ;
  assign n11666 = n3325 ^ n416 ^ 1'b0 ;
  assign n11667 = n6523 & n7847 ;
  assign n11668 = n3139 ^ n3006 ^ 1'b0 ;
  assign n11669 = n11668 ^ n1236 ^ 1'b0 ;
  assign n11670 = n8298 ^ n6925 ^ n2160 ;
  assign n11671 = ~n11669 & n11670 ;
  assign n11672 = n10729 ^ n10288 ^ 1'b0 ;
  assign n11673 = n10855 & n11672 ;
  assign n11675 = ( n1309 & n2464 ) | ( n1309 & ~n2589 ) | ( n2464 & ~n2589 ) ;
  assign n11676 = ( n2503 & ~n7345 ) | ( n2503 & n11675 ) | ( ~n7345 & n11675 ) ;
  assign n11674 = ~n2642 & n4660 ;
  assign n11677 = n11676 ^ n11674 ^ 1'b0 ;
  assign n11678 = n2726 | n3325 ;
  assign n11679 = n4292 | n11678 ;
  assign n11680 = n11679 ^ n7762 ^ n5330 ;
  assign n11681 = n4850 ^ n4620 ^ n3155 ;
  assign n11682 = n5256 ^ x73 ^ 1'b0 ;
  assign n11683 = n3904 & ~n11682 ;
  assign n11684 = ~n3681 & n7918 ;
  assign n11685 = n11684 ^ x17 ^ 1'b0 ;
  assign n11686 = n11387 ^ n1869 ^ 1'b0 ;
  assign n11687 = n3192 & n11686 ;
  assign n11688 = n5922 & n11687 ;
  assign n11689 = n1451 | n3193 ;
  assign n11690 = n11689 ^ n516 ^ 1'b0 ;
  assign n11691 = ( ~n3380 & n9110 ) | ( ~n3380 & n11690 ) | ( n9110 & n11690 ) ;
  assign n11692 = n4915 ^ n4211 ^ 1'b0 ;
  assign n11693 = n11691 | n11692 ;
  assign n11694 = n11693 ^ n10002 ^ 1'b0 ;
  assign n11699 = ( n1269 & n4440 ) | ( n1269 & n10549 ) | ( n4440 & n10549 ) ;
  assign n11696 = n5548 | n6363 ;
  assign n11697 = n11696 ^ n265 ^ 1'b0 ;
  assign n11698 = n7962 & n11697 ;
  assign n11695 = n2837 | n3538 ;
  assign n11700 = n11699 ^ n11698 ^ n11695 ;
  assign n11701 = n5027 & ~n6182 ;
  assign n11702 = n1566 ^ n486 ^ 1'b0 ;
  assign n11703 = n11702 ^ x118 ^ 1'b0 ;
  assign n11704 = n6251 & ~n11703 ;
  assign n11705 = n3063 & ~n9821 ;
  assign n11706 = n5548 & n11705 ;
  assign n11707 = ( ~n3366 & n10530 ) | ( ~n3366 & n11706 ) | ( n10530 & n11706 ) ;
  assign n11708 = n2505 & n4164 ;
  assign n11709 = ~n5437 & n11708 ;
  assign n11710 = n5802 ^ n663 ^ 1'b0 ;
  assign n11711 = n944 & n11710 ;
  assign n11712 = n11711 ^ n1693 ^ 1'b0 ;
  assign n11713 = ( n1869 & ~n2551 ) | ( n1869 & n9144 ) | ( ~n2551 & n9144 ) ;
  assign n11714 = ~n469 & n11713 ;
  assign n11715 = ( n3697 & n11712 ) | ( n3697 & n11714 ) | ( n11712 & n11714 ) ;
  assign n11716 = n11709 & n11715 ;
  assign n11717 = n7003 ^ n5528 ^ 1'b0 ;
  assign n11718 = n8768 | n11717 ;
  assign n11719 = ( n3958 & n8389 ) | ( n3958 & n11486 ) | ( n8389 & n11486 ) ;
  assign n11720 = n11432 ^ n9747 ^ 1'b0 ;
  assign n11721 = n6335 | n11720 ;
  assign n11722 = n387 & ~n840 ;
  assign n11723 = n1291 & n11722 ;
  assign n11724 = ~n5255 & n11569 ;
  assign n11725 = n11723 & n11724 ;
  assign n11726 = ~n2484 & n9276 ;
  assign n11727 = n2484 & n11726 ;
  assign n11728 = n1387 ^ n167 ^ 1'b0 ;
  assign n11729 = n6979 & ~n11728 ;
  assign n11730 = n11729 ^ n8150 ^ 1'b0 ;
  assign n11731 = n5680 | n11730 ;
  assign n11732 = n5410 & ~n11731 ;
  assign n11733 = n11727 & n11732 ;
  assign n11734 = n11733 ^ n7713 ^ 1'b0 ;
  assign n11735 = ~x13 & n11734 ;
  assign n11736 = n1504 & n8960 ;
  assign n11737 = n11165 ^ n765 ^ 1'b0 ;
  assign n11738 = n11737 ^ n8991 ^ 1'b0 ;
  assign n11739 = n11736 | n11738 ;
  assign n11740 = n11739 ^ n4113 ^ 1'b0 ;
  assign n11741 = ~n3842 & n11740 ;
  assign n11742 = n5680 & n9617 ;
  assign n11743 = ~n5118 & n11742 ;
  assign n11744 = n3892 | n4919 ;
  assign n11745 = n11744 ^ x70 ^ 1'b0 ;
  assign n11746 = n11745 ^ n4466 ^ 1'b0 ;
  assign n11747 = ~n6063 & n7318 ;
  assign n11748 = ( n314 & n2165 ) | ( n314 & ~n5737 ) | ( n2165 & ~n5737 ) ;
  assign n11749 = n3754 ^ n197 ^ 1'b0 ;
  assign n11750 = ~n8720 & n9999 ;
  assign n11751 = ( ~n4760 & n11207 ) | ( ~n4760 & n11750 ) | ( n11207 & n11750 ) ;
  assign n11752 = n9926 ^ n1677 ^ 1'b0 ;
  assign n11753 = n11752 ^ n8009 ^ n2389 ;
  assign n11754 = n1605 | n6868 ;
  assign n11755 = n7461 & ~n11754 ;
  assign n11756 = ~n10266 & n11755 ;
  assign n11757 = n10504 ^ x48 ^ 1'b0 ;
  assign n11758 = n3835 & ~n11757 ;
  assign n11759 = n11087 ^ n4257 ^ 1'b0 ;
  assign n11760 = n9335 ^ n8441 ^ n5573 ;
  assign n11761 = n1017 | n2313 ;
  assign n11762 = ~n5101 & n6245 ;
  assign n11763 = n882 | n1658 ;
  assign n11764 = n11763 ^ n812 ^ 1'b0 ;
  assign n11765 = n11762 & n11764 ;
  assign n11766 = n4813 ^ n2658 ^ 1'b0 ;
  assign n11767 = ~n6719 & n11766 ;
  assign n11768 = ( n1394 & n3551 ) | ( n1394 & n11767 ) | ( n3551 & n11767 ) ;
  assign n11769 = n10356 & n11768 ;
  assign n11770 = n11769 ^ n5765 ^ 1'b0 ;
  assign n11771 = n509 & ~n11770 ;
  assign n11772 = n3438 | n3950 ;
  assign n11773 = ~n8479 & n9344 ;
  assign n11774 = n2956 & n11773 ;
  assign n11782 = n5382 ^ n335 ^ 1'b0 ;
  assign n11783 = n3195 & n11782 ;
  assign n11775 = n4095 & n9513 ;
  assign n11776 = n4966 & n11775 ;
  assign n11777 = n4654 & n11217 ;
  assign n11778 = n11777 ^ n10293 ^ 1'b0 ;
  assign n11779 = n11778 ^ n10751 ^ 1'b0 ;
  assign n11780 = n2206 & n11779 ;
  assign n11781 = n11776 & n11780 ;
  assign n11784 = n11783 ^ n11781 ^ 1'b0 ;
  assign n11785 = ~n7347 & n11784 ;
  assign n11786 = n1327 & n1342 ;
  assign n11787 = n5010 ^ x60 ^ 1'b0 ;
  assign n11788 = n4331 | n11787 ;
  assign n11789 = n11786 | n11788 ;
  assign n11790 = n6353 ^ n4655 ^ 1'b0 ;
  assign n11791 = n3113 | n11790 ;
  assign n11792 = n3178 | n3797 ;
  assign n11793 = n1243 & ~n8512 ;
  assign n11794 = ~n1083 & n11793 ;
  assign n11795 = n11794 ^ n2980 ^ 1'b0 ;
  assign n11796 = n1251 & ~n11795 ;
  assign n11797 = n4237 & n11796 ;
  assign n11798 = n11797 ^ n4820 ^ 1'b0 ;
  assign n11799 = n9374 ^ n4625 ^ n3439 ;
  assign n11800 = n6422 & n11799 ;
  assign n11801 = n11800 ^ n633 ^ 1'b0 ;
  assign n11802 = n10961 & ~n11801 ;
  assign n11803 = n2104 & ~n3934 ;
  assign n11804 = ( n3073 & n3185 ) | ( n3073 & ~n8050 ) | ( n3185 & ~n8050 ) ;
  assign n11805 = n1596 & ~n1943 ;
  assign n11806 = n897 & ~n11805 ;
  assign n11807 = n11804 & n11806 ;
  assign n11813 = ~n3948 & n5486 ;
  assign n11808 = n2253 ^ n895 ^ 1'b0 ;
  assign n11809 = ( n785 & ~n917 ) | ( n785 & n11808 ) | ( ~n917 & n11808 ) ;
  assign n11810 = n11809 ^ n5355 ^ 1'b0 ;
  assign n11811 = ~n8645 & n11810 ;
  assign n11812 = ~n10145 & n11811 ;
  assign n11814 = n11813 ^ n11812 ^ n10219 ;
  assign n11815 = n4594 | n6868 ;
  assign n11816 = n9476 ^ n1791 ^ 1'b0 ;
  assign n11817 = n7979 | n11816 ;
  assign n11818 = ~n975 & n2463 ;
  assign n11819 = n7200 & ~n8289 ;
  assign n11820 = n10738 & n11819 ;
  assign n11821 = n5963 & n11820 ;
  assign n11822 = ~n1122 & n10628 ;
  assign n11823 = n8332 & n11822 ;
  assign n11824 = x126 & n2823 ;
  assign n11825 = n4055 & n11824 ;
  assign n11826 = n11825 ^ n3609 ^ 1'b0 ;
  assign n11827 = n7181 | n11826 ;
  assign n11828 = n10978 ^ n4165 ^ 1'b0 ;
  assign n11829 = ( n474 & n5573 ) | ( n474 & ~n10200 ) | ( n5573 & ~n10200 ) ;
  assign n11830 = n7123 & ~n8035 ;
  assign n11831 = n190 | n2125 ;
  assign n11832 = n11831 ^ n9477 ^ n1746 ;
  assign n11833 = n11830 & n11832 ;
  assign n11834 = n3288 & ~n11833 ;
  assign n11835 = n11834 ^ n8729 ^ 1'b0 ;
  assign n11836 = n5420 ^ n4102 ^ 1'b0 ;
  assign n11837 = n7729 ^ n6728 ^ 1'b0 ;
  assign n11838 = n11836 & ~n11837 ;
  assign n11839 = ~n6257 & n10996 ;
  assign n11840 = n11839 ^ n11817 ^ 1'b0 ;
  assign n11841 = n8055 ^ n3317 ^ 1'b0 ;
  assign n11842 = ~n10750 & n11841 ;
  assign n11843 = n4498 & ~n5485 ;
  assign n11844 = ( n8512 & n8776 ) | ( n8512 & ~n9972 ) | ( n8776 & ~n9972 ) ;
  assign n11845 = n4164 & n5960 ;
  assign n11846 = n11845 ^ n4510 ^ 1'b0 ;
  assign n11847 = ( n1044 & n1427 ) | ( n1044 & n11846 ) | ( n1427 & n11846 ) ;
  assign n11848 = ~n3393 & n11847 ;
  assign n11849 = ~n8994 & n11848 ;
  assign n11850 = ( n3412 & n6452 ) | ( n3412 & ~n8005 ) | ( n6452 & ~n8005 ) ;
  assign n11851 = n11850 ^ n7389 ^ n4459 ;
  assign n11853 = n4898 ^ n871 ^ 1'b0 ;
  assign n11854 = n7850 | n11853 ;
  assign n11852 = ( n513 & n778 ) | ( n513 & n1108 ) | ( n778 & n1108 ) ;
  assign n11855 = n11854 ^ n11852 ^ 1'b0 ;
  assign n11856 = n5059 | n11855 ;
  assign n11859 = n6134 ^ n944 ^ 1'b0 ;
  assign n11857 = n11180 ^ n4553 ^ 1'b0 ;
  assign n11858 = n8862 & ~n11857 ;
  assign n11860 = n11859 ^ n11858 ^ n3199 ;
  assign n11861 = n11860 ^ n3379 ^ 1'b0 ;
  assign n11866 = n5834 ^ n5603 ^ n5535 ;
  assign n11867 = n2775 & n11866 ;
  assign n11868 = ~n8956 & n11867 ;
  assign n11862 = n4915 & n5790 ;
  assign n11863 = ~n336 & n11862 ;
  assign n11864 = n11863 ^ n6566 ^ 1'b0 ;
  assign n11865 = n505 & n11864 ;
  assign n11869 = n11868 ^ n11865 ^ 1'b0 ;
  assign n11870 = n1849 & ~n11869 ;
  assign n11871 = n11870 ^ n4050 ^ 1'b0 ;
  assign n11872 = n11861 & ~n11871 ;
  assign n11873 = n8427 ^ n8107 ^ 1'b0 ;
  assign n11874 = x52 & ~n11873 ;
  assign n11875 = n8044 ^ n1710 ^ 1'b0 ;
  assign n11876 = x126 & ~n762 ;
  assign n11877 = ~n5785 & n11876 ;
  assign n11878 = ~n1229 & n7120 ;
  assign n11879 = n11878 ^ n8141 ^ 1'b0 ;
  assign n11880 = n9056 | n11879 ;
  assign n11882 = ~n4839 & n7434 ;
  assign n11881 = n5606 ^ n3886 ^ 1'b0 ;
  assign n11883 = n11882 ^ n11881 ^ n6900 ;
  assign n11884 = ~n5067 & n11883 ;
  assign n11885 = n11884 ^ n5396 ^ 1'b0 ;
  assign n11886 = n11530 ^ n1796 ^ 1'b0 ;
  assign n11887 = ~n1459 & n4023 ;
  assign n11888 = n11887 ^ n6118 ^ 1'b0 ;
  assign n11889 = n4216 | n11888 ;
  assign n11890 = n11889 ^ n11469 ^ 1'b0 ;
  assign n11892 = n1739 & n2214 ;
  assign n11893 = n11892 ^ n3668 ^ 1'b0 ;
  assign n11891 = n10455 & n10959 ;
  assign n11894 = n11893 ^ n11891 ^ 1'b0 ;
  assign n11895 = n7958 & n10701 ;
  assign n11896 = n11895 ^ n8966 ^ 1'b0 ;
  assign n11897 = n2927 | n4122 ;
  assign n11898 = n11897 ^ n654 ^ 1'b0 ;
  assign n11899 = n2317 & n2605 ;
  assign n11900 = n11898 & n11899 ;
  assign n11901 = ~n8425 & n11900 ;
  assign n11902 = n11901 ^ n418 ^ 1'b0 ;
  assign n11903 = x122 & n11203 ;
  assign n11904 = n7489 ^ n1617 ^ 1'b0 ;
  assign n11905 = n11903 & n11904 ;
  assign n11906 = n575 & ~n8378 ;
  assign n11907 = n11905 & n11906 ;
  assign n11908 = ~n6333 & n11907 ;
  assign n11909 = n2956 | n11908 ;
  assign n11910 = n11909 ^ n5031 ^ 1'b0 ;
  assign n11911 = n11910 ^ n7506 ^ 1'b0 ;
  assign n11912 = n910 & n11911 ;
  assign n11913 = n262 & n5190 ;
  assign n11914 = n11913 ^ n3619 ^ 1'b0 ;
  assign n11915 = n4670 | n11914 ;
  assign n11916 = n7521 ^ n6461 ^ 1'b0 ;
  assign n11917 = ~n11436 & n11916 ;
  assign n11918 = n5058 ^ n3424 ^ 1'b0 ;
  assign n11919 = ~n1044 & n11918 ;
  assign n11920 = ~n2014 & n11919 ;
  assign n11921 = n2379 & ~n2860 ;
  assign n11922 = ( n8512 & ~n10583 ) | ( n8512 & n11921 ) | ( ~n10583 & n11921 ) ;
  assign n11923 = n5169 | n11330 ;
  assign n11924 = n4559 & ~n11923 ;
  assign n11925 = ~n1542 & n2678 ;
  assign n11928 = n2443 ^ n1853 ^ 1'b0 ;
  assign n11929 = n1186 & n11928 ;
  assign n11930 = n3617 | n11929 ;
  assign n11931 = n11930 ^ n3961 ^ 1'b0 ;
  assign n11932 = n11931 ^ n8584 ^ 1'b0 ;
  assign n11933 = n593 & ~n11932 ;
  assign n11926 = ~n2219 & n6909 ;
  assign n11927 = ~n7174 & n11926 ;
  assign n11934 = n11933 ^ n11927 ^ n1435 ;
  assign n11935 = n11934 ^ n510 ^ 1'b0 ;
  assign n11936 = n4667 ^ n1589 ^ 1'b0 ;
  assign n11937 = n11935 & n11936 ;
  assign n11938 = n11066 ^ n10772 ^ 1'b0 ;
  assign n11939 = n2981 & ~n11938 ;
  assign n11940 = ( n3455 & n9908 ) | ( n3455 & ~n11939 ) | ( n9908 & ~n11939 ) ;
  assign n11941 = n2809 ^ n381 ^ 1'b0 ;
  assign n11942 = n3291 & n11872 ;
  assign n11948 = n2605 ^ x66 ^ 1'b0 ;
  assign n11949 = ( n5118 & n7416 ) | ( n5118 & ~n11948 ) | ( n7416 & ~n11948 ) ;
  assign n11943 = n6257 ^ n1308 ^ 1'b0 ;
  assign n11944 = n4327 & n11943 ;
  assign n11945 = n11944 ^ n5755 ^ n2969 ;
  assign n11946 = n11945 ^ n5089 ^ 1'b0 ;
  assign n11947 = n7368 & ~n11946 ;
  assign n11950 = n11949 ^ n11947 ^ 1'b0 ;
  assign n11951 = n8927 ^ n7988 ^ 1'b0 ;
  assign n11953 = n8185 ^ n7103 ^ 1'b0 ;
  assign n11952 = n2676 & ~n7044 ;
  assign n11954 = n11953 ^ n11952 ^ 1'b0 ;
  assign n11955 = ~n2349 & n11954 ;
  assign n11956 = n10772 ^ n3732 ^ 1'b0 ;
  assign n11957 = n3366 | n11956 ;
  assign n11958 = n8032 & ~n11957 ;
  assign n11959 = n11958 ^ n9489 ^ 1'b0 ;
  assign n11960 = n10138 ^ n3808 ^ 1'b0 ;
  assign n11961 = n4601 & n4669 ;
  assign n11962 = n7103 ^ n1044 ^ 1'b0 ;
  assign n11963 = n11962 ^ n11635 ^ 1'b0 ;
  assign n11964 = n7615 & n11963 ;
  assign n11966 = ( ~n265 & n1637 ) | ( ~n265 & n1944 ) | ( n1637 & n1944 ) ;
  assign n11965 = ~n1854 & n4394 ;
  assign n11967 = n11966 ^ n11965 ^ 1'b0 ;
  assign n11968 = n9153 ^ n1846 ^ 1'b0 ;
  assign n11969 = ~n5665 & n11968 ;
  assign n11970 = n11969 ^ n2940 ^ 1'b0 ;
  assign n11971 = n5274 ^ n935 ^ x97 ;
  assign n11972 = ( ~n7177 & n11364 ) | ( ~n7177 & n11971 ) | ( n11364 & n11971 ) ;
  assign n11973 = n4948 ^ n2551 ^ 1'b0 ;
  assign n11974 = ~n3785 & n6026 ;
  assign n11975 = n11973 & n11974 ;
  assign n11976 = n10010 ^ n6279 ^ 1'b0 ;
  assign n11977 = n1000 | n3297 ;
  assign n11978 = n9822 ^ n6667 ^ 1'b0 ;
  assign n11979 = ~n633 & n8572 ;
  assign n11980 = n11978 & n11979 ;
  assign n11981 = n11980 ^ n256 ^ 1'b0 ;
  assign n11982 = n11284 ^ n217 ^ 1'b0 ;
  assign n11985 = ( n2107 & n4054 ) | ( n2107 & ~n8295 ) | ( n4054 & ~n8295 ) ;
  assign n11986 = n4812 & n11985 ;
  assign n11983 = n4721 ^ n1033 ^ 1'b0 ;
  assign n11984 = n4376 | n11983 ;
  assign n11987 = n11986 ^ n11984 ^ 1'b0 ;
  assign n11988 = ~n7583 & n9684 ;
  assign n11989 = n7808 ^ n7420 ^ 1'b0 ;
  assign n11990 = ~n2506 & n11989 ;
  assign n11991 = n7361 ^ n4453 ^ 1'b0 ;
  assign n11992 = n5096 | n11991 ;
  assign n11993 = n8977 ^ n6253 ^ 1'b0 ;
  assign n11994 = n5376 ^ n3977 ^ 1'b0 ;
  assign n11995 = ~n11993 & n11994 ;
  assign n11996 = n2295 & ~n7101 ;
  assign n11997 = n11996 ^ n4285 ^ 1'b0 ;
  assign n11998 = ( n9814 & ~n11995 ) | ( n9814 & n11997 ) | ( ~n11995 & n11997 ) ;
  assign n12000 = n5539 ^ n1871 ^ n461 ;
  assign n11999 = n7085 & ~n10517 ;
  assign n12001 = n12000 ^ n11999 ^ 1'b0 ;
  assign n12002 = ~n696 & n12001 ;
  assign n12003 = ~n438 & n8120 ;
  assign n12004 = n1628 & ~n11079 ;
  assign n12005 = n3786 ^ n842 ^ 1'b0 ;
  assign n12006 = n1251 | n12005 ;
  assign n12007 = n12006 ^ n1944 ^ 1'b0 ;
  assign n12008 = n3721 & n12007 ;
  assign n12009 = n1246 & n7462 ;
  assign n12010 = n6248 ^ n4255 ^ 1'b0 ;
  assign n12011 = n5051 & ~n12010 ;
  assign n12012 = n5218 ^ x41 ^ 1'b0 ;
  assign n12013 = ~n12011 & n12012 ;
  assign n12014 = n8156 ^ n1258 ^ 1'b0 ;
  assign n12015 = n2915 | n9409 ;
  assign n12016 = n12015 ^ n11423 ^ 1'b0 ;
  assign n12017 = n558 | n5419 ;
  assign n12018 = n10198 ^ n9722 ^ 1'b0 ;
  assign n12019 = n5598 ^ n2933 ^ 1'b0 ;
  assign n12020 = n2540 & ~n3143 ;
  assign n12021 = ~n12019 & n12020 ;
  assign n12022 = n5730 & n12021 ;
  assign n12023 = n8615 ^ n5937 ^ 1'b0 ;
  assign n12024 = n11241 ^ n4197 ^ 1'b0 ;
  assign n12025 = n5281 ^ n588 ^ 1'b0 ;
  assign n12026 = ~n8084 & n12025 ;
  assign n12027 = n1181 & n12026 ;
  assign n12028 = n4876 & n6016 ;
  assign n12029 = n12027 & n12028 ;
  assign n12033 = n6195 & ~n6695 ;
  assign n12034 = ~x11 & n12033 ;
  assign n12031 = n1521 ^ n1374 ^ 1'b0 ;
  assign n12032 = ~n1461 & n12031 ;
  assign n12030 = n2280 & ~n4793 ;
  assign n12035 = n12034 ^ n12032 ^ n12030 ;
  assign n12036 = n11490 ^ n7707 ^ n2229 ;
  assign n12042 = n1312 & ~n6134 ;
  assign n12043 = n12042 ^ n1627 ^ 1'b0 ;
  assign n12037 = n5950 & ~n9682 ;
  assign n12038 = n9774 ^ n2083 ^ 1'b0 ;
  assign n12039 = ~n5530 & n12038 ;
  assign n12040 = ~n4111 & n12039 ;
  assign n12041 = n12037 | n12040 ;
  assign n12044 = n12043 ^ n12041 ^ 1'b0 ;
  assign n12045 = n5497 ^ n1775 ^ 1'b0 ;
  assign n12046 = n7497 ^ n3228 ^ 1'b0 ;
  assign n12047 = n4767 & ~n11031 ;
  assign n12048 = n12047 ^ n717 ^ 1'b0 ;
  assign n12049 = n12048 ^ n8340 ^ n7325 ;
  assign n12050 = n361 | n4570 ;
  assign n12051 = n12050 ^ n12034 ^ n182 ;
  assign n12053 = ~n3617 & n4020 ;
  assign n12054 = n12053 ^ n908 ^ 1'b0 ;
  assign n12052 = ~n5610 & n7896 ;
  assign n12055 = n12054 ^ n12052 ^ 1'b0 ;
  assign n12056 = n9589 ^ n2368 ^ 1'b0 ;
  assign n12057 = n12055 & n12056 ;
  assign n12058 = ~n3121 & n12057 ;
  assign n12059 = n794 ^ n399 ^ 1'b0 ;
  assign n12060 = n12058 & n12059 ;
  assign n12061 = n4448 ^ n1265 ^ n503 ;
  assign n12062 = n5475 ^ n450 ^ 1'b0 ;
  assign n12063 = n6816 & ~n12062 ;
  assign n12064 = x14 & ~n4867 ;
  assign n12065 = n12064 ^ n2994 ^ 1'b0 ;
  assign n12066 = n6698 | n9819 ;
  assign n12067 = ~n3431 & n12066 ;
  assign n12068 = ~n4146 & n4163 ;
  assign n12069 = n2755 ^ n1413 ^ 1'b0 ;
  assign n12070 = ~n12068 & n12069 ;
  assign n12071 = n11316 ^ n7425 ^ 1'b0 ;
  assign n12072 = n9209 ^ n1943 ^ 1'b0 ;
  assign n12073 = n4572 & ~n12072 ;
  assign n12074 = n2199 ^ n1998 ^ 1'b0 ;
  assign n12075 = n12074 ^ n10121 ^ 1'b0 ;
  assign n12076 = n12073 & n12075 ;
  assign n12077 = n8054 ^ n7930 ^ 1'b0 ;
  assign n12078 = ~n3020 & n3056 ;
  assign n12079 = ( n2932 & n9968 ) | ( n2932 & n12078 ) | ( n9968 & n12078 ) ;
  assign n12081 = n1689 & n3614 ;
  assign n12082 = n12081 ^ n11300 ^ n2485 ;
  assign n12080 = n5064 | n9896 ;
  assign n12083 = n12082 ^ n12080 ^ 1'b0 ;
  assign n12084 = n3519 & ~n4504 ;
  assign n12085 = n9630 ^ n2304 ^ n1860 ;
  assign n12086 = n4693 | n7692 ;
  assign n12087 = n1222 & n12086 ;
  assign n12088 = n190 & n12087 ;
  assign n12089 = n12088 ^ n2066 ^ 1'b0 ;
  assign n12090 = n3999 & n4988 ;
  assign n12091 = n2268 ^ n1440 ^ 1'b0 ;
  assign n12092 = n808 ^ n483 ^ 1'b0 ;
  assign n12093 = n12092 ^ n7806 ^ 1'b0 ;
  assign n12094 = n12091 & n12093 ;
  assign n12095 = ~n10464 & n12094 ;
  assign n12096 = ~n12090 & n12095 ;
  assign n12097 = n5565 | n9773 ;
  assign n12098 = n4368 ^ n3662 ^ x84 ;
  assign n12099 = n12098 ^ n2814 ^ 1'b0 ;
  assign n12100 = n4502 | n10854 ;
  assign n12101 = n9424 & ~n12100 ;
  assign n12106 = n6428 ^ n1952 ^ 1'b0 ;
  assign n12102 = n1703 & ~n2768 ;
  assign n12103 = n12102 ^ n2200 ^ 1'b0 ;
  assign n12104 = ~n9010 & n12103 ;
  assign n12105 = ~n4398 & n12104 ;
  assign n12107 = n12106 ^ n12105 ^ 1'b0 ;
  assign n12108 = n6878 & ~n8256 ;
  assign n12109 = n12108 ^ n10758 ^ 1'b0 ;
  assign n12110 = ( n796 & ~n11765 ) | ( n796 & n12109 ) | ( ~n11765 & n12109 ) ;
  assign n12111 = n6629 & n6849 ;
  assign n12112 = n12111 ^ n9514 ^ 1'b0 ;
  assign n12113 = n9466 ^ n1393 ^ 1'b0 ;
  assign n12114 = n6076 ^ n5371 ^ n176 ;
  assign n12115 = n9062 & ~n12114 ;
  assign n12116 = n4990 ^ n1724 ^ 1'b0 ;
  assign n12117 = ~n3328 & n12116 ;
  assign n12118 = n12117 ^ n7085 ^ 1'b0 ;
  assign n12119 = ~n9703 & n12118 ;
  assign n12120 = n1789 & ~n4358 ;
  assign n12121 = n8313 & n10032 ;
  assign n12122 = n9972 ^ n8157 ^ n6811 ;
  assign n12123 = n4050 | n10136 ;
  assign n12124 = n12123 ^ n1561 ^ 1'b0 ;
  assign n12125 = n1316 ^ n1021 ^ n642 ;
  assign n12126 = ( n3509 & n7114 ) | ( n3509 & ~n7186 ) | ( n7114 & ~n7186 ) ;
  assign n12127 = n327 | n8150 ;
  assign n12128 = n2299 & n12127 ;
  assign n12129 = n12128 ^ n2258 ^ 1'b0 ;
  assign n12130 = n9607 ^ n1660 ^ 1'b0 ;
  assign n12131 = x73 & n4000 ;
  assign n12132 = n12131 ^ n4915 ^ 1'b0 ;
  assign n12133 = n6996 | n9667 ;
  assign n12134 = ~n2956 & n7126 ;
  assign n12135 = ~n12133 & n12134 ;
  assign n12136 = n6778 ^ n2634 ^ 1'b0 ;
  assign n12137 = n5391 ^ n1075 ^ n1033 ;
  assign n12138 = n4886 | n5746 ;
  assign n12139 = n12138 ^ n9766 ^ 1'b0 ;
  assign n12140 = ( ~n452 & n3279 ) | ( ~n452 & n12139 ) | ( n3279 & n12139 ) ;
  assign n12141 = n1159 & ~n6555 ;
  assign n12142 = n3105 | n5770 ;
  assign n12143 = n12142 ^ n9412 ^ 1'b0 ;
  assign n12144 = n8295 & ~n9388 ;
  assign n12145 = ~n12143 & n12144 ;
  assign n12148 = n1373 & ~n4935 ;
  assign n12149 = n12148 ^ n1323 ^ 1'b0 ;
  assign n12150 = ~n4285 & n12149 ;
  assign n12146 = ~n5651 & n10384 ;
  assign n12147 = n12146 ^ n3710 ^ 1'b0 ;
  assign n12151 = n12150 ^ n12147 ^ 1'b0 ;
  assign n12152 = n2522 & ~n12151 ;
  assign n12156 = x77 & ~n403 ;
  assign n12157 = ~n2766 & n12156 ;
  assign n12153 = n9889 ^ n7163 ^ 1'b0 ;
  assign n12154 = n9090 | n12153 ;
  assign n12155 = n7819 & ~n12154 ;
  assign n12158 = n12157 ^ n12155 ^ 1'b0 ;
  assign n12161 = n3249 | n6641 ;
  assign n12162 = n6641 & ~n12161 ;
  assign n12159 = ~n2839 & n3083 ;
  assign n12160 = ~n6193 & n12159 ;
  assign n12163 = n12162 ^ n12160 ^ 1'b0 ;
  assign n12164 = ~n12158 & n12163 ;
  assign n12165 = n8835 ^ n8407 ^ 1'b0 ;
  assign n12166 = n1981 | n9754 ;
  assign n12167 = ( n1525 & ~n6357 ) | ( n1525 & n12166 ) | ( ~n6357 & n12166 ) ;
  assign n12168 = ( n1684 & n3399 ) | ( n1684 & n4955 ) | ( n3399 & n4955 ) ;
  assign n12170 = ~n4235 & n4936 ;
  assign n12171 = n12170 ^ n486 ^ 1'b0 ;
  assign n12172 = n12171 ^ n7720 ^ 1'b0 ;
  assign n12169 = n7763 ^ n7558 ^ n5548 ;
  assign n12173 = n12172 ^ n12169 ^ n7032 ;
  assign n12179 = n5656 ^ n4631 ^ 1'b0 ;
  assign n12174 = n884 | n4509 ;
  assign n12175 = n9515 & ~n12174 ;
  assign n12176 = n2772 & ~n12175 ;
  assign n12177 = n12176 ^ n7196 ^ 1'b0 ;
  assign n12178 = n373 & n12177 ;
  assign n12180 = n12179 ^ n12178 ^ 1'b0 ;
  assign n12181 = n1182 | n9341 ;
  assign n12182 = n2099 | n12181 ;
  assign n12183 = n11464 ^ n3811 ^ 1'b0 ;
  assign n12184 = n12182 & ~n12183 ;
  assign n12185 = n493 & n10962 ;
  assign n12186 = n12185 ^ n6658 ^ 1'b0 ;
  assign n12187 = ~n5898 & n12186 ;
  assign n12188 = ~n3005 & n11836 ;
  assign n12189 = n6149 & ~n12188 ;
  assign n12190 = n12189 ^ n5641 ^ 1'b0 ;
  assign n12191 = ~n10161 & n12190 ;
  assign n12192 = ~n242 & n12191 ;
  assign n12193 = n3830 & n6384 ;
  assign n12194 = n9572 & ~n12193 ;
  assign n12195 = n6674 ^ n510 ^ 1'b0 ;
  assign n12196 = ~n2435 & n10445 ;
  assign n12197 = n12196 ^ n8577 ^ 1'b0 ;
  assign n12198 = ( ~n2007 & n6993 ) | ( ~n2007 & n12197 ) | ( n6993 & n12197 ) ;
  assign n12199 = n5797 & ~n5962 ;
  assign n12200 = n2021 & n10005 ;
  assign n12201 = n5391 & n12200 ;
  assign n12202 = n10428 ^ n4644 ^ 1'b0 ;
  assign n12203 = n3900 & ~n5918 ;
  assign n12204 = n12202 & n12203 ;
  assign n12205 = n565 & n5859 ;
  assign n12206 = n5527 & n12205 ;
  assign n12207 = n8539 ^ n5050 ^ 1'b0 ;
  assign n12208 = n11323 ^ n2295 ^ 1'b0 ;
  assign n12209 = n5621 & n12208 ;
  assign n12210 = n12207 & ~n12209 ;
  assign n12211 = ~n2777 & n6251 ;
  assign n12212 = n12211 ^ n4457 ^ 1'b0 ;
  assign n12213 = n12212 ^ n5324 ^ 1'b0 ;
  assign n12214 = ~n3607 & n12213 ;
  assign n12215 = ~n5079 & n12214 ;
  assign n12216 = ~n12210 & n12215 ;
  assign n12217 = n2310 ^ n1347 ^ 1'b0 ;
  assign n12218 = n1634 | n12217 ;
  assign n12219 = x21 & n773 ;
  assign n12220 = n5781 | n11391 ;
  assign n12226 = n2222 & ~n6169 ;
  assign n12224 = n2622 | n3836 ;
  assign n12225 = ~n3203 & n12224 ;
  assign n12227 = n12226 ^ n12225 ^ 1'b0 ;
  assign n12221 = ~x27 & n8317 ;
  assign n12222 = n12221 ^ n6097 ^ n2802 ;
  assign n12223 = n567 & n12222 ;
  assign n12228 = n12227 ^ n12223 ^ 1'b0 ;
  assign n12229 = n12228 ^ n9786 ^ n2419 ;
  assign n12230 = n3901 & ~n10921 ;
  assign n12231 = n8547 ^ n4419 ^ 1'b0 ;
  assign n12232 = n665 | n3208 ;
  assign n12233 = n6327 & ~n12232 ;
  assign n12234 = n5706 ^ n2600 ^ 1'b0 ;
  assign n12235 = n12233 | n12234 ;
  assign n12237 = n6135 ^ n319 ^ 1'b0 ;
  assign n12238 = n7627 & n12237 ;
  assign n12236 = n5121 & ~n10868 ;
  assign n12239 = n12238 ^ n12236 ^ 1'b0 ;
  assign n12240 = n5051 & n8020 ;
  assign n12241 = ~n1254 & n12240 ;
  assign n12242 = ( n2549 & n2888 ) | ( n2549 & ~n8934 ) | ( n2888 & ~n8934 ) ;
  assign n12243 = n8730 ^ n7773 ^ 1'b0 ;
  assign n12244 = ~n7263 & n12243 ;
  assign n12245 = n2634 | n7251 ;
  assign n12246 = n12245 ^ n5030 ^ 1'b0 ;
  assign n12247 = n3793 & n3825 ;
  assign n12248 = n12246 & n12247 ;
  assign n12249 = n9591 ^ n7790 ^ n1578 ;
  assign n12250 = n1521 ^ n361 ^ 1'b0 ;
  assign n12251 = n12249 & n12250 ;
  assign n12252 = ( n635 & n1849 ) | ( n635 & ~n3805 ) | ( n1849 & ~n3805 ) ;
  assign n12253 = ( ~n369 & n11109 ) | ( ~n369 & n12252 ) | ( n11109 & n12252 ) ;
  assign n12254 = n7804 ^ n2640 ^ 1'b0 ;
  assign n12255 = n12254 ^ n1586 ^ 1'b0 ;
  assign n12256 = n12255 ^ n7866 ^ 1'b0 ;
  assign n12257 = x83 & ~n7613 ;
  assign n12258 = ~n3281 & n12257 ;
  assign n12259 = n1379 | n7103 ;
  assign n12260 = n12258 | n12259 ;
  assign n12261 = n12260 ^ n2199 ^ 1'b0 ;
  assign n12262 = n1999 & ~n12261 ;
  assign n12263 = ~n12256 & n12262 ;
  assign n12264 = n3297 | n3480 ;
  assign n12265 = ~n2793 & n4904 ;
  assign n12266 = n12265 ^ n10454 ^ 1'b0 ;
  assign n12267 = n3849 ^ n1203 ^ 1'b0 ;
  assign n12268 = n4975 | n5030 ;
  assign n12269 = n12268 ^ n4492 ^ 1'b0 ;
  assign n12270 = n2661 ^ n1168 ^ 1'b0 ;
  assign n12271 = n4472 & ~n12270 ;
  assign n12272 = n12271 ^ x3 ^ 1'b0 ;
  assign n12273 = ~n6717 & n12272 ;
  assign n12274 = n3417 | n8200 ;
  assign n12275 = n12274 ^ n7734 ^ 1'b0 ;
  assign n12278 = n4670 & ~n8860 ;
  assign n12279 = n12278 ^ n1627 ^ 1'b0 ;
  assign n12280 = n6923 & ~n12279 ;
  assign n12281 = n12280 ^ n3590 ^ 1'b0 ;
  assign n12276 = n4100 & ~n7099 ;
  assign n12277 = n12276 ^ n1682 ^ 1'b0 ;
  assign n12282 = n12281 ^ n12277 ^ 1'b0 ;
  assign n12283 = x86 & n4613 ;
  assign n12284 = n3268 & n12283 ;
  assign n12285 = n9275 & n11903 ;
  assign n12286 = n12284 & n12285 ;
  assign n12287 = n5526 ^ n5476 ^ n4044 ;
  assign n12288 = n12287 ^ n5875 ^ 1'b0 ;
  assign n12289 = n9686 | n12288 ;
  assign n12290 = n10959 ^ n2157 ^ 1'b0 ;
  assign n12291 = n10868 | n12290 ;
  assign n12295 = n4065 ^ n824 ^ 1'b0 ;
  assign n12296 = n6156 & n12295 ;
  assign n12297 = n3365 & n12296 ;
  assign n12298 = ~n6311 & n12297 ;
  assign n12299 = n4285 | n12298 ;
  assign n12292 = n2622 ^ n1372 ^ 1'b0 ;
  assign n12293 = ( ~n454 & n4097 ) | ( ~n454 & n10689 ) | ( n4097 & n10689 ) ;
  assign n12294 = ~n12292 & n12293 ;
  assign n12300 = n12299 ^ n12294 ^ 1'b0 ;
  assign n12301 = n6573 ^ n1582 ^ 1'b0 ;
  assign n12302 = n12300 & ~n12301 ;
  assign n12303 = n6974 & n12302 ;
  assign n12304 = n6039 ^ n5581 ^ 1'b0 ;
  assign n12305 = ( ~n4599 & n11531 ) | ( ~n4599 & n12304 ) | ( n11531 & n12304 ) ;
  assign n12306 = n5589 ^ n3307 ^ 1'b0 ;
  assign n12307 = n12305 & ~n12306 ;
  assign n12308 = ~n7935 & n12307 ;
  assign n12309 = n12308 ^ n4644 ^ n1829 ;
  assign n12310 = n12116 ^ n7514 ^ n836 ;
  assign n12311 = n3287 & ~n6705 ;
  assign n12312 = ~n2483 & n12311 ;
  assign n12313 = n3269 & ~n12312 ;
  assign n12314 = ~n7562 & n12313 ;
  assign n12315 = n7255 | n11794 ;
  assign n12316 = n12314 & ~n12315 ;
  assign n12317 = n8673 ^ n7906 ^ n2399 ;
  assign n12318 = n2970 & n8069 ;
  assign n12319 = ~n1979 & n3070 ;
  assign n12320 = n4948 | n8277 ;
  assign n12321 = n9817 ^ n5637 ^ 1'b0 ;
  assign n12322 = n381 & ~n12321 ;
  assign n12323 = n7924 ^ n6219 ^ 1'b0 ;
  assign n12324 = n381 | n8058 ;
  assign n12325 = n12324 ^ n6157 ^ 1'b0 ;
  assign n12326 = n12325 ^ n276 ^ 1'b0 ;
  assign n12327 = n9182 & n10200 ;
  assign n12328 = n12327 ^ n1022 ^ 1'b0 ;
  assign n12329 = ( n5834 & n10673 ) | ( n5834 & n12328 ) | ( n10673 & n12328 ) ;
  assign n12332 = ~n6350 & n12081 ;
  assign n12330 = x60 & ~n6101 ;
  assign n12331 = n12330 ^ n3105 ^ 1'b0 ;
  assign n12333 = n12332 ^ n12331 ^ 1'b0 ;
  assign n12334 = n4025 & ~n6991 ;
  assign n12335 = ~n4602 & n6155 ;
  assign n12336 = n940 & n12335 ;
  assign n12337 = n2244 & ~n6903 ;
  assign n12338 = n12337 ^ n3758 ^ 1'b0 ;
  assign n12339 = n9167 | n12338 ;
  assign n12340 = n12339 ^ n12107 ^ 1'b0 ;
  assign n12341 = n2668 & n12340 ;
  assign n12342 = n7813 | n9368 ;
  assign n12343 = n337 & ~n12342 ;
  assign n12345 = n3098 | n3964 ;
  assign n12346 = n12345 ^ n1938 ^ 1'b0 ;
  assign n12347 = ( n1191 & n7156 ) | ( n1191 & ~n12346 ) | ( n7156 & ~n12346 ) ;
  assign n12344 = ~n4355 & n5118 ;
  assign n12348 = n12347 ^ n12344 ^ 1'b0 ;
  assign n12349 = ( ~n954 & n3156 ) | ( ~n954 & n5142 ) | ( n3156 & n5142 ) ;
  assign n12350 = n12349 ^ n1930 ^ n939 ;
  assign n12351 = n1373 & n12350 ;
  assign n12352 = n3048 & ~n4238 ;
  assign n12353 = n12352 ^ n4335 ^ 1'b0 ;
  assign n12354 = n5600 & ~n12353 ;
  assign n12355 = n12354 ^ n1913 ^ 1'b0 ;
  assign n12356 = n4708 ^ n3371 ^ 1'b0 ;
  assign n12357 = n10592 | n12356 ;
  assign n12358 = n594 & ~n9735 ;
  assign n12359 = n3869 ^ n2741 ^ 1'b0 ;
  assign n12360 = n5516 & n12359 ;
  assign n12361 = ~n8994 & n12360 ;
  assign n12362 = ~n1012 & n5351 ;
  assign n12363 = n4094 | n12362 ;
  assign n12364 = n12363 ^ n8126 ^ 1'b0 ;
  assign n12365 = n373 & n11618 ;
  assign n12366 = n12365 ^ n1854 ^ 1'b0 ;
  assign n12368 = n503 & n5836 ;
  assign n12367 = n4481 | n5581 ;
  assign n12369 = n12368 ^ n12367 ^ n791 ;
  assign n12370 = ~n2611 & n3297 ;
  assign n12371 = n12370 ^ n6166 ^ 1'b0 ;
  assign n12372 = n12371 ^ n4041 ^ 1'b0 ;
  assign n12373 = n5916 & n12372 ;
  assign n12374 = ( n1171 & ~n1332 ) | ( n1171 & n2535 ) | ( ~n1332 & n2535 ) ;
  assign n12375 = n6013 & n7878 ;
  assign n12376 = n12375 ^ n1236 ^ 1'b0 ;
  assign n12377 = n594 & n1798 ;
  assign n12378 = n12377 ^ n1637 ^ 1'b0 ;
  assign n12379 = ~n1638 & n6528 ;
  assign n12380 = n12379 ^ n9574 ^ 1'b0 ;
  assign n12382 = n5318 ^ n1869 ^ n895 ;
  assign n12381 = ~n6899 & n7872 ;
  assign n12383 = n12382 ^ n12381 ^ 1'b0 ;
  assign n12384 = n12118 & n12383 ;
  assign n12385 = ~n403 & n5852 ;
  assign n12386 = ~n1479 & n2313 ;
  assign n12387 = n12386 ^ n909 ^ 1'b0 ;
  assign n12388 = ( n2647 & n4025 ) | ( n2647 & n6564 ) | ( n4025 & n6564 ) ;
  assign n12389 = n9263 | n12388 ;
  assign n12390 = n1000 & ~n12389 ;
  assign n12391 = n944 | n10977 ;
  assign n12392 = x100 & ~n3911 ;
  assign n12393 = n1848 & n12392 ;
  assign n12394 = n2897 | n12353 ;
  assign n12395 = n12394 ^ n4672 ^ 1'b0 ;
  assign n12396 = ~n12393 & n12395 ;
  assign n12397 = n12396 ^ n3627 ^ 1'b0 ;
  assign n12401 = n6511 ^ n2244 ^ 1'b0 ;
  assign n12398 = n2099 & ~n6308 ;
  assign n12399 = n4500 | n12398 ;
  assign n12400 = n3696 | n12399 ;
  assign n12402 = n12401 ^ n12400 ^ 1'b0 ;
  assign n12403 = n645 & ~n5717 ;
  assign n12404 = n12403 ^ n4097 ^ 1'b0 ;
  assign n12407 = n3995 & ~n7893 ;
  assign n12405 = n5208 ^ n2734 ^ 1'b0 ;
  assign n12406 = n4449 & n12405 ;
  assign n12408 = n12407 ^ n12406 ^ 1'b0 ;
  assign n12409 = n4802 & ~n10504 ;
  assign n12410 = ~n12408 & n12409 ;
  assign n12411 = n621 & ~n6700 ;
  assign n12412 = n12410 | n12411 ;
  assign n12413 = n3476 | n12412 ;
  assign n12414 = n7605 | n12413 ;
  assign n12415 = n8543 & ~n12414 ;
  assign n12416 = n7056 & ~n7604 ;
  assign n12417 = n2728 & n4880 ;
  assign n12418 = n11819 ^ n6052 ^ n3811 ;
  assign n12419 = n4779 ^ n4564 ^ 1'b0 ;
  assign n12420 = ( n1074 & ~n1482 ) | ( n1074 & n7027 ) | ( ~n1482 & n7027 ) ;
  assign n12421 = ~n6217 & n6399 ;
  assign n12422 = n12421 ^ n6634 ^ 1'b0 ;
  assign n12423 = n12422 ^ n6365 ^ 1'b0 ;
  assign n12424 = n1036 & ~n10372 ;
  assign n12425 = n11739 & n12424 ;
  assign n12426 = n4291 & n6516 ;
  assign n12427 = n1847 & n3558 ;
  assign n12428 = n1318 & n12427 ;
  assign n12429 = n11263 | n12428 ;
  assign n12430 = n12429 ^ n452 ^ 1'b0 ;
  assign n12431 = n4510 ^ n3516 ^ 1'b0 ;
  assign n12432 = ~n4246 & n12431 ;
  assign n12433 = n7296 | n10497 ;
  assign n12434 = n5227 & ~n6853 ;
  assign n12435 = n12434 ^ x9 ^ 1'b0 ;
  assign n12436 = n12435 ^ n8694 ^ n7172 ;
  assign n12437 = ~n2291 & n9710 ;
  assign n12438 = ( ~n11331 & n12436 ) | ( ~n11331 & n12437 ) | ( n12436 & n12437 ) ;
  assign n12439 = ( ~n832 & n1842 ) | ( ~n832 & n8357 ) | ( n1842 & n8357 ) ;
  assign n12440 = ( n5854 & n9880 ) | ( n5854 & n12439 ) | ( n9880 & n12439 ) ;
  assign n12441 = n12440 ^ n1894 ^ n1868 ;
  assign n12442 = ~n498 & n1206 ;
  assign n12443 = ~n2827 & n12442 ;
  assign n12444 = n5573 ^ n2675 ^ 1'b0 ;
  assign n12445 = n12443 | n12444 ;
  assign n12446 = n2258 & ~n12445 ;
  assign n12447 = n12446 ^ n2622 ^ 1'b0 ;
  assign n12448 = n5706 ^ n2577 ^ 1'b0 ;
  assign n12449 = n5736 & n12448 ;
  assign n12450 = n12449 ^ n2558 ^ 1'b0 ;
  assign n12451 = n2595 ^ n1017 ^ 1'b0 ;
  assign n12452 = n12451 ^ n8902 ^ 1'b0 ;
  assign n12453 = ~n12450 & n12452 ;
  assign n12455 = ( n4165 & ~n5925 ) | ( n4165 & n11418 ) | ( ~n5925 & n11418 ) ;
  assign n12454 = n1779 & n7619 ;
  assign n12456 = n12455 ^ n12454 ^ 1'b0 ;
  assign n12457 = n6457 ^ n4000 ^ 1'b0 ;
  assign n12458 = n12457 ^ n202 ^ 1'b0 ;
  assign n12459 = n12458 ^ n193 ^ 1'b0 ;
  assign n12460 = ~n933 & n1876 ;
  assign n12461 = ~n10134 & n12460 ;
  assign n12462 = n9932 & ~n12461 ;
  assign n12463 = n12462 ^ n10428 ^ 1'b0 ;
  assign n12464 = n1888 & n3243 ;
  assign n12465 = n10282 | n12464 ;
  assign n12466 = n12088 ^ n1775 ^ n1504 ;
  assign n12467 = n2622 & ~n10951 ;
  assign n12468 = n3093 & ~n5291 ;
  assign n12469 = n12468 ^ n3334 ^ 1'b0 ;
  assign n12470 = ( n6146 & n12467 ) | ( n6146 & n12469 ) | ( n12467 & n12469 ) ;
  assign n12471 = n7983 & n12470 ;
  assign n12472 = n635 & n1299 ;
  assign n12473 = n7744 ^ n7556 ^ 1'b0 ;
  assign n12474 = n12472 & ~n12473 ;
  assign n12475 = ~n671 & n1724 ;
  assign n12477 = n9486 & ~n10233 ;
  assign n12478 = n12477 ^ n2705 ^ 1'b0 ;
  assign n12479 = n8699 | n12478 ;
  assign n12476 = x88 & ~n8204 ;
  assign n12480 = n12479 ^ n12476 ^ 1'b0 ;
  assign n12481 = n7814 & ~n7945 ;
  assign n12482 = n12481 ^ n2938 ^ 1'b0 ;
  assign n12483 = n2945 & n4865 ;
  assign n12484 = n12483 ^ n4911 ^ 1'b0 ;
  assign n12485 = n12482 & n12484 ;
  assign n12486 = n910 & ~n12485 ;
  assign n12490 = n1257 ^ n872 ^ 1'b0 ;
  assign n12487 = n3803 ^ n1044 ^ x27 ;
  assign n12488 = ~n2802 & n12487 ;
  assign n12489 = ~n10095 & n12488 ;
  assign n12491 = n12490 ^ n12489 ^ 1'b0 ;
  assign n12492 = ~n752 & n12491 ;
  assign n12493 = ( x97 & n3664 ) | ( x97 & n11763 ) | ( n3664 & n11763 ) ;
  assign n12494 = ( n1521 & n2493 ) | ( n1521 & ~n3031 ) | ( n2493 & ~n3031 ) ;
  assign n12495 = n11198 | n12494 ;
  assign n12496 = n5895 ^ n4819 ^ 1'b0 ;
  assign n12497 = n673 & n12496 ;
  assign n12498 = ( x126 & n7400 ) | ( x126 & n7789 ) | ( n7400 & n7789 ) ;
  assign n12499 = n6874 & ~n11557 ;
  assign n12500 = ~n2419 & n9039 ;
  assign n12501 = n1506 & ~n7654 ;
  assign n12502 = ( n2051 & ~n12500 ) | ( n2051 & n12501 ) | ( ~n12500 & n12501 ) ;
  assign n12503 = n3006 & ~n12502 ;
  assign n12504 = n973 | n12401 ;
  assign n12505 = n4025 ^ n725 ^ 1'b0 ;
  assign n12506 = n10397 | n12505 ;
  assign n12507 = n3199 | n12015 ;
  assign n12508 = n3297 | n12507 ;
  assign n12509 = n5734 ^ n2433 ^ 1'b0 ;
  assign n12510 = ~n3411 & n6095 ;
  assign n12511 = ( x111 & ~n1586 ) | ( x111 & n3766 ) | ( ~n1586 & n3766 ) ;
  assign n12512 = n471 & ~n12511 ;
  assign n12513 = n8382 & ~n12512 ;
  assign n12514 = n12513 ^ n3788 ^ 1'b0 ;
  assign n12515 = n5964 & ~n12348 ;
  assign n12516 = n9936 ^ n2151 ^ 1'b0 ;
  assign n12519 = n3827 ^ n2328 ^ 1'b0 ;
  assign n12520 = n4160 & n12519 ;
  assign n12517 = n9223 ^ n2146 ^ 1'b0 ;
  assign n12518 = n871 | n12517 ;
  assign n12521 = n12520 ^ n12518 ^ n499 ;
  assign n12522 = n11128 ^ n7988 ^ n7893 ;
  assign n12523 = n4547 & ~n5093 ;
  assign n12524 = n4271 | n11550 ;
  assign n12525 = n3156 & ~n7367 ;
  assign n12526 = n12525 ^ n6896 ^ 1'b0 ;
  assign n12527 = n6002 & n12526 ;
  assign n12528 = n12527 ^ n691 ^ 1'b0 ;
  assign n12529 = n2956 | n4136 ;
  assign n12530 = n521 | n3132 ;
  assign n12531 = n12530 ^ n4948 ^ 1'b0 ;
  assign n12532 = n12531 ^ n6541 ^ 1'b0 ;
  assign n12533 = n12529 & ~n12532 ;
  assign n12534 = n12533 ^ n10061 ^ n9331 ;
  assign n12536 = x39 & ~n1766 ;
  assign n12535 = x93 & ~n1286 ;
  assign n12537 = n12536 ^ n12535 ^ n9674 ;
  assign n12538 = n778 & n2462 ;
  assign n12539 = n12538 ^ n3386 ^ 1'b0 ;
  assign n12540 = n8623 & n12539 ;
  assign n12541 = n8002 ^ n7452 ^ 1'b0 ;
  assign n12542 = n9599 ^ n6215 ^ 1'b0 ;
  assign n12543 = n10860 & n12542 ;
  assign n12544 = n12543 ^ n9657 ^ 1'b0 ;
  assign n12545 = n1106 | n8676 ;
  assign n12546 = n4606 & ~n12545 ;
  assign n12547 = n1879 | n12546 ;
  assign n12548 = n1911 | n12547 ;
  assign n12549 = ( n3947 & ~n8849 ) | ( n3947 & n12548 ) | ( ~n8849 & n12548 ) ;
  assign n12550 = n12549 ^ n4124 ^ 1'b0 ;
  assign n12551 = n1966 & n2205 ;
  assign n12552 = n7099 & n12551 ;
  assign n12553 = n2172 & ~n5098 ;
  assign n12554 = ~n322 & n12553 ;
  assign n12555 = ( n1452 & n7504 ) | ( n1452 & n8938 ) | ( n7504 & n8938 ) ;
  assign n12556 = ~n341 & n12555 ;
  assign n12557 = n1075 & ~n7984 ;
  assign n12558 = n4745 & n12557 ;
  assign n12559 = n2804 & n9320 ;
  assign n12560 = ( n3250 & n12558 ) | ( n3250 & ~n12559 ) | ( n12558 & ~n12559 ) ;
  assign n12561 = n8345 & ~n12560 ;
  assign n12562 = n7850 ^ n4270 ^ n1983 ;
  assign n12563 = ( n5052 & ~n8425 ) | ( n5052 & n12562 ) | ( ~n8425 & n12562 ) ;
  assign n12564 = n12563 ^ n8108 ^ 1'b0 ;
  assign n12565 = n674 & ~n12564 ;
  assign n12566 = n12565 ^ n3859 ^ 1'b0 ;
  assign n12567 = ~n1811 & n4985 ;
  assign n12568 = n12567 ^ n202 ^ 1'b0 ;
  assign n12569 = ~n2656 & n8385 ;
  assign n12570 = n7656 & n12569 ;
  assign n12571 = n1802 & ~n3011 ;
  assign n12572 = n12571 ^ n9008 ^ n1587 ;
  assign n12573 = n3947 & ~n9514 ;
  assign n12574 = n452 & n1741 ;
  assign n12575 = n2693 & n12574 ;
  assign n12576 = x47 & n7565 ;
  assign n12577 = n9979 & n12576 ;
  assign n12578 = n5107 | n12577 ;
  assign n12579 = n1840 & ~n12578 ;
  assign n12580 = n3947 | n12579 ;
  assign n12581 = n4761 & n5458 ;
  assign n12582 = ~n8813 & n12581 ;
  assign n12583 = ~n1332 & n2312 ;
  assign n12584 = n12583 ^ n3883 ^ 1'b0 ;
  assign n12585 = n12584 ^ n2159 ^ 1'b0 ;
  assign n12586 = n10937 ^ n4351 ^ 1'b0 ;
  assign n12587 = ~n1108 & n2917 ;
  assign n12588 = n2923 ^ n2596 ^ 1'b0 ;
  assign n12589 = n4400 & n12588 ;
  assign n12590 = ~n299 & n5669 ;
  assign n12591 = n12590 ^ n8526 ^ 1'b0 ;
  assign n12592 = n1840 & ~n5633 ;
  assign n12593 = n2608 & n12592 ;
  assign n12594 = n6446 | n10035 ;
  assign n12595 = n730 & n11061 ;
  assign n12596 = ~n7632 & n7759 ;
  assign n12597 = n12317 ^ n8776 ^ 1'b0 ;
  assign n12598 = n1846 & ~n12597 ;
  assign n12599 = ~n8567 & n9343 ;
  assign n12600 = n12599 ^ n5495 ^ 1'b0 ;
  assign n12601 = n1139 | n4186 ;
  assign n12602 = n2691 & ~n10061 ;
  assign n12603 = n12602 ^ n12505 ^ 1'b0 ;
  assign n12606 = n2703 & n7012 ;
  assign n12607 = ~n7012 & n12606 ;
  assign n12604 = n3172 & n6424 ;
  assign n12605 = n12604 ^ n6617 ^ 1'b0 ;
  assign n12608 = n12607 ^ n12605 ^ n1974 ;
  assign n12609 = n928 | n1821 ;
  assign n12610 = n12609 ^ n7930 ^ 1'b0 ;
  assign n12611 = n12610 ^ n5815 ^ 1'b0 ;
  assign n12612 = n9743 ^ n972 ^ 1'b0 ;
  assign n12613 = x70 | n3814 ;
  assign n12614 = n12613 ^ n5925 ^ 1'b0 ;
  assign n12615 = n12614 ^ n676 ^ 1'b0 ;
  assign n12616 = n12612 | n12615 ;
  assign n12617 = ( n815 & n9989 ) | ( n815 & ~n10878 ) | ( n9989 & ~n10878 ) ;
  assign n12618 = n12617 ^ n12023 ^ 1'b0 ;
  assign n12619 = ~n2839 & n8966 ;
  assign n12620 = n4712 | n9472 ;
  assign n12621 = ( n2554 & n3845 ) | ( n2554 & n3960 ) | ( n3845 & n3960 ) ;
  assign n12622 = n10491 & ~n12621 ;
  assign n12623 = n12622 ^ n6735 ^ 1'b0 ;
  assign n12624 = n3638 ^ n1079 ^ 1'b0 ;
  assign n12625 = n3204 | n12624 ;
  assign n12626 = ( n3744 & ~n5681 ) | ( n3744 & n8233 ) | ( ~n5681 & n8233 ) ;
  assign n12627 = n12626 ^ n7165 ^ 1'b0 ;
  assign n12628 = ~n12625 & n12627 ;
  assign n12629 = n9904 ^ n6519 ^ n764 ;
  assign n12630 = n1794 & n5800 ;
  assign n12631 = ~n5093 & n8279 ;
  assign n12632 = n12631 ^ n282 ^ 1'b0 ;
  assign n12633 = ~n10985 & n12632 ;
  assign n12634 = n828 | n4359 ;
  assign n12635 = n12634 ^ n11130 ^ n6141 ;
  assign n12636 = n148 | n8360 ;
  assign n12637 = ~n4319 & n12133 ;
  assign n12638 = n12637 ^ n7685 ^ 1'b0 ;
  assign n12639 = n129 & ~n8692 ;
  assign n12640 = n2582 ^ n1387 ^ 1'b0 ;
  assign n12641 = ~n2846 & n9210 ;
  assign n12642 = n9667 ^ n8732 ^ n6135 ;
  assign n12643 = ~n1408 & n1998 ;
  assign n12644 = ~n6908 & n12643 ;
  assign n12645 = ~n7750 & n8766 ;
  assign n12646 = n4052 ^ n2207 ^ 1'b0 ;
  assign n12647 = ~n5618 & n12646 ;
  assign n12648 = n3516 & n12647 ;
  assign n12649 = n2870 & ~n3995 ;
  assign n12650 = ~n2069 & n12649 ;
  assign n12651 = n5091 ^ n818 ^ 1'b0 ;
  assign n12653 = n462 ^ x1 ^ 1'b0 ;
  assign n12652 = x104 & ~n8197 ;
  assign n12654 = n12653 ^ n12652 ^ 1'b0 ;
  assign n12655 = ~n12651 & n12654 ;
  assign n12656 = ~n12650 & n12655 ;
  assign n12657 = n12656 ^ n2957 ^ 1'b0 ;
  assign n12658 = n5950 ^ n2866 ^ 1'b0 ;
  assign n12659 = n4740 ^ n2850 ^ 1'b0 ;
  assign n12660 = n12659 ^ n2694 ^ 1'b0 ;
  assign n12661 = ( n1599 & n3080 ) | ( n1599 & n12660 ) | ( n3080 & n12660 ) ;
  assign n12662 = n2622 & n12661 ;
  assign n12663 = n12662 ^ n3396 ^ 1'b0 ;
  assign n12664 = n7368 ^ n3456 ^ n2065 ;
  assign n12665 = n4279 | n6159 ;
  assign n12666 = n12665 ^ n9007 ^ 1'b0 ;
  assign n12667 = n654 | n12666 ;
  assign n12668 = n12667 ^ n804 ^ 1'b0 ;
  assign n12669 = n12664 & ~n12668 ;
  assign n12670 = n3339 ^ n2306 ^ 1'b0 ;
  assign n12671 = x86 & n12670 ;
  assign n12672 = n12669 & ~n12671 ;
  assign n12673 = n330 & ~n9029 ;
  assign n12674 = n5383 ^ n331 ^ 1'b0 ;
  assign n12675 = n2525 & ~n3869 ;
  assign n12676 = n12675 ^ n6408 ^ 1'b0 ;
  assign n12677 = n12676 ^ n1172 ^ 1'b0 ;
  assign n12678 = n11474 ^ n7909 ^ 1'b0 ;
  assign n12679 = n7101 & ~n12660 ;
  assign n12681 = n134 & ~n933 ;
  assign n12682 = n3147 & n12681 ;
  assign n12683 = n12682 ^ n4428 ^ n1869 ;
  assign n12684 = n4950 | n12683 ;
  assign n12680 = n2930 & ~n7311 ;
  assign n12685 = n12684 ^ n12680 ^ 1'b0 ;
  assign n12686 = ~n2806 & n6501 ;
  assign n12687 = n9268 & ~n12686 ;
  assign n12689 = ~n5910 & n12127 ;
  assign n12690 = n8042 & n12689 ;
  assign n12688 = n2888 ^ x95 ^ 1'b0 ;
  assign n12691 = n12690 ^ n12688 ^ 1'b0 ;
  assign n12692 = n2906 ^ n2173 ^ n2098 ;
  assign n12693 = n1427 ^ n1312 ^ 1'b0 ;
  assign n12694 = n4124 | n12693 ;
  assign n12695 = n11927 & n12694 ;
  assign n12696 = n10426 ^ n8231 ^ 1'b0 ;
  assign n12697 = n12696 ^ x91 ^ 1'b0 ;
  assign n12698 = n1938 & ~n2591 ;
  assign n12699 = n9638 & n12698 ;
  assign n12700 = ~n1410 & n12699 ;
  assign n12701 = n9052 | n12700 ;
  assign n12702 = n12701 ^ n8678 ^ 1'b0 ;
  assign n12703 = n12410 ^ n2605 ^ 1'b0 ;
  assign n12704 = n7857 | n9760 ;
  assign n12705 = n2570 & n9494 ;
  assign n12706 = n12705 ^ n7887 ^ 1'b0 ;
  assign n12707 = n8603 ^ n5366 ^ 1'b0 ;
  assign n12708 = n12707 ^ n6225 ^ 1'b0 ;
  assign n12709 = ~n2715 & n12708 ;
  assign n12710 = n678 | n1868 ;
  assign n12711 = n6629 | n12710 ;
  assign n12712 = n12682 & n12711 ;
  assign n12713 = n8113 ^ n5948 ^ 1'b0 ;
  assign n12714 = n3453 & n6874 ;
  assign n12715 = n10434 ^ n4091 ^ 1'b0 ;
  assign n12716 = ~n5517 & n12715 ;
  assign n12717 = n12716 ^ n5536 ^ n229 ;
  assign n12718 = n12717 ^ n8376 ^ 1'b0 ;
  assign n12719 = ~n2622 & n12205 ;
  assign n12720 = x22 & n2577 ;
  assign n12721 = n12720 ^ n6903 ^ 1'b0 ;
  assign n12722 = n11404 & n12721 ;
  assign n12723 = n2043 & n5183 ;
  assign n12724 = n1329 | n8966 ;
  assign n12725 = n12724 ^ n4959 ^ 1'b0 ;
  assign n12726 = n11921 ^ n2649 ^ n1860 ;
  assign n12727 = n6779 ^ n3623 ^ n1700 ;
  assign n12728 = n12727 ^ n5603 ^ 1'b0 ;
  assign n12729 = n12150 ^ n4230 ^ 1'b0 ;
  assign n12730 = n4964 | n12729 ;
  assign n12731 = n12728 & ~n12730 ;
  assign n12732 = n1511 ^ n1109 ^ 1'b0 ;
  assign n12733 = ~n2860 & n6998 ;
  assign n12734 = ~n2305 & n12733 ;
  assign n12735 = n6711 & ~n12734 ;
  assign n12736 = n12734 & n12735 ;
  assign n12737 = ~n2956 & n10198 ;
  assign n12738 = n12737 ^ n7109 ^ 1'b0 ;
  assign n12739 = ~n690 & n1100 ;
  assign n12740 = n12739 ^ n10260 ^ 1'b0 ;
  assign n12741 = n12738 & ~n12740 ;
  assign n12743 = n4611 ^ n1573 ^ 1'b0 ;
  assign n12744 = n6157 | n12743 ;
  assign n12745 = n2300 & ~n12744 ;
  assign n12746 = n12745 ^ n701 ^ 1'b0 ;
  assign n12747 = n12746 ^ n12434 ^ 1'b0 ;
  assign n12742 = n2507 | n12695 ;
  assign n12748 = n12747 ^ n12742 ^ 1'b0 ;
  assign n12749 = ~n2523 & n3910 ;
  assign n12750 = n4863 | n12749 ;
  assign n12751 = n8122 ^ n4440 ^ 1'b0 ;
  assign n12752 = n3404 | n12751 ;
  assign n12753 = n12750 | n12752 ;
  assign n12754 = n6786 & ~n11012 ;
  assign n12755 = ~n372 & n9532 ;
  assign n12756 = n12755 ^ n2209 ^ 1'b0 ;
  assign n12757 = n12754 & ~n12756 ;
  assign n12758 = ( n2611 & n9221 ) | ( n2611 & ~n11008 ) | ( n9221 & ~n11008 ) ;
  assign n12759 = n12758 ^ n5915 ^ 1'b0 ;
  assign n12760 = n3958 & ~n12759 ;
  assign n12761 = ~n6001 & n12760 ;
  assign n12762 = n829 & n1749 ;
  assign n12763 = n12761 & n12762 ;
  assign n12764 = n2703 & ~n3208 ;
  assign n12765 = n4923 & n12764 ;
  assign n12766 = n4717 | n12765 ;
  assign n12767 = ~n7301 & n7990 ;
  assign n12768 = n11684 & ~n12767 ;
  assign n12769 = n8582 & n12768 ;
  assign n12770 = n12221 ^ x88 ^ 1'b0 ;
  assign n12771 = n2074 & ~n12770 ;
  assign n12772 = n12771 ^ n1777 ^ n1580 ;
  assign n12773 = n12772 ^ n8531 ^ 1'b0 ;
  assign n12774 = n2679 ^ n2119 ^ 1'b0 ;
  assign n12775 = ~n2702 & n12774 ;
  assign n12776 = n12775 ^ n8534 ^ 1'b0 ;
  assign n12777 = ( ~n2465 & n10081 ) | ( ~n2465 & n12776 ) | ( n10081 & n12776 ) ;
  assign n12779 = ( ~n463 & n1809 ) | ( ~n463 & n1933 ) | ( n1809 & n1933 ) ;
  assign n12780 = n1572 ^ n510 ^ 1'b0 ;
  assign n12781 = ~n12779 & n12780 ;
  assign n12778 = x77 & n7131 ;
  assign n12782 = n12781 ^ n12778 ^ 1'b0 ;
  assign n12783 = x85 & ~n998 ;
  assign n12784 = n4053 & n12783 ;
  assign n12785 = n5307 & ~n12784 ;
  assign n12786 = n5967 & ~n12785 ;
  assign n12787 = n12786 ^ n5242 ^ 1'b0 ;
  assign n12788 = n4224 ^ n2180 ^ 1'b0 ;
  assign n12789 = n12788 ^ n2787 ^ n1526 ;
  assign n12790 = n12789 ^ n8991 ^ 1'b0 ;
  assign n12791 = ~n1081 & n5824 ;
  assign n12792 = ~n806 & n1436 ;
  assign n12793 = ~n1436 & n12792 ;
  assign n12794 = ~n1893 & n12793 ;
  assign n12795 = ~n1350 & n12794 ;
  assign n12796 = n12795 ^ n3861 ^ 1'b0 ;
  assign n12797 = ~n6763 & n12796 ;
  assign n12798 = n5447 & ~n12797 ;
  assign n12799 = ~n12791 & n12798 ;
  assign n12800 = n9645 | n11559 ;
  assign n12801 = ~n10895 & n12800 ;
  assign n12802 = ~n6049 & n12395 ;
  assign n12803 = ~n2962 & n6202 ;
  assign n12804 = n12073 ^ n4545 ^ 1'b0 ;
  assign n12805 = n2052 & n12804 ;
  assign n12806 = n5908 ^ n2408 ^ 1'b0 ;
  assign n12807 = n3108 & ~n12806 ;
  assign n12808 = x123 & n1633 ;
  assign n12809 = n12808 ^ n2034 ^ 1'b0 ;
  assign n12810 = n12809 ^ n4525 ^ n1893 ;
  assign n12811 = n3966 & ~n6196 ;
  assign n12812 = n12811 ^ n159 ^ 1'b0 ;
  assign n12813 = n12812 ^ n8605 ^ 1'b0 ;
  assign n12814 = ( x47 & n4382 ) | ( x47 & n4662 ) | ( n4382 & n4662 ) ;
  assign n12815 = ~n5296 & n12814 ;
  assign n12816 = ~n5175 & n12815 ;
  assign n12817 = n12813 | n12816 ;
  assign n12818 = n7666 & n11096 ;
  assign n12819 = ~n2619 & n12818 ;
  assign n12820 = n8389 & ~n12819 ;
  assign n12821 = n12817 & n12820 ;
  assign n12822 = n1581 & ~n8288 ;
  assign n12823 = n8832 | n12822 ;
  assign n12824 = n3223 & ~n7403 ;
  assign n12825 = n12824 ^ n1835 ^ 1'b0 ;
  assign n12826 = n4915 | n10403 ;
  assign n12827 = ( n770 & n2340 ) | ( n770 & ~n2472 ) | ( n2340 & ~n2472 ) ;
  assign n12828 = n12827 ^ n5463 ^ 1'b0 ;
  assign n12829 = n2193 & ~n12828 ;
  assign n12830 = n7286 ^ n892 ^ 1'b0 ;
  assign n12831 = n12830 ^ n826 ^ 1'b0 ;
  assign n12832 = n12831 ^ n579 ^ 1'b0 ;
  assign n12833 = n4983 | n12832 ;
  assign n12834 = n3631 & ~n7288 ;
  assign n12835 = ~n2087 & n12834 ;
  assign n12836 = n4917 & ~n12835 ;
  assign n12837 = n10356 & n11440 ;
  assign n12838 = n1610 & n12837 ;
  assign n12842 = ~x91 & n2198 ;
  assign n12843 = n12842 ^ x51 ^ 1'b0 ;
  assign n12839 = n4422 ^ n3983 ^ 1'b0 ;
  assign n12840 = n11130 & n12839 ;
  assign n12841 = n3946 & ~n12840 ;
  assign n12844 = n12843 ^ n12841 ^ 1'b0 ;
  assign n12845 = ~n4702 & n12844 ;
  assign n12850 = n1000 | n4229 ;
  assign n12851 = n12850 ^ n3212 ^ 1'b0 ;
  assign n12852 = ~n6820 & n12851 ;
  assign n12853 = n12852 ^ n5141 ^ 1'b0 ;
  assign n12846 = x112 & n3012 ;
  assign n12847 = n335 & ~n3172 ;
  assign n12848 = n12847 ^ n1138 ^ n258 ;
  assign n12849 = n12846 | n12848 ;
  assign n12854 = n12853 ^ n12849 ^ 1'b0 ;
  assign n12855 = ~n707 & n11454 ;
  assign n12856 = ~n720 & n12855 ;
  assign n12857 = n2957 ^ n1390 ^ 1'b0 ;
  assign n12858 = n6259 | n12857 ;
  assign n12859 = n5269 | n12858 ;
  assign n12860 = n1036 & n12859 ;
  assign n12861 = n389 & ~n6135 ;
  assign n12862 = ~n12860 & n12861 ;
  assign n12863 = n3353 & n10194 ;
  assign n12864 = ( n4605 & n5141 ) | ( n4605 & ~n12863 ) | ( n5141 & ~n12863 ) ;
  assign n12865 = n12864 ^ n7303 ^ 1'b0 ;
  assign n12866 = n1503 & n9350 ;
  assign n12867 = n11355 ^ n1703 ^ 1'b0 ;
  assign n12868 = n8667 & ~n12867 ;
  assign n12869 = n1481 & n3203 ;
  assign n12870 = n3580 & n12869 ;
  assign n12871 = n12870 ^ n2103 ^ 1'b0 ;
  assign n12872 = ~n182 & n12871 ;
  assign n12873 = ( n2067 & ~n4042 ) | ( n2067 & n12872 ) | ( ~n4042 & n12872 ) ;
  assign n12874 = n12873 ^ n6251 ^ 1'b0 ;
  assign n12875 = n8130 & ~n12874 ;
  assign n12876 = ~n1405 & n4335 ;
  assign n12877 = ~n4651 & n12876 ;
  assign n12878 = ( n309 & ~n673 ) | ( n309 & n12877 ) | ( ~n673 & n12877 ) ;
  assign n12879 = n1765 | n3428 ;
  assign n12880 = n9292 | n12879 ;
  assign n12881 = ~n7792 & n12880 ;
  assign n12882 = n5920 ^ n3288 ^ 1'b0 ;
  assign n12883 = ~n3901 & n12882 ;
  assign n12884 = n794 & n12883 ;
  assign n12885 = n12881 | n12884 ;
  assign n12886 = x75 & n12885 ;
  assign n12887 = n12878 & n12886 ;
  assign n12888 = n4225 & n11277 ;
  assign n12889 = ~n10583 & n12888 ;
  assign n12890 = n5520 & n7888 ;
  assign n12891 = n12037 & n12890 ;
  assign n12893 = n4382 ^ n2647 ^ 1'b0 ;
  assign n12892 = n8038 & n10228 ;
  assign n12894 = n12893 ^ n12892 ^ 1'b0 ;
  assign n12895 = n5361 ^ n4292 ^ 1'b0 ;
  assign n12896 = n1677 & ~n12895 ;
  assign n12897 = n12896 ^ n1599 ^ 1'b0 ;
  assign n12898 = n324 | n12897 ;
  assign n12904 = n6833 ^ x104 ^ 1'b0 ;
  assign n12905 = n4946 | n12904 ;
  assign n12903 = n7936 ^ n6609 ^ 1'b0 ;
  assign n12899 = n7403 ^ n3836 ^ 1'b0 ;
  assign n12900 = n3457 & n12899 ;
  assign n12901 = ~n7576 & n12900 ;
  assign n12902 = n5760 & n12901 ;
  assign n12906 = n12905 ^ n12903 ^ n12902 ;
  assign n12907 = n7491 & n12906 ;
  assign n12908 = n12907 ^ n4439 ^ n250 ;
  assign n12909 = n1522 & ~n3533 ;
  assign n12910 = ~n3149 & n12909 ;
  assign n12911 = n3123 & ~n12910 ;
  assign n12912 = n1680 | n9227 ;
  assign n12913 = n10922 & ~n12912 ;
  assign n12914 = n2847 ^ n1041 ^ 1'b0 ;
  assign n12915 = n7487 & ~n12914 ;
  assign n12916 = n12915 ^ n8344 ^ 1'b0 ;
  assign n12917 = n12916 ^ n5402 ^ 1'b0 ;
  assign n12918 = n8849 ^ n4988 ^ 1'b0 ;
  assign n12919 = n5278 ^ n1085 ^ 1'b0 ;
  assign n12920 = n6391 & n12919 ;
  assign n12921 = n12920 ^ n7840 ^ n5389 ;
  assign n12922 = n11179 ^ n3304 ^ 1'b0 ;
  assign n12924 = ~n2607 & n3268 ;
  assign n12923 = n12775 ^ n9691 ^ n9591 ;
  assign n12925 = n12924 ^ n12923 ^ 1'b0 ;
  assign n12926 = ~n11607 & n12925 ;
  assign n12927 = ~n7530 & n12926 ;
  assign n12928 = n4059 | n7936 ;
  assign n12929 = n1660 & ~n12928 ;
  assign n12930 = n12929 ^ n4325 ^ 1'b0 ;
  assign n12931 = ~n9593 & n12930 ;
  assign n12933 = n404 | n1511 ;
  assign n12934 = n12933 ^ n9446 ^ 1'b0 ;
  assign n12932 = n4942 & n5875 ;
  assign n12935 = n12934 ^ n12932 ^ n7478 ;
  assign n12936 = n1122 & n2738 ;
  assign n12937 = n1835 | n10924 ;
  assign n12938 = ~n567 & n1738 ;
  assign n12939 = n3755 & ~n12938 ;
  assign n12940 = n12939 ^ n7571 ^ 1'b0 ;
  assign n12941 = n3562 | n7859 ;
  assign n12942 = n12941 ^ n2852 ^ 1'b0 ;
  assign n12943 = n12942 ^ n7272 ^ n996 ;
  assign n12952 = x63 & n210 ;
  assign n12953 = ~n210 & n12952 ;
  assign n12954 = n612 & n12953 ;
  assign n12955 = n513 & n566 ;
  assign n12956 = ~n513 & n12955 ;
  assign n12957 = n1461 | n12956 ;
  assign n12958 = n12956 & ~n12957 ;
  assign n12959 = n5535 | n12958 ;
  assign n12960 = n12954 & ~n12959 ;
  assign n12944 = n285 & ~n1994 ;
  assign n12945 = ~n285 & n12944 ;
  assign n12946 = x12 & n12945 ;
  assign n12947 = n1399 | n8536 ;
  assign n12948 = n12946 & ~n12947 ;
  assign n12949 = x123 & ~n12948 ;
  assign n12950 = n12948 & n12949 ;
  assign n12951 = n10293 | n12950 ;
  assign n12961 = n12960 ^ n12951 ^ n6534 ;
  assign n12962 = n12500 ^ n5204 ^ 1'b0 ;
  assign n12963 = n5045 ^ n4315 ^ 1'b0 ;
  assign n12964 = n6688 & ~n12963 ;
  assign n12965 = ~n250 & n12964 ;
  assign n12966 = ~n10190 & n10783 ;
  assign n12967 = n1706 | n6040 ;
  assign n12968 = n3803 & ~n12967 ;
  assign n12969 = n12968 ^ n10768 ^ 1'b0 ;
  assign n12970 = ~n5816 & n12750 ;
  assign n12971 = n6257 ^ n3631 ^ x77 ;
  assign n12972 = n5743 | n12971 ;
  assign n12973 = n7204 ^ n6684 ^ 1'b0 ;
  assign n12974 = n12972 | n12973 ;
  assign n12975 = ~x20 & n2819 ;
  assign n12976 = n11240 ^ n5434 ^ 1'b0 ;
  assign n12977 = n4181 ^ n3437 ^ 1'b0 ;
  assign n12978 = n12977 ^ n1567 ^ 1'b0 ;
  assign n12979 = n8681 ^ n7604 ^ 1'b0 ;
  assign n12980 = ~n3265 & n12979 ;
  assign n12981 = n12980 ^ n3223 ^ 1'b0 ;
  assign n12982 = n640 | n4819 ;
  assign n12983 = n12982 ^ n442 ^ 1'b0 ;
  assign n12984 = n12983 ^ n5517 ^ 1'b0 ;
  assign n12985 = n386 & ~n12984 ;
  assign n12986 = n12985 ^ n6691 ^ 1'b0 ;
  assign n12987 = ~n6284 & n12986 ;
  assign n12988 = n5840 ^ n5785 ^ 1'b0 ;
  assign n12989 = ~n320 & n12988 ;
  assign n12990 = ~n1872 & n12989 ;
  assign n12991 = n10637 & n12990 ;
  assign n12992 = n3070 ^ n1360 ^ 1'b0 ;
  assign n12993 = n3767 | n12992 ;
  assign n12994 = ( n5545 & ~n5695 ) | ( n5545 & n7177 ) | ( ~n5695 & n7177 ) ;
  assign n12995 = n12994 ^ n3755 ^ 1'b0 ;
  assign n12996 = n7032 & ~n12399 ;
  assign n12997 = ~n4812 & n12679 ;
  assign n12998 = n2824 & n5941 ;
  assign n12999 = n827 & n12998 ;
  assign n13000 = n12999 ^ n865 ^ 1'b0 ;
  assign n13001 = n2451 | n6426 ;
  assign n13002 = n375 | n13001 ;
  assign n13003 = n13002 ^ n1033 ^ 1'b0 ;
  assign n13004 = ( ~n2980 & n9162 ) | ( ~n2980 & n13003 ) | ( n9162 & n13003 ) ;
  assign n13005 = n10152 ^ n8900 ^ 1'b0 ;
  assign n13006 = n2510 ^ n2282 ^ 1'b0 ;
  assign n13007 = n7567 & n13006 ;
  assign n13008 = n13007 ^ n3499 ^ 1'b0 ;
  assign n13009 = n7111 & n13008 ;
  assign n13010 = ~n8256 & n13009 ;
  assign n13011 = ~n5714 & n13010 ;
  assign n13012 = ( n3619 & ~n6536 ) | ( n3619 & n9950 ) | ( ~n6536 & n9950 ) ;
  assign n13013 = n9321 ^ n1739 ^ 1'b0 ;
  assign n13014 = n13012 | n13013 ;
  assign n13015 = x126 & n2366 ;
  assign n13016 = n353 & n13015 ;
  assign n13017 = n9658 ^ n8128 ^ 1'b0 ;
  assign n13021 = n681 | n1512 ;
  assign n13018 = n2479 ^ x121 ^ 1'b0 ;
  assign n13019 = n482 & ~n13018 ;
  assign n13020 = ( n668 & n4832 ) | ( n668 & ~n13019 ) | ( n4832 & ~n13019 ) ;
  assign n13022 = n13021 ^ n13020 ^ 1'b0 ;
  assign n13023 = n3347 | n7008 ;
  assign n13024 = n13022 & ~n13023 ;
  assign n13027 = n1609 & ~n1850 ;
  assign n13028 = n4393 & n13027 ;
  assign n13025 = ( n783 & n1682 ) | ( n783 & ~n4084 ) | ( n1682 & ~n4084 ) ;
  assign n13026 = ~n204 & n13025 ;
  assign n13029 = n13028 ^ n13026 ^ 1'b0 ;
  assign n13030 = ~n5802 & n11865 ;
  assign n13031 = ~n9140 & n13030 ;
  assign n13032 = n3838 & n12975 ;
  assign n13033 = n6023 ^ n5034 ^ 1'b0 ;
  assign n13034 = n6675 & ~n13033 ;
  assign n13035 = n13034 ^ n1393 ^ 1'b0 ;
  assign n13036 = n9565 & ~n10930 ;
  assign n13037 = n13036 ^ n4144 ^ 1'b0 ;
  assign n13038 = ( n1184 & n3178 ) | ( n1184 & n5291 ) | ( n3178 & n5291 ) ;
  assign n13039 = n13038 ^ n4597 ^ 1'b0 ;
  assign n13040 = n6996 & n9984 ;
  assign n13041 = n13040 ^ n5572 ^ n1230 ;
  assign n13042 = ~n9110 & n9307 ;
  assign n13043 = n4135 & n13042 ;
  assign n13044 = n13043 ^ n9346 ^ 1'b0 ;
  assign n13045 = ~n6735 & n9045 ;
  assign n13046 = n13045 ^ n2656 ^ 1'b0 ;
  assign n13047 = n6346 ^ n4839 ^ n1940 ;
  assign n13048 = n13047 ^ n12772 ^ 1'b0 ;
  assign n13049 = n13048 ^ n10780 ^ 1'b0 ;
  assign n13050 = ~n1920 & n2702 ;
  assign n13051 = n6547 | n12034 ;
  assign n13052 = n13050 | n13051 ;
  assign n13053 = n2980 & n11399 ;
  assign n13054 = n13053 ^ n6470 ^ 1'b0 ;
  assign n13055 = n13052 & ~n13054 ;
  assign n13056 = ~n5165 & n13055 ;
  assign n13057 = n3259 | n4348 ;
  assign n13058 = n707 | n13057 ;
  assign n13059 = n13058 ^ n7632 ^ n3698 ;
  assign n13060 = ~n5721 & n10811 ;
  assign n13061 = ( ~n10418 & n13059 ) | ( ~n10418 & n13060 ) | ( n13059 & n13060 ) ;
  assign n13066 = n2987 & ~n12501 ;
  assign n13062 = x79 & n5381 ;
  assign n13063 = n13062 ^ n8378 ^ 1'b0 ;
  assign n13064 = n5675 & ~n13063 ;
  assign n13065 = n6655 & n13064 ;
  assign n13067 = n13066 ^ n13065 ^ 1'b0 ;
  assign n13068 = ~n6311 & n8413 ;
  assign n13069 = n1198 | n13068 ;
  assign n13070 = n13069 ^ n1329 ^ 1'b0 ;
  assign n13071 = n4315 & ~n13070 ;
  assign n13072 = n13071 ^ n2661 ^ 1'b0 ;
  assign n13073 = n5749 & ~n10890 ;
  assign n13074 = n7595 & n13073 ;
  assign n13075 = n13074 ^ n4219 ^ 1'b0 ;
  assign n13076 = n13040 ^ n6617 ^ n5177 ;
  assign n13077 = ~n7560 & n13076 ;
  assign n13078 = x16 & ~n544 ;
  assign n13079 = n13078 ^ n11179 ^ n9999 ;
  assign n13082 = n1963 ^ n1044 ^ 1'b0 ;
  assign n13083 = ~n3995 & n13082 ;
  assign n13080 = n760 & ~n4820 ;
  assign n13081 = n3703 | n13080 ;
  assign n13084 = n13083 ^ n13081 ^ 1'b0 ;
  assign n13085 = n4065 & ~n8774 ;
  assign n13086 = n13084 & n13085 ;
  assign n13087 = n2355 & ~n11344 ;
  assign n13088 = n13087 ^ n8733 ^ 1'b0 ;
  assign n13089 = n530 & n10126 ;
  assign n13090 = n6988 & n13089 ;
  assign n13091 = n7503 & ~n13090 ;
  assign n13092 = n1041 & n13091 ;
  assign n13093 = n9090 ^ n7461 ^ n5920 ;
  assign n13094 = n13093 ^ n8545 ^ 1'b0 ;
  assign n13096 = n765 & n7487 ;
  assign n13097 = n13096 ^ n11017 ^ 1'b0 ;
  assign n13095 = ~n6450 & n9492 ;
  assign n13098 = n13097 ^ n13095 ^ n12650 ;
  assign n13099 = n2023 & ~n6687 ;
  assign n13100 = ~n3489 & n13099 ;
  assign n13101 = x58 & n10266 ;
  assign n13102 = n4974 & ~n5259 ;
  assign n13103 = n1266 & n13102 ;
  assign n13104 = n2208 | n5746 ;
  assign n13105 = n12034 & n13104 ;
  assign n13106 = n12650 ^ n1193 ^ 1'b0 ;
  assign n13107 = n2886 & n13106 ;
  assign n13108 = n13107 ^ n9502 ^ 1'b0 ;
  assign n13109 = n11297 & n13108 ;
  assign n13110 = n474 & ~n7872 ;
  assign n13111 = n13110 ^ n4254 ^ 1'b0 ;
  assign n13112 = n8512 ^ n8190 ^ n1083 ;
  assign n13113 = n2399 | n13112 ;
  assign n13114 = n13113 ^ n5413 ^ n3349 ;
  assign n13115 = n13114 ^ n8753 ^ 1'b0 ;
  assign n13116 = n13111 | n13115 ;
  assign n13117 = n4420 & n6936 ;
  assign n13118 = ~n3788 & n5371 ;
  assign n13119 = ~n13117 & n13118 ;
  assign n13123 = n2748 ^ n925 ^ 1'b0 ;
  assign n13124 = ~n642 & n13123 ;
  assign n13120 = n425 | n3638 ;
  assign n13121 = n13120 ^ n1266 ^ 1'b0 ;
  assign n13122 = ~n4005 & n13121 ;
  assign n13125 = n13124 ^ n13122 ^ n10377 ;
  assign n13126 = n12212 & n13125 ;
  assign n13127 = n726 & n13126 ;
  assign n13128 = n6337 & n13127 ;
  assign n13129 = n13128 ^ n11549 ^ 1'b0 ;
  assign n13130 = n13119 | n13129 ;
  assign n13131 = n4336 ^ n1050 ^ 1'b0 ;
  assign n13132 = n6751 & ~n13131 ;
  assign n13133 = ( n1319 & n2217 ) | ( n1319 & n4851 ) | ( n2217 & n4851 ) ;
  assign n13134 = ~n9496 & n13133 ;
  assign n13135 = n13134 ^ n1492 ^ 1'b0 ;
  assign n13136 = n6705 & n13135 ;
  assign n13137 = n8984 & ~n12318 ;
  assign n13138 = n10376 ^ n1607 ^ 1'b0 ;
  assign n13139 = n6097 ^ n1762 ^ 1'b0 ;
  assign n13140 = n8196 ^ n3281 ^ 1'b0 ;
  assign n13141 = ~n13139 & n13140 ;
  assign n13142 = n8231 ^ n5463 ^ 1'b0 ;
  assign n13143 = ~n3428 & n12659 ;
  assign n13144 = ~n1133 & n13143 ;
  assign n13145 = ( n539 & n13142 ) | ( n539 & n13144 ) | ( n13142 & n13144 ) ;
  assign n13146 = ~n7457 & n12971 ;
  assign n13147 = ~n5085 & n13146 ;
  assign n13148 = ~n1403 & n5763 ;
  assign n13149 = n13148 ^ n6040 ^ 1'b0 ;
  assign n13150 = ~n2399 & n13149 ;
  assign n13151 = ~n8925 & n13150 ;
  assign n13152 = ~n449 & n487 ;
  assign n13153 = ~n4004 & n13152 ;
  assign n13154 = n13153 ^ n1509 ^ 1'b0 ;
  assign n13155 = n1079 & ~n11962 ;
  assign n13156 = ~n13154 & n13155 ;
  assign n13157 = n2148 ^ n1234 ^ 1'b0 ;
  assign n13158 = n12207 & n13157 ;
  assign n13159 = ~n4732 & n5356 ;
  assign n13160 = n8134 & ~n13159 ;
  assign n13161 = n5446 | n7522 ;
  assign n13162 = n2052 | n13161 ;
  assign n13166 = n1236 ^ n742 ^ 1'b0 ;
  assign n13167 = n3670 & ~n13166 ;
  assign n13163 = n1257 & ~n4204 ;
  assign n13164 = n2287 & n13163 ;
  assign n13165 = n13164 ^ n9953 ^ 1'b0 ;
  assign n13168 = n13167 ^ n13165 ^ n12139 ;
  assign n13169 = n6359 | n8537 ;
  assign n13170 = n5409 & ~n11384 ;
  assign n13171 = n12659 ^ n1067 ^ 1'b0 ;
  assign n13172 = ( x70 & n6521 ) | ( x70 & ~n13171 ) | ( n6521 & ~n13171 ) ;
  assign n13173 = ~x7 & n13172 ;
  assign n13174 = n7646 ^ n6199 ^ 1'b0 ;
  assign n13175 = ( n1067 & ~n3066 ) | ( n1067 & n9426 ) | ( ~n3066 & n9426 ) ;
  assign n13176 = n13175 ^ n5468 ^ n1877 ;
  assign n13177 = n5352 & ~n8720 ;
  assign n13178 = n13177 ^ n12132 ^ 1'b0 ;
  assign n13186 = n3166 ^ n1641 ^ 1'b0 ;
  assign n13187 = n3103 & n13186 ;
  assign n13188 = n13187 ^ n11442 ^ 1'b0 ;
  assign n13179 = n3267 & ~n3455 ;
  assign n13180 = n5378 & n13179 ;
  assign n13181 = n13180 ^ n379 ^ 1'b0 ;
  assign n13182 = ~n277 & n2283 ;
  assign n13183 = n655 | n10058 ;
  assign n13184 = n13182 & ~n13183 ;
  assign n13185 = n13181 & ~n13184 ;
  assign n13189 = n13188 ^ n13185 ^ 1'b0 ;
  assign n13190 = n819 | n6872 ;
  assign n13191 = n13190 ^ n12880 ^ 1'b0 ;
  assign n13192 = ~n3208 & n13191 ;
  assign n13193 = ( n2910 & n4119 ) | ( n2910 & ~n13192 ) | ( n4119 & ~n13192 ) ;
  assign n13194 = n2618 | n9963 ;
  assign n13195 = n1549 | n13194 ;
  assign n13196 = n13195 ^ n11547 ^ n8687 ;
  assign n13197 = n771 | n1706 ;
  assign n13198 = n13197 ^ n3041 ^ 1'b0 ;
  assign n13199 = n8526 & ~n13198 ;
  assign n13200 = ~n7520 & n13199 ;
  assign n13201 = n13200 ^ n9201 ^ 1'b0 ;
  assign n13202 = n13196 & n13201 ;
  assign n13203 = n1700 | n3525 ;
  assign n13204 = n4909 & n13203 ;
  assign n13206 = n5717 | n11645 ;
  assign n13207 = n13206 ^ n1641 ^ 1'b0 ;
  assign n13205 = n830 & ~n3066 ;
  assign n13208 = n13207 ^ n13205 ^ 1'b0 ;
  assign n13209 = n2070 & n5790 ;
  assign n13210 = ( n10611 & n13208 ) | ( n10611 & n13209 ) | ( n13208 & n13209 ) ;
  assign n13211 = ~n3117 & n10783 ;
  assign n13212 = n13211 ^ n9268 ^ 1'b0 ;
  assign n13213 = n13212 ^ n8212 ^ 1'b0 ;
  assign n13214 = n10472 ^ n149 ^ 1'b0 ;
  assign n13215 = n13214 ^ n9625 ^ n5785 ;
  assign n13216 = n13215 ^ n8790 ^ 1'b0 ;
  assign n13217 = n760 | n1758 ;
  assign n13218 = n1413 | n9575 ;
  assign n13219 = n13218 ^ n379 ^ 1'b0 ;
  assign n13220 = ~n5297 & n10471 ;
  assign n13221 = n11272 & n13220 ;
  assign n13222 = n4041 & ~n13221 ;
  assign n13223 = n13219 & n13222 ;
  assign n13224 = n13223 ^ n9686 ^ n8776 ;
  assign n13233 = ~n1929 & n2827 ;
  assign n13232 = n5667 ^ n590 ^ 1'b0 ;
  assign n13225 = n3351 & ~n4502 ;
  assign n13226 = ~n1674 & n13225 ;
  assign n13227 = n13226 ^ n5342 ^ 1'b0 ;
  assign n13228 = ~n1111 & n13227 ;
  assign n13229 = n13228 ^ n6670 ^ n3110 ;
  assign n13230 = n9024 ^ n2461 ^ 1'b0 ;
  assign n13231 = n13229 & n13230 ;
  assign n13234 = n13233 ^ n13232 ^ n13231 ;
  assign n13237 = n12977 ^ n3446 ^ n1277 ;
  assign n13238 = n13237 ^ n892 ^ 1'b0 ;
  assign n13239 = n12045 | n13238 ;
  assign n13240 = n13239 ^ n6390 ^ 1'b0 ;
  assign n13235 = n1182 | n6197 ;
  assign n13236 = n7025 | n13235 ;
  assign n13241 = n13240 ^ n13236 ^ 1'b0 ;
  assign n13242 = n1608 & ~n7473 ;
  assign n13243 = n13242 ^ n6584 ^ 1'b0 ;
  assign n13244 = n1423 ^ n990 ^ n752 ;
  assign n13245 = n13244 ^ n3281 ^ 1'b0 ;
  assign n13246 = n13245 ^ n12692 ^ n4197 ;
  assign n13247 = n5459 ^ n2456 ^ 1'b0 ;
  assign n13248 = ~n1765 & n7851 ;
  assign n13249 = n13247 | n13248 ;
  assign n13250 = n13246 & ~n13249 ;
  assign n13251 = n5533 ^ n2429 ^ 1'b0 ;
  assign n13252 = n1722 & ~n13251 ;
  assign n13253 = ( n3591 & ~n4975 ) | ( n3591 & n13252 ) | ( ~n4975 & n13252 ) ;
  assign n13254 = n3344 & ~n6874 ;
  assign n13255 = n13254 ^ n9093 ^ n7973 ;
  assign n13256 = n6497 ^ n4829 ^ 1'b0 ;
  assign n13257 = n8623 ^ n7599 ^ 1'b0 ;
  assign n13258 = n8637 ^ n2189 ^ 1'b0 ;
  assign n13259 = ~n2081 & n6610 ;
  assign n13262 = n673 ^ n257 ^ 1'b0 ;
  assign n13263 = ~n9176 & n13262 ;
  assign n13264 = n5056 & n13263 ;
  assign n13265 = ( n7546 & ~n10569 ) | ( n7546 & n13264 ) | ( ~n10569 & n13264 ) ;
  assign n13260 = n5669 ^ n3518 ^ n1641 ;
  assign n13261 = ~n2642 & n13260 ;
  assign n13266 = n13265 ^ n13261 ^ 1'b0 ;
  assign n13267 = n975 | n13266 ;
  assign n13268 = n1711 & n2818 ;
  assign n13269 = n1765 & n13268 ;
  assign n13270 = ( n7225 & n7496 ) | ( n7225 & n13269 ) | ( n7496 & n13269 ) ;
  assign n13271 = n11420 & ~n13270 ;
  assign n13272 = n13271 ^ n12472 ^ 1'b0 ;
  assign n13273 = n1720 & ~n5366 ;
  assign n13274 = n2521 & n13273 ;
  assign n13275 = n1339 | n3033 ;
  assign n13276 = n13275 ^ n856 ^ 1'b0 ;
  assign n13277 = n13274 | n13276 ;
  assign n13278 = n10355 ^ n470 ^ 1'b0 ;
  assign n13279 = n6027 & ~n13278 ;
  assign n13280 = n10729 ^ n1034 ^ 1'b0 ;
  assign n13281 = n5509 ^ n888 ^ 1'b0 ;
  assign n13282 = n10414 | n13281 ;
  assign n13283 = n11854 ^ n11699 ^ 1'b0 ;
  assign n13284 = n5606 & ~n8311 ;
  assign n13285 = n12711 ^ n8759 ^ n8317 ;
  assign n13286 = n6425 | n6617 ;
  assign n13287 = n13286 ^ n9874 ^ 1'b0 ;
  assign n13288 = n3525 | n6470 ;
  assign n13289 = n13287 & ~n13288 ;
  assign n13290 = n13289 ^ n1504 ^ 1'b0 ;
  assign n13291 = n11477 & n13290 ;
  assign n13292 = n13291 ^ n9489 ^ 1'b0 ;
  assign n13293 = n8038 ^ n6763 ^ n5528 ;
  assign n13294 = n9936 ^ n9814 ^ 1'b0 ;
  assign n13295 = ~n639 & n9925 ;
  assign n13296 = n13295 ^ n1627 ^ 1'b0 ;
  assign n13297 = n648 & ~n13296 ;
  assign n13298 = n5201 ^ n2287 ^ 1'b0 ;
  assign n13299 = n9315 | n13298 ;
  assign n13300 = n13297 & ~n13299 ;
  assign n13301 = n7280 & n13300 ;
  assign n13304 = n194 | n247 ;
  assign n13302 = n4686 ^ n4494 ^ n1067 ;
  assign n13303 = n9200 & ~n13302 ;
  assign n13305 = n13304 ^ n13303 ^ 1'b0 ;
  assign n13306 = n6157 ^ n5686 ^ n3214 ;
  assign n13307 = n10104 ^ n8138 ^ 1'b0 ;
  assign n13308 = ( x93 & n196 ) | ( x93 & ~n13307 ) | ( n196 & ~n13307 ) ;
  assign n13309 = ( n10661 & n13306 ) | ( n10661 & n13308 ) | ( n13306 & n13308 ) ;
  assign n13310 = n9884 ^ n9072 ^ 1'b0 ;
  assign n13311 = n4650 ^ n185 ^ 1'b0 ;
  assign n13312 = ( ~n13219 & n13310 ) | ( ~n13219 & n13311 ) | ( n13310 & n13311 ) ;
  assign n13313 = n4584 ^ n3249 ^ 1'b0 ;
  assign n13314 = n9278 & n13313 ;
  assign n13315 = n7881 ^ n3979 ^ 1'b0 ;
  assign n13316 = n12853 ^ n3258 ^ 1'b0 ;
  assign n13317 = n1406 & ~n8478 ;
  assign n13318 = n13316 & n13317 ;
  assign n13319 = n3639 & ~n9320 ;
  assign n13320 = n13319 ^ n6612 ^ 1'b0 ;
  assign n13321 = n13320 ^ n3036 ^ 1'b0 ;
  assign n13322 = n11026 ^ n10463 ^ 1'b0 ;
  assign n13323 = n3411 ^ n3066 ^ 1'b0 ;
  assign n13324 = n4355 | n9035 ;
  assign n13325 = n13324 ^ n1567 ^ 1'b0 ;
  assign n13326 = n9800 ^ n8058 ^ 1'b0 ;
  assign n13327 = n2241 & ~n12430 ;
  assign n13328 = n1906 ^ n712 ^ 1'b0 ;
  assign n13329 = ~n4130 & n13328 ;
  assign n13330 = ~n13002 & n13329 ;
  assign n13331 = n13330 ^ n11466 ^ 1'b0 ;
  assign n13332 = n1341 | n2706 ;
  assign n13333 = n13332 ^ n2900 ^ 1'b0 ;
  assign n13334 = n7688 | n10106 ;
  assign n13335 = n1311 & ~n11633 ;
  assign n13336 = n3985 | n13335 ;
  assign n13337 = n11985 & ~n13336 ;
  assign n13338 = n701 | n9527 ;
  assign n13339 = n5178 ^ n4439 ^ n532 ;
  assign n13340 = n13339 ^ n869 ^ 1'b0 ;
  assign n13341 = n2345 | n13340 ;
  assign n13342 = n1578 & ~n13341 ;
  assign n13343 = n8067 | n9918 ;
  assign n13344 = ( n6048 & ~n13342 ) | ( n6048 & n13343 ) | ( ~n13342 & n13343 ) ;
  assign n13345 = n6590 | n7547 ;
  assign n13346 = n3446 & ~n13345 ;
  assign n13347 = n6805 & ~n13346 ;
  assign n13348 = n4180 | n13347 ;
  assign n13349 = ( n3639 & n3882 ) | ( n3639 & n4739 ) | ( n3882 & n4739 ) ;
  assign n13350 = ~n2788 & n13349 ;
  assign n13351 = ~n2229 & n7410 ;
  assign n13352 = ~n884 & n2353 ;
  assign n13353 = ( n2431 & n13351 ) | ( n2431 & ~n13352 ) | ( n13351 & ~n13352 ) ;
  assign n13354 = n7271 ^ x41 ^ 1'b0 ;
  assign n13355 = n12535 ^ n5790 ^ 1'b0 ;
  assign n13356 = n13153 | n13355 ;
  assign n13357 = n13354 | n13356 ;
  assign n13358 = n13357 ^ n3135 ^ 1'b0 ;
  assign n13359 = n2461 & ~n7229 ;
  assign n13360 = ~x36 & n13359 ;
  assign n13361 = n2692 & n13360 ;
  assign n13362 = n5330 & ~n13361 ;
  assign n13363 = n13362 ^ n259 ^ 1'b0 ;
  assign n13364 = n13363 ^ n8619 ^ n2510 ;
  assign n13365 = n758 & ~n8334 ;
  assign n13366 = ~n1222 & n13365 ;
  assign n13367 = n13366 ^ n13207 ^ 1'b0 ;
  assign n13368 = n3648 & ~n8581 ;
  assign n13369 = ( n10456 & n12752 ) | ( n10456 & ~n13368 ) | ( n12752 & ~n13368 ) ;
  assign n13370 = n3708 ^ n2020 ^ n1320 ;
  assign n13371 = ~n8371 & n13370 ;
  assign n13372 = n13371 ^ n6937 ^ 1'b0 ;
  assign n13373 = ~n6576 & n9008 ;
  assign n13374 = ~n6004 & n13373 ;
  assign n13375 = ( ~n6655 & n13372 ) | ( ~n6655 & n13374 ) | ( n13372 & n13374 ) ;
  assign n13376 = n631 & ~n9703 ;
  assign n13377 = n6705 | n8872 ;
  assign n13378 = n13377 ^ n8341 ^ 1'b0 ;
  assign n13379 = n3424 & ~n11017 ;
  assign n13380 = n6117 & n13379 ;
  assign n13381 = n3351 ^ n672 ^ 1'b0 ;
  assign n13382 = n1909 & n13381 ;
  assign n13383 = n12246 ^ n6209 ^ n703 ;
  assign n13384 = n13383 ^ n6815 ^ 1'b0 ;
  assign n13385 = n8377 & ~n13384 ;
  assign n13386 = ~n5536 & n7726 ;
  assign n13387 = n13386 ^ n11833 ^ 1'b0 ;
  assign n13388 = n10650 & n12185 ;
  assign n13389 = n5967 ^ n1019 ^ 1'b0 ;
  assign n13390 = n1439 ^ n438 ^ 1'b0 ;
  assign n13391 = ~n8212 & n13390 ;
  assign n13392 = n5687 ^ x70 ^ 1'b0 ;
  assign n13393 = n4534 ^ x120 ^ 1'b0 ;
  assign n13394 = n10613 & n13393 ;
  assign n13395 = n13394 ^ n7430 ^ 1'b0 ;
  assign n13396 = n4446 & ~n4773 ;
  assign n13397 = ~n4446 & n13396 ;
  assign n13398 = n13397 ^ n835 ^ 1'b0 ;
  assign n13399 = n2285 ^ n2005 ^ 1'b0 ;
  assign n13400 = n13399 ^ n2011 ^ 1'b0 ;
  assign n13401 = n13400 ^ n5324 ^ 1'b0 ;
  assign n13402 = n13398 & n13401 ;
  assign n13403 = n935 ^ n726 ^ 1'b0 ;
  assign n13404 = n901 & n13403 ;
  assign n13405 = ~n425 & n13404 ;
  assign n13406 = n9562 & ~n13200 ;
  assign n13407 = n10544 ^ n7776 ^ 1'b0 ;
  assign n13408 = n1650 & ~n13407 ;
  assign n13409 = n13048 ^ n6264 ^ n5041 ;
  assign n13411 = x119 & ~n4157 ;
  assign n13412 = n13411 ^ n4430 ^ 1'b0 ;
  assign n13410 = n7416 ^ n6976 ^ n3879 ;
  assign n13413 = n13412 ^ n13410 ^ 1'b0 ;
  assign n13414 = n7471 ^ n2933 ^ 1'b0 ;
  assign n13415 = n13414 ^ n11894 ^ n3738 ;
  assign n13416 = x2 & n7223 ;
  assign n13417 = ~n11504 & n13416 ;
  assign n13418 = ~n2459 & n6808 ;
  assign n13419 = n13418 ^ n8085 ^ 1'b0 ;
  assign n13420 = n1671 ^ n771 ^ 1'b0 ;
  assign n13421 = n13419 | n13420 ;
  assign n13422 = n2976 & ~n10588 ;
  assign n13424 = n1818 & n3179 ;
  assign n13423 = n461 & ~n7799 ;
  assign n13425 = n13424 ^ n13423 ^ 1'b0 ;
  assign n13426 = ( n5881 & n7920 ) | ( n5881 & ~n13425 ) | ( n7920 & ~n13425 ) ;
  assign n13427 = n13426 ^ n12402 ^ n8024 ;
  assign n13428 = n8515 ^ n7402 ^ 1'b0 ;
  assign n13429 = ~n1765 & n7653 ;
  assign n13430 = ( n12023 & n13428 ) | ( n12023 & ~n13429 ) | ( n13428 & ~n13429 ) ;
  assign n13431 = n3975 & n5156 ;
  assign n13432 = n5487 ^ n1953 ^ n703 ;
  assign n13433 = n13432 ^ n5211 ^ n3986 ;
  assign n13434 = ( ~n2930 & n8983 ) | ( ~n2930 & n13433 ) | ( n8983 & n13433 ) ;
  assign n13435 = n4017 & ~n5072 ;
  assign n13436 = n370 & ~n2259 ;
  assign n13437 = n13436 ^ n2529 ^ 1'b0 ;
  assign n13438 = n1014 | n11402 ;
  assign n13439 = n13437 | n13438 ;
  assign n13440 = ~n5304 & n8924 ;
  assign n13441 = ~n13439 & n13440 ;
  assign n13442 = n2751 | n9653 ;
  assign n13443 = n2751 & ~n13442 ;
  assign n13444 = n2391 & n13443 ;
  assign n13445 = ~n2608 & n3602 ;
  assign n13446 = n3625 & n13445 ;
  assign n13447 = ~n13444 & n13446 ;
  assign n13448 = n11111 ^ n672 ^ 1'b0 ;
  assign n13449 = n13448 ^ n6833 ^ n1275 ;
  assign n13450 = n10649 ^ n9773 ^ 1'b0 ;
  assign n13451 = n13450 ^ n11868 ^ 1'b0 ;
  assign n13452 = n13449 & ~n13451 ;
  assign n13453 = n2543 & ~n3672 ;
  assign n13454 = n13453 ^ n264 ^ 1'b0 ;
  assign n13455 = n13454 ^ n2665 ^ 1'b0 ;
  assign n13456 = n1677 & ~n3741 ;
  assign n13457 = n13456 ^ n5692 ^ 1'b0 ;
  assign n13458 = ~n2897 & n13457 ;
  assign n13464 = n2999 ^ n1323 ^ 1'b0 ;
  assign n13459 = n1380 ^ n919 ^ 1'b0 ;
  assign n13460 = ~n1410 & n13459 ;
  assign n13461 = n9887 ^ n8820 ^ 1'b0 ;
  assign n13462 = n13460 & ~n13461 ;
  assign n13463 = ~n9328 & n13462 ;
  assign n13465 = n13464 ^ n13463 ^ 1'b0 ;
  assign n13466 = x61 & ~n10424 ;
  assign n13467 = ~n6496 & n13466 ;
  assign n13468 = n13467 ^ n6575 ^ 1'b0 ;
  assign n13469 = n1291 | n13468 ;
  assign n13471 = n4205 | n10286 ;
  assign n13470 = ~n159 & n7626 ;
  assign n13472 = n13471 ^ n13470 ^ 1'b0 ;
  assign n13473 = n8510 ^ n7218 ^ n4462 ;
  assign n13480 = ~n7495 & n10747 ;
  assign n13481 = n13480 ^ n10066 ^ 1'b0 ;
  assign n13482 = ~n606 & n13481 ;
  assign n13483 = n13482 ^ n7167 ^ 1'b0 ;
  assign n13484 = ( n708 & n5394 ) | ( n708 & ~n13483 ) | ( n5394 & ~n13483 ) ;
  assign n13485 = n6243 ^ n6073 ^ 1'b0 ;
  assign n13486 = n9348 | n13485 ;
  assign n13487 = n3253 & ~n13486 ;
  assign n13488 = ~n13484 & n13487 ;
  assign n13474 = n4320 | n7178 ;
  assign n13475 = n1668 | n5163 ;
  assign n13476 = n13474 & ~n13475 ;
  assign n13477 = n4410 ^ n1861 ^ 1'b0 ;
  assign n13478 = ~n13476 & n13477 ;
  assign n13479 = n10064 & n13478 ;
  assign n13489 = n13488 ^ n13479 ^ 1'b0 ;
  assign n13495 = n4070 | n7452 ;
  assign n13496 = n6816 | n13495 ;
  assign n13491 = n2836 & ~n3025 ;
  assign n13490 = n7021 & ~n11985 ;
  assign n13492 = n13491 ^ n13490 ^ 1'b0 ;
  assign n13493 = n13492 ^ n11531 ^ n1111 ;
  assign n13494 = n7756 & n13493 ;
  assign n13497 = n13496 ^ n13494 ^ 1'b0 ;
  assign n13498 = n2806 & ~n8652 ;
  assign n13499 = n13498 ^ n11562 ^ 1'b0 ;
  assign n13500 = n13499 ^ n6168 ^ 1'b0 ;
  assign n13501 = n13497 | n13500 ;
  assign n13502 = n1337 | n1811 ;
  assign n13503 = n8444 & ~n13502 ;
  assign n13504 = n13503 ^ n4281 ^ 1'b0 ;
  assign n13505 = n13504 ^ n3776 ^ 1'b0 ;
  assign n13506 = ~n4942 & n10971 ;
  assign n13507 = n6824 & n10583 ;
  assign n13508 = n13507 ^ n1624 ^ 1'b0 ;
  assign n13509 = n11199 ^ n3199 ^ 1'b0 ;
  assign n13510 = n12420 ^ n7666 ^ 1'b0 ;
  assign n13511 = n2106 & ~n3152 ;
  assign n13512 = n13511 ^ n3067 ^ 1'b0 ;
  assign n13513 = n13512 ^ n8761 ^ 1'b0 ;
  assign n13514 = n3488 | n13513 ;
  assign n13515 = ~n5387 & n9278 ;
  assign n13516 = n13515 ^ n3933 ^ 1'b0 ;
  assign n13517 = n5953 & ~n10306 ;
  assign n13518 = n13517 ^ n6617 ^ 1'b0 ;
  assign n13519 = n1677 | n1768 ;
  assign n13520 = n5731 & ~n13519 ;
  assign n13521 = n5986 | n13520 ;
  assign n13522 = n13521 ^ n12938 ^ 1'b0 ;
  assign n13523 = n13275 ^ n4076 ^ 1'b0 ;
  assign n13524 = n12195 & n13523 ;
  assign n13525 = n399 & n6580 ;
  assign n13526 = n337 ^ x13 ^ 1'b0 ;
  assign n13527 = n8903 ^ n269 ^ 1'b0 ;
  assign n13528 = n8512 | n13527 ;
  assign n13529 = ~n12079 & n13528 ;
  assign n13530 = n6439 ^ n4760 ^ n3468 ;
  assign n13531 = n7490 & n13530 ;
  assign n13532 = n13531 ^ n11414 ^ 1'b0 ;
  assign n13533 = n13532 ^ n9863 ^ n5265 ;
  assign n13534 = n3652 | n10387 ;
  assign n13535 = n13533 | n13534 ;
  assign n13537 = n6317 ^ n4300 ^ 1'b0 ;
  assign n13538 = n1308 | n13537 ;
  assign n13536 = ~n134 & n2609 ;
  assign n13539 = n13538 ^ n13536 ^ 1'b0 ;
  assign n13540 = n13535 & n13539 ;
  assign n13541 = ~n2323 & n3476 ;
  assign n13542 = n13541 ^ n7615 ^ 1'b0 ;
  assign n13543 = ~n4230 & n8678 ;
  assign n13544 = n13543 ^ n1000 ^ x96 ;
  assign n13549 = ( n603 & n1521 ) | ( n603 & n4757 ) | ( n1521 & n4757 ) ;
  assign n13548 = ( n425 & n1542 ) | ( n425 & n4420 ) | ( n1542 & n4420 ) ;
  assign n13550 = n13549 ^ n13548 ^ n2526 ;
  assign n13545 = x63 | n3828 ;
  assign n13546 = n1051 | n12610 ;
  assign n13547 = n13545 & ~n13546 ;
  assign n13551 = n13550 ^ n13547 ^ 1'b0 ;
  assign n13552 = ( n8281 & ~n12845 ) | ( n8281 & n13551 ) | ( ~n12845 & n13551 ) ;
  assign n13553 = n4821 ^ n2036 ^ 1'b0 ;
  assign n13554 = n13047 ^ n758 ^ 1'b0 ;
  assign n13555 = n1424 ^ n632 ^ 1'b0 ;
  assign n13556 = n13554 & ~n13555 ;
  assign n13557 = ~n1880 & n5554 ;
  assign n13558 = n13557 ^ n3533 ^ 1'b0 ;
  assign n13559 = n1578 ^ x110 ^ 1'b0 ;
  assign n13560 = n10325 & ~n13559 ;
  assign n13561 = n13560 ^ n8657 ^ 1'b0 ;
  assign n13562 = ~n1774 & n13561 ;
  assign n13563 = ~n8520 & n13562 ;
  assign n13564 = n6051 & n12384 ;
  assign n13565 = ~n1968 & n3339 ;
  assign n13566 = ~x22 & n13565 ;
  assign n13567 = n12610 ^ n10637 ^ 1'b0 ;
  assign n13568 = n13567 ^ n2569 ^ 1'b0 ;
  assign n13569 = n1041 ^ n159 ^ 1'b0 ;
  assign n13570 = n1766 & ~n13569 ;
  assign n13571 = ~n1540 & n6546 ;
  assign n13572 = ~n13570 & n13571 ;
  assign n13573 = n5031 | n12546 ;
  assign n13575 = ~n6860 & n12977 ;
  assign n13576 = n13575 ^ n9889 ^ 1'b0 ;
  assign n13577 = n13576 ^ x14 ^ 1'b0 ;
  assign n13578 = n5629 ^ n1692 ^ 1'b0 ;
  assign n13579 = ~n2255 & n13578 ;
  assign n13580 = n13577 & n13579 ;
  assign n13574 = ~n6450 & n12198 ;
  assign n13581 = n13580 ^ n13574 ^ 1'b0 ;
  assign n13582 = n11890 ^ n7988 ^ 1'b0 ;
  assign n13583 = n2940 & n13582 ;
  assign n13584 = n6095 ^ n3113 ^ 1'b0 ;
  assign n13585 = ( ~n4204 & n8913 ) | ( ~n4204 & n13584 ) | ( n8913 & n13584 ) ;
  assign n13586 = n13467 ^ n8856 ^ n8706 ;
  assign n13587 = n12995 & n13586 ;
  assign n13588 = n2369 | n3085 ;
  assign n13589 = n2414 & ~n13588 ;
  assign n13590 = n13589 ^ n1311 ^ 1'b0 ;
  assign n13591 = n3590 & ~n13590 ;
  assign n13592 = n13591 ^ n1760 ^ 1'b0 ;
  assign n13593 = n7579 ^ n2461 ^ n2282 ;
  assign n13594 = n13593 ^ n8914 ^ 1'b0 ;
  assign n13595 = n3542 ^ n1808 ^ 1'b0 ;
  assign n13596 = n6264 ^ n828 ^ 1'b0 ;
  assign n13597 = n2107 ^ n1913 ^ 1'b0 ;
  assign n13598 = n1186 & ~n13597 ;
  assign n13599 = n13598 ^ n7119 ^ 1'b0 ;
  assign n13600 = ~n1420 & n7497 ;
  assign n13601 = n4122 & n13600 ;
  assign n13602 = n2983 & ~n3703 ;
  assign n13603 = n1021 & n11866 ;
  assign n13604 = ~n690 & n13603 ;
  assign n13605 = n2160 & ~n13604 ;
  assign n13606 = n13605 ^ n8253 ^ 1'b0 ;
  assign n13607 = n13565 ^ n5432 ^ 1'b0 ;
  assign n13608 = n13606 & ~n13607 ;
  assign n13609 = n1345 & n7383 ;
  assign n13610 = ~n6468 & n13609 ;
  assign n13611 = ~n877 & n1513 ;
  assign n13612 = ~n676 & n13611 ;
  assign n13613 = n1269 | n13612 ;
  assign n13614 = n3336 | n13613 ;
  assign n13615 = n5916 ^ n2173 ^ 1'b0 ;
  assign n13616 = n13615 ^ n3811 ^ 1'b0 ;
  assign n13617 = n2956 & ~n7032 ;
  assign n13618 = ( x47 & n1069 ) | ( x47 & n1257 ) | ( n1069 & n1257 ) ;
  assign n13619 = ~n11957 & n13618 ;
  assign n13620 = n13619 ^ n7987 ^ 1'b0 ;
  assign n13621 = n3377 & n8146 ;
  assign n13622 = n4817 & n13621 ;
  assign n13623 = n4880 & ~n13622 ;
  assign n13624 = n13620 & n13623 ;
  assign n13625 = n4465 & ~n5043 ;
  assign n13626 = ~n6068 & n13625 ;
  assign n13627 = n13626 ^ n10215 ^ 1'b0 ;
  assign n13628 = n11604 & n13627 ;
  assign n13629 = n393 & ~n11656 ;
  assign n13634 = n2256 & n2443 ;
  assign n13635 = n3625 & n13634 ;
  assign n13630 = n4932 & ~n6970 ;
  assign n13631 = ( ~n606 & n3624 ) | ( ~n606 & n13630 ) | ( n3624 & n13630 ) ;
  assign n13632 = n4254 ^ n2109 ^ 1'b0 ;
  assign n13633 = n13631 & ~n13632 ;
  assign n13636 = n13635 ^ n13633 ^ 1'b0 ;
  assign n13637 = n4263 & ~n13636 ;
  assign n13638 = n1472 & n8106 ;
  assign n13639 = n13638 ^ n9615 ^ n2643 ;
  assign n13640 = n11940 ^ n11340 ^ 1'b0 ;
  assign n13641 = n954 & n13640 ;
  assign n13642 = ~n5480 & n7382 ;
  assign n13643 = n8804 & n13642 ;
  assign n13645 = n2751 | n3340 ;
  assign n13644 = n4881 ^ n3113 ^ 1'b0 ;
  assign n13646 = n13645 ^ n13644 ^ 1'b0 ;
  assign n13647 = ~n1517 & n5363 ;
  assign n13648 = n13647 ^ n1698 ^ 1'b0 ;
  assign n13649 = n4136 ^ n869 ^ x38 ;
  assign n13650 = n561 & ~n13649 ;
  assign n13651 = n13648 & n13650 ;
  assign n13652 = n13651 ^ n13391 ^ 1'b0 ;
  assign n13653 = ~n984 & n4455 ;
  assign n13654 = n1089 & ~n6787 ;
  assign n13655 = n5288 & n13654 ;
  assign n13656 = ( n2291 & ~n13653 ) | ( n2291 & n13655 ) | ( ~n13653 & n13655 ) ;
  assign n13657 = n10650 ^ n7827 ^ 1'b0 ;
  assign n13658 = n3849 & n13657 ;
  assign n13659 = n10281 ^ n4489 ^ n1306 ;
  assign n13660 = ( n4581 & n5165 ) | ( n4581 & n10312 ) | ( n5165 & n10312 ) ;
  assign n13661 = ( n1139 & ~n3803 ) | ( n1139 & n4987 ) | ( ~n3803 & n4987 ) ;
  assign n13662 = n13661 ^ n706 ^ 1'b0 ;
  assign n13663 = n5858 & ~n13662 ;
  assign n13665 = n2870 & n4231 ;
  assign n13666 = n13665 ^ n4648 ^ 1'b0 ;
  assign n13667 = n13666 ^ n12647 ^ n11966 ;
  assign n13664 = x55 | n6283 ;
  assign n13668 = n13667 ^ n13664 ^ 1'b0 ;
  assign n13669 = n13668 ^ n1688 ^ 1'b0 ;
  assign n13670 = n4180 | n11474 ;
  assign n13671 = n939 & n10751 ;
  assign n13672 = n13671 ^ n2634 ^ n210 ;
  assign n13673 = n12319 ^ n7368 ^ n4827 ;
  assign n13674 = ( ~n1559 & n1589 ) | ( ~n1559 & n5671 ) | ( n1589 & n5671 ) ;
  assign n13675 = n13674 ^ n7733 ^ 1'b0 ;
  assign n13676 = n6327 & n10420 ;
  assign n13677 = n5401 & n9602 ;
  assign n13678 = n13677 ^ n2952 ^ 1'b0 ;
  assign n13679 = ( n9910 & ~n11046 ) | ( n9910 & n13678 ) | ( ~n11046 & n13678 ) ;
  assign n13680 = n6284 & ~n8877 ;
  assign n13681 = n13680 ^ n6087 ^ n2364 ;
  assign n13682 = ( n1841 & n6741 ) | ( n1841 & n11836 ) | ( n6741 & n11836 ) ;
  assign n13683 = ~n12435 & n13682 ;
  assign n13684 = n13683 ^ n12371 ^ 1'b0 ;
  assign n13685 = ~n740 & n13684 ;
  assign n13691 = ( n6623 & n7311 ) | ( n6623 & ~n9137 ) | ( n7311 & ~n9137 ) ;
  assign n13688 = n3981 ^ x57 ^ 1'b0 ;
  assign n13689 = n5250 & ~n13688 ;
  assign n13690 = n6558 & ~n13689 ;
  assign n13692 = n13691 ^ n13690 ^ 1'b0 ;
  assign n13686 = n12942 ^ n8739 ^ 1'b0 ;
  assign n13687 = n11905 & ~n13686 ;
  assign n13693 = n13692 ^ n13687 ^ 1'b0 ;
  assign n13694 = n764 & ~n10538 ;
  assign n13695 = n4677 ^ n2934 ^ 1'b0 ;
  assign n13698 = ~n1765 & n4012 ;
  assign n13697 = n551 | n8422 ;
  assign n13699 = n13698 ^ n13697 ^ 1'b0 ;
  assign n13700 = n4707 | n13699 ;
  assign n13701 = n13700 ^ n6753 ^ n5123 ;
  assign n13702 = ~n3664 & n13701 ;
  assign n13703 = n13702 ^ n10364 ^ 1'b0 ;
  assign n13696 = n1467 & ~n7616 ;
  assign n13704 = n13703 ^ n13696 ^ 1'b0 ;
  assign n13705 = n5763 & n8258 ;
  assign n13706 = n4285 & n13705 ;
  assign n13707 = n7090 & ~n13706 ;
  assign n13708 = n11298 ^ n10173 ^ n8545 ;
  assign n13709 = n4508 | n11446 ;
  assign n13710 = n13709 ^ n12883 ^ n1308 ;
  assign n13711 = n7953 | n11645 ;
  assign n13712 = n4837 & ~n13711 ;
  assign n13713 = ~n3957 & n11556 ;
  assign n13714 = n13713 ^ n8528 ^ 1'b0 ;
  assign n13715 = n13712 & n13714 ;
  assign n13716 = n1181 | n6023 ;
  assign n13717 = n10762 | n13716 ;
  assign n13718 = n2944 ^ n1111 ^ 1'b0 ;
  assign n13719 = n2325 | n3906 ;
  assign n13720 = n13719 ^ n7295 ^ 1'b0 ;
  assign n13721 = n6689 ^ n3319 ^ 1'b0 ;
  assign n13722 = ~n10424 & n13721 ;
  assign n13723 = ( n5833 & n13720 ) | ( n5833 & n13722 ) | ( n13720 & n13722 ) ;
  assign n13724 = n7550 ^ n7100 ^ 1'b0 ;
  assign n13725 = ( ~n4907 & n11366 ) | ( ~n4907 & n13724 ) | ( n11366 & n13724 ) ;
  assign n13726 = n4684 ^ x102 ^ 1'b0 ;
  assign n13727 = n3254 | n7135 ;
  assign n13728 = n13727 ^ n9929 ^ 1'b0 ;
  assign n13729 = n12060 & ~n13377 ;
  assign n13730 = n10060 ^ n8909 ^ 1'b0 ;
  assign n13731 = n10168 & ~n13730 ;
  assign n13732 = n11102 & n13731 ;
  assign n13733 = n1365 & n1533 ;
  assign n13734 = n4429 & ~n13733 ;
  assign n13735 = ~n13732 & n13734 ;
  assign n13736 = n3585 & n10626 ;
  assign n13737 = ~n3046 & n13736 ;
  assign n13738 = n9167 ^ n5468 ^ n1630 ;
  assign n13739 = n13738 ^ n6281 ^ 1'b0 ;
  assign n13740 = n10188 ^ n4208 ^ n3156 ;
  assign n13741 = n13740 ^ n9237 ^ 1'b0 ;
  assign n13744 = n4034 ^ n3043 ^ 1'b0 ;
  assign n13742 = n1870 & ~n13112 ;
  assign n13743 = n13742 ^ n8355 ^ 1'b0 ;
  assign n13745 = n13744 ^ n13743 ^ 1'b0 ;
  assign n13746 = n6701 & ~n13745 ;
  assign n13747 = n11691 ^ n5687 ^ 1'b0 ;
  assign n13748 = n3831 ^ n1008 ^ 1'b0 ;
  assign n13749 = n13747 & ~n13748 ;
  assign n13750 = ~n196 & n13749 ;
  assign n13751 = n13671 & n13750 ;
  assign n13752 = n3387 ^ n1887 ^ n740 ;
  assign n13753 = n13751 | n13752 ;
  assign n13754 = ~n1086 & n12405 ;
  assign n13755 = n7632 & n13754 ;
  assign n13756 = n8048 ^ n4806 ^ 1'b0 ;
  assign n13757 = ~n5415 & n5477 ;
  assign n13758 = n7602 & n13757 ;
  assign n13759 = n4522 & ~n13758 ;
  assign n13760 = n13526 ^ n1519 ^ 1'b0 ;
  assign n13761 = n13760 ^ n2903 ^ 1'b0 ;
  assign n13762 = n6154 & n13761 ;
  assign n13763 = n442 | n5752 ;
  assign n13764 = n13763 ^ n366 ^ 1'b0 ;
  assign n13765 = n5613 ^ n4933 ^ n2900 ;
  assign n13766 = ~n3470 & n5715 ;
  assign n13767 = n13765 & n13766 ;
  assign n13768 = n13767 ^ n7654 ^ 1'b0 ;
  assign n13769 = ~n3067 & n13768 ;
  assign n13770 = n13764 & n13769 ;
  assign n13771 = n13770 ^ n5497 ^ 1'b0 ;
  assign n13772 = n6770 ^ n3056 ^ 1'b0 ;
  assign n13773 = n12814 & ~n13772 ;
  assign n13774 = n3447 ^ n1277 ^ 1'b0 ;
  assign n13775 = n730 & n13275 ;
  assign n13776 = n13775 ^ n3859 ^ 1'b0 ;
  assign n13777 = n11097 | n13776 ;
  assign n13780 = n1630 | n3105 ;
  assign n13778 = ~n3811 & n13124 ;
  assign n13779 = n3158 & ~n13778 ;
  assign n13781 = n13780 ^ n13779 ^ 1'b0 ;
  assign n13783 = n755 | n2839 ;
  assign n13784 = n13783 ^ n7461 ^ 1'b0 ;
  assign n13782 = n4472 & n5589 ;
  assign n13785 = n13784 ^ n13782 ^ 1'b0 ;
  assign n13786 = ~x40 & n11190 ;
  assign n13787 = ( ~n2673 & n8878 ) | ( ~n2673 & n10530 ) | ( n8878 & n10530 ) ;
  assign n13788 = n13787 ^ n13554 ^ 1'b0 ;
  assign n13789 = n13786 | n13788 ;
  assign n13794 = n5785 ^ n1752 ^ 1'b0 ;
  assign n13795 = ~n3066 & n13794 ;
  assign n13792 = n2498 | n6046 ;
  assign n13793 = n5499 & ~n13792 ;
  assign n13796 = n13795 ^ n13793 ^ 1'b0 ;
  assign n13790 = n2260 & ~n9751 ;
  assign n13791 = n7420 & n13790 ;
  assign n13797 = n13796 ^ n13791 ^ n10780 ;
  assign n13798 = n3441 & ~n4946 ;
  assign n13799 = n13798 ^ n3739 ^ 1'b0 ;
  assign n13801 = n8697 ^ n6151 ^ n2489 ;
  assign n13800 = n1734 & ~n3452 ;
  assign n13802 = n13801 ^ n13800 ^ 1'b0 ;
  assign n13803 = ( n5600 & n13799 ) | ( n5600 & n13802 ) | ( n13799 & n13802 ) ;
  assign n13804 = n13803 ^ n5517 ^ 1'b0 ;
  assign n13805 = n3284 & n13804 ;
  assign n13806 = n13526 ^ n1450 ^ 1'b0 ;
  assign n13807 = ~n4309 & n13806 ;
  assign n13808 = n13807 ^ n9031 ^ 1'b0 ;
  assign n13813 = n808 | n2836 ;
  assign n13814 = n1165 | n13813 ;
  assign n13809 = n2151 & ~n3896 ;
  assign n13810 = n2720 & n13809 ;
  assign n13811 = n7578 & n13810 ;
  assign n13812 = n9524 & ~n13811 ;
  assign n13815 = n13814 ^ n13812 ^ 1'b0 ;
  assign n13816 = ( n4962 & ~n13808 ) | ( n4962 & n13815 ) | ( ~n13808 & n13815 ) ;
  assign n13817 = n1802 | n8835 ;
  assign n13818 = n2671 & ~n13816 ;
  assign n13819 = n368 | n13190 ;
  assign n13820 = n4757 & ~n10387 ;
  assign n13821 = n13224 & n13820 ;
  assign n13822 = n13821 ^ n422 ^ 1'b0 ;
  assign n13823 = ~n3403 & n4272 ;
  assign n13824 = n13823 ^ n4199 ^ 1'b0 ;
  assign n13825 = ( n10610 & n12277 ) | ( n10610 & n13824 ) | ( n12277 & n13824 ) ;
  assign n13827 = n11178 ^ n1680 ^ 1'b0 ;
  assign n13828 = ( n9175 & n12228 ) | ( n9175 & n13827 ) | ( n12228 & n13827 ) ;
  assign n13826 = n1841 & n7806 ;
  assign n13829 = n13828 ^ n13826 ^ 1'b0 ;
  assign n13830 = n13829 ^ n4769 ^ 1'b0 ;
  assign n13831 = ~n4113 & n10395 ;
  assign n13832 = n13831 ^ n12847 ^ 1'b0 ;
  assign n13833 = n8455 ^ n3639 ^ 1'b0 ;
  assign n13834 = ~n937 & n13833 ;
  assign n13835 = n261 & ~n13834 ;
  assign n13836 = n6969 ^ n6297 ^ n2277 ;
  assign n13837 = n740 & ~n6169 ;
  assign n13838 = n7123 ^ n5057 ^ n703 ;
  assign n13839 = ( n1154 & n7231 ) | ( n1154 & n13838 ) | ( n7231 & n13838 ) ;
  assign n13840 = ~n4561 & n7230 ;
  assign n13841 = n1034 ^ x40 ^ 1'b0 ;
  assign n13842 = n1564 & ~n13841 ;
  assign n13843 = n461 & ~n13842 ;
  assign n13844 = n13843 ^ n6003 ^ 1'b0 ;
  assign n13845 = n10847 ^ n1971 ^ 1'b0 ;
  assign n13846 = n9610 ^ n7575 ^ 1'b0 ;
  assign n13847 = n10619 & n11881 ;
  assign n13848 = n13846 & n13847 ;
  assign n13849 = n8085 & n11396 ;
  assign n13850 = n13849 ^ n4851 ^ 1'b0 ;
  assign n13851 = n8107 & n13850 ;
  assign n13852 = n10469 ^ n1645 ^ 1'b0 ;
  assign n13853 = n9039 | n13852 ;
  assign n13854 = x24 & ~n2770 ;
  assign n13855 = n13854 ^ n4441 ^ 1'b0 ;
  assign n13856 = n13855 ^ n5865 ^ 1'b0 ;
  assign n13857 = ~n1475 & n10788 ;
  assign n13858 = n177 & n13857 ;
  assign n13859 = ( n2994 & ~n13476 ) | ( n2994 & n13641 ) | ( ~n13476 & n13641 ) ;
  assign n13860 = ( ~n9334 & n10262 ) | ( ~n9334 & n11401 ) | ( n10262 & n11401 ) ;
  assign n13861 = n1162 & n1758 ;
  assign n13862 = ~n13860 & n13861 ;
  assign n13863 = n3376 ^ n1974 ^ 1'b0 ;
  assign n13864 = ~n3597 & n13863 ;
  assign n13865 = ( n8169 & n12767 ) | ( n8169 & n13864 ) | ( n12767 & n13864 ) ;
  assign n13866 = n10125 ^ n2195 ^ 1'b0 ;
  assign n13867 = ~n13865 & n13866 ;
  assign n13868 = n5013 ^ n2827 ^ n868 ;
  assign n13869 = n4317 | n13868 ;
  assign n13870 = n13869 ^ n11115 ^ n10623 ;
  assign n13871 = n13867 & ~n13870 ;
  assign n13872 = n13871 ^ n6208 ^ 1'b0 ;
  assign n13873 = n13872 ^ n7806 ^ 1'b0 ;
  assign n13874 = n8946 & ~n13873 ;
  assign n13875 = n2307 & ~n13874 ;
  assign n13876 = n2696 | n10240 ;
  assign n13877 = n11115 & ~n13876 ;
  assign n13878 = n8748 & n10554 ;
  assign n13879 = n13878 ^ n8752 ^ 1'b0 ;
  assign n13880 = n13879 ^ n11426 ^ 1'b0 ;
  assign n13881 = n11327 ^ n3143 ^ 1'b0 ;
  assign n13882 = ~n5539 & n13881 ;
  assign n13883 = n6996 ^ n1726 ^ 1'b0 ;
  assign n13884 = ~n10300 & n13883 ;
  assign n13885 = ~n7949 & n13884 ;
  assign n13886 = ~n13882 & n13885 ;
  assign n13887 = ~n6202 & n13886 ;
  assign n13888 = n196 & n12370 ;
  assign n13889 = n8609 & ~n13776 ;
  assign n13890 = n13889 ^ x51 ^ 1'b0 ;
  assign n13891 = n13474 ^ n259 ^ 1'b0 ;
  assign n13893 = x45 & ~n5875 ;
  assign n13894 = n13893 ^ n3343 ^ 1'b0 ;
  assign n13895 = ( n595 & n4468 ) | ( n595 & ~n13894 ) | ( n4468 & ~n13894 ) ;
  assign n13892 = n7173 & ~n9450 ;
  assign n13896 = n13895 ^ n13892 ^ n3181 ;
  assign n13897 = n1931 ^ n1720 ^ 1'b0 ;
  assign n13898 = ( n1658 & ~n3084 ) | ( n1658 & n10581 ) | ( ~n3084 & n10581 ) ;
  assign n13899 = n4836 ^ n1106 ^ 1'b0 ;
  assign n13900 = n1275 | n13899 ;
  assign n13901 = n884 | n3365 ;
  assign n13902 = n13901 ^ n1899 ^ 1'b0 ;
  assign n13903 = n3858 & ~n13902 ;
  assign n13904 = n3669 | n13903 ;
  assign n13905 = ( ~n4237 & n8776 ) | ( ~n4237 & n10125 ) | ( n8776 & n10125 ) ;
  assign n13906 = ~n1016 & n6118 ;
  assign n13907 = n13906 ^ n11077 ^ 1'b0 ;
  assign n13908 = n1562 ^ n1208 ^ n1041 ;
  assign n13909 = n13908 ^ n5879 ^ 1'b0 ;
  assign n13910 = n11595 & n13909 ;
  assign n13911 = n6787 | n9263 ;
  assign n13912 = n9927 & ~n13911 ;
  assign n13913 = n4502 ^ n176 ^ 1'b0 ;
  assign n13914 = n3419 | n13913 ;
  assign n13915 = n13914 ^ n3244 ^ n1462 ;
  assign n13916 = n13915 ^ n8790 ^ n337 ;
  assign n13917 = ~n13912 & n13916 ;
  assign n13919 = x107 & n6701 ;
  assign n13920 = ~n6936 & n13919 ;
  assign n13918 = n3703 ^ n2083 ^ 1'b0 ;
  assign n13921 = n13920 ^ n13918 ^ 1'b0 ;
  assign n13922 = n13801 ^ n5584 ^ 1'b0 ;
  assign n13923 = n8279 | n13922 ;
  assign n13924 = ( n997 & n13921 ) | ( n997 & ~n13923 ) | ( n13921 & ~n13923 ) ;
  assign n13925 = ~n2440 & n4255 ;
  assign n13926 = n13925 ^ n1440 ^ 1'b0 ;
  assign n13927 = n13926 ^ n3568 ^ 1'b0 ;
  assign n13928 = n615 | n13927 ;
  assign n13929 = n5539 & ~n6915 ;
  assign n13930 = ( ~n4545 & n13928 ) | ( ~n4545 & n13929 ) | ( n13928 & n13929 ) ;
  assign n13931 = n13930 ^ n1428 ^ 1'b0 ;
  assign n13932 = n6202 | n9409 ;
  assign n13933 = n13931 & ~n13932 ;
  assign n13934 = n10837 ^ n10019 ^ 1'b0 ;
  assign n13935 = n4670 & n9020 ;
  assign n13936 = n2432 ^ n1939 ^ 1'b0 ;
  assign n13937 = n3189 & n13936 ;
  assign n13938 = n13937 ^ n1077 ^ 1'b0 ;
  assign n13939 = n10293 & ~n13938 ;
  assign n13940 = n2498 & n12983 ;
  assign n13941 = n9635 ^ n5308 ^ 1'b0 ;
  assign n13942 = ~n13940 & n13941 ;
  assign n13943 = n4289 ^ n3664 ^ 1'b0 ;
  assign n13944 = n13943 ^ n3594 ^ 1'b0 ;
  assign n13945 = n13942 & n13944 ;
  assign n13946 = n1184 & n2170 ;
  assign n13947 = ~n5107 & n13946 ;
  assign n13948 = n6240 ^ n4108 ^ n929 ;
  assign n13949 = n744 ^ n730 ^ 1'b0 ;
  assign n13950 = n1042 & ~n13949 ;
  assign n13951 = n13950 ^ n11043 ^ n4886 ;
  assign n13952 = ( n4293 & n13948 ) | ( n4293 & ~n13951 ) | ( n13948 & ~n13951 ) ;
  assign n13953 = ( n6333 & n13947 ) | ( n6333 & n13952 ) | ( n13947 & n13952 ) ;
  assign n13954 = n1788 & ~n2837 ;
  assign n13955 = n13954 ^ n4902 ^ 1'b0 ;
  assign n13956 = n7662 | n13955 ;
  assign n13957 = n361 & ~n13956 ;
  assign n13958 = n5199 ^ n1362 ^ 1'b0 ;
  assign n13959 = n2654 & ~n2814 ;
  assign n13960 = ( ~n3964 & n13958 ) | ( ~n3964 & n13959 ) | ( n13958 & n13959 ) ;
  assign n13961 = n10741 | n10981 ;
  assign n13962 = n13960 & ~n13961 ;
  assign n13963 = n7705 ^ n6023 ^ 1'b0 ;
  assign n13964 = n4432 & n10834 ;
  assign n13965 = n13964 ^ n3886 ^ 1'b0 ;
  assign n13966 = n8534 | n10204 ;
  assign n13967 = n13966 ^ n11399 ^ 1'b0 ;
  assign n13968 = n12496 ^ n6950 ^ 1'b0 ;
  assign n13969 = n1884 & ~n13968 ;
  assign n13970 = n11376 ^ n11122 ^ n4088 ;
  assign n13971 = n13969 & n13970 ;
  assign n13972 = n1858 | n11118 ;
  assign n13974 = n7887 & n8390 ;
  assign n13975 = ~n13807 & n13974 ;
  assign n13976 = ~n6671 & n13975 ;
  assign n13973 = n7455 ^ n5504 ^ n1666 ;
  assign n13977 = n13976 ^ n13973 ^ n10785 ;
  assign n13978 = n2703 & n3242 ;
  assign n13979 = n13978 ^ n1669 ^ 1'b0 ;
  assign n13980 = n5482 | n13979 ;
  assign n13981 = n13980 ^ n7473 ^ 1'b0 ;
  assign n13982 = ~n1196 & n13981 ;
  assign n13983 = n13982 ^ n11162 ^ 1'b0 ;
  assign n13984 = n5486 | n13983 ;
  assign n13985 = n3386 | n9528 ;
  assign n13986 = n10668 & ~n12535 ;
  assign n13987 = n6905 & n10318 ;
  assign n13988 = n1127 | n2770 ;
  assign n13989 = n13987 & ~n13988 ;
  assign n13990 = n3623 & ~n13989 ;
  assign n13995 = n6629 & ~n10106 ;
  assign n13994 = n11739 ^ n10576 ^ 1'b0 ;
  assign n13991 = n6616 ^ n5240 ^ 1'b0 ;
  assign n13992 = n7658 | n13991 ;
  assign n13993 = n1212 & n13992 ;
  assign n13996 = n13995 ^ n13994 ^ n13993 ;
  assign n13997 = ~n1923 & n13996 ;
  assign n13998 = ( n2958 & n4620 ) | ( n2958 & n13997 ) | ( n4620 & n13997 ) ;
  assign n13999 = n13216 ^ n6442 ^ 1'b0 ;
  assign n14000 = n3453 & ~n13999 ;
  assign n14001 = n7906 ^ n1860 ^ 1'b0 ;
  assign n14002 = ~n2011 & n14001 ;
  assign n14003 = ~n1458 & n14002 ;
  assign n14004 = n9314 & ~n14003 ;
  assign n14005 = ~n2276 & n6237 ;
  assign n14006 = n3155 & n14005 ;
  assign n14007 = n10486 & n11096 ;
  assign n14008 = ~n2528 & n14007 ;
  assign n14009 = ( n10778 & n14006 ) | ( n10778 & n14008 ) | ( n14006 & n14008 ) ;
  assign n14010 = n9915 & ~n11394 ;
  assign n14011 = ~n13019 & n14010 ;
  assign n14012 = n6281 | n11597 ;
  assign n14013 = n3718 & ~n14012 ;
  assign n14014 = n4759 ^ n3625 ^ 1'b0 ;
  assign n14015 = ~n1690 & n8545 ;
  assign n14016 = ( n946 & n3135 ) | ( n946 & ~n14015 ) | ( n3135 & ~n14015 ) ;
  assign n14017 = ~n14014 & n14016 ;
  assign n14018 = n14017 ^ n11930 ^ 1'b0 ;
  assign n14019 = n2393 & ~n4903 ;
  assign n14020 = n14019 ^ n4757 ^ 1'b0 ;
  assign n14021 = n14020 ^ n243 ^ 1'b0 ;
  assign n14022 = ~n3580 & n5409 ;
  assign n14023 = ~n6993 & n10060 ;
  assign n14024 = n14023 ^ n2748 ^ 1'b0 ;
  assign n14025 = ( x64 & n7370 ) | ( x64 & ~n11287 ) | ( n7370 & ~n11287 ) ;
  assign n14026 = n14025 ^ n13872 ^ n10487 ;
  assign n14027 = ~n621 & n1794 ;
  assign n14028 = n3940 & ~n4520 ;
  assign n14029 = ~n2694 & n14028 ;
  assign n14030 = ( n895 & ~n3476 ) | ( n895 & n7649 ) | ( ~n3476 & n7649 ) ;
  assign n14031 = n895 | n1366 ;
  assign n14032 = n14031 ^ n429 ^ 1'b0 ;
  assign n14033 = n14032 ^ n3756 ^ 1'b0 ;
  assign n14034 = n7113 & ~n14033 ;
  assign n14035 = n6407 ^ n5526 ^ 1'b0 ;
  assign n14036 = n10658 | n14035 ;
  assign n14037 = n1887 & n12402 ;
  assign n14039 = n1157 | n11787 ;
  assign n14040 = n3791 & ~n14039 ;
  assign n14038 = ~n3476 & n11997 ;
  assign n14041 = n14040 ^ n14038 ^ 1'b0 ;
  assign n14042 = n6109 ^ n2928 ^ 1'b0 ;
  assign n14043 = n10799 ^ n4833 ^ 1'b0 ;
  assign n14044 = n3166 & ~n4247 ;
  assign n14045 = n6430 ^ n5203 ^ 1'b0 ;
  assign n14046 = ~n6058 & n14045 ;
  assign n14047 = n338 & n14046 ;
  assign n14048 = ~x83 & n9395 ;
  assign n14049 = n6408 | n14048 ;
  assign n14050 = n914 | n14049 ;
  assign n14051 = n4957 ^ n1139 ^ 1'b0 ;
  assign n14052 = ~n12157 & n14051 ;
  assign n14053 = n14052 ^ n8190 ^ 1'b0 ;
  assign n14054 = n2384 & n4307 ;
  assign n14055 = n14054 ^ n11865 ^ 1'b0 ;
  assign n14056 = ~n12127 & n14055 ;
  assign n14057 = n3298 & n14056 ;
  assign n14058 = n14053 & n14057 ;
  assign n14059 = ( ~n6157 & n6909 ) | ( ~n6157 & n9889 ) | ( n6909 & n9889 ) ;
  assign n14060 = n14059 ^ n4133 ^ 1'b0 ;
  assign n14061 = n14060 ^ n833 ^ 1'b0 ;
  assign n14062 = ~n1203 & n14061 ;
  assign n14063 = n877 | n4466 ;
  assign n14064 = n14063 ^ n6870 ^ 1'b0 ;
  assign n14065 = n14062 & ~n14064 ;
  assign n14066 = n14058 & n14065 ;
  assign n14067 = ~n2223 & n10412 ;
  assign n14068 = n6206 ^ n1048 ^ 1'b0 ;
  assign n14069 = n6482 ^ n1684 ^ 1'b0 ;
  assign n14070 = n13749 & ~n14069 ;
  assign n14071 = ~n12287 & n14070 ;
  assign n14072 = n5620 & n9005 ;
  assign n14073 = n14072 ^ n12484 ^ 1'b0 ;
  assign n14074 = n10594 ^ n5339 ^ 1'b0 ;
  assign n14075 = n4904 & ~n14074 ;
  assign n14076 = n14075 ^ n2048 ^ 1'b0 ;
  assign n14077 = n14073 & n14076 ;
  assign n14078 = ( n612 & n14071 ) | ( n612 & n14077 ) | ( n14071 & n14077 ) ;
  assign n14079 = x120 & ~n12854 ;
  assign n14080 = n858 ^ n502 ^ 1'b0 ;
  assign n14081 = ~n838 & n14080 ;
  assign n14082 = n1775 & n12653 ;
  assign n14083 = ~n14081 & n14082 ;
  assign n14084 = n9046 & ~n14083 ;
  assign n14085 = n5326 ^ n4720 ^ 1'b0 ;
  assign n14086 = n4255 & ~n14085 ;
  assign n14087 = n14086 ^ n700 ^ 1'b0 ;
  assign n14088 = n8178 ^ n1761 ^ 1'b0 ;
  assign n14089 = ( n3763 & ~n9326 ) | ( n3763 & n14088 ) | ( ~n9326 & n14088 ) ;
  assign n14090 = n608 & n14089 ;
  assign n14091 = n14090 ^ n7691 ^ 1'b0 ;
  assign n14092 = n1603 | n1629 ;
  assign n14093 = n14092 ^ n3006 ^ 1'b0 ;
  assign n14094 = n7171 ^ n2176 ^ 1'b0 ;
  assign n14095 = ~n13223 & n14094 ;
  assign n14096 = n4292 | n7881 ;
  assign n14097 = n1205 & ~n8308 ;
  assign n14098 = n6707 & n14097 ;
  assign n14099 = n14098 ^ n8768 ^ 1'b0 ;
  assign n14100 = ~n14096 & n14099 ;
  assign n14101 = n3374 ^ n1837 ^ n711 ;
  assign n14105 = n9956 ^ n406 ^ 1'b0 ;
  assign n14102 = n4822 ^ n2705 ^ 1'b0 ;
  assign n14103 = n6171 | n14102 ;
  assign n14104 = n1017 & n14103 ;
  assign n14106 = n14105 ^ n14104 ^ 1'b0 ;
  assign n14107 = ( n9687 & ~n9733 ) | ( n9687 & n10379 ) | ( ~n9733 & n10379 ) ;
  assign n14108 = n14106 & ~n14107 ;
  assign n14109 = n13803 ^ n9315 ^ 1'b0 ;
  assign n14110 = n14108 & ~n14109 ;
  assign n14111 = ~n10108 & n11339 ;
  assign n14112 = n6135 | n13927 ;
  assign n14113 = n12451 ^ n3249 ^ 1'b0 ;
  assign n14114 = n11910 ^ n4555 ^ 1'b0 ;
  assign n14115 = n6131 & ~n11911 ;
  assign n14116 = n8911 ^ n3583 ^ 1'b0 ;
  assign n14117 = n3767 ^ n2408 ^ n1085 ;
  assign n14118 = ~n2330 & n14117 ;
  assign n14119 = n14116 & n14118 ;
  assign n14120 = ~n2280 & n14119 ;
  assign n14121 = ( n2637 & ~n8499 ) | ( n2637 & n12809 ) | ( ~n8499 & n12809 ) ;
  assign n14122 = n11826 ^ n1162 ^ 1'b0 ;
  assign n14123 = n454 & n14122 ;
  assign n14124 = n2570 | n7298 ;
  assign n14125 = ( n5218 & n12139 ) | ( n5218 & n14124 ) | ( n12139 & n14124 ) ;
  assign n14126 = ~n466 & n2503 ;
  assign n14127 = n14126 ^ n6455 ^ n2359 ;
  assign n14128 = n11492 ^ n1631 ^ 1'b0 ;
  assign n14129 = n12486 | n14128 ;
  assign n14130 = n14129 ^ n7114 ^ 1'b0 ;
  assign n14131 = n7670 & ~n14130 ;
  assign n14132 = n3310 & ~n13483 ;
  assign n14133 = n7592 | n14132 ;
  assign n14134 = n13796 & ~n14133 ;
  assign n14135 = n14134 ^ n4560 ^ 1'b0 ;
  assign n14136 = n842 & ~n14135 ;
  assign n14137 = n6148 ^ n6051 ^ n2038 ;
  assign n14138 = n3554 & n9438 ;
  assign n14139 = n4090 & ~n4745 ;
  assign n14140 = n8677 & n14139 ;
  assign n14141 = n13853 ^ n5413 ^ 1'b0 ;
  assign n14147 = n2692 ^ n1081 ^ 1'b0 ;
  assign n14148 = ~n2846 & n14147 ;
  assign n14142 = ~n5437 & n10879 ;
  assign n14143 = ~n150 & n14142 ;
  assign n14144 = n7526 | n14143 ;
  assign n14145 = n14144 ^ n8605 ^ 1'b0 ;
  assign n14146 = ~n9702 & n14145 ;
  assign n14149 = n14148 ^ n14146 ^ n708 ;
  assign n14150 = ~n7924 & n12865 ;
  assign n14154 = ( n179 & n1758 ) | ( n179 & n3008 ) | ( n1758 & n3008 ) ;
  assign n14151 = n10066 ^ n3181 ^ 1'b0 ;
  assign n14152 = ( n6812 & n8121 ) | ( n6812 & ~n10710 ) | ( n8121 & ~n10710 ) ;
  assign n14153 = n14151 | n14152 ;
  assign n14155 = n14154 ^ n14153 ^ 1'b0 ;
  assign n14156 = n13287 | n14155 ;
  assign n14158 = n398 & n1025 ;
  assign n14157 = ~n7850 & n11101 ;
  assign n14159 = n14158 ^ n14157 ^ 1'b0 ;
  assign n14160 = n8107 & n11058 ;
  assign n14161 = n3468 & n14160 ;
  assign n14162 = n3411 & n14161 ;
  assign n14163 = ( ~n1459 & n1861 ) | ( ~n1459 & n12408 ) | ( n1861 & n12408 ) ;
  assign n14164 = ~n12802 & n14163 ;
  assign n14165 = n14164 ^ n9093 ^ 1'b0 ;
  assign n14166 = n3634 | n9591 ;
  assign n14167 = ~n3259 & n14166 ;
  assign n14168 = ( n199 & n2640 ) | ( n199 & ~n13970 ) | ( n2640 & ~n13970 ) ;
  assign n14169 = n9464 ^ n8140 ^ 1'b0 ;
  assign n14170 = n14168 | n14169 ;
  assign n14171 = n14170 ^ n1848 ^ 1'b0 ;
  assign n14172 = n6456 & n7620 ;
  assign n14173 = ~n13803 & n14172 ;
  assign n14174 = n4466 | n5050 ;
  assign n14175 = ~n785 & n4115 ;
  assign n14176 = ~n8680 & n14175 ;
  assign n14177 = n11567 ^ n8681 ^ 1'b0 ;
  assign n14178 = n9011 & ~n14177 ;
  assign n14179 = n14178 ^ n9176 ^ 1'b0 ;
  assign n14180 = n14179 ^ n7851 ^ 1'b0 ;
  assign n14181 = ~n5822 & n11288 ;
  assign n14182 = ( n153 & n9963 ) | ( n153 & ~n14181 ) | ( n9963 & ~n14181 ) ;
  assign n14183 = n4715 | n7649 ;
  assign n14184 = n14182 | n14183 ;
  assign n14185 = ~n1123 & n6840 ;
  assign n14186 = n14069 ^ n510 ^ 1'b0 ;
  assign n14187 = n1637 & n2599 ;
  assign n14188 = n4678 & n14187 ;
  assign n14189 = n14186 & ~n14188 ;
  assign n14190 = n14185 | n14189 ;
  assign n14191 = n14190 ^ n4266 ^ 1'b0 ;
  assign n14192 = n2329 & n8505 ;
  assign n14193 = n14143 & n14192 ;
  assign n14194 = n4451 ^ n3343 ^ 1'b0 ;
  assign n14195 = n8885 ^ n5459 ^ 1'b0 ;
  assign n14196 = n5567 & ~n6951 ;
  assign n14197 = ~n3319 & n14196 ;
  assign n14198 = ~n3995 & n8395 ;
  assign n14199 = n398 & n14198 ;
  assign n14200 = n14199 ^ n6048 ^ n823 ;
  assign n14201 = n8965 ^ n7481 ^ n7064 ;
  assign n14202 = ~n14200 & n14201 ;
  assign n14203 = n9795 | n11653 ;
  assign n14204 = n4929 & n14203 ;
  assign n14205 = n5662 & n14204 ;
  assign n14207 = ( ~n2389 & n6287 ) | ( ~n2389 & n6678 ) | ( n6287 & n6678 ) ;
  assign n14206 = n2788 | n12906 ;
  assign n14208 = n14207 ^ n14206 ^ 1'b0 ;
  assign n14209 = n4394 ^ n661 ^ 1'b0 ;
  assign n14210 = n7514 & n14209 ;
  assign n14211 = ( n373 & n8730 ) | ( n373 & ~n9950 ) | ( n8730 & ~n9950 ) ;
  assign n14212 = n1794 ^ n1364 ^ 1'b0 ;
  assign n14213 = n14212 ^ n7627 ^ 1'b0 ;
  assign n14214 = n4409 ^ n1601 ^ 1'b0 ;
  assign n14215 = n308 & ~n6726 ;
  assign n14216 = n4516 & n8132 ;
  assign n14217 = ~n6079 & n14216 ;
  assign n14218 = n14217 ^ n2670 ^ 1'b0 ;
  assign n14219 = n12142 ^ n11084 ^ 1'b0 ;
  assign n14220 = n8081 ^ n8021 ^ n5154 ;
  assign n14221 = n3624 & ~n5908 ;
  assign n14222 = ~n2985 & n5733 ;
  assign n14223 = n13474 | n14222 ;
  assign n14224 = n14221 & ~n14223 ;
  assign n14225 = n5404 | n8498 ;
  assign n14226 = n14225 ^ n3922 ^ 1'b0 ;
  assign n14227 = n14226 ^ n5483 ^ 1'b0 ;
  assign n14228 = ~n1449 & n5089 ;
  assign n14229 = n8945 ^ n5139 ^ 1'b0 ;
  assign n14230 = x45 & ~n14229 ;
  assign n14231 = n5862 ^ n1044 ^ 1'b0 ;
  assign n14232 = n1021 & ~n10776 ;
  assign n14233 = n14232 ^ n7461 ^ 1'b0 ;
  assign n14234 = n510 & ~n1002 ;
  assign n14235 = ~n6791 & n14234 ;
  assign n14236 = n10472 & n14235 ;
  assign n14237 = ~n4573 & n4622 ;
  assign n14238 = n14237 ^ n1207 ^ 1'b0 ;
  assign n14239 = n14238 ^ n4771 ^ 1'b0 ;
  assign n14240 = ~n6337 & n14239 ;
  assign n14241 = n1362 | n14240 ;
  assign n14242 = n12430 ^ n10609 ^ n4819 ;
  assign n14243 = n14241 | n14242 ;
  assign n14244 = n12386 ^ n7142 ^ x125 ;
  assign n14245 = n2022 | n3291 ;
  assign n14246 = n14245 ^ n1239 ^ 1'b0 ;
  assign n14247 = ( n2642 & ~n4357 ) | ( n2642 & n14246 ) | ( ~n4357 & n14246 ) ;
  assign n14248 = n12116 ^ x110 ^ 1'b0 ;
  assign n14249 = n4217 | n14248 ;
  assign n14250 = n14247 & ~n14249 ;
  assign n14251 = n14250 ^ n8085 ^ n4217 ;
  assign n14252 = ~n7723 & n9787 ;
  assign n14253 = n873 ^ x59 ^ 1'b0 ;
  assign n14254 = ~n8867 & n14253 ;
  assign n14255 = ~n14252 & n14254 ;
  assign n14257 = n654 | n7909 ;
  assign n14256 = n6001 & ~n8491 ;
  assign n14258 = n14257 ^ n14256 ^ 1'b0 ;
  assign n14259 = x80 & ~n11122 ;
  assign n14260 = ~n4490 & n14259 ;
  assign n14261 = n9777 ^ n3838 ^ 1'b0 ;
  assign n14267 = n3999 & ~n9921 ;
  assign n14268 = n12650 | n14267 ;
  assign n14269 = n975 & ~n14268 ;
  assign n14262 = n342 | n1193 ;
  assign n14263 = n1833 & ~n14262 ;
  assign n14264 = n920 ^ x84 ^ 1'b0 ;
  assign n14265 = ~n1150 & n14264 ;
  assign n14266 = ~n14263 & n14265 ;
  assign n14270 = n14269 ^ n14266 ^ 1'b0 ;
  assign n14271 = n13598 ^ n11059 ^ 1'b0 ;
  assign n14273 = n11330 ^ n4371 ^ 1'b0 ;
  assign n14274 = ~n3625 & n14273 ;
  assign n14272 = n8873 | n12388 ;
  assign n14275 = n14274 ^ n14272 ^ 1'b0 ;
  assign n14276 = n4340 ^ n240 ^ 1'b0 ;
  assign n14277 = n10033 & ~n14276 ;
  assign n14278 = ( ~x76 & n4902 ) | ( ~x76 & n14277 ) | ( n4902 & n14277 ) ;
  assign n14279 = n452 & n4420 ;
  assign n14280 = n14279 ^ x95 ^ 1'b0 ;
  assign n14281 = n14280 ^ n10094 ^ n1220 ;
  assign n14282 = n10031 ^ n6811 ^ 1'b0 ;
  assign n14283 = ~n7328 & n14282 ;
  assign n14284 = n8705 ^ n6506 ^ 1'b0 ;
  assign n14285 = ~n5585 & n14284 ;
  assign n14286 = n1181 | n14285 ;
  assign n14287 = n4428 ^ n828 ^ n515 ;
  assign n14288 = ~n4204 & n14287 ;
  assign n14289 = n14288 ^ n10963 ^ 1'b0 ;
  assign n14290 = n1724 | n14289 ;
  assign n14291 = n11210 ^ n10267 ^ n4288 ;
  assign n14293 = ~n3386 & n4001 ;
  assign n14294 = n14293 ^ n8341 ^ 1'b0 ;
  assign n14292 = n2032 ^ n563 ^ 1'b0 ;
  assign n14295 = n14294 ^ n14292 ^ 1'b0 ;
  assign n14296 = n8397 & ~n14295 ;
  assign n14297 = n9777 ^ n8999 ^ 1'b0 ;
  assign n14298 = ~n11084 & n14297 ;
  assign n14299 = n9322 ^ n9198 ^ n1777 ;
  assign n14300 = n6073 ^ n1326 ^ 1'b0 ;
  assign n14301 = n4528 & ~n9145 ;
  assign n14302 = n14301 ^ n639 ^ 1'b0 ;
  assign n14305 = ~n3448 & n3922 ;
  assign n14303 = n1169 | n1739 ;
  assign n14304 = n14303 ^ n9463 ^ n2682 ;
  assign n14306 = n14305 ^ n14304 ^ 1'b0 ;
  assign n14307 = ( n1364 & n1702 ) | ( n1364 & ~n5538 ) | ( n1702 & ~n5538 ) ;
  assign n14308 = n311 & ~n14307 ;
  assign n14309 = ( n5565 & ~n6338 ) | ( n5565 & n14308 ) | ( ~n6338 & n14308 ) ;
  assign n14310 = n4683 ^ n4123 ^ 1'b0 ;
  assign n14311 = ~n6241 & n14310 ;
  assign n14312 = n5551 & n14311 ;
  assign n14313 = ( n1465 & n14309 ) | ( n1465 & ~n14312 ) | ( n14309 & ~n14312 ) ;
  assign n14314 = n2547 ^ n420 ^ 1'b0 ;
  assign n14315 = ~n5369 & n14314 ;
  assign n14316 = n14315 ^ n4131 ^ 1'b0 ;
  assign n14317 = n4270 & n14316 ;
  assign n14318 = ( n1168 & n6826 ) | ( n1168 & ~n14317 ) | ( n6826 & ~n14317 ) ;
  assign n14319 = n13709 ^ n6002 ^ x8 ;
  assign n14320 = n6394 & ~n10796 ;
  assign n14321 = n3618 ^ n2880 ^ 1'b0 ;
  assign n14322 = n6914 & n14321 ;
  assign n14323 = n14322 ^ n5002 ^ 1'b0 ;
  assign n14324 = n4846 & ~n14323 ;
  assign n14325 = n14324 ^ n654 ^ 1'b0 ;
  assign n14326 = n13492 ^ n10006 ^ 1'b0 ;
  assign n14327 = n14326 ^ n10136 ^ n5119 ;
  assign n14328 = n10395 ^ n6071 ^ 1'b0 ;
  assign n14329 = n8337 & n14328 ;
  assign n14330 = n14329 ^ n2334 ^ 1'b0 ;
  assign n14331 = n12977 ^ n1805 ^ 1'b0 ;
  assign n14332 = n14331 ^ n5771 ^ 1'b0 ;
  assign n14333 = n14332 ^ n330 ^ 1'b0 ;
  assign n14334 = x22 & ~n14333 ;
  assign n14335 = n8974 & n14334 ;
  assign n14336 = ~n1371 & n14335 ;
  assign n14337 = n1420 ^ x57 ^ 1'b0 ;
  assign n14338 = n2234 & ~n14337 ;
  assign n14339 = ~n3882 & n14338 ;
  assign n14340 = n7632 & n14339 ;
  assign n14341 = n6792 | n14340 ;
  assign n14342 = n14341 ^ n4498 ^ 1'b0 ;
  assign n14343 = n10048 & n14342 ;
  assign n14344 = n4391 & ~n8029 ;
  assign n14345 = n14343 & n14344 ;
  assign n14346 = n3914 & ~n13544 ;
  assign n14350 = n10008 ^ n9647 ^ 1'b0 ;
  assign n14348 = n10856 ^ n3191 ^ 1'b0 ;
  assign n14349 = n7981 & n14348 ;
  assign n14347 = n3516 ^ n3167 ^ 1'b0 ;
  assign n14351 = n14350 ^ n14349 ^ n14347 ;
  assign n14352 = n2541 | n7355 ;
  assign n14353 = n1479 ^ n1443 ^ 1'b0 ;
  assign n14354 = ~n3999 & n14353 ;
  assign n14355 = n14354 ^ n2786 ^ 1'b0 ;
  assign n14356 = n14355 ^ n8106 ^ 1'b0 ;
  assign n14357 = ( n2091 & n14352 ) | ( n2091 & ~n14356 ) | ( n14352 & ~n14356 ) ;
  assign n14358 = n1248 | n1418 ;
  assign n14359 = n14358 ^ n4489 ^ 1'b0 ;
  assign n14360 = n14359 ^ n3494 ^ x83 ;
  assign n14361 = ~n508 & n8942 ;
  assign n14362 = n10109 ^ n2705 ^ 1'b0 ;
  assign n14363 = n5783 ^ n2005 ^ 1'b0 ;
  assign n14364 = ~n283 & n14363 ;
  assign n14365 = n2572 | n5107 ;
  assign n14366 = n14365 ^ n10277 ^ n6070 ;
  assign n14367 = n13439 ^ n8745 ^ 1'b0 ;
  assign n14368 = n4097 ^ x56 ^ 1'b0 ;
  assign n14369 = n11075 & ~n14368 ;
  assign n14370 = n11589 ^ n7226 ^ 1'b0 ;
  assign n14371 = n7934 ^ n3856 ^ 1'b0 ;
  assign n14372 = n14371 ^ n8759 ^ n6584 ;
  assign n14373 = n4120 ^ x81 ^ 1'b0 ;
  assign n14374 = n14373 ^ n5255 ^ 1'b0 ;
  assign n14375 = n12721 ^ n9708 ^ n4612 ;
  assign n14376 = n14375 ^ n4479 ^ 1'b0 ;
  assign n14377 = n14374 & n14376 ;
  assign n14378 = ~n8981 & n14377 ;
  assign n14379 = n14372 & n14378 ;
  assign n14381 = ~n1860 & n13034 ;
  assign n14382 = ~n1254 & n14381 ;
  assign n14380 = n3265 ^ n527 ^ 1'b0 ;
  assign n14383 = n14382 ^ n14380 ^ n12037 ;
  assign n14384 = n1938 & n5824 ;
  assign n14385 = n4690 & n14384 ;
  assign n14386 = n7046 ^ n5973 ^ 1'b0 ;
  assign n14387 = n817 & n14386 ;
  assign n14388 = n14387 ^ n4573 ^ 1'b0 ;
  assign n14389 = n14385 | n14388 ;
  assign n14390 = n4605 & n6030 ;
  assign n14391 = n14390 ^ n3126 ^ x104 ;
  assign n14392 = n1116 | n14391 ;
  assign n14395 = ~n3119 & n3192 ;
  assign n14396 = n206 & n14395 ;
  assign n14397 = n8259 & ~n14396 ;
  assign n14398 = ~n2409 & n14397 ;
  assign n14393 = n7258 | n13526 ;
  assign n14394 = n14393 ^ n3369 ^ 1'b0 ;
  assign n14399 = n14398 ^ n14394 ^ n9659 ;
  assign n14400 = n2789 ^ x49 ^ 1'b0 ;
  assign n14401 = n1185 & ~n14400 ;
  assign n14402 = n14401 ^ n1407 ^ 1'b0 ;
  assign n14403 = n1251 & n2030 ;
  assign n14404 = n10257 & n14403 ;
  assign n14405 = n2507 ^ n1371 ^ n872 ;
  assign n14406 = ( ~n314 & n4730 ) | ( ~n314 & n14405 ) | ( n4730 & n14405 ) ;
  assign n14407 = n14406 ^ n4498 ^ 1'b0 ;
  assign n14408 = n14407 ^ n2964 ^ 1'b0 ;
  assign n14409 = n14404 | n14408 ;
  assign n14410 = ( n642 & n939 ) | ( n642 & n4915 ) | ( n939 & n4915 ) ;
  assign n14411 = n2639 | n14410 ;
  assign n14412 = n1684 | n14411 ;
  assign n14413 = ~n2190 & n14412 ;
  assign n14414 = ~n7103 & n14413 ;
  assign n14415 = n8006 ^ n6534 ^ 1'b0 ;
  assign n14416 = ( ~n555 & n10170 ) | ( ~n555 & n14415 ) | ( n10170 & n14415 ) ;
  assign n14418 = ~n3528 & n12408 ;
  assign n14417 = n1734 & ~n9733 ;
  assign n14419 = n14418 ^ n14417 ^ n11185 ;
  assign n14420 = n13708 & n14419 ;
  assign n14421 = n11683 ^ n6729 ^ 1'b0 ;
  assign n14422 = n5282 ^ n1465 ^ n1423 ;
  assign n14423 = n14422 ^ n13529 ^ n6308 ;
  assign n14424 = n2057 & n11919 ;
  assign n14425 = n6046 ^ n142 ^ 1'b0 ;
  assign n14426 = ~n7408 & n14425 ;
  assign n14427 = ( ~n764 & n7332 ) | ( ~n764 & n14426 ) | ( n7332 & n14426 ) ;
  assign n14428 = ~n1189 & n11683 ;
  assign n14429 = n14428 ^ n10616 ^ 1'b0 ;
  assign n14430 = n8086 ^ n2846 ^ 1'b0 ;
  assign n14431 = n2411 & ~n14430 ;
  assign n14432 = n6198 & ~n14431 ;
  assign n14434 = n1236 & n5185 ;
  assign n14433 = n8441 & n11698 ;
  assign n14435 = n14434 ^ n14433 ^ 1'b0 ;
  assign n14439 = ( n1578 & n1600 ) | ( n1578 & n3743 ) | ( n1600 & n3743 ) ;
  assign n14440 = ( ~n1345 & n3861 ) | ( ~n1345 & n14439 ) | ( n3861 & n14439 ) ;
  assign n14436 = n1869 ^ n830 ^ 1'b0 ;
  assign n14437 = n3479 & ~n14436 ;
  assign n14438 = ( n2705 & n12405 ) | ( n2705 & n14437 ) | ( n12405 & n14437 ) ;
  assign n14441 = n14440 ^ n14438 ^ n3480 ;
  assign n14442 = n14441 ^ n6661 ^ n1853 ;
  assign n14443 = ~n2389 & n5946 ;
  assign n14444 = n13545 & n14443 ;
  assign n14445 = n311 | n11899 ;
  assign n14447 = ( n5897 & ~n6868 ) | ( n5897 & n7075 ) | ( ~n6868 & n7075 ) ;
  assign n14446 = ( n1118 & n4121 ) | ( n1118 & n14160 ) | ( n4121 & n14160 ) ;
  assign n14448 = n14447 ^ n14446 ^ n2605 ;
  assign n14449 = n14448 ^ n254 ^ 1'b0 ;
  assign n14450 = x65 & ~n6770 ;
  assign n14451 = n14450 ^ n3475 ^ 1'b0 ;
  assign n14452 = ( n7353 & n7827 ) | ( n7353 & n14451 ) | ( n7827 & n14451 ) ;
  assign n14453 = n9069 ^ n3342 ^ 1'b0 ;
  assign n14454 = n4261 ^ n1171 ^ 1'b0 ;
  assign n14455 = ~n14453 & n14454 ;
  assign n14456 = n5123 | n9072 ;
  assign n14457 = ~n7679 & n8594 ;
  assign n14458 = ~n14456 & n14457 ;
  assign n14459 = n14455 & ~n14458 ;
  assign n14460 = n8769 ^ n8095 ^ x22 ;
  assign n14461 = n13142 ^ n610 ^ 1'b0 ;
  assign n14462 = n4025 & n14461 ;
  assign n14463 = n6441 | n14058 ;
  assign n14464 = n14462 | n14463 ;
  assign n14465 = n3521 ^ x31 ^ 1'b0 ;
  assign n14466 = ~n13501 & n14465 ;
  assign n14467 = n5623 | n6337 ;
  assign n14468 = ( n779 & n4281 ) | ( n779 & n14188 ) | ( n4281 & n14188 ) ;
  assign n14469 = ~n5227 & n6798 ;
  assign n14470 = ~n3116 & n3590 ;
  assign n14471 = n2997 | n9104 ;
  assign n14472 = n2997 & ~n14471 ;
  assign n14473 = n248 & ~n8185 ;
  assign n14474 = n8185 & n14473 ;
  assign n14475 = x37 & ~n790 ;
  assign n14476 = ~x37 & n14475 ;
  assign n14477 = n2091 & n4399 ;
  assign n14478 = n14476 & n14477 ;
  assign n14479 = n14474 | n14478 ;
  assign n14480 = n14474 & ~n14479 ;
  assign n14481 = n14472 | n14480 ;
  assign n14482 = n14472 & ~n14481 ;
  assign n14483 = n14482 ^ n2190 ^ 1'b0 ;
  assign n14484 = n14483 ^ n4280 ^ 1'b0 ;
  assign n14485 = n14470 & n14484 ;
  assign n14486 = n3842 ^ n1387 ^ 1'b0 ;
  assign n14487 = ( n5012 & n5373 ) | ( n5012 & n8220 ) | ( n5373 & n8220 ) ;
  assign n14488 = n14487 ^ n12292 ^ 1'b0 ;
  assign n14489 = n14486 & ~n14488 ;
  assign n14490 = ~n859 & n11162 ;
  assign n14491 = n1535 & n14490 ;
  assign n14492 = n1108 ^ n984 ^ 1'b0 ;
  assign n14495 = n3476 & n7323 ;
  assign n14496 = ~n11055 & n14495 ;
  assign n14493 = n6753 | n9172 ;
  assign n14494 = n8391 | n14493 ;
  assign n14497 = n14496 ^ n14494 ^ n9216 ;
  assign n14498 = ~n5749 & n14426 ;
  assign n14499 = n14498 ^ n8419 ^ 1'b0 ;
  assign n14500 = n4875 & n5898 ;
  assign n14501 = n7131 ^ n5304 ^ 1'b0 ;
  assign n14502 = n6248 | n14501 ;
  assign n14503 = n2496 ^ n529 ^ 1'b0 ;
  assign n14504 = n4640 & n14503 ;
  assign n14505 = n496 | n14504 ;
  assign n14506 = ~n239 & n614 ;
  assign n14507 = ~n1870 & n14506 ;
  assign n14508 = n6432 | n14507 ;
  assign n14509 = n815 | n14508 ;
  assign n14510 = ( n2165 & n4725 ) | ( n2165 & n14509 ) | ( n4725 & n14509 ) ;
  assign n14511 = n12712 ^ n3153 ^ 1'b0 ;
  assign n14512 = ( n3814 & n14510 ) | ( n3814 & n14511 ) | ( n14510 & n14511 ) ;
  assign n14513 = n1929 | n3553 ;
  assign n14514 = n11800 | n14513 ;
  assign n14515 = n910 & n4064 ;
  assign n14516 = n14515 ^ n461 ^ 1'b0 ;
  assign n14517 = n9391 ^ n5632 ^ 1'b0 ;
  assign n14518 = n4369 & n14517 ;
  assign n14520 = n3767 | n5625 ;
  assign n14519 = ~n7776 & n11528 ;
  assign n14521 = n14520 ^ n14519 ^ 1'b0 ;
  assign n14522 = ( ~n4817 & n6429 ) | ( ~n4817 & n14521 ) | ( n6429 & n14521 ) ;
  assign n14523 = n5937 & n14522 ;
  assign n14524 = n5875 & n14523 ;
  assign n14525 = n11101 ^ n9525 ^ n3249 ;
  assign n14526 = n12205 & n12405 ;
  assign n14527 = n14526 ^ n5706 ^ 1'b0 ;
  assign n14528 = n398 & n14527 ;
  assign n14529 = n7582 ^ n6986 ^ n2871 ;
  assign n14530 = n14529 ^ n12717 ^ n745 ;
  assign n14531 = n12789 ^ n10841 ^ n1012 ;
  assign n14532 = n13133 ^ n3644 ^ 1'b0 ;
  assign n14533 = ~n1368 & n14532 ;
  assign n14534 = n8491 ^ n1088 ^ 1'b0 ;
  assign n14535 = n11731 | n14534 ;
  assign n14536 = n6182 | n14535 ;
  assign n14537 = n14533 | n14536 ;
  assign n14538 = n8299 & n11046 ;
  assign n14539 = n14537 | n14538 ;
  assign n14540 = n4531 & ~n8124 ;
  assign n14541 = n1666 & ~n4990 ;
  assign n14542 = n9773 & n14541 ;
  assign n14543 = n6363 ^ n3761 ^ 1'b0 ;
  assign n14544 = ~n753 & n3800 ;
  assign n14545 = n11266 ^ n10454 ^ n9086 ;
  assign n14546 = ( n1506 & n2411 ) | ( n1506 & ~n3594 ) | ( n2411 & ~n3594 ) ;
  assign n14547 = n3210 & n14546 ;
  assign n14548 = n8471 ^ n6937 ^ n1909 ;
  assign n14549 = n628 | n13197 ;
  assign n14550 = n14549 ^ n2309 ^ 1'b0 ;
  assign n14551 = n4499 ^ n4057 ^ 1'b0 ;
  assign n14552 = n14550 & n14551 ;
  assign n14553 = n221 | n3878 ;
  assign n14554 = ( n9587 & ~n14552 ) | ( n9587 & n14553 ) | ( ~n14552 & n14553 ) ;
  assign n14555 = n12305 ^ n11587 ^ n1372 ;
  assign n14556 = n3340 & ~n12347 ;
  assign n14557 = n14556 ^ n4408 ^ 1'b0 ;
  assign n14558 = n13076 & n13641 ;
  assign n14559 = ~n14557 & n14558 ;
  assign n14560 = ~n2929 & n10856 ;
  assign n14561 = n942 & n14560 ;
  assign n14562 = ( n2535 & ~n7781 ) | ( n2535 & n7818 ) | ( ~n7781 & n7818 ) ;
  assign n14563 = n14562 ^ n9018 ^ 1'b0 ;
  assign n14564 = ( n1072 & ~n3738 ) | ( n1072 & n12398 ) | ( ~n3738 & n12398 ) ;
  assign n14565 = n5274 & n6981 ;
  assign n14566 = n1939 & n4896 ;
  assign n14567 = ~n12851 & n14566 ;
  assign n14568 = n14567 ^ n13867 ^ 1'b0 ;
  assign n14569 = n10910 | n14568 ;
  assign n14570 = n9350 | n12647 ;
  assign n14571 = n386 & n2804 ;
  assign n14572 = n14571 ^ n9743 ^ 1'b0 ;
  assign n14573 = n14572 ^ n2431 ^ 1'b0 ;
  assign n14574 = n9816 & n14573 ;
  assign n14575 = ( n3035 & n3299 ) | ( n3035 & ~n4584 ) | ( n3299 & ~n4584 ) ;
  assign n14576 = ~n1079 & n14575 ;
  assign n14577 = n14455 ^ n12848 ^ n1803 ;
  assign n14578 = n12487 ^ n11326 ^ 1'b0 ;
  assign n14579 = n1504 | n14578 ;
  assign n14580 = ( n1681 & ~n4426 ) | ( n1681 & n6354 ) | ( ~n4426 & n6354 ) ;
  assign n14581 = n14580 ^ n2198 ^ 1'b0 ;
  assign n14582 = n2735 ^ n1738 ^ 1'b0 ;
  assign n14583 = n14582 ^ n2467 ^ 1'b0 ;
  assign n14584 = n3117 | n13737 ;
  assign n14585 = n14584 ^ n6190 ^ 1'b0 ;
  assign n14586 = n595 & n2737 ;
  assign n14587 = n14586 ^ n4376 ^ 1'b0 ;
  assign n14589 = ( n1610 & ~n4833 ) | ( n1610 & n14287 ) | ( ~n4833 & n14287 ) ;
  assign n14588 = n4640 ^ n3209 ^ 1'b0 ;
  assign n14590 = n14589 ^ n14588 ^ 1'b0 ;
  assign n14591 = n14587 & n14590 ;
  assign n14593 = n1669 & n1944 ;
  assign n14594 = ~n1140 & n14593 ;
  assign n14592 = x125 & n5693 ;
  assign n14595 = n14594 ^ n14592 ^ 1'b0 ;
  assign n14596 = n6083 ^ n2694 ^ 1'b0 ;
  assign n14597 = ~n3409 & n14596 ;
  assign n14598 = n8344 ^ n6428 ^ n4983 ;
  assign n14599 = n14557 ^ n9388 ^ 1'b0 ;
  assign n14600 = n3869 ^ n311 ^ 1'b0 ;
  assign n14602 = n2985 ^ n978 ^ 1'b0 ;
  assign n14603 = n755 | n14602 ;
  assign n14601 = n2198 & ~n4963 ;
  assign n14604 = n14603 ^ n14601 ^ n7583 ;
  assign n14605 = ~n14600 & n14604 ;
  assign n14606 = ~n11226 & n14605 ;
  assign n14607 = n819 & ~n5682 ;
  assign n14608 = n14607 ^ n3145 ^ 1'b0 ;
  assign n14609 = n14608 ^ n4467 ^ 1'b0 ;
  assign n14610 = ~n3896 & n14609 ;
  assign n14611 = ( n469 & n1927 ) | ( n469 & n14610 ) | ( n1927 & n14610 ) ;
  assign n14612 = n7616 | n8381 ;
  assign n14613 = n1841 & ~n14612 ;
  assign n14614 = n3625 & ~n14613 ;
  assign n14615 = ~n14611 & n14614 ;
  assign n14616 = n2760 & ~n7295 ;
  assign n14617 = ~n11298 & n14616 ;
  assign n14618 = n2380 | n5836 ;
  assign n14619 = n14618 ^ n8555 ^ 1'b0 ;
  assign n14620 = n14619 ^ n3137 ^ 1'b0 ;
  assign n14621 = n1379 & ~n6146 ;
  assign n14622 = ~n527 & n1136 ;
  assign n14623 = x30 & n9323 ;
  assign n14624 = n14623 ^ n13047 ^ 1'b0 ;
  assign n14625 = n5866 & n7564 ;
  assign n14626 = ~n14624 & n14625 ;
  assign n14627 = n1212 & n14626 ;
  assign n14628 = n12173 & ~n14627 ;
  assign n14629 = n12601 & n14628 ;
  assign n14630 = n9947 ^ n6392 ^ 1'b0 ;
  assign n14631 = n9840 & ~n14630 ;
  assign n14632 = n6963 ^ n2184 ^ 1'b0 ;
  assign n14633 = n14631 & n14632 ;
  assign n14634 = n728 | n6490 ;
  assign n14635 = n11699 ^ n8887 ^ n3845 ;
  assign n14636 = ~n1901 & n3716 ;
  assign n14641 = ~n986 & n5705 ;
  assign n14637 = n3476 ^ n2636 ^ 1'b0 ;
  assign n14638 = n670 | n1203 ;
  assign n14639 = n3102 | n14638 ;
  assign n14640 = ( n11460 & n14637 ) | ( n11460 & ~n14639 ) | ( n14637 & ~n14639 ) ;
  assign n14642 = n14641 ^ n14640 ^ n1892 ;
  assign n14643 = n14642 ^ n1893 ^ 1'b0 ;
  assign n14644 = n14636 | n14643 ;
  assign n14645 = n5156 & ~n13990 ;
  assign n14646 = n5328 & n9586 ;
  assign n14647 = n3244 & n14646 ;
  assign n14648 = ~n2535 & n13807 ;
  assign n14649 = n2668 | n14648 ;
  assign n14650 = n9481 | n14649 ;
  assign n14651 = n642 & ~n2413 ;
  assign n14652 = n2804 & n14651 ;
  assign n14653 = n14652 ^ n13584 ^ 1'b0 ;
  assign n14654 = n11105 ^ n2639 ^ 1'b0 ;
  assign n14655 = n11934 ^ n6031 ^ 1'b0 ;
  assign n14656 = n9686 ^ n6961 ^ 1'b0 ;
  assign n14657 = ~n6403 & n14656 ;
  assign n14658 = n6701 ^ n5656 ^ 1'b0 ;
  assign n14659 = n3224 & n14658 ;
  assign n14660 = n4204 & ~n14659 ;
  assign n14661 = n14660 ^ n11269 ^ 1'b0 ;
  assign n14662 = ( n4514 & n6680 ) | ( n4514 & n11043 ) | ( n6680 & n11043 ) ;
  assign n14663 = n9686 ^ n3838 ^ n2750 ;
  assign n14664 = n9942 | n14663 ;
  assign n14665 = ( ~n1931 & n6546 ) | ( ~n1931 & n10943 ) | ( n6546 & n10943 ) ;
  assign n14666 = n14665 ^ n276 ^ 1'b0 ;
  assign n14667 = n4594 & ~n13237 ;
  assign n14668 = n2643 & ~n9466 ;
  assign n14669 = n14668 ^ n8956 ^ 1'b0 ;
  assign n14670 = ( n404 & ~n7851 ) | ( n404 & n14669 ) | ( ~n7851 & n14669 ) ;
  assign n14671 = n2873 & n5410 ;
  assign n14672 = n14671 ^ n2065 ^ 1'b0 ;
  assign n14673 = x84 & n1811 ;
  assign n14674 = n14672 | n14673 ;
  assign n14675 = n7458 ^ n2583 ^ 1'b0 ;
  assign n14676 = n7916 & n14675 ;
  assign n14677 = n14674 & n14676 ;
  assign n14678 = n7386 | n9938 ;
  assign n14683 = ( ~n2441 & n4095 ) | ( ~n2441 & n5858 ) | ( n4095 & n5858 ) ;
  assign n14679 = n2192 & n4400 ;
  assign n14680 = n14679 ^ n1504 ^ 1'b0 ;
  assign n14681 = n3023 & ~n14680 ;
  assign n14682 = n6350 | n14681 ;
  assign n14684 = n14683 ^ n14682 ^ 1'b0 ;
  assign n14685 = n2668 | n7234 ;
  assign n14686 = n14685 ^ n4597 ^ 1'b0 ;
  assign n14687 = n4398 | n13778 ;
  assign n14688 = n14687 ^ n3542 ^ 1'b0 ;
  assign n14689 = n10028 ^ n2462 ^ 1'b0 ;
  assign n14690 = ( n1961 & n10305 ) | ( n1961 & ~n14149 ) | ( n10305 & ~n14149 ) ;
  assign n14691 = x21 & ~n14690 ;
  assign n14692 = n4952 & ~n10888 ;
  assign n14693 = n13250 ^ n8571 ^ 1'b0 ;
  assign n14694 = n14664 ^ n646 ^ 1'b0 ;
  assign n14696 = n2443 ^ n561 ^ 1'b0 ;
  assign n14697 = n6406 & n14696 ;
  assign n14695 = n1671 & n7199 ;
  assign n14698 = n14697 ^ n14695 ^ 1'b0 ;
  assign n14699 = ~n8260 & n14698 ;
  assign n14700 = n3083 & n6527 ;
  assign n14701 = ~n14166 & n14700 ;
  assign n14702 = ( ~n3488 & n5417 ) | ( ~n3488 & n14701 ) | ( n5417 & n14701 ) ;
  assign n14703 = n9651 | n10480 ;
  assign n14704 = ~n2811 & n6614 ;
  assign n14705 = n12722 & ~n14704 ;
  assign n14706 = ~n11101 & n14705 ;
  assign n14708 = n7304 ^ n760 ^ 1'b0 ;
  assign n14707 = n275 | n2469 ;
  assign n14709 = n14708 ^ n14707 ^ 1'b0 ;
  assign n14710 = n2175 & n2599 ;
  assign n14711 = n3664 & n14710 ;
  assign n14712 = ( n4651 & n4876 ) | ( n4651 & ~n10554 ) | ( n4876 & ~n10554 ) ;
  assign n14713 = ~n7315 & n14712 ;
  assign n14715 = ~n5032 & n13943 ;
  assign n14716 = n14715 ^ n1106 ^ 1'b0 ;
  assign n14714 = n9909 & ~n10032 ;
  assign n14717 = n14716 ^ n14714 ^ 1'b0 ;
  assign n14718 = n2198 & ~n2535 ;
  assign n14719 = ( ~x50 & n4745 ) | ( ~x50 & n14718 ) | ( n4745 & n14718 ) ;
  assign n14720 = n615 & n8935 ;
  assign n14721 = n2927 & n14720 ;
  assign n14722 = n14719 & ~n14721 ;
  assign n14723 = n9677 ^ n1903 ^ 1'b0 ;
  assign n14724 = n14723 ^ n12011 ^ n6440 ;
  assign n14725 = n8632 ^ n1800 ^ 1'b0 ;
  assign n14726 = ~n4044 & n7074 ;
  assign n14727 = ~n2933 & n14726 ;
  assign n14728 = n865 | n14727 ;
  assign n14729 = n10218 & ~n14728 ;
  assign n14730 = n14725 | n14729 ;
  assign n14731 = ~n1636 & n2007 ;
  assign n14732 = n2774 ^ n2667 ^ 1'b0 ;
  assign n14733 = n3503 & ~n14732 ;
  assign n14734 = n14733 ^ n11266 ^ n9398 ;
  assign n14735 = n10195 ^ n5901 ^ 1'b0 ;
  assign n14736 = n10228 ^ n9134 ^ n9085 ;
  assign n14737 = n3836 ^ n3738 ^ n1123 ;
  assign n14738 = ( n1374 & n9743 ) | ( n1374 & ~n14737 ) | ( n9743 & ~n14737 ) ;
  assign n14739 = n12766 ^ n630 ^ 1'b0 ;
  assign n14740 = n14738 | n14739 ;
  assign n14741 = n1309 | n3582 ;
  assign n14742 = ~n330 & n14601 ;
  assign n14743 = ~x95 & n13799 ;
  assign n14744 = n2800 ^ n2063 ^ n457 ;
  assign n14745 = n4307 & n6346 ;
  assign n14746 = ~n4854 & n14745 ;
  assign n14747 = n14744 & n14746 ;
  assign n14748 = n14747 ^ n401 ^ 1'b0 ;
  assign n14749 = n5395 ^ n3208 ^ 1'b0 ;
  assign n14750 = n3654 & n4865 ;
  assign n14751 = ~n14749 & n14750 ;
  assign n14752 = n14749 & n14751 ;
  assign n14753 = n11111 | n14752 ;
  assign n14754 = n6487 & ~n14753 ;
  assign n14755 = n7990 ^ n6027 ^ 1'b0 ;
  assign n14756 = x45 & n14755 ;
  assign n14757 = n4524 & ~n9035 ;
  assign n14758 = n9733 ^ n2663 ^ 1'b0 ;
  assign n14759 = ~n6040 & n14758 ;
  assign n14760 = n13701 ^ n11147 ^ n3434 ;
  assign n14761 = ( n7207 & ~n10025 ) | ( n7207 & n11751 ) | ( ~n10025 & n11751 ) ;
  assign n14762 = n7731 ^ n3383 ^ 1'b0 ;
  assign n14763 = n9827 ^ n7796 ^ 1'b0 ;
  assign n14764 = n317 | n14763 ;
  assign n14765 = n5145 ^ n3857 ^ 1'b0 ;
  assign n14766 = n3990 & n14765 ;
  assign n14767 = n3037 | n14766 ;
  assign n14768 = ~n3993 & n12368 ;
  assign n14769 = ( n185 & ~n1316 ) | ( n185 & n11941 ) | ( ~n1316 & n11941 ) ;
  assign n14774 = n1191 & ~n10186 ;
  assign n14770 = n1191 & ~n5722 ;
  assign n14771 = n14770 ^ n1952 ^ 1'b0 ;
  assign n14772 = n5573 | n10333 ;
  assign n14773 = n14771 | n14772 ;
  assign n14775 = n14774 ^ n14773 ^ 1'b0 ;
  assign n14776 = n2912 | n12091 ;
  assign n14777 = n6315 & n11945 ;
  assign n14778 = ~n14776 & n14777 ;
  assign n14779 = n7234 ^ n6412 ^ 1'b0 ;
  assign n14782 = ~n7309 & n12487 ;
  assign n14783 = n8713 & n14782 ;
  assign n14780 = n2403 | n7567 ;
  assign n14781 = ( n636 & ~n6991 ) | ( n636 & n14780 ) | ( ~n6991 & n14780 ) ;
  assign n14784 = n14783 ^ n14781 ^ n1583 ;
  assign n14785 = n3050 | n14784 ;
  assign n14786 = n6247 & ~n14785 ;
  assign n14788 = n5581 & n8750 ;
  assign n14789 = n2817 & n14788 ;
  assign n14787 = n5718 | n10393 ;
  assign n14790 = n14789 ^ n14787 ^ 1'b0 ;
  assign n14791 = n14790 ^ n11476 ^ 1'b0 ;
  assign n14793 = n2866 ^ n932 ^ 1'b0 ;
  assign n14794 = ( n387 & n4254 ) | ( n387 & ~n14793 ) | ( n4254 & ~n14793 ) ;
  assign n14795 = n14794 ^ n413 ^ 1'b0 ;
  assign n14796 = n9839 | n14795 ;
  assign n14792 = ( ~n7046 & n9625 ) | ( ~n7046 & n11234 ) | ( n9625 & n11234 ) ;
  assign n14797 = n14796 ^ n14792 ^ n5486 ;
  assign n14799 = n3684 ^ n1582 ^ 1'b0 ;
  assign n14798 = ( n3658 & n5203 ) | ( n3658 & n9821 ) | ( n5203 & n9821 ) ;
  assign n14800 = n14799 ^ n14798 ^ n11668 ;
  assign n14801 = n4081 & n5356 ;
  assign n14802 = ~n12573 & n14801 ;
  assign n14803 = n14802 ^ n1399 ^ 1'b0 ;
  assign n14804 = n5836 & n9858 ;
  assign n14805 = n14804 ^ n13540 ^ 1'b0 ;
  assign n14807 = ( ~n2117 & n2625 ) | ( ~n2117 & n3967 ) | ( n2625 & n3967 ) ;
  assign n14808 = n14807 ^ n8181 ^ 1'b0 ;
  assign n14806 = n2945 & ~n8783 ;
  assign n14809 = n14808 ^ n14806 ^ 1'b0 ;
  assign n14810 = n6303 & n14809 ;
  assign n14811 = n14810 ^ n8249 ^ n1560 ;
  assign n14812 = ~n2377 & n2878 ;
  assign n14813 = ~n341 & n14812 ;
  assign n14814 = n14813 ^ n14740 ^ n11042 ;
  assign n14815 = n8608 ^ n6168 ^ 1'b0 ;
  assign n14816 = n5501 & ~n8582 ;
  assign n14817 = n14816 ^ n12413 ^ 1'b0 ;
  assign n14818 = n4122 & ~n8086 ;
  assign n14819 = n9679 | n13948 ;
  assign n14820 = n6122 ^ n1741 ^ 1'b0 ;
  assign n14821 = n3712 & n14820 ;
  assign n14822 = n14821 ^ n7189 ^ 1'b0 ;
  assign n14823 = ~n14819 & n14822 ;
  assign n14824 = n13953 ^ n2346 ^ 1'b0 ;
  assign n14825 = n2383 | n14824 ;
  assign n14826 = n3285 ^ n804 ^ 1'b0 ;
  assign n14827 = n169 | n534 ;
  assign n14828 = n2865 | n14827 ;
  assign n14829 = ~n14826 & n14828 ;
  assign n14830 = n14642 & ~n14829 ;
  assign n14831 = n405 & n10686 ;
  assign n14832 = n14831 ^ n12328 ^ 1'b0 ;
  assign n14833 = n14832 ^ n5059 ^ 1'b0 ;
  assign n14836 = n4827 | n7256 ;
  assign n14837 = n9593 ^ n7182 ^ n4575 ;
  assign n14838 = ~n14836 & n14837 ;
  assign n14834 = x95 | n6295 ;
  assign n14835 = n14834 ^ n1410 ^ 1'b0 ;
  assign n14839 = n14838 ^ n14835 ^ 1'b0 ;
  assign n14840 = x56 & n14839 ;
  assign n14841 = n138 & n10223 ;
  assign n14842 = ~n1461 & n13200 ;
  assign n14843 = ~n14841 & n14842 ;
  assign n14844 = n1451 | n10647 ;
  assign n14845 = n14844 ^ n2574 ^ n612 ;
  assign n14846 = n5815 ^ n323 ^ 1'b0 ;
  assign n14847 = n1372 | n14846 ;
  assign n14848 = n12893 & ~n14847 ;
  assign n14849 = n7004 & n12115 ;
  assign n14850 = n14849 ^ n9724 ^ 1'b0 ;
  assign n14851 = n13339 ^ n886 ^ 1'b0 ;
  assign n14852 = n4796 ^ n484 ^ 1'b0 ;
  assign n14853 = n11368 ^ n6686 ^ n1907 ;
  assign n14854 = ( n14077 & ~n14852 ) | ( n14077 & n14853 ) | ( ~n14852 & n14853 ) ;
  assign n14855 = n7117 & ~n7933 ;
  assign n14856 = n14855 ^ n13450 ^ 1'b0 ;
  assign n14857 = n6999 ^ n3946 ^ 1'b0 ;
  assign n14858 = ~n1397 & n10954 ;
  assign n14859 = n13701 ^ n3313 ^ 1'b0 ;
  assign n14860 = n2937 | n11458 ;
  assign n14861 = ~n628 & n11263 ;
  assign n14862 = n13653 & n14861 ;
  assign n14864 = n5043 ^ n4702 ^ 1'b0 ;
  assign n14865 = n4120 & n14864 ;
  assign n14863 = n5581 & ~n7653 ;
  assign n14866 = n14865 ^ n14863 ^ 1'b0 ;
  assign n14867 = n889 | n3593 ;
  assign n14868 = n4292 ^ n1033 ^ n582 ;
  assign n14869 = n7538 ^ n6030 ^ 1'b0 ;
  assign n14870 = n5623 ^ n683 ^ 1'b0 ;
  assign n14871 = ~n13958 & n14870 ;
  assign n14872 = n7806 ^ n4497 ^ 1'b0 ;
  assign n14873 = ~n5255 & n12536 ;
  assign n14874 = ( n1090 & ~n14872 ) | ( n1090 & n14873 ) | ( ~n14872 & n14873 ) ;
  assign n14875 = n4272 & n4292 ;
  assign n14876 = n7089 & n14875 ;
  assign n14877 = n13233 & ~n14876 ;
  assign n14878 = ~n7604 & n8861 ;
  assign n14879 = n14878 ^ n13997 ^ 1'b0 ;
  assign n14880 = ( x123 & n14877 ) | ( x123 & n14879 ) | ( n14877 & n14879 ) ;
  assign n14881 = n10901 ^ x107 ^ 1'b0 ;
  assign n14882 = n14880 & ~n14881 ;
  assign n14883 = n6093 & n12497 ;
  assign n14884 = n5099 & n14883 ;
  assign n14885 = n7587 ^ n5211 ^ 1'b0 ;
  assign n14886 = ~n4512 & n5916 ;
  assign n14887 = n14885 & n14886 ;
  assign n14888 = n7347 & ~n10372 ;
  assign n14890 = n3358 & n3781 ;
  assign n14889 = ( n806 & n6116 ) | ( n806 & ~n9067 ) | ( n6116 & ~n9067 ) ;
  assign n14891 = n14890 ^ n14889 ^ n6802 ;
  assign n14892 = ~n4457 & n5267 ;
  assign n14893 = ~n11589 & n14892 ;
  assign n14896 = n492 & ~n9381 ;
  assign n14897 = n14896 ^ n2841 ^ 1'b0 ;
  assign n14894 = ~n4250 & n4264 ;
  assign n14895 = ~n1627 & n14894 ;
  assign n14898 = n14897 ^ n14895 ^ 1'b0 ;
  assign n14899 = x124 & n671 ;
  assign n14900 = ~n8036 & n14899 ;
  assign n14901 = n8113 ^ n2007 ^ 1'b0 ;
  assign n14902 = ~n14900 & n14901 ;
  assign n14903 = n14902 ^ n7491 ^ n3832 ;
  assign n14904 = n2135 | n12601 ;
  assign n14905 = n14904 ^ n655 ^ 1'b0 ;
  assign n14906 = n4992 ^ n2821 ^ 1'b0 ;
  assign n14907 = ~n3299 & n14906 ;
  assign n14908 = n14439 ^ n5541 ^ n3317 ;
  assign n14909 = n14907 & ~n14908 ;
  assign n14910 = n4761 & ~n5027 ;
  assign n14911 = n6190 & n14910 ;
  assign n14912 = n13592 ^ n6299 ^ 1'b0 ;
  assign n14913 = n14911 | n14912 ;
  assign n14914 = n14913 ^ n4977 ^ 1'b0 ;
  assign n14915 = ~n7930 & n14914 ;
  assign n14916 = n14915 ^ n4518 ^ 1'b0 ;
  assign n14917 = n14916 ^ n6233 ^ n3221 ;
  assign n14918 = n13882 ^ n1196 ^ 1'b0 ;
  assign n14919 = n10645 & ~n14918 ;
  assign n14920 = n1002 ^ n174 ^ 1'b0 ;
  assign n14921 = n3889 | n14920 ;
  assign n14922 = n1950 & n14921 ;
  assign n14923 = ( ~n6629 & n9340 ) | ( ~n6629 & n14081 ) | ( n9340 & n14081 ) ;
  assign n14924 = n4796 ^ n2409 ^ n505 ;
  assign n14925 = n14924 ^ n2751 ^ 1'b0 ;
  assign n14926 = n2254 | n14925 ;
  assign n14927 = ~n8367 & n14926 ;
  assign n14930 = n4563 ^ n3952 ^ 1'b0 ;
  assign n14931 = ( n1970 & n2419 ) | ( n1970 & n14930 ) | ( n2419 & n14930 ) ;
  assign n14928 = ( x78 & n4806 ) | ( x78 & n5897 ) | ( n4806 & n5897 ) ;
  assign n14929 = x108 & ~n14928 ;
  assign n14932 = n14931 ^ n14929 ^ 1'b0 ;
  assign n14933 = ( n5464 & n9686 ) | ( n5464 & ~n12090 ) | ( n9686 & ~n12090 ) ;
  assign n14934 = n7592 ^ n7176 ^ 1'b0 ;
  assign n14935 = n14933 | n14934 ;
  assign n14936 = n431 & ~n10366 ;
  assign n14937 = n6837 & n14936 ;
  assign n14938 = ( n1034 & n10317 ) | ( n1034 & n14937 ) | ( n10317 & n14937 ) ;
  assign n14939 = n14835 ^ n1517 ^ 1'b0 ;
  assign n14940 = n9327 ^ n5737 ^ 1'b0 ;
  assign n14941 = n14940 ^ n1669 ^ 1'b0 ;
  assign n14942 = n980 & ~n14941 ;
  assign n14943 = n5432 | n8882 ;
  assign n14944 = n10697 & ~n14943 ;
  assign n14945 = n11276 ^ n3556 ^ 1'b0 ;
  assign n14946 = ~n9791 & n14945 ;
  assign n14947 = ~n5889 & n14946 ;
  assign n14948 = ~n299 & n14947 ;
  assign n14949 = n4520 | n14627 ;
  assign n14950 = n8140 ^ n6241 ^ 1'b0 ;
  assign n14951 = n3267 ^ n1307 ^ 1'b0 ;
  assign n14952 = ~n13504 & n14951 ;
  assign n14953 = n5001 ^ x97 ^ 1'b0 ;
  assign n14954 = ~n8009 & n14953 ;
  assign n14955 = n14952 & ~n14954 ;
  assign n14956 = n14955 ^ n1794 ^ 1'b0 ;
  assign n14957 = n2151 & ~n5221 ;
  assign n14958 = n3842 ^ n1798 ^ 1'b0 ;
  assign n14959 = n14958 ^ n8680 ^ 1'b0 ;
  assign n14960 = n717 | n1554 ;
  assign n14961 = n12744 ^ n9522 ^ n4767 ;
  assign n14962 = ( ~n2634 & n14960 ) | ( ~n2634 & n14961 ) | ( n14960 & n14961 ) ;
  assign n14963 = n10096 ^ n5883 ^ 1'b0 ;
  assign n14964 = n9962 ^ n2529 ^ 1'b0 ;
  assign n14965 = n7420 ^ n6027 ^ n3939 ;
  assign n14966 = n129 & ~n1410 ;
  assign n14967 = ~n2896 & n14966 ;
  assign n14968 = n14967 ^ n5365 ^ 1'b0 ;
  assign n14969 = n9564 & n14968 ;
  assign n14970 = ~n14806 & n14969 ;
  assign n14971 = n9968 & n14970 ;
  assign n14972 = n8377 & n10847 ;
  assign n14973 = n1085 & n14972 ;
  assign n14974 = ~n13053 & n14973 ;
  assign n14975 = n7395 ^ n1661 ^ 1'b0 ;
  assign n14976 = n14975 ^ n6761 ^ n5122 ;
  assign n14978 = ( ~n3741 & n4727 ) | ( ~n3741 & n13767 ) | ( n4727 & n13767 ) ;
  assign n14977 = n1776 ^ n1631 ^ 1'b0 ;
  assign n14979 = n14978 ^ n14977 ^ n1208 ;
  assign n14980 = n681 & n4770 ;
  assign n14981 = n14979 & n14980 ;
  assign n14982 = n14976 & ~n14981 ;
  assign n14983 = ~n2691 & n14982 ;
  assign n14984 = n10381 ^ n938 ^ 1'b0 ;
  assign n14985 = n3610 ^ n2346 ^ 1'b0 ;
  assign n14986 = x68 & ~n12711 ;
  assign n14987 = n5407 ^ n891 ^ 1'b0 ;
  assign n14988 = n2740 & n14987 ;
  assign n14989 = n6157 ^ x126 ^ 1'b0 ;
  assign n14990 = n3184 & ~n14989 ;
  assign n14991 = ~n12199 & n14990 ;
  assign n14992 = n13845 ^ n4439 ^ 1'b0 ;
  assign n14993 = n4115 & n14992 ;
  assign n14994 = n14424 & n14993 ;
  assign n14995 = n1189 & n14994 ;
  assign n14996 = ~n3999 & n12103 ;
  assign n14997 = n5687 & n14996 ;
  assign n14998 = n10719 | n14162 ;
  assign n14999 = n14997 & ~n14998 ;
  assign n15000 = ( n2341 & ~n11329 ) | ( n2341 & n12979 ) | ( ~n11329 & n12979 ) ;
  assign n15001 = n14037 ^ n6097 ^ 1'b0 ;
  assign n15002 = n2940 & ~n15001 ;
  assign n15003 = ~n177 & n15002 ;
  assign n15004 = n7971 & n15003 ;
  assign n15005 = n6828 ^ n5923 ^ n4111 ;
  assign n15006 = n2090 & n8723 ;
  assign n15007 = n7232 & n15006 ;
  assign n15008 = n7857 & ~n15007 ;
  assign n15009 = n15008 ^ n857 ^ 1'b0 ;
  assign n15010 = ( n2860 & n10298 ) | ( n2860 & n15009 ) | ( n10298 & n15009 ) ;
  assign n15018 = n6789 & ~n12683 ;
  assign n15019 = n15018 ^ n9220 ^ 1'b0 ;
  assign n15012 = n5132 | n10057 ;
  assign n15013 = n5039 & ~n15012 ;
  assign n15014 = n14222 | n15013 ;
  assign n15015 = n4371 & ~n15014 ;
  assign n15011 = ~n1034 & n2198 ;
  assign n15016 = n15015 ^ n15011 ^ 1'b0 ;
  assign n15017 = n373 & n15016 ;
  assign n15020 = n15019 ^ n15017 ^ 1'b0 ;
  assign n15021 = n2958 & n7514 ;
  assign n15022 = ~n1765 & n4124 ;
  assign n15023 = n1765 | n15022 ;
  assign n15024 = n1843 & ~n4727 ;
  assign n15025 = n15024 ^ n6547 ^ n909 ;
  assign n15026 = n1649 & n15025 ;
  assign n15027 = n15026 ^ n9402 ^ 1'b0 ;
  assign n15028 = n15027 ^ n912 ^ 1'b0 ;
  assign n15029 = n12660 ^ n6199 ^ 1'b0 ;
  assign n15030 = n5078 ^ n4195 ^ 1'b0 ;
  assign n15031 = n13135 & n15030 ;
  assign n15032 = n15029 & n15031 ;
  assign n15033 = n3751 ^ n129 ^ 1'b0 ;
  assign n15034 = n1844 ^ n785 ^ n381 ;
  assign n15035 = ~n1286 & n15034 ;
  assign n15036 = ~n15033 & n15035 ;
  assign n15037 = n8828 & n13233 ;
  assign n15038 = n15037 ^ n3204 ^ 1'b0 ;
  assign n15039 = n12098 ^ n5927 ^ 1'b0 ;
  assign n15040 = n15038 & ~n15039 ;
  assign n15041 = n3529 | n13492 ;
  assign n15042 = n15041 ^ n10716 ^ 1'b0 ;
  assign n15043 = n13855 ^ n7079 ^ n2219 ;
  assign n15044 = n15043 ^ n9144 ^ 1'b0 ;
  assign n15045 = n15042 & ~n15044 ;
  assign n15046 = n14979 & n15045 ;
  assign n15047 = n6140 ^ x102 ^ 1'b0 ;
  assign n15048 = n12091 ^ n3970 ^ 1'b0 ;
  assign n15049 = n1597 | n15048 ;
  assign n15050 = n3770 & ~n15049 ;
  assign n15051 = n14240 ^ n1423 ^ 1'b0 ;
  assign n15052 = n15050 | n15051 ;
  assign n15053 = n10224 & n14587 ;
  assign n15054 = n1571 & n15007 ;
  assign n15055 = n7475 ^ n1703 ^ 1'b0 ;
  assign n15056 = ( n930 & n9434 ) | ( n930 & ~n12931 ) | ( n9434 & ~n12931 ) ;
  assign n15057 = n13532 ^ n7482 ^ n7195 ;
  assign n15058 = n9426 & ~n10136 ;
  assign n15059 = n7032 ^ n1879 ^ 1'b0 ;
  assign n15060 = ~n15058 & n15059 ;
  assign n15061 = n1428 & ~n8948 ;
  assign n15062 = n15061 ^ n12531 ^ 1'b0 ;
  assign n15063 = n1760 & ~n8624 ;
  assign n15064 = n15063 ^ n3728 ^ 1'b0 ;
  assign n15065 = ( n10303 & ~n10495 ) | ( n10303 & n15064 ) | ( ~n10495 & n15064 ) ;
  assign n15066 = n14531 ^ n9209 ^ 1'b0 ;
  assign n15067 = n15065 & ~n15066 ;
  assign n15068 = n854 & ~n11294 ;
  assign n15069 = n14895 ^ n12653 ^ 1'b0 ;
  assign n15070 = n1246 & n2586 ;
  assign n15071 = n15070 ^ n4420 ^ 1'b0 ;
  assign n15072 = n14257 ^ n4384 ^ 1'b0 ;
  assign n15073 = n15071 | n15072 ;
  assign n15074 = ~n2932 & n8354 ;
  assign n15075 = n7156 & n15074 ;
  assign n15076 = n9880 ^ n7709 ^ 1'b0 ;
  assign n15077 = n191 & n15076 ;
  assign n15078 = n5747 | n15077 ;
  assign n15083 = n3067 | n7971 ;
  assign n15084 = n15083 ^ n4261 ^ 1'b0 ;
  assign n15080 = n2979 & n6940 ;
  assign n15081 = ~n1154 & n15080 ;
  assign n15082 = n15081 ^ n8331 ^ n1094 ;
  assign n15079 = n9643 ^ n7497 ^ n2612 ;
  assign n15085 = n15084 ^ n15082 ^ n15079 ;
  assign n15086 = ~n331 & n2219 ;
  assign n15087 = n15086 ^ n11690 ^ 1'b0 ;
  assign n15088 = n4133 | n7488 ;
  assign n15089 = n2147 | n5256 ;
  assign n15090 = n15089 ^ n11230 ^ 1'b0 ;
  assign n15091 = n5237 & n14086 ;
  assign n15092 = n15091 ^ n10691 ^ 1'b0 ;
  assign n15093 = ~n2022 & n8684 ;
  assign n15094 = n15093 ^ n630 ^ 1'b0 ;
  assign n15095 = n10448 ^ n7808 ^ n7251 ;
  assign n15096 = n4041 & ~n10733 ;
  assign n15097 = ~n15095 & n15096 ;
  assign n15098 = n5927 ^ n3681 ^ 1'b0 ;
  assign n15099 = n10272 ^ n6586 ^ n3706 ;
  assign n15100 = n15099 ^ n13917 ^ n2017 ;
  assign n15101 = n11061 ^ n6729 ^ 1'b0 ;
  assign n15102 = n9336 | n15101 ;
  assign n15103 = n11939 & ~n13698 ;
  assign n15104 = n14166 ^ n2849 ^ 1'b0 ;
  assign n15105 = ~n8905 & n15104 ;
  assign n15106 = n3113 | n4716 ;
  assign n15107 = n1182 | n12895 ;
  assign n15108 = n15106 & ~n15107 ;
  assign n15109 = n391 & ~n15108 ;
  assign n15110 = n15109 ^ n13195 ^ 1'b0 ;
  assign n15111 = n13981 ^ n11044 ^ 1'b0 ;
  assign n15112 = n3429 ^ x53 ^ 1'b0 ;
  assign n15113 = n888 & ~n15112 ;
  assign n15114 = ~n5487 & n10096 ;
  assign n15115 = n4303 & n15114 ;
  assign n15116 = n5219 & ~n15115 ;
  assign n15117 = n15116 ^ n5107 ^ 1'b0 ;
  assign n15118 = ~n11632 & n15117 ;
  assign n15119 = n6287 ^ n3684 ^ 1'b0 ;
  assign n15120 = n15118 & n15119 ;
  assign n15121 = n2138 & n10339 ;
  assign n15122 = ~n10735 & n15121 ;
  assign n15123 = ( ~n1621 & n5900 ) | ( ~n1621 & n11444 ) | ( n5900 & n11444 ) ;
  assign n15124 = n2081 | n15123 ;
  assign n15125 = n15124 ^ n442 ^ 1'b0 ;
  assign n15126 = n15125 ^ n4815 ^ 1'b0 ;
  assign n15127 = n663 & ~n5918 ;
  assign n15128 = n11280 & ~n15127 ;
  assign n15129 = n5428 ^ n5344 ^ 1'b0 ;
  assign n15130 = n9819 ^ n2622 ^ 1'b0 ;
  assign n15131 = n7949 & n9881 ;
  assign n15132 = n681 & ~n3158 ;
  assign n15133 = n3435 & n15132 ;
  assign n15134 = n15133 ^ n7391 ^ 1'b0 ;
  assign n15135 = ~n1089 & n8425 ;
  assign n15136 = n15135 ^ x126 ^ 1'b0 ;
  assign n15137 = n8289 ^ n7872 ^ 1'b0 ;
  assign n15138 = n1796 | n15137 ;
  assign n15139 = n7380 | n8641 ;
  assign n15140 = n15139 ^ n279 ^ 1'b0 ;
  assign n15141 = n9868 ^ n805 ^ 1'b0 ;
  assign n15142 = ~n640 & n671 ;
  assign n15143 = n15142 ^ n7573 ^ 1'b0 ;
  assign n15144 = n7877 ^ n1009 ^ 1'b0 ;
  assign n15145 = n1991 & ~n15144 ;
  assign n15146 = n12814 ^ n1623 ^ 1'b0 ;
  assign n15147 = ( n2605 & n3725 ) | ( n2605 & n9294 ) | ( n3725 & n9294 ) ;
  assign n15148 = n1353 & n2258 ;
  assign n15149 = ~n282 & n15148 ;
  assign n15150 = n15149 ^ n9591 ^ 1'b0 ;
  assign n15151 = n8771 ^ n305 ^ 1'b0 ;
  assign n15152 = n6024 & ~n15151 ;
  assign n15153 = n15150 | n15152 ;
  assign n15154 = n5579 & ~n13043 ;
  assign n15155 = n3221 ^ n2065 ^ n1154 ;
  assign n15156 = n420 | n15155 ;
  assign n15157 = n3214 & ~n5628 ;
  assign n15158 = n15157 ^ n1485 ^ 1'b0 ;
  assign n15159 = ~n6420 & n6545 ;
  assign n15160 = n15159 ^ n4672 ^ 1'b0 ;
  assign n15161 = n13573 ^ n5389 ^ 1'b0 ;
  assign n15162 = n12614 ^ n3724 ^ 1'b0 ;
  assign n15163 = ~n9243 & n15162 ;
  assign n15164 = n15163 ^ n1250 ^ 1'b0 ;
  assign n15167 = n8325 | n8798 ;
  assign n15165 = x108 & n14968 ;
  assign n15166 = n15165 ^ n7344 ^ 1'b0 ;
  assign n15168 = n15167 ^ n15166 ^ 1'b0 ;
  assign n15169 = n12411 & n15168 ;
  assign n15170 = n15169 ^ n14115 ^ n11884 ;
  assign n15171 = n1568 & ~n13979 ;
  assign n15172 = n1408 & n15171 ;
  assign n15173 = n4259 | n12443 ;
  assign n15174 = n15172 & ~n15173 ;
  assign n15175 = n12396 & n15174 ;
  assign n15176 = n2115 | n10089 ;
  assign n15177 = n15176 ^ n10104 ^ 1'b0 ;
  assign n15178 = n5758 ^ x13 ^ 1'b0 ;
  assign n15179 = n15177 & ~n15178 ;
  assign n15180 = n15179 ^ n13228 ^ 1'b0 ;
  assign n15181 = n5401 & n15180 ;
  assign n15182 = n7178 ^ n3999 ^ n1765 ;
  assign n15183 = n3279 & ~n15182 ;
  assign n15184 = n833 & n15183 ;
  assign n15185 = ~n605 & n6829 ;
  assign n15186 = n15185 ^ n869 ^ 1'b0 ;
  assign n15187 = n5747 | n9545 ;
  assign n15188 = n15187 ^ n11432 ^ 1'b0 ;
  assign n15189 = ( ~n4532 & n15186 ) | ( ~n4532 & n15188 ) | ( n15186 & n15188 ) ;
  assign n15190 = n4518 | n5355 ;
  assign n15191 = n3033 & ~n15190 ;
  assign n15192 = n1477 | n1828 ;
  assign n15193 = ( n1746 & n1782 ) | ( n1746 & n3485 ) | ( n1782 & n3485 ) ;
  assign n15194 = n15193 ^ n4454 ^ 1'b0 ;
  assign n15195 = n3935 | n15194 ;
  assign n15196 = n15192 | n15195 ;
  assign n15198 = n1477 | n10815 ;
  assign n15199 = n4599 & ~n15198 ;
  assign n15197 = n10971 & n14520 ;
  assign n15200 = n15199 ^ n15197 ^ 1'b0 ;
  assign n15201 = n4030 & ~n6847 ;
  assign n15202 = n11944 ^ n11467 ^ n938 ;
  assign n15203 = ( ~n6003 & n15201 ) | ( ~n6003 & n15202 ) | ( n15201 & n15202 ) ;
  assign n15204 = n2690 | n4755 ;
  assign n15205 = n15203 & n15204 ;
  assign n15209 = n5190 & n9903 ;
  assign n15210 = ~x100 & n15209 ;
  assign n15211 = n15210 ^ n5965 ^ 1'b0 ;
  assign n15206 = n12905 ^ x21 ^ 1'b0 ;
  assign n15207 = n14059 | n15206 ;
  assign n15208 = n11481 | n15207 ;
  assign n15212 = n15211 ^ n15208 ^ 1'b0 ;
  assign n15213 = n9519 & n13892 ;
  assign n15214 = n4593 & n15213 ;
  assign n15215 = ~n1705 & n10709 ;
  assign n15216 = n3332 ^ n1628 ^ 1'b0 ;
  assign n15217 = ( ~n3247 & n7713 ) | ( ~n3247 & n15216 ) | ( n7713 & n15216 ) ;
  assign n15218 = n10466 & n15217 ;
  assign n15219 = n15215 | n15218 ;
  assign n15220 = n15214 & n15219 ;
  assign n15221 = n15211 ^ n11071 ^ n1500 ;
  assign n15222 = n11761 ^ n10270 ^ n7506 ;
  assign n15223 = n14310 ^ n10229 ^ n8586 ;
  assign n15224 = n9670 & n10449 ;
  assign n15225 = n15224 ^ n7601 ^ 1'b0 ;
  assign n15226 = n2775 | n3678 ;
  assign n15227 = n15226 ^ n4138 ^ n2523 ;
  assign n15228 = n15227 ^ n1786 ^ 1'b0 ;
  assign n15229 = n6668 & ~n15228 ;
  assign n15230 = n15229 ^ n8273 ^ 1'b0 ;
  assign n15231 = ~n4574 & n13107 ;
  assign n15232 = n15231 ^ n2672 ^ 1'b0 ;
  assign n15233 = n857 & ~n15081 ;
  assign n15234 = n15233 ^ n5625 ^ 1'b0 ;
  assign n15235 = n15234 ^ n6629 ^ 1'b0 ;
  assign n15236 = n3138 & ~n15235 ;
  assign n15237 = n7142 ^ n4122 ^ 1'b0 ;
  assign n15238 = n4038 & n15237 ;
  assign n15239 = ~n3315 & n15238 ;
  assign n15240 = n539 & ~n4285 ;
  assign n15241 = n8471 ^ n513 ^ 1'b0 ;
  assign n15242 = ( ~n4620 & n10361 ) | ( ~n4620 & n11066 ) | ( n10361 & n11066 ) ;
  assign n15243 = ~n15241 & n15242 ;
  assign n15244 = n15243 ^ n6516 ^ 1'b0 ;
  assign n15245 = n13044 & n13729 ;
  assign n15246 = n5963 ^ n3252 ^ n2700 ;
  assign n15247 = n4757 ^ n1592 ^ 1'b0 ;
  assign n15248 = ( n3729 & ~n8677 ) | ( n3729 & n15247 ) | ( ~n8677 & n15247 ) ;
  assign n15249 = n15248 ^ n5396 ^ n1292 ;
  assign n15250 = n4247 | n6768 ;
  assign n15252 = n5206 & ~n9328 ;
  assign n15251 = n6550 & ~n9388 ;
  assign n15253 = n15252 ^ n15251 ^ 1'b0 ;
  assign n15254 = n15253 ^ n3568 ^ 1'b0 ;
  assign n15255 = n13903 & n15254 ;
  assign n15256 = n429 & n12226 ;
  assign n15257 = ~n8856 & n15256 ;
  assign n15258 = n4589 ^ n3728 ^ 1'b0 ;
  assign n15259 = n7046 ^ n5519 ^ n2069 ;
  assign n15260 = n6931 ^ n2178 ^ 1'b0 ;
  assign n15261 = ( n7067 & n15259 ) | ( n7067 & ~n15260 ) | ( n15259 & ~n15260 ) ;
  assign n15262 = n9384 | n15261 ;
  assign n15263 = n15258 & ~n15262 ;
  assign n15264 = x13 & ~n15263 ;
  assign n15265 = n5712 ^ n2715 ^ n566 ;
  assign n15266 = n3061 ^ n2285 ^ 1'b0 ;
  assign n15267 = n2117 & n4169 ;
  assign n15268 = n5310 | n15267 ;
  assign n15269 = n15266 | n15268 ;
  assign n15273 = n8953 & n12858 ;
  assign n15274 = n484 & ~n15273 ;
  assign n15275 = n7960 & n15274 ;
  assign n15270 = n2594 ^ n383 ^ 1'b0 ;
  assign n15271 = x6 & ~n15270 ;
  assign n15272 = ~n8441 & n15271 ;
  assign n15276 = n15275 ^ n15272 ^ 1'b0 ;
  assign n15277 = n15276 ^ n13671 ^ n9841 ;
  assign n15278 = n6007 & ~n6738 ;
  assign n15279 = ~n2325 & n15278 ;
  assign n15280 = n413 | n988 ;
  assign n15281 = n7992 | n11574 ;
  assign n15282 = n14214 ^ n5070 ^ 1'b0 ;
  assign n15283 = n12935 & n15282 ;
  assign n15284 = ~n399 & n2760 ;
  assign n15285 = ~n13233 & n15284 ;
  assign n15286 = n7320 & ~n15285 ;
  assign n15287 = n15286 ^ n3406 ^ 1'b0 ;
  assign n15289 = n6219 & ~n8534 ;
  assign n15290 = n15289 ^ n7575 ^ 1'b0 ;
  assign n15288 = n6171 & n7416 ;
  assign n15291 = n15290 ^ n15288 ^ 1'b0 ;
  assign n15292 = ( x54 & n4132 ) | ( x54 & ~n6830 ) | ( n4132 & ~n6830 ) ;
  assign n15293 = ~n2371 & n3946 ;
  assign n15294 = n15293 ^ n1624 ^ 1'b0 ;
  assign n15295 = n2603 ^ n788 ^ 1'b0 ;
  assign n15296 = n13950 & n15295 ;
  assign n15297 = n2690 & n15296 ;
  assign n15298 = ~n12092 & n15297 ;
  assign n15299 = n12018 | n15298 ;
  assign n15300 = n312 & n11504 ;
  assign n15301 = n15300 ^ n341 ^ 1'b0 ;
  assign n15302 = n8200 | n10195 ;
  assign n15303 = n15302 ^ x36 ^ 1'b0 ;
  assign n15304 = ~n648 & n9489 ;
  assign n15305 = ~n15303 & n15304 ;
  assign n15306 = n3376 ^ n1743 ^ n1217 ;
  assign n15307 = n15306 ^ n4030 ^ 1'b0 ;
  assign n15308 = n6271 & n11686 ;
  assign n15309 = ( n1420 & n5810 ) | ( n1420 & n8351 ) | ( n5810 & n8351 ) ;
  assign n15310 = n541 | n635 ;
  assign n15311 = x9 | n15310 ;
  assign n15312 = n8187 & n15311 ;
  assign n15313 = n7972 & n15312 ;
  assign n15314 = n15313 ^ n5199 ^ 1'b0 ;
  assign n15315 = ~n2896 & n15314 ;
  assign n15316 = n15315 ^ n14718 ^ 1'b0 ;
  assign n15317 = n188 & n1892 ;
  assign n15318 = n15317 ^ n4847 ^ 1'b0 ;
  assign n15320 = ~n229 & n2464 ;
  assign n15319 = n2940 & n8503 ;
  assign n15321 = n15320 ^ n15319 ^ 1'b0 ;
  assign n15322 = n14455 ^ n3791 ^ 1'b0 ;
  assign n15323 = n846 & ~n12934 ;
  assign n15324 = ~n15322 & n15323 ;
  assign n15325 = ( ~n7772 & n11518 ) | ( ~n7772 & n13126 ) | ( n11518 & n13126 ) ;
  assign n15326 = n15325 ^ n240 ^ 1'b0 ;
  assign n15327 = n15324 | n15326 ;
  assign n15328 = n15327 ^ n3977 ^ 1'b0 ;
  assign n15329 = ~n9138 & n13570 ;
  assign n15330 = n6599 & ~n11772 ;
  assign n15332 = n2937 ^ n2888 ^ x48 ;
  assign n15333 = ( n2841 & n13706 ) | ( n2841 & ~n15332 ) | ( n13706 & ~n15332 ) ;
  assign n15331 = n3922 & n8300 ;
  assign n15334 = n15333 ^ n15331 ^ 1'b0 ;
  assign n15337 = n6243 ^ n299 ^ 1'b0 ;
  assign n15335 = n6933 ^ n375 ^ 1'b0 ;
  assign n15336 = n593 & ~n15335 ;
  assign n15338 = n15337 ^ n15336 ^ 1'b0 ;
  assign n15339 = n6826 & n14257 ;
  assign n15340 = n1669 & n3415 ;
  assign n15341 = n7837 | n15340 ;
  assign n15342 = n14349 ^ n9172 ^ 1'b0 ;
  assign n15343 = n5810 & ~n15342 ;
  assign n15350 = n4406 | n7376 ;
  assign n15344 = n9161 ^ n4363 ^ 1'b0 ;
  assign n15345 = n15344 ^ n5785 ^ n1265 ;
  assign n15346 = n15345 ^ n3922 ^ 1'b0 ;
  assign n15347 = n15346 ^ n3831 ^ 1'b0 ;
  assign n15348 = n3408 & ~n4489 ;
  assign n15349 = n15347 & n15348 ;
  assign n15351 = n15350 ^ n15349 ^ n9786 ;
  assign n15352 = n15351 ^ n7451 ^ 1'b0 ;
  assign n15353 = n10609 & ~n15352 ;
  assign n15354 = ( ~n6806 & n9860 ) | ( ~n6806 & n15353 ) | ( n9860 & n15353 ) ;
  assign n15355 = n15081 ^ n9823 ^ n2752 ;
  assign n15356 = ~n646 & n10700 ;
  assign n15357 = ( n5774 & n12727 ) | ( n5774 & n15356 ) | ( n12727 & n15356 ) ;
  assign n15358 = n9562 & ~n12932 ;
  assign n15359 = n9334 ^ n4205 ^ 1'b0 ;
  assign n15360 = n12125 ^ n3887 ^ 1'b0 ;
  assign n15361 = n5291 | n6855 ;
  assign n15362 = n15361 ^ n987 ^ 1'b0 ;
  assign n15363 = n15362 ^ n2375 ^ 1'b0 ;
  assign n15364 = n9400 & ~n15363 ;
  assign n15365 = n15364 ^ n4952 ^ 1'b0 ;
  assign n15366 = n6742 | n15365 ;
  assign n15367 = n6506 ^ n3277 ^ n338 ;
  assign n15368 = n271 & n11813 ;
  assign n15369 = n15368 ^ n7669 ^ 1'b0 ;
  assign n15370 = n4651 ^ x3 ^ 1'b0 ;
  assign n15371 = ~n6815 & n15370 ;
  assign n15372 = ~n5866 & n15371 ;
  assign n15373 = n13618 ^ n953 ^ 1'b0 ;
  assign n15374 = n1526 | n15373 ;
  assign n15375 = ~n3989 & n7048 ;
  assign n15376 = ( ~n10517 & n15374 ) | ( ~n10517 & n15375 ) | ( n15374 & n15375 ) ;
  assign n15377 = n5778 ^ n3167 ^ 1'b0 ;
  assign n15378 = n15377 ^ n13471 ^ 1'b0 ;
  assign n15379 = n10950 ^ n8967 ^ 1'b0 ;
  assign n15380 = n1734 & n3746 ;
  assign n15381 = ~n1734 & n15380 ;
  assign n15382 = n15381 ^ n8740 ^ 1'b0 ;
  assign n15383 = n14435 | n15382 ;
  assign n15384 = n129 & n210 ;
  assign n15385 = n7462 & n15384 ;
  assign n15386 = n15385 ^ n12612 ^ 1'b0 ;
  assign n15387 = ~n3674 & n15386 ;
  assign n15388 = n15387 ^ n13306 ^ 1'b0 ;
  assign n15389 = ~n734 & n7666 ;
  assign n15390 = ~n12691 & n15389 ;
  assign n15391 = n13681 ^ n3151 ^ 1'b0 ;
  assign n15392 = n3143 & ~n15391 ;
  assign n15393 = n8946 ^ n3756 ^ n1892 ;
  assign n15394 = n8924 ^ n7891 ^ 1'b0 ;
  assign n15395 = n6643 ^ n4049 ^ 1'b0 ;
  assign n15396 = n7790 & n9492 ;
  assign n15397 = n3585 ^ n2721 ^ n2291 ;
  assign n15398 = n7567 ^ n6266 ^ 1'b0 ;
  assign n15399 = ~n15397 & n15398 ;
  assign n15400 = n954 ^ n276 ^ 1'b0 ;
  assign n15401 = n282 | n15400 ;
  assign n15402 = n2154 & ~n4010 ;
  assign n15403 = n13807 ^ n3385 ^ 1'b0 ;
  assign n15404 = ~n15402 & n15403 ;
  assign n15405 = n10006 & n15404 ;
  assign n15406 = n15401 & n15405 ;
  assign n15407 = n12964 ^ n11042 ^ n10588 ;
  assign n15408 = n9225 ^ n7759 ^ n3268 ;
  assign n15409 = ~n975 & n10978 ;
  assign n15410 = ~n15408 & n15409 ;
  assign n15411 = n9322 & n10062 ;
  assign n15412 = n15411 ^ n11273 ^ 1'b0 ;
  assign n15413 = n6849 ^ n2364 ^ 1'b0 ;
  assign n15414 = ~n974 & n15413 ;
  assign n15415 = n3135 & ~n15414 ;
  assign n15416 = n14470 ^ n8052 ^ n7029 ;
  assign n15417 = ~n1784 & n10855 ;
  assign n15418 = ~n10855 & n15417 ;
  assign n15419 = ~n4895 & n14158 ;
  assign n15420 = n4895 & n15419 ;
  assign n15421 = n467 | n686 ;
  assign n15422 = n467 & ~n15421 ;
  assign n15423 = n692 & n1940 ;
  assign n15424 = ~n1560 & n15423 ;
  assign n15425 = n215 | n5057 ;
  assign n15426 = n15425 ^ n2749 ^ 1'b0 ;
  assign n15427 = n15424 | n15426 ;
  assign n15428 = n15424 & ~n15427 ;
  assign n15429 = n15422 | n15428 ;
  assign n15430 = n15420 & ~n15429 ;
  assign n15431 = ~n15418 & n15430 ;
  assign n15432 = ~n2694 & n10719 ;
  assign n15433 = n688 & ~n15432 ;
  assign n15434 = n15433 ^ n14535 ^ n3815 ;
  assign n15435 = n4246 ^ n3249 ^ 1'b0 ;
  assign n15436 = n15434 & n15435 ;
  assign n15437 = n9357 & ~n12418 ;
  assign n15439 = n620 & n1089 ;
  assign n15440 = n15439 ^ n5288 ^ 1'b0 ;
  assign n15438 = n6958 ^ n3578 ^ n2440 ;
  assign n15441 = n15440 ^ n15438 ^ 1'b0 ;
  assign n15443 = n14552 ^ n9968 ^ 1'b0 ;
  assign n15442 = ~n2531 & n13233 ;
  assign n15444 = n15443 ^ n15442 ^ 1'b0 ;
  assign n15445 = n2007 | n9939 ;
  assign n15446 = n15445 ^ n12791 ^ 1'b0 ;
  assign n15447 = n4527 & ~n5616 ;
  assign n15448 = ~n3336 & n15447 ;
  assign n15449 = n1413 & n15448 ;
  assign n15450 = n1212 & n1430 ;
  assign n15451 = n15450 ^ n3861 ^ 1'b0 ;
  assign n15452 = n8969 ^ n3831 ^ 1'b0 ;
  assign n15453 = n1183 & ~n15452 ;
  assign n15454 = n15453 ^ n10107 ^ 1'b0 ;
  assign n15455 = n3065 & n15454 ;
  assign n15456 = n5191 & n15455 ;
  assign n15457 = n15456 ^ n5842 ^ 1'b0 ;
  assign n15458 = n13846 ^ n992 ^ 1'b0 ;
  assign n15459 = n1734 & n15458 ;
  assign n15460 = ~n4749 & n15459 ;
  assign n15461 = n9425 ^ n7939 ^ 1'b0 ;
  assign n15462 = n15461 ^ n3376 ^ 1'b0 ;
  assign n15463 = n2857 ^ n2166 ^ 1'b0 ;
  assign n15464 = ~n1106 & n15463 ;
  assign n15465 = ~n3582 & n12457 ;
  assign n15466 = n15465 ^ n10459 ^ 1'b0 ;
  assign n15467 = ~n6694 & n15466 ;
  assign n15468 = n4230 & ~n15174 ;
  assign n15469 = n6415 | n7153 ;
  assign n15470 = n7962 | n15469 ;
  assign n15471 = ( n1198 & ~n8753 ) | ( n1198 & n15470 ) | ( ~n8753 & n15470 ) ;
  assign n15472 = ( n11756 & n14374 ) | ( n11756 & ~n15057 ) | ( n14374 & ~n15057 ) ;
  assign n15473 = ~n5043 & n14030 ;
  assign n15474 = n11184 ^ n5925 ^ n2661 ;
  assign n15475 = ~n12487 & n15474 ;
  assign n15476 = ( ~n4782 & n7683 ) | ( ~n4782 & n8842 ) | ( n7683 & n8842 ) ;
  assign n15479 = n6332 ^ n3249 ^ 1'b0 ;
  assign n15480 = n3931 & n15479 ;
  assign n15481 = n11368 | n15480 ;
  assign n15477 = n8743 ^ n4667 ^ 1'b0 ;
  assign n15478 = ~n8749 & n15477 ;
  assign n15482 = n15481 ^ n15478 ^ 1'b0 ;
  assign n15483 = n1089 & ~n8401 ;
  assign n15484 = ~n9492 & n15483 ;
  assign n15485 = n744 & n10962 ;
  assign n15488 = n2339 | n4937 ;
  assign n15486 = n3036 ^ n1550 ^ 1'b0 ;
  assign n15487 = ~n10770 & n15486 ;
  assign n15489 = n15488 ^ n15487 ^ 1'b0 ;
  assign n15490 = ( ~n6866 & n12489 ) | ( ~n6866 & n15489 ) | ( n12489 & n15489 ) ;
  assign n15491 = n4110 & n11764 ;
  assign n15492 = n2581 & n4630 ;
  assign n15493 = n1006 & n5556 ;
  assign n15494 = n1135 & n15493 ;
  assign n15495 = n4538 & ~n15494 ;
  assign n15496 = n15495 ^ n1655 ^ 1'b0 ;
  assign n15497 = n12707 ^ n1451 ^ 1'b0 ;
  assign n15498 = n11338 & ~n15497 ;
  assign n15499 = n15498 ^ n8967 ^ 1'b0 ;
  assign n15500 = n5610 | n15499 ;
  assign n15501 = n7676 ^ n264 ^ 1'b0 ;
  assign n15502 = n306 & ~n3432 ;
  assign n15503 = n15502 ^ n640 ^ 1'b0 ;
  assign n15504 = n7265 & n12068 ;
  assign n15505 = n5742 & ~n5902 ;
  assign n15506 = n15504 & n15505 ;
  assign n15507 = n4044 & ~n9096 ;
  assign n15508 = n2535 | n2964 ;
  assign n15509 = n12754 & n15508 ;
  assign n15510 = n9630 ^ n9067 ^ 1'b0 ;
  assign n15511 = ~n3366 & n15510 ;
  assign n15512 = n15511 ^ n13182 ^ 1'b0 ;
  assign n15513 = ( n167 & n8613 ) | ( n167 & ~n15512 ) | ( n8613 & ~n15512 ) ;
  assign n15514 = n10001 ^ n8481 ^ n821 ;
  assign n15515 = n10624 ^ n7685 ^ 1'b0 ;
  assign n15516 = n3792 & ~n5816 ;
  assign n15517 = n15516 ^ n868 ^ 1'b0 ;
  assign n15518 = n10006 & ~n14928 ;
  assign n15519 = n15518 ^ n1669 ^ 1'b0 ;
  assign n15520 = n1159 ^ n1056 ^ 1'b0 ;
  assign n15521 = n9315 | n15520 ;
  assign n15522 = ~n6036 & n8178 ;
  assign n15523 = n3480 | n5910 ;
  assign n15524 = n5824 | n15523 ;
  assign n15525 = ~n7238 & n15524 ;
  assign n15526 = n12331 ^ n5876 ^ 1'b0 ;
  assign n15527 = ~n15525 & n15526 ;
  assign n15528 = n1868 ^ n1670 ^ n1372 ;
  assign n15529 = ~n9063 & n15528 ;
  assign n15530 = n13652 ^ n9387 ^ 1'b0 ;
  assign n15531 = ( n12395 & n15529 ) | ( n12395 & n15530 ) | ( n15529 & n15530 ) ;
  assign n15532 = n15296 ^ n4648 ^ 1'b0 ;
  assign n15533 = n15531 & ~n15532 ;
  assign n15534 = n1111 & ~n11241 ;
  assign n15535 = n15534 ^ n2717 ^ 1'b0 ;
  assign n15539 = ~n193 & n3631 ;
  assign n15540 = ~n1870 & n15539 ;
  assign n15536 = n671 & ~n2329 ;
  assign n15537 = n8526 & n12038 ;
  assign n15538 = ~n15536 & n15537 ;
  assign n15541 = n15540 ^ n15538 ^ 1'b0 ;
  assign n15542 = n4451 | n8885 ;
  assign n15543 = n15073 ^ n10313 ^ 1'b0 ;
  assign n15544 = n4612 ^ n2091 ^ 1'b0 ;
  assign n15545 = n7230 | n15544 ;
  assign n15546 = n14686 ^ n1072 ^ 1'b0 ;
  assign n15547 = n1803 ^ n1089 ^ 1'b0 ;
  assign n15548 = n332 & ~n937 ;
  assign n15549 = ~n2322 & n15548 ;
  assign n15550 = ( ~n1376 & n3871 ) | ( ~n1376 & n11024 ) | ( n3871 & n11024 ) ;
  assign n15551 = n15550 ^ n7031 ^ 1'b0 ;
  assign n15552 = n15549 | n15551 ;
  assign n15553 = ~n1392 & n4390 ;
  assign n15554 = n15553 ^ n7002 ^ 1'b0 ;
  assign n15555 = n5493 & n15554 ;
  assign n15556 = n15199 | n15555 ;
  assign n15557 = ~n7056 & n8440 ;
  assign n15558 = n15557 ^ n4230 ^ 1'b0 ;
  assign n15559 = n2432 & ~n9677 ;
  assign n15560 = n6806 & n15559 ;
  assign n15561 = ~n374 & n3091 ;
  assign n15562 = n11441 ^ n3126 ^ 1'b0 ;
  assign n15563 = n15561 & ~n15562 ;
  assign n15567 = n6786 & ~n10707 ;
  assign n15568 = n15567 ^ n4323 ^ 1'b0 ;
  assign n15566 = ~n1034 & n1800 ;
  assign n15569 = n15568 ^ n15566 ^ 1'b0 ;
  assign n15570 = n6806 | n15569 ;
  assign n15564 = n6849 ^ n6625 ^ 1'b0 ;
  assign n15565 = ~n12458 & n15564 ;
  assign n15571 = n15570 ^ n15565 ^ 1'b0 ;
  assign n15572 = n1017 | n6338 ;
  assign n15573 = ~n4537 & n6464 ;
  assign n15574 = n8353 ^ n502 ^ 1'b0 ;
  assign n15575 = n9779 | n15574 ;
  assign n15576 = n10517 ^ n10208 ^ 1'b0 ;
  assign n15577 = n2590 & ~n13112 ;
  assign n15578 = ~n1364 & n15577 ;
  assign n15582 = ~n452 & n3840 ;
  assign n15583 = n15582 ^ n8539 ^ 1'b0 ;
  assign n15579 = n3496 ^ n1585 ^ 1'b0 ;
  assign n15580 = n1722 | n15579 ;
  assign n15581 = n14355 & ~n15580 ;
  assign n15584 = n15583 ^ n15581 ^ 1'b0 ;
  assign n15587 = n1724 & ~n7022 ;
  assign n15588 = ~n1788 & n15587 ;
  assign n15585 = ( n1309 & n6308 ) | ( n1309 & ~n8311 ) | ( n6308 & ~n8311 ) ;
  assign n15586 = n2472 & n15585 ;
  assign n15589 = n15588 ^ n15586 ^ 1'b0 ;
  assign n15590 = n2756 ^ n2676 ^ 1'b0 ;
  assign n15591 = n7513 ^ n4327 ^ n576 ;
  assign n15592 = n2060 & n12386 ;
  assign n15593 = ( ~n2756 & n15591 ) | ( ~n2756 & n15592 ) | ( n15591 & n15592 ) ;
  assign n15594 = n15590 & n15593 ;
  assign n15595 = n633 & ~n12043 ;
  assign n15596 = ~n1099 & n14800 ;
  assign n15597 = n15595 & n15596 ;
  assign n15598 = n8345 ^ n2268 ^ 1'b0 ;
  assign n15600 = n13894 ^ n9226 ^ 1'b0 ;
  assign n15601 = ~n346 & n15600 ;
  assign n15599 = n990 & ~n9422 ;
  assign n15602 = n15601 ^ n15599 ^ 1'b0 ;
  assign n15603 = ~n6214 & n7303 ;
  assign n15604 = n15603 ^ n6023 ^ 1'b0 ;
  assign n15605 = n12333 ^ n2798 ^ 1'b0 ;
  assign n15606 = n3494 & ~n15605 ;
  assign n15607 = ~n15604 & n15606 ;
  assign n15608 = n10355 ^ n612 ^ 1'b0 ;
  assign n15609 = n2159 | n15608 ;
  assign n15610 = n15609 ^ n6631 ^ n5041 ;
  assign n15611 = n8046 & ~n9228 ;
  assign n15612 = n15610 & n15611 ;
  assign n15613 = ( ~n10435 & n10495 ) | ( ~n10435 & n15612 ) | ( n10495 & n15612 ) ;
  assign n15614 = n15578 ^ n417 ^ 1'b0 ;
  assign n15615 = n15217 | n15614 ;
  assign n15616 = ~n1487 & n4380 ;
  assign n15617 = n6930 & n15616 ;
  assign n15618 = ( n745 & n4181 ) | ( n745 & ~n4651 ) | ( n4181 & ~n4651 ) ;
  assign n15619 = n5209 | n15618 ;
  assign n15620 = n15619 ^ n6717 ^ 1'b0 ;
  assign n15621 = n15620 ^ n3062 ^ 1'b0 ;
  assign n15622 = ~n3324 & n15621 ;
  assign n15623 = ( x3 & ~n14864 ) | ( x3 & n15622 ) | ( ~n14864 & n15622 ) ;
  assign n15624 = ~n4376 & n4948 ;
  assign n15625 = n15624 ^ n3202 ^ n1573 ;
  assign n15626 = ~n12054 & n12753 ;
  assign n15627 = n3953 & n15626 ;
  assign n15628 = ~n8437 & n13178 ;
  assign n15629 = n10563 ^ n5514 ^ 1'b0 ;
  assign n15630 = n15629 ^ n7259 ^ 1'b0 ;
  assign n15631 = n4348 | n10387 ;
  assign n15632 = n15631 ^ n8776 ^ 1'b0 ;
  assign n15633 = n11123 ^ n4429 ^ n3055 ;
  assign n15634 = n15633 ^ n12910 ^ n8220 ;
  assign n15635 = ~n1131 & n15634 ;
  assign n15636 = ~n15632 & n15635 ;
  assign n15637 = n9703 & ~n10801 ;
  assign n15638 = n15637 ^ n11944 ^ 1'b0 ;
  assign n15639 = ( n1843 & n8813 ) | ( n1843 & ~n15638 ) | ( n8813 & ~n15638 ) ;
  assign n15640 = n529 | n9927 ;
  assign n15641 = ~n11490 & n15640 ;
  assign n15642 = n15491 ^ n2081 ^ 1'b0 ;
  assign n15643 = ~n8547 & n15642 ;
  assign n15644 = n276 & n7265 ;
  assign n15645 = n15644 ^ n1013 ^ 1'b0 ;
  assign n15646 = n4911 & n15645 ;
  assign n15647 = n11129 & n14574 ;
  assign n15648 = ~n15646 & n15647 ;
  assign n15649 = n13863 ^ n612 ^ 1'b0 ;
  assign n15653 = n385 & ~n3653 ;
  assign n15654 = n15653 ^ n1529 ^ 1'b0 ;
  assign n15650 = n2137 | n2692 ;
  assign n15651 = n15650 ^ n1948 ^ 1'b0 ;
  assign n15652 = n7999 & ~n15651 ;
  assign n15655 = n15654 ^ n15652 ^ 1'b0 ;
  assign n15656 = n10707 | n15655 ;
  assign n15657 = n15656 ^ n10921 ^ 1'b0 ;
  assign n15658 = n1384 ^ n374 ^ n361 ;
  assign n15659 = n15658 ^ n11445 ^ 1'b0 ;
  assign n15660 = n11288 & ~n15659 ;
  assign n15661 = n8953 ^ n7724 ^ 1'b0 ;
  assign n15662 = n15385 ^ n8799 ^ x84 ;
  assign n15664 = ( n301 & n2209 ) | ( n301 & ~n9348 ) | ( n2209 & ~n9348 ) ;
  assign n15663 = n6073 ^ x110 ^ x37 ;
  assign n15665 = n15664 ^ n15663 ^ 1'b0 ;
  assign n15666 = n1856 | n15665 ;
  assign n15667 = n5633 ^ n4010 ^ 1'b0 ;
  assign n15668 = n5468 | n15667 ;
  assign n15669 = n1580 & ~n15668 ;
  assign n15670 = n15668 & n15669 ;
  assign n15671 = n527 | n3617 ;
  assign n15672 = n3617 & ~n15671 ;
  assign n15673 = n15672 ^ n7251 ^ 1'b0 ;
  assign n15674 = n15670 | n15673 ;
  assign n15675 = n15674 ^ n7201 ^ 1'b0 ;
  assign n15676 = ( ~n4689 & n8572 ) | ( ~n4689 & n15675 ) | ( n8572 & n15675 ) ;
  assign n15677 = x64 & ~n2089 ;
  assign n15678 = n2089 & n15677 ;
  assign n15679 = n2396 & n2525 ;
  assign n15680 = ~n2396 & n15679 ;
  assign n15681 = n15680 ^ n3994 ^ 1'b0 ;
  assign n15682 = n691 & n15681 ;
  assign n15683 = n15678 & n15682 ;
  assign n15684 = n15683 ^ n9192 ^ 1'b0 ;
  assign n15685 = n12190 & ~n15684 ;
  assign n15686 = n1819 & n8226 ;
  assign n15687 = n15261 ^ n7274 ^ 1'b0 ;
  assign n15688 = n241 & n12631 ;
  assign n15689 = n15688 ^ n4305 ^ 1'b0 ;
  assign n15690 = n7005 & ~n13168 ;
  assign n15691 = n381 & n15690 ;
  assign n15692 = ~n886 & n1029 ;
  assign n15693 = ~n1036 & n15692 ;
  assign n15694 = n3563 & n15031 ;
  assign n15695 = n15694 ^ n746 ^ 1'b0 ;
  assign n15696 = n3938 & n15695 ;
  assign n15697 = n9496 ^ n1540 ^ 1'b0 ;
  assign n15698 = n15697 ^ n13478 ^ n3706 ;
  assign n15699 = n7499 ^ n1675 ^ 1'b0 ;
  assign n15700 = n15699 ^ n7504 ^ 1'b0 ;
  assign n15701 = n5082 & n14539 ;
  assign n15702 = n15701 ^ n4614 ^ 1'b0 ;
  assign n15705 = x120 & ~n7163 ;
  assign n15706 = n15705 ^ n5840 ^ 1'b0 ;
  assign n15707 = n1785 | n15706 ;
  assign n15708 = n15707 ^ n4288 ^ 1'b0 ;
  assign n15703 = n13667 ^ n588 ^ 1'b0 ;
  assign n15704 = x20 & ~n15703 ;
  assign n15709 = n15708 ^ n15704 ^ 1'b0 ;
  assign n15715 = n3734 ^ n1193 ^ 1'b0 ;
  assign n15716 = n2810 | n15715 ;
  assign n15710 = n2348 ^ n674 ^ 1'b0 ;
  assign n15711 = n857 & n15710 ;
  assign n15712 = n15711 ^ n7272 ^ 1'b0 ;
  assign n15713 = n4344 | n15712 ;
  assign n15714 = ( n8252 & n15601 ) | ( n8252 & ~n15713 ) | ( n15601 & ~n15713 ) ;
  assign n15717 = n15716 ^ n15714 ^ n842 ;
  assign n15718 = ~n707 & n12598 ;
  assign n15719 = n856 & n15718 ;
  assign n15720 = n593 & ~n15719 ;
  assign n15721 = n4443 | n8437 ;
  assign n15722 = ( ~n2998 & n4594 ) | ( ~n2998 & n15721 ) | ( n4594 & n15721 ) ;
  assign n15723 = n15722 ^ n1462 ^ n703 ;
  assign n15724 = ~x13 & n1045 ;
  assign n15725 = n15724 ^ n4048 ^ 1'b0 ;
  assign n15726 = ( n5183 & ~n11102 ) | ( n5183 & n13332 ) | ( ~n11102 & n13332 ) ;
  assign n15727 = n15726 ^ n11579 ^ n8652 ;
  assign n15728 = n5683 ^ n3491 ^ n2376 ;
  assign n15729 = n15727 & ~n15728 ;
  assign n15730 = ~n15725 & n15729 ;
  assign n15731 = n15730 ^ n13746 ^ 1'b0 ;
  assign n15732 = ~n1980 & n15731 ;
  assign n15733 = n8587 ^ x19 ^ 1'b0 ;
  assign n15734 = n1920 | n7837 ;
  assign n15735 = n15734 ^ n12103 ^ n5645 ;
  assign n15736 = n6823 & n15735 ;
  assign n15737 = n3453 ^ n2108 ^ n275 ;
  assign n15738 = n15737 ^ n10469 ^ 1'b0 ;
  assign n15748 = ~n2395 & n5433 ;
  assign n15741 = n4662 ^ n1777 ^ 1'b0 ;
  assign n15742 = n2178 & n15741 ;
  assign n15743 = n15742 ^ n3301 ^ 1'b0 ;
  assign n15744 = n3675 & n15743 ;
  assign n15745 = ~n8358 & n15744 ;
  assign n15746 = n11149 & n15745 ;
  assign n15739 = n9745 ^ n2325 ^ 1'b0 ;
  assign n15740 = n6844 & n15739 ;
  assign n15747 = n15746 ^ n15740 ^ 1'b0 ;
  assign n15749 = n15748 ^ n15747 ^ n372 ;
  assign n15750 = n3865 & ~n11753 ;
  assign n15751 = n4749 ^ n2647 ^ 1'b0 ;
  assign n15752 = n13724 & ~n15751 ;
  assign n15753 = n8187 & ~n12393 ;
  assign n15754 = n11382 | n15753 ;
  assign n15755 = n15754 ^ n9307 ^ 1'b0 ;
  assign n15756 = ~n8515 & n15755 ;
  assign n15757 = ~n869 & n10318 ;
  assign n15758 = n14958 ^ n6182 ^ 1'b0 ;
  assign n15759 = n3937 | n15758 ;
  assign n15760 = n5888 & ~n15759 ;
  assign n15761 = n14194 ^ n2947 ^ 1'b0 ;
  assign n15762 = n1658 & ~n9569 ;
  assign n15763 = ( n5125 & n14006 ) | ( n5125 & ~n15762 ) | ( n14006 & ~n15762 ) ;
  assign n15764 = n12319 ^ n557 ^ 1'b0 ;
  assign n15765 = ~n4845 & n5585 ;
  assign n15766 = n12193 ^ n2246 ^ 1'b0 ;
  assign n15767 = n1375 | n15766 ;
  assign n15768 = n15767 ^ n14086 ^ 1'b0 ;
  assign n15769 = n15768 ^ n14201 ^ n12106 ;
  assign n15770 = n15769 ^ n2159 ^ 1'b0 ;
  assign n15771 = n2712 | n15770 ;
  assign n15772 = n7717 ^ n3444 ^ 1'b0 ;
  assign n15773 = n2203 & ~n15772 ;
  assign n15774 = ( n2998 & n3497 ) | ( n2998 & n15773 ) | ( n3497 & n15773 ) ;
  assign n15775 = n9096 ^ n7147 ^ 1'b0 ;
  assign n15776 = n1414 & n4136 ;
  assign n15777 = ~n4136 & n15776 ;
  assign n15778 = n3861 | n7509 ;
  assign n15779 = n3861 & ~n15778 ;
  assign n15780 = n5300 | n15779 ;
  assign n15781 = n15777 & ~n15780 ;
  assign n15782 = n5330 ^ n4837 ^ 1'b0 ;
  assign n15783 = n3842 | n15782 ;
  assign n15784 = n2357 & ~n15783 ;
  assign n15785 = n15784 ^ n8895 ^ 1'b0 ;
  assign n15786 = n1514 ^ n1228 ^ 1'b0 ;
  assign n15787 = n620 & ~n15786 ;
  assign n15788 = n15787 ^ n12397 ^ 1'b0 ;
  assign n15789 = ~n15785 & n15788 ;
  assign n15790 = n7850 ^ n199 ^ 1'b0 ;
  assign n15793 = x118 | n2104 ;
  assign n15794 = n15793 ^ n3340 ^ 1'b0 ;
  assign n15795 = n15794 ^ n6415 ^ 1'b0 ;
  assign n15796 = n3851 | n15795 ;
  assign n15791 = n4811 & ~n8691 ;
  assign n15792 = n15791 ^ n13289 ^ 1'b0 ;
  assign n15797 = n15796 ^ n15792 ^ 1'b0 ;
  assign n15798 = ( n5243 & ~n13870 ) | ( n5243 & n15797 ) | ( ~n13870 & n15797 ) ;
  assign n15799 = n12535 ^ n12143 ^ 1'b0 ;
  assign n15800 = n7113 & n15799 ;
  assign n15802 = x67 | n1122 ;
  assign n15801 = n2945 ^ n337 ^ 1'b0 ;
  assign n15803 = n15802 ^ n15801 ^ 1'b0 ;
  assign n15804 = n15803 ^ n901 ^ 1'b0 ;
  assign n15805 = ~n182 & n15196 ;
  assign n15806 = n15805 ^ n13492 ^ 1'b0 ;
  assign n15807 = n5806 & ~n15340 ;
  assign n15808 = n15807 ^ n4625 ^ 1'b0 ;
  assign n15809 = n5920 ^ n3724 ^ 1'b0 ;
  assign n15810 = n2012 & ~n15809 ;
  assign n15811 = n1320 & n5110 ;
  assign n15812 = n15811 ^ n811 ^ 1'b0 ;
  assign n15813 = n15812 ^ n13342 ^ 1'b0 ;
  assign n15814 = n11327 & n15813 ;
  assign n15815 = ~n2380 & n2677 ;
  assign n15816 = ~n9366 & n15815 ;
  assign n15817 = ~n8980 & n15816 ;
  assign n15818 = n15817 ^ n4331 ^ 1'b0 ;
  assign n15819 = ( x117 & n3557 ) | ( x117 & ~n3562 ) | ( n3557 & ~n3562 ) ;
  assign n15820 = n13691 ^ n7476 ^ 1'b0 ;
  assign n15821 = n1244 | n15820 ;
  assign n15822 = n11129 ^ n6047 ^ 1'b0 ;
  assign n15823 = n15822 ^ n895 ^ 1'b0 ;
  assign n15824 = n5203 | n6657 ;
  assign n15825 = n2554 | n7953 ;
  assign n15826 = n15825 ^ n3878 ^ 1'b0 ;
  assign n15827 = n15824 | n15826 ;
  assign n15828 = ~n5216 & n7660 ;
  assign n15829 = n5466 | n15828 ;
  assign n15830 = n15827 | n15829 ;
  assign n15831 = n13983 ^ n8775 ^ n3977 ;
  assign n15832 = n15831 ^ n13499 ^ 1'b0 ;
  assign n15833 = n1261 | n15832 ;
  assign n15834 = n11017 ^ n1560 ^ 1'b0 ;
  assign n15835 = ( n4108 & n4757 ) | ( n4108 & n15834 ) | ( n4757 & n15834 ) ;
  assign n15836 = n8745 & n15835 ;
  assign n15837 = n1048 & n15836 ;
  assign n15838 = n13544 ^ n1243 ^ 1'b0 ;
  assign n15839 = n15837 | n15838 ;
  assign n15840 = n517 & ~n10237 ;
  assign n15841 = n15840 ^ n5581 ^ 1'b0 ;
  assign n15842 = x48 & n4584 ;
  assign n15843 = ( ~n473 & n3036 ) | ( ~n473 & n3647 ) | ( n3036 & n3647 ) ;
  assign n15844 = n15843 ^ n6560 ^ 1'b0 ;
  assign n15845 = n15842 & n15844 ;
  assign n15846 = ~n856 & n6599 ;
  assign n15847 = ~n8357 & n15846 ;
  assign n15848 = n14968 ^ n4553 ^ 1'b0 ;
  assign n15849 = ~n15847 & n15848 ;
  assign n15850 = n3304 & n15849 ;
  assign n15851 = n12853 ^ n8227 ^ 1'b0 ;
  assign n15852 = n4079 & n15851 ;
  assign n15853 = n2066 | n6541 ;
  assign n15854 = n15853 ^ n6712 ^ 1'b0 ;
  assign n15855 = ~n3511 & n15854 ;
  assign n15856 = n7197 ^ n6280 ^ n2371 ;
  assign n15857 = n15855 & ~n15856 ;
  assign n15858 = n15857 ^ n13060 ^ n6007 ;
  assign n15859 = n10617 ^ n7116 ^ 1'b0 ;
  assign n15860 = n10381 ^ n8935 ^ 1'b0 ;
  assign n15861 = n6524 | n15860 ;
  assign n15862 = n8313 ^ n5805 ^ 1'b0 ;
  assign n15863 = n15861 | n15862 ;
  assign n15864 = n5475 | n9474 ;
  assign n15865 = n6279 & ~n15864 ;
  assign n15866 = n245 & n8343 ;
  assign n15867 = n12871 & n15866 ;
  assign n15868 = n15867 ^ n9534 ^ 1'b0 ;
  assign n15869 = ~n1408 & n15868 ;
  assign n15870 = n13047 ^ n11978 ^ 1'b0 ;
  assign n15871 = n10758 & ~n13441 ;
  assign n15872 = n15871 ^ n15504 ^ 1'b0 ;
  assign n15873 = n10374 | n13471 ;
  assign n15874 = n15057 ^ n12550 ^ 1'b0 ;
  assign n15875 = n12612 | n15874 ;
  assign n15876 = n8455 ^ n4795 ^ 1'b0 ;
  assign n15877 = n14453 | n15876 ;
  assign n15878 = ~n3516 & n15877 ;
  assign n15879 = n2231 ^ n1131 ^ 1'b0 ;
  assign n15880 = n6872 | n8681 ;
  assign n15881 = n15144 | n15880 ;
  assign n15882 = n15879 & ~n15881 ;
  assign n15883 = n141 & ~n4346 ;
  assign n15884 = n10900 & n15883 ;
  assign n15885 = n7850 ^ n6663 ^ 1'b0 ;
  assign n15886 = n771 | n9751 ;
  assign n15887 = n7385 & ~n9090 ;
  assign n15888 = n8956 & ~n15887 ;
  assign n15889 = n7476 ^ n2782 ^ 1'b0 ;
  assign n15890 = n15888 & ~n15889 ;
  assign n15891 = n3684 & ~n9786 ;
  assign n15892 = n616 & n15891 ;
  assign n15893 = n9900 & ~n15892 ;
  assign n15894 = n15893 ^ n12848 ^ 1'b0 ;
  assign n15895 = n2621 & ~n7158 ;
  assign n15896 = x126 & n15895 ;
  assign n15897 = n13133 & ~n13197 ;
  assign n15898 = n11706 & n15897 ;
  assign n15899 = n2087 ^ n299 ^ 1'b0 ;
  assign n15900 = ~n10315 & n15899 ;
  assign n15901 = ~n15898 & n15900 ;
  assign n15902 = n15901 ^ n524 ^ 1'b0 ;
  assign n15903 = ( n2907 & n5129 ) | ( n2907 & n6898 ) | ( n5129 & n6898 ) ;
  assign n15904 = n2549 ^ n1684 ^ 1'b0 ;
  assign n15905 = n8854 & n15904 ;
  assign n15906 = ( ~n6367 & n8480 ) | ( ~n6367 & n15905 ) | ( n8480 & n15905 ) ;
  assign n15907 = n11190 ^ n3012 ^ n2728 ;
  assign n15908 = n10341 ^ n7160 ^ 1'b0 ;
  assign n15909 = n15907 & n15908 ;
  assign n15910 = n5747 | n6339 ;
  assign n15911 = n5993 & ~n15910 ;
  assign n15912 = ~n6003 & n15911 ;
  assign n15913 = n1694 & ~n15912 ;
  assign n15914 = n14888 | n15913 ;
  assign n15916 = n2106 & ~n8919 ;
  assign n15917 = n15916 ^ n6293 ^ 1'b0 ;
  assign n15915 = n4091 & n10686 ;
  assign n15918 = n15917 ^ n15915 ^ 1'b0 ;
  assign n15919 = n2692 | n15918 ;
  assign n15920 = n15919 ^ n2605 ^ 1'b0 ;
  assign n15921 = n10034 ^ n9669 ^ 1'b0 ;
  assign n15922 = n15920 & n15921 ;
  assign n15923 = n1139 & ~n12741 ;
  assign n15924 = n3213 & n3277 ;
  assign n15925 = n15924 ^ n912 ^ 1'b0 ;
  assign n15926 = n15925 ^ n15029 ^ 1'b0 ;
  assign n15927 = n15926 ^ n6670 ^ 1'b0 ;
  assign n15928 = ~n10060 & n15927 ;
  assign n15929 = n11365 ^ n3056 ^ 1'b0 ;
  assign n15930 = n3975 & ~n15929 ;
  assign n15931 = n15930 ^ n4832 ^ 1'b0 ;
  assign n15932 = n5545 | n15504 ;
  assign n15933 = n9074 | n15932 ;
  assign n15937 = n461 & n1965 ;
  assign n15938 = n5330 & ~n15937 ;
  assign n15939 = n15938 ^ n3028 ^ 1'b0 ;
  assign n15934 = n2149 & n8895 ;
  assign n15935 = n15934 ^ n2866 ^ 1'b0 ;
  assign n15936 = n10900 | n15935 ;
  assign n15940 = n15939 ^ n15936 ^ 1'b0 ;
  assign n15941 = n13439 ^ n10971 ^ 1'b0 ;
  assign n15942 = n1958 ^ n849 ^ 1'b0 ;
  assign n15943 = ( n3366 & ~n9875 ) | ( n3366 & n15942 ) | ( ~n9875 & n15942 ) ;
  assign n15944 = ~n5878 & n7639 ;
  assign n15945 = n15944 ^ n15588 ^ 1'b0 ;
  assign n15948 = n4576 ^ n4071 ^ 1'b0 ;
  assign n15949 = ~n937 & n15948 ;
  assign n15946 = n1605 ^ n485 ^ n239 ;
  assign n15947 = n1408 & n15946 ;
  assign n15950 = n15949 ^ n15947 ^ n9584 ;
  assign n15951 = n14432 ^ n3076 ^ 1'b0 ;
  assign n15953 = n15663 ^ n4645 ^ n673 ;
  assign n15954 = n1347 & ~n7365 ;
  assign n15955 = n15954 ^ n2194 ^ 1'b0 ;
  assign n15956 = ~n15953 & n15955 ;
  assign n15952 = ~n1224 & n6755 ;
  assign n15957 = n15956 ^ n15952 ^ 1'b0 ;
  assign n15959 = n863 & ~n6490 ;
  assign n15958 = n452 | n2677 ;
  assign n15960 = n15959 ^ n15958 ^ 1'b0 ;
  assign n15962 = n2437 & ~n6102 ;
  assign n15961 = n2464 & ~n8233 ;
  assign n15963 = n15962 ^ n15961 ^ 1'b0 ;
  assign n15964 = n3244 ^ n306 ^ 1'b0 ;
  assign n15965 = ~n1430 & n3055 ;
  assign n15966 = ~n15964 & n15965 ;
  assign n15967 = n9474 ^ n7818 ^ 1'b0 ;
  assign n15968 = n11708 & ~n15967 ;
  assign n15969 = n1861 & ~n8548 ;
  assign n15970 = n594 & n15969 ;
  assign n15971 = n15968 & n15970 ;
  assign n15973 = ( n2355 & ~n6212 ) | ( n2355 & n12158 ) | ( ~n6212 & n12158 ) ;
  assign n15972 = n10700 & ~n12631 ;
  assign n15974 = n15973 ^ n15972 ^ 1'b0 ;
  assign n15975 = n3983 ^ n3773 ^ 1'b0 ;
  assign n15976 = n1674 & n15842 ;
  assign n15977 = ~n7380 & n15976 ;
  assign n15978 = n8056 & ~n15977 ;
  assign n15979 = n3036 & n15978 ;
  assign n15980 = n6739 & n6860 ;
  assign n15981 = n15980 ^ n14073 ^ 1'b0 ;
  assign n15982 = n14236 ^ n4293 ^ 1'b0 ;
  assign n15983 = ~n306 & n1056 ;
  assign n15984 = n15983 ^ n6421 ^ n5725 ;
  assign n15985 = n9333 ^ n9183 ^ 1'b0 ;
  assign n15986 = n15985 ^ n10071 ^ 1'b0 ;
  assign n15988 = n488 & n2840 ;
  assign n15989 = ~n11174 & n15988 ;
  assign n15992 = ~n2239 & n3472 ;
  assign n15993 = ~n3472 & n15992 ;
  assign n15990 = n129 & n3434 ;
  assign n15991 = ~n3434 & n15990 ;
  assign n15994 = n15993 ^ n15991 ^ 1'b0 ;
  assign n15995 = ~n15989 & n15994 ;
  assign n15987 = ~n4186 & n7782 ;
  assign n15996 = n15995 ^ n15987 ^ n10688 ;
  assign n15997 = ~n994 & n3542 ;
  assign n15998 = n6367 & ~n15997 ;
  assign n15999 = ~x72 & n15998 ;
  assign n16000 = n3723 ^ n3003 ^ 1'b0 ;
  assign n16001 = n2373 & ~n16000 ;
  assign n16002 = n1472 & ~n6661 ;
  assign n16003 = n16002 ^ n3882 ^ 1'b0 ;
  assign n16004 = n3047 & n16003 ;
  assign n16005 = n16004 ^ n2915 ^ 1'b0 ;
  assign n16006 = n3298 & n16005 ;
  assign n16007 = n16006 ^ n756 ^ 1'b0 ;
  assign n16008 = n630 | n7434 ;
  assign n16009 = n659 | n16008 ;
  assign n16010 = n748 | n12936 ;
  assign n16011 = n1967 ^ n450 ^ 1'b0 ;
  assign n16012 = n6927 & n16011 ;
  assign n16013 = n14048 | n14170 ;
  assign n16014 = n16013 ^ n8618 ^ 1'b0 ;
  assign n16015 = n4323 & n16014 ;
  assign n16016 = ~n16012 & n16015 ;
  assign n16017 = n6063 & ~n9956 ;
  assign n16018 = n9052 & n16017 ;
  assign n16019 = n4068 & n5224 ;
  assign n16020 = ~n11647 & n16019 ;
  assign n16021 = n10996 ^ n5122 ^ 1'b0 ;
  assign n16022 = n10982 ^ n5772 ^ 1'b0 ;
  assign n16023 = ( n2958 & n5933 ) | ( n2958 & ~n16022 ) | ( n5933 & ~n16022 ) ;
  assign n16024 = n12091 ^ n3205 ^ 1'b0 ;
  assign n16025 = n3574 & n16024 ;
  assign n16026 = n8510 ^ n1202 ^ 1'b0 ;
  assign n16027 = n16025 & ~n16026 ;
  assign n16028 = ~n3476 & n16027 ;
  assign n16029 = n14404 ^ n3618 ^ 1'b0 ;
  assign n16030 = n1800 & n16029 ;
  assign n16031 = n15022 ^ n6364 ^ 1'b0 ;
  assign n16032 = ~n11688 & n16031 ;
  assign n16033 = ~n9653 & n11611 ;
  assign n16034 = n16033 ^ n469 ^ 1'b0 ;
  assign n16035 = ( n4752 & ~n12212 ) | ( n4752 & n16034 ) | ( ~n12212 & n16034 ) ;
  assign n16036 = n9495 | n16035 ;
  assign n16037 = n2138 & n12789 ;
  assign n16038 = n10460 ^ n6549 ^ 1'b0 ;
  assign n16039 = n4118 & ~n13977 ;
  assign n16040 = n16039 ^ n14137 ^ 1'b0 ;
  assign n16041 = ~n3964 & n6076 ;
  assign n16042 = n7151 ^ n2886 ^ 1'b0 ;
  assign n16043 = n2980 & n16042 ;
  assign n16044 = n16043 ^ n12665 ^ 1'b0 ;
  assign n16045 = ~n5274 & n6936 ;
  assign n16046 = n16045 ^ n1611 ^ 1'b0 ;
  assign n16047 = ~n6457 & n16046 ;
  assign n16048 = n2034 & n16047 ;
  assign n16049 = n15050 ^ n8903 ^ n6632 ;
  assign n16050 = n16049 ^ n5127 ^ 1'b0 ;
  assign n16051 = n10097 & n16050 ;
  assign n16052 = n1230 & ~n1306 ;
  assign n16053 = ~n2511 & n7218 ;
  assign n16054 = n16052 & n16053 ;
  assign n16055 = n477 & n16054 ;
  assign n16056 = n15917 ^ n1189 ^ 1'b0 ;
  assign n16057 = n8471 & ~n16056 ;
  assign n16058 = n16057 ^ n15084 ^ 1'b0 ;
  assign n16059 = n16055 | n16058 ;
  assign n16060 = n5479 ^ n519 ^ 1'b0 ;
  assign n16061 = n9461 & ~n16060 ;
  assign n16062 = n4344 ^ n3178 ^ 1'b0 ;
  assign n16063 = ( n6807 & n7563 ) | ( n6807 & n13666 ) | ( n7563 & n13666 ) ;
  assign n16064 = n8713 ^ n6327 ^ n1999 ;
  assign n16065 = n16063 & n16064 ;
  assign n16066 = ~n16062 & n16065 ;
  assign n16067 = n1920 & ~n16066 ;
  assign n16068 = n15019 & n16067 ;
  assign n16069 = n4224 | n15404 ;
  assign n16072 = ~n4025 & n12370 ;
  assign n16073 = n16072 ^ n3946 ^ 1'b0 ;
  assign n16070 = n5189 | n10156 ;
  assign n16071 = n1382 & n16070 ;
  assign n16074 = n16073 ^ n16071 ^ 1'b0 ;
  assign n16075 = n5327 | n15332 ;
  assign n16076 = n16075 ^ n12917 ^ 1'b0 ;
  assign n16077 = n13838 ^ x82 ^ 1'b0 ;
  assign n16078 = n9867 | n16077 ;
  assign n16079 = n14354 ^ n2151 ^ 1'b0 ;
  assign n16080 = n13604 ^ n4354 ^ 1'b0 ;
  assign n16081 = ( n3156 & n16079 ) | ( n3156 & n16080 ) | ( n16079 & n16080 ) ;
  assign n16086 = n12086 ^ n10580 ^ n4665 ;
  assign n16082 = n3714 & n7138 ;
  assign n16083 = ~n7761 & n16082 ;
  assign n16084 = n16083 ^ n10376 ^ 1'b0 ;
  assign n16085 = n3298 & ~n16084 ;
  assign n16087 = n16086 ^ n16085 ^ 1'b0 ;
  assign n16088 = ( n3958 & n5175 ) | ( n3958 & ~n9760 ) | ( n5175 & ~n9760 ) ;
  assign n16089 = ~n7455 & n16088 ;
  assign n16090 = n3793 & ~n14165 ;
  assign n16091 = n14727 & n16090 ;
  assign n16092 = n7428 | n7920 ;
  assign n16093 = n3202 | n14851 ;
  assign n16094 = ~n5909 & n12771 ;
  assign n16095 = n5942 | n7386 ;
  assign n16096 = n16095 ^ n295 ^ 1'b0 ;
  assign n16097 = n4455 | n16096 ;
  assign n16098 = n16097 ^ n7665 ^ 1'b0 ;
  assign n16099 = n6868 ^ n3943 ^ 1'b0 ;
  assign n16100 = ~n2985 & n4044 ;
  assign n16101 = ~n1658 & n8835 ;
  assign n16102 = ( n7222 & n10975 ) | ( n7222 & n13722 ) | ( n10975 & n13722 ) ;
  assign n16103 = n3608 ^ n2463 ^ 1'b0 ;
  assign n16104 = x101 & n16103 ;
  assign n16105 = ~n312 & n3091 ;
  assign n16106 = n2551 & n5562 ;
  assign n16107 = ~n2786 & n16106 ;
  assign n16108 = n4125 & n5661 ;
  assign n16109 = ( n1765 & n3181 ) | ( n1765 & n12371 ) | ( n3181 & n12371 ) ;
  assign n16110 = n11463 ^ n3012 ^ 1'b0 ;
  assign n16111 = n498 & n8455 ;
  assign n16112 = n16111 ^ n5029 ^ 1'b0 ;
  assign n16113 = n10796 & ~n16112 ;
  assign n16114 = ~n4374 & n9484 ;
  assign n16115 = n1903 | n8005 ;
  assign n16116 = n16115 ^ n11370 ^ n5389 ;
  assign n16117 = n14210 & n16116 ;
  assign n16118 = n16114 & n16117 ;
  assign n16119 = ~n2291 & n2582 ;
  assign n16120 = n7458 ^ n1034 ^ 1'b0 ;
  assign n16121 = n2206 & n5546 ;
  assign n16122 = n16121 ^ n2102 ^ 1'b0 ;
  assign n16123 = n16122 ^ n3684 ^ 1'b0 ;
  assign n16124 = n16120 & n16123 ;
  assign n16125 = n16119 & n16124 ;
  assign n16126 = n16125 ^ n5813 ^ 1'b0 ;
  assign n16127 = n3330 & ~n9615 ;
  assign n16128 = n16126 & n16127 ;
  assign n16129 = n2414 | n9069 ;
  assign n16130 = n7836 & ~n16129 ;
  assign n16131 = ( n6729 & n12281 ) | ( n6729 & n16130 ) | ( n12281 & n16130 ) ;
  assign n16132 = ~n12731 & n16131 ;
  assign n16133 = n15190 ^ n14020 ^ n7299 ;
  assign n16134 = n5263 & n10081 ;
  assign n16135 = n16134 ^ n10161 ^ 1'b0 ;
  assign n16136 = n659 & ~n16135 ;
  assign n16137 = n4822 & n8317 ;
  assign n16138 = n14774 ^ n12184 ^ 1'b0 ;
  assign n16139 = n13543 & ~n16138 ;
  assign n16140 = n3345 | n7891 ;
  assign n16141 = n9719 ^ n9656 ^ 1'b0 ;
  assign n16142 = n8660 ^ n7716 ^ 1'b0 ;
  assign n16143 = ~n16141 & n16142 ;
  assign n16144 = n10833 ^ n5996 ^ 1'b0 ;
  assign n16145 = ( ~n6739 & n9894 ) | ( ~n6739 & n12906 ) | ( n9894 & n12906 ) ;
  assign n16146 = ( n8361 & n16144 ) | ( n8361 & n16145 ) | ( n16144 & n16145 ) ;
  assign n16147 = n14323 ^ n8619 ^ 1'b0 ;
  assign n16148 = ~n5928 & n14494 ;
  assign n16149 = n5057 & n16148 ;
  assign n16150 = n13307 ^ n7776 ^ n4052 ;
  assign n16151 = n9969 & ~n16150 ;
  assign n16152 = n16149 & n16151 ;
  assign n16153 = n182 | n13012 ;
  assign n16154 = n4602 | n14092 ;
  assign n16155 = n2494 | n16154 ;
  assign n16156 = n16155 ^ n9781 ^ 1'b0 ;
  assign n16157 = n1583 & n16156 ;
  assign n16158 = n1055 & n16157 ;
  assign n16159 = ~n7853 & n16158 ;
  assign n16160 = n1256 & ~n11436 ;
  assign n16161 = n2297 | n2783 ;
  assign n16162 = n16161 ^ x56 ^ 1'b0 ;
  assign n16163 = n16162 ^ n7794 ^ 1'b0 ;
  assign n16164 = ~n13078 & n16163 ;
  assign n16165 = n7739 & ~n8727 ;
  assign n16166 = n16165 ^ n8067 ^ 1'b0 ;
  assign n16167 = n6747 ^ n5930 ^ 1'b0 ;
  assign n16168 = n12470 ^ n7229 ^ 1'b0 ;
  assign n16169 = n1532 & n10422 ;
  assign n16170 = ~n4181 & n16169 ;
  assign n16171 = n16170 ^ n7347 ^ 1'b0 ;
  assign n16172 = ~n3876 & n16171 ;
  assign n16173 = n10577 ^ n2909 ^ 1'b0 ;
  assign n16174 = n6635 ^ n1746 ^ 1'b0 ;
  assign n16175 = n3291 | n4606 ;
  assign n16176 = n16175 ^ n5004 ^ 1'b0 ;
  assign n16177 = n10350 ^ n3361 ^ 1'b0 ;
  assign n16178 = n2893 & ~n16177 ;
  assign n16179 = ~n16176 & n16178 ;
  assign n16180 = n16174 & ~n16179 ;
  assign n16181 = n16173 & n16180 ;
  assign n16182 = n748 | n1680 ;
  assign n16183 = n1864 & ~n10559 ;
  assign n16184 = n3686 ^ n1843 ^ 1'b0 ;
  assign n16185 = n1428 & ~n16184 ;
  assign n16186 = ~n8842 & n16185 ;
  assign n16187 = n16186 ^ n9175 ^ 1'b0 ;
  assign n16188 = n16183 & n16187 ;
  assign n16189 = n14675 ^ n10649 ^ n6402 ;
  assign n16190 = n16189 ^ n12497 ^ 1'b0 ;
  assign n16191 = n14042 & n16190 ;
  assign n16192 = n9791 ^ n4474 ^ 1'b0 ;
  assign n16193 = ~n2195 & n16192 ;
  assign n16194 = n4529 ^ n691 ^ 1'b0 ;
  assign n16195 = n1434 & n16194 ;
  assign n16196 = n16195 ^ n13243 ^ n6139 ;
  assign n16197 = ~n5549 & n8751 ;
  assign n16199 = n7156 ^ n6126 ^ n5092 ;
  assign n16198 = ~n9584 & n10943 ;
  assign n16200 = n16199 ^ n16198 ^ 1'b0 ;
  assign n16201 = n9931 ^ n7012 ^ n4893 ;
  assign n16202 = n2487 | n2830 ;
  assign n16203 = n6922 & ~n16202 ;
  assign n16204 = n16203 ^ n9499 ^ 1'b0 ;
  assign n16205 = n319 | n16204 ;
  assign n16206 = ( n1427 & ~n4578 ) | ( n1427 & n16205 ) | ( ~n4578 & n16205 ) ;
  assign n16207 = n10094 ^ n2618 ^ 1'b0 ;
  assign n16208 = n2579 & n16207 ;
  assign n16209 = ~n5725 & n12518 ;
  assign n16210 = ~n2770 & n3351 ;
  assign n16211 = n4466 & n16210 ;
  assign n16212 = n16211 ^ n2930 ^ 1'b0 ;
  assign n16213 = ~n3881 & n13905 ;
  assign n16214 = n15374 ^ n12921 ^ 1'b0 ;
  assign n16215 = n1590 | n7362 ;
  assign n16216 = ~n6159 & n7928 ;
  assign n16217 = ( n5288 & n16215 ) | ( n5288 & n16216 ) | ( n16215 & n16216 ) ;
  assign n16219 = n8300 ^ n5620 ^ 1'b0 ;
  assign n16218 = ~n884 & n13793 ;
  assign n16220 = n16219 ^ n16218 ^ n3424 ;
  assign n16221 = ~n5296 & n5902 ;
  assign n16222 = n3689 ^ n2622 ^ 1'b0 ;
  assign n16223 = n16222 ^ n6683 ^ 1'b0 ;
  assign n16224 = n411 | n16223 ;
  assign n16226 = n1471 ^ n1434 ^ 1'b0 ;
  assign n16225 = n1086 | n4650 ;
  assign n16227 = n16226 ^ n16225 ^ 1'b0 ;
  assign n16229 = n2052 & n5697 ;
  assign n16230 = n16229 ^ n4715 ^ 1'b0 ;
  assign n16228 = ~n632 & n9041 ;
  assign n16231 = n16230 ^ n16228 ^ 1'b0 ;
  assign n16232 = n3540 & ~n16231 ;
  assign n16233 = n5805 ^ n3946 ^ n2092 ;
  assign n16234 = n6243 ^ n5841 ^ n1627 ;
  assign n16235 = n16234 ^ n3396 ^ 1'b0 ;
  assign n16236 = n9162 ^ n8447 ^ n7652 ;
  assign n16237 = n8260 | n16236 ;
  assign n16238 = n9035 & ~n16237 ;
  assign n16239 = ( ~n9141 & n16235 ) | ( ~n9141 & n16238 ) | ( n16235 & n16238 ) ;
  assign n16240 = n13538 ^ n301 ^ 1'b0 ;
  assign n16241 = ~n8523 & n12074 ;
  assign n16242 = n9880 & n16241 ;
  assign n16243 = n9464 ^ n7305 ^ n3607 ;
  assign n16244 = n5217 ^ n2246 ^ 1'b0 ;
  assign n16245 = ~n15826 & n16244 ;
  assign n16246 = n5585 & n16245 ;
  assign n16247 = n7682 & ~n13799 ;
  assign n16248 = n16247 ^ n1736 ^ 1'b0 ;
  assign n16249 = n4050 | n16248 ;
  assign n16250 = ( ~n403 & n7471 ) | ( ~n403 & n10598 ) | ( n7471 & n10598 ) ;
  assign n16251 = n4820 ^ n4487 ^ n2485 ;
  assign n16252 = n16251 ^ n13020 ^ 1'b0 ;
  assign n16253 = n1624 & n16252 ;
  assign n16254 = n12166 ^ n3554 ^ 1'b0 ;
  assign n16255 = n449 | n16254 ;
  assign n16256 = n16255 ^ n1485 ^ n477 ;
  assign n16257 = n14398 ^ n8199 ^ n6893 ;
  assign n16258 = n16256 & ~n16257 ;
  assign n16259 = ~n16253 & n16258 ;
  assign n16260 = n16150 ^ n5788 ^ 1'b0 ;
  assign n16261 = n16260 ^ n12971 ^ n374 ;
  assign n16266 = n671 & n13855 ;
  assign n16264 = n196 | n10800 ;
  assign n16265 = n16264 ^ n1153 ^ 1'b0 ;
  assign n16262 = n5046 & n6927 ;
  assign n16263 = n16262 ^ n8068 ^ 1'b0 ;
  assign n16267 = n16266 ^ n16265 ^ n16263 ;
  assign n16268 = ( n1055 & n3460 ) | ( n1055 & ~n16267 ) | ( n3460 & ~n16267 ) ;
  assign n16269 = n5669 ^ n1774 ^ n1151 ;
  assign n16270 = n16269 ^ n14619 ^ n9615 ;
  assign n16271 = n7992 ^ n7125 ^ 1'b0 ;
  assign n16272 = ~n11312 & n16271 ;
  assign n16273 = n4446 & n7453 ;
  assign n16274 = n16273 ^ x116 ^ 1'b0 ;
  assign n16275 = n1924 | n16274 ;
  assign n16276 = ~n806 & n14265 ;
  assign n16277 = ~n9854 & n16276 ;
  assign n16278 = n1242 | n12168 ;
  assign n16279 = n5433 | n16278 ;
  assign n16280 = n173 | n8271 ;
  assign n16281 = n16280 ^ n12261 ^ n5283 ;
  assign n16282 = n593 & n1529 ;
  assign n16283 = ( n7709 & ~n15340 ) | ( n7709 & n16282 ) | ( ~n15340 & n16282 ) ;
  assign n16284 = n8021 ^ n1496 ^ 1'b0 ;
  assign n16285 = n5281 ^ x32 ^ 1'b0 ;
  assign n16286 = n16285 ^ n5675 ^ 1'b0 ;
  assign n16287 = n14186 | n16286 ;
  assign n16292 = ( ~n2926 & n9017 ) | ( ~n2926 & n13586 ) | ( n9017 & n13586 ) ;
  assign n16290 = n2192 & n2825 ;
  assign n16289 = ( n2099 & ~n3142 ) | ( n2099 & n7520 ) | ( ~n3142 & n7520 ) ;
  assign n16288 = ( n1435 & n4247 ) | ( n1435 & ~n11865 ) | ( n4247 & ~n11865 ) ;
  assign n16291 = n16290 ^ n16289 ^ n16288 ;
  assign n16293 = n16292 ^ n16291 ^ 1'b0 ;
  assign n16294 = n12386 ^ n8748 ^ 1'b0 ;
  assign n16295 = n262 & ~n2457 ;
  assign n16296 = n16005 ^ n12338 ^ 1'b0 ;
  assign n16297 = ~n13576 & n16296 ;
  assign n16298 = ( ~n601 & n12368 ) | ( ~n601 & n14738 ) | ( n12368 & n14738 ) ;
  assign n16299 = n7579 ^ n3591 ^ 1'b0 ;
  assign n16300 = n3109 | n15540 ;
  assign n16301 = n16300 ^ n9939 ^ 1'b0 ;
  assign n16302 = n16301 ^ n15704 ^ 1'b0 ;
  assign n16303 = n6555 & n15455 ;
  assign n16304 = ~n5909 & n16303 ;
  assign n16305 = n14813 ^ n6361 ^ n1101 ;
  assign n16306 = n6200 ^ n2489 ^ 1'b0 ;
  assign n16307 = n6501 & n8328 ;
  assign n16308 = n2871 ^ n2178 ^ 1'b0 ;
  assign n16309 = ~n10439 & n16308 ;
  assign n16310 = n374 & ~n5631 ;
  assign n16311 = n16310 ^ n1484 ^ 1'b0 ;
  assign n16312 = n888 & ~n13586 ;
  assign n16313 = n8310 ^ n5796 ^ 1'b0 ;
  assign n16314 = n4456 & ~n5567 ;
  assign n16315 = ~n16313 & n16314 ;
  assign n16316 = n14073 ^ n1765 ^ 1'b0 ;
  assign n16317 = n2926 | n7602 ;
  assign n16318 = ~n16316 & n16317 ;
  assign n16319 = n6735 ^ n5584 ^ n3892 ;
  assign n16320 = n10057 ^ n9153 ^ 1'b0 ;
  assign n16321 = ( ~n4984 & n7391 ) | ( ~n4984 & n16320 ) | ( n7391 & n16320 ) ;
  assign n16322 = n13238 | n14269 ;
  assign n16323 = n14438 | n16322 ;
  assign n16324 = n14580 & n16323 ;
  assign n16325 = ~n2249 & n16324 ;
  assign n16326 = n4562 | n9210 ;
  assign n16327 = n11935 ^ n10444 ^ 1'b0 ;
  assign n16328 = n3428 | n16327 ;
  assign n16329 = n3080 ^ n1968 ^ 1'b0 ;
  assign n16330 = n16251 | n16329 ;
  assign n16331 = n4025 & n10303 ;
  assign n16332 = n16330 & n16331 ;
  assign n16333 = n380 & ~n16332 ;
  assign n16334 = ~n3789 & n7862 ;
  assign n16335 = n6898 & n8655 ;
  assign n16336 = n2819 | n9583 ;
  assign n16337 = n6787 | n16336 ;
  assign n16338 = n996 | n16337 ;
  assign n16339 = n946 & ~n8425 ;
  assign n16340 = ~n1385 & n16339 ;
  assign n16341 = n6921 | n15015 ;
  assign n16342 = n3325 & ~n11505 ;
  assign n16343 = n4596 & ~n16342 ;
  assign n16344 = n1874 & n16343 ;
  assign n16345 = n2321 | n16344 ;
  assign n16346 = n2112 & ~n16345 ;
  assign n16347 = n3791 & n13316 ;
  assign n16348 = ( n2335 & ~n3429 ) | ( n2335 & n16347 ) | ( ~n3429 & n16347 ) ;
  assign n16349 = n4837 ^ n3253 ^ 1'b0 ;
  assign n16350 = n4343 & ~n16349 ;
  assign n16351 = ~n306 & n16350 ;
  assign n16352 = n15022 & n16351 ;
  assign n16353 = n10609 & ~n16352 ;
  assign n16354 = ~n12687 & n16353 ;
  assign n16355 = n13057 ^ n3011 ^ 1'b0 ;
  assign n16356 = n6555 & ~n16355 ;
  assign n16357 = n15202 ^ n5890 ^ 1'b0 ;
  assign n16358 = n6539 ^ n5538 ^ 1'b0 ;
  assign n16359 = n16357 | n16358 ;
  assign n16360 = ~n2010 & n4064 ;
  assign n16361 = n16360 ^ n5357 ^ 1'b0 ;
  assign n16362 = n2728 & ~n16361 ;
  assign n16363 = n1851 ^ n1800 ^ 1'b0 ;
  assign n16364 = n16362 & n16363 ;
  assign n16365 = n2162 & ~n7872 ;
  assign n16366 = ~n16364 & n16365 ;
  assign n16367 = n12304 ^ n11948 ^ 1'b0 ;
  assign n16368 = n7897 ^ n199 ^ 1'b0 ;
  assign n16369 = n7277 & ~n16368 ;
  assign n16370 = n2933 ^ n1762 ^ n1619 ;
  assign n16371 = n1529 | n6482 ;
  assign n16372 = n16371 ^ n4992 ^ 1'b0 ;
  assign n16373 = n16372 ^ n2292 ^ 1'b0 ;
  assign n16374 = n16370 & n16373 ;
  assign n16375 = n16374 ^ n9198 ^ n6547 ;
  assign n16376 = n16375 ^ n4789 ^ 1'b0 ;
  assign n16377 = n1500 & ~n10498 ;
  assign n16378 = n10498 & n16377 ;
  assign n16379 = n643 & ~n972 ;
  assign n16380 = n972 & n16379 ;
  assign n16381 = n786 | n1761 ;
  assign n16382 = n786 & ~n16381 ;
  assign n16383 = n1573 | n16382 ;
  assign n16384 = n16382 & ~n16383 ;
  assign n16385 = n16380 | n16384 ;
  assign n16386 = n16378 | n16385 ;
  assign n16387 = n16386 ^ n9615 ^ 1'b0 ;
  assign n16388 = n8978 ^ n3728 ^ 1'b0 ;
  assign n16389 = n12716 | n16214 ;
  assign n16390 = ~n1276 & n7012 ;
  assign n16391 = n6376 & n8106 ;
  assign n16392 = ~n16390 & n16391 ;
  assign n16393 = n6916 & n8792 ;
  assign n16394 = n5683 & ~n16393 ;
  assign n16395 = n9795 ^ n3462 ^ 1'b0 ;
  assign n16396 = n2809 | n9265 ;
  assign n16397 = n1568 & ~n13928 ;
  assign n16398 = n16397 ^ n12025 ^ n6638 ;
  assign n16403 = n6051 ^ n4230 ^ n1504 ;
  assign n16400 = n135 & n2652 ;
  assign n16399 = n2401 & ~n3399 ;
  assign n16401 = n16400 ^ n16399 ^ 1'b0 ;
  assign n16402 = n421 & ~n16401 ;
  assign n16404 = n16403 ^ n16402 ^ n9578 ;
  assign n16405 = n691 & n1273 ;
  assign n16406 = n9424 ^ n1337 ^ 1'b0 ;
  assign n16407 = n16336 ^ n990 ^ 1'b0 ;
  assign n16408 = n9580 & n16407 ;
  assign n16410 = n697 | n764 ;
  assign n16411 = n16410 ^ n9091 ^ 1'b0 ;
  assign n16409 = ( ~n2749 & n6698 ) | ( ~n2749 & n9867 ) | ( n6698 & n9867 ) ;
  assign n16412 = n16411 ^ n16409 ^ 1'b0 ;
  assign n16413 = ( n7955 & n8385 ) | ( n7955 & n14222 ) | ( n8385 & n14222 ) ;
  assign n16414 = n3903 ^ n415 ^ 1'b0 ;
  assign n16415 = n13068 | n16414 ;
  assign n16416 = n1621 & ~n16415 ;
  assign n16417 = ~n16413 & n16416 ;
  assign n16418 = n13880 & ~n16417 ;
  assign n16419 = n5936 | n16418 ;
  assign n16420 = n11714 ^ n8070 ^ n5247 ;
  assign n16421 = n2511 & ~n3289 ;
  assign n16422 = n16421 ^ n3412 ^ 1'b0 ;
  assign n16423 = n16420 & n16422 ;
  assign n16427 = n7268 ^ n6977 ^ 1'b0 ;
  assign n16426 = n7312 ^ n5464 ^ n4707 ;
  assign n16424 = n15324 ^ n9619 ^ 1'b0 ;
  assign n16425 = n12331 & ~n16424 ;
  assign n16428 = n16427 ^ n16426 ^ n16425 ;
  assign n16429 = n16428 ^ n5077 ^ n1321 ;
  assign n16433 = n6688 ^ n2212 ^ 1'b0 ;
  assign n16434 = ~n6848 & n16433 ;
  assign n16435 = ~n1959 & n16434 ;
  assign n16430 = n718 & ~n11275 ;
  assign n16431 = n10281 | n16430 ;
  assign n16432 = n16431 ^ n1511 ^ 1'b0 ;
  assign n16436 = n16435 ^ n16432 ^ n2519 ;
  assign n16437 = n9565 ^ n4096 ^ 1'b0 ;
  assign n16438 = n8555 & n16437 ;
  assign n16439 = n15162 ^ n8669 ^ 1'b0 ;
  assign n16440 = n12364 & n16439 ;
  assign n16441 = n6588 ^ n4084 ^ n3480 ;
  assign n16442 = n4246 ^ n3673 ^ n1284 ;
  assign n16443 = n4561 ^ n3916 ^ 1'b0 ;
  assign n16444 = ( x78 & ~n16442 ) | ( x78 & n16443 ) | ( ~n16442 & n16443 ) ;
  assign n16445 = ( n612 & n5223 ) | ( n612 & n16444 ) | ( n5223 & n16444 ) ;
  assign n16454 = ~n4612 & n4948 ;
  assign n16447 = n5352 & ~n7489 ;
  assign n16448 = ~n5352 & n16447 ;
  assign n16449 = n16448 ^ n403 ^ 1'b0 ;
  assign n16450 = ~n439 & n1006 ;
  assign n16451 = n439 & n16450 ;
  assign n16452 = n16449 | n16451 ;
  assign n16453 = n16449 & ~n16452 ;
  assign n16446 = n12281 ^ n8983 ^ 1'b0 ;
  assign n16455 = n16454 ^ n16453 ^ n16446 ;
  assign n16456 = n4213 & ~n11502 ;
  assign n16457 = ~n16455 & n16456 ;
  assign n16458 = n2463 | n4552 ;
  assign n16459 = n13057 ^ n12374 ^ n5144 ;
  assign n16460 = n12098 ^ n11079 ^ 1'b0 ;
  assign n16461 = n2833 | n16460 ;
  assign n16462 = n13243 | n16461 ;
  assign n16463 = n4026 & ~n16462 ;
  assign n16464 = n15490 ^ n13659 ^ 1'b0 ;
  assign n16465 = n16463 | n16464 ;
  assign n16469 = n1973 | n11847 ;
  assign n16466 = n11905 ^ n9268 ^ 1'b0 ;
  assign n16467 = n11457 | n16466 ;
  assign n16468 = n3351 & ~n16467 ;
  assign n16470 = n16469 ^ n16468 ^ 1'b0 ;
  assign n16471 = n12411 ^ n2554 ^ 1'b0 ;
  assign n16472 = n11825 | n16471 ;
  assign n16473 = n16472 ^ n3882 ^ 1'b0 ;
  assign n16474 = n3102 & n16473 ;
  assign n16475 = n9830 ^ n8185 ^ n3373 ;
  assign n16476 = n10823 ^ n8036 ^ 1'b0 ;
  assign n16477 = n2927 | n16476 ;
  assign n16478 = n6661 ^ n5520 ^ 1'b0 ;
  assign n16479 = n13987 | n16478 ;
  assign n16480 = n14426 | n16479 ;
  assign n16481 = n422 & n7448 ;
  assign n16482 = n4294 & n16481 ;
  assign n16483 = n165 & n13884 ;
  assign n16484 = n4443 | n14665 ;
  assign n16485 = ( ~n2098 & n7022 ) | ( ~n2098 & n9489 ) | ( n7022 & n9489 ) ;
  assign n16486 = n16485 ^ n3413 ^ 1'b0 ;
  assign n16487 = n4216 | n16486 ;
  assign n16488 = n16487 ^ n890 ^ 1'b0 ;
  assign n16489 = n2438 ^ n1384 ^ 1'b0 ;
  assign n16490 = n8492 ^ n3058 ^ 1'b0 ;
  assign n16491 = n5945 | n16490 ;
  assign n16492 = x110 | n2169 ;
  assign n16493 = n16492 ^ n2800 ^ 1'b0 ;
  assign n16494 = ~n840 & n1353 ;
  assign n16495 = ~n630 & n13683 ;
  assign n16496 = n6927 & n11168 ;
  assign n16497 = n16496 ^ n6013 ^ 1'b0 ;
  assign n16498 = n3117 | n9450 ;
  assign n16499 = n8156 | n16498 ;
  assign n16500 = n16499 ^ n12943 ^ n10626 ;
  assign n16501 = n8308 ^ n1010 ^ n677 ;
  assign n16502 = n16500 & ~n16501 ;
  assign n16503 = n16156 ^ n8927 ^ 1'b0 ;
  assign n16504 = n5051 ^ x23 ^ 1'b0 ;
  assign n16505 = ( n190 & n620 ) | ( n190 & ~n16504 ) | ( n620 & ~n16504 ) ;
  assign n16506 = n8100 | n16505 ;
  assign n16507 = n5983 & ~n13265 ;
  assign n16508 = ~n2052 & n16507 ;
  assign n16509 = ( n980 & n5475 ) | ( n980 & ~n16508 ) | ( n5475 & ~n16508 ) ;
  assign n16510 = n16509 ^ n13865 ^ n13715 ;
  assign n16511 = n6288 ^ n5648 ^ 1'b0 ;
  assign n16512 = n9235 & n16511 ;
  assign n16513 = n16512 ^ n14084 ^ 1'b0 ;
  assign n16514 = n3712 & ~n16513 ;
  assign n16515 = n11329 | n16514 ;
  assign n16516 = n2706 ^ n427 ^ 1'b0 ;
  assign n16517 = n3143 ^ n1095 ^ 1'b0 ;
  assign n16518 = n16517 ^ n535 ^ 1'b0 ;
  assign n16519 = n15520 ^ n395 ^ 1'b0 ;
  assign n16520 = n16519 ^ n8296 ^ 1'b0 ;
  assign n16521 = ~n4123 & n15169 ;
  assign n16522 = n16520 & n16521 ;
  assign n16523 = n7703 ^ n2599 ^ 1'b0 ;
  assign n16524 = n16522 | n16523 ;
  assign n16525 = n4358 ^ n1781 ^ 1'b0 ;
  assign n16526 = n12722 & n16525 ;
  assign n16527 = n15062 ^ x116 ^ 1'b0 ;
  assign n16528 = n9349 ^ n4785 ^ n3972 ;
  assign n16529 = n2409 & ~n15226 ;
  assign n16530 = n16529 ^ n5063 ^ 1'b0 ;
  assign n16531 = ~n16528 & n16530 ;
  assign n16532 = n2805 | n3728 ;
  assign n16533 = n16532 ^ n5526 ^ 1'b0 ;
  assign n16534 = n16533 ^ n16245 ^ 1'b0 ;
  assign n16535 = n16230 & n16534 ;
  assign n16536 = ~n9542 & n16535 ;
  assign n16537 = n4850 ^ n4820 ^ 1'b0 ;
  assign n16538 = n12814 & n16537 ;
  assign n16539 = n16538 ^ n5840 ^ 1'b0 ;
  assign n16540 = n3946 & n8347 ;
  assign n16541 = n5791 & n7918 ;
  assign n16542 = n16541 ^ n892 ^ 1'b0 ;
  assign n16543 = n16542 ^ x80 ^ 1'b0 ;
  assign n16545 = n3124 & ~n4105 ;
  assign n16544 = ( n1010 & n4481 ) | ( n1010 & ~n9449 ) | ( n4481 & ~n9449 ) ;
  assign n16546 = n16545 ^ n16544 ^ n742 ;
  assign n16547 = n6381 | n8090 ;
  assign n16548 = n16547 ^ n14199 ^ 1'b0 ;
  assign n16549 = n11875 & n16548 ;
  assign n16550 = n8046 & n15565 ;
  assign n16551 = n12546 & n16550 ;
  assign n16552 = n7479 ^ n2316 ^ 1'b0 ;
  assign n16553 = ~n9092 & n16552 ;
  assign n16554 = ~n1184 & n16553 ;
  assign n16557 = n4097 & ~n4254 ;
  assign n16558 = n16557 ^ n6860 ^ 1'b0 ;
  assign n16555 = n691 & ~n8599 ;
  assign n16556 = ~n1130 & n16555 ;
  assign n16559 = n16558 ^ n16556 ^ n2845 ;
  assign n16560 = n14611 ^ n13167 ^ n3391 ;
  assign n16561 = n14194 ^ n6747 ^ 1'b0 ;
  assign n16562 = n4532 & n16561 ;
  assign n16563 = n6841 & ~n11172 ;
  assign n16564 = n16563 ^ n4394 ^ 1'b0 ;
  assign n16565 = n2200 ^ n1649 ^ 1'b0 ;
  assign n16566 = n7467 | n7520 ;
  assign n16567 = n16566 ^ n553 ^ 1'b0 ;
  assign n16568 = ~n6819 & n16567 ;
  assign n16569 = n1143 | n13679 ;
  assign n16570 = n1324 | n16569 ;
  assign n16571 = n16332 ^ n305 ^ 1'b0 ;
  assign n16572 = ~n4361 & n16571 ;
  assign n16573 = n9765 ^ n6251 ^ 1'b0 ;
  assign n16574 = ~n6146 & n16573 ;
  assign n16576 = n8496 ^ n1482 ^ 1'b0 ;
  assign n16577 = n12577 | n16576 ;
  assign n16575 = n6781 & n13403 ;
  assign n16578 = n16577 ^ n16575 ^ 1'b0 ;
  assign n16579 = ( ~n2824 & n3228 ) | ( ~n2824 & n10583 ) | ( n3228 & n10583 ) ;
  assign n16581 = n11550 ^ n6102 ^ 1'b0 ;
  assign n16582 = ~n10248 & n16581 ;
  assign n16583 = n16582 ^ n1791 ^ n1758 ;
  assign n16580 = n1462 | n7758 ;
  assign n16584 = n16583 ^ n16580 ^ n14511 ;
  assign n16585 = ( ~n1484 & n1840 ) | ( ~n1484 & n15801 ) | ( n1840 & n15801 ) ;
  assign n16586 = n3151 | n15519 ;
  assign n16587 = n16585 & ~n16586 ;
  assign n16588 = n7723 & n7962 ;
  assign n16589 = n16588 ^ n6131 ^ 1'b0 ;
  assign n16590 = n6517 ^ n247 ^ 1'b0 ;
  assign n16591 = n11460 & n16590 ;
  assign n16592 = n13596 ^ n1953 ^ 1'b0 ;
  assign n16596 = n551 & ~n670 ;
  assign n16597 = n670 & n16596 ;
  assign n16598 = n671 & ~n16597 ;
  assign n16593 = n2720 | n14340 ;
  assign n16594 = n14340 & ~n16593 ;
  assign n16595 = n2755 | n16594 ;
  assign n16599 = n16598 ^ n16595 ^ n3849 ;
  assign n16600 = n7553 ^ n2447 ^ 1'b0 ;
  assign n16601 = n10738 & n16600 ;
  assign n16602 = n12360 ^ n355 ^ 1'b0 ;
  assign n16603 = ( n16599 & n16601 ) | ( n16599 & n16602 ) | ( n16601 & n16602 ) ;
  assign n16604 = n1708 & n13104 ;
  assign n16605 = n16604 ^ n9507 ^ 1'b0 ;
  assign n16606 = n6075 | n6834 ;
  assign n16607 = n15320 ^ n14673 ^ 1'b0 ;
  assign n16608 = n4844 & ~n16607 ;
  assign n16609 = n16608 ^ n962 ^ 1'b0 ;
  assign n16610 = n8505 & n16609 ;
  assign n16611 = ~n8929 & n16610 ;
  assign n16612 = n1461 | n9204 ;
  assign n16613 = n11085 & ~n16612 ;
  assign n16614 = n3232 | n16613 ;
  assign n16615 = n16614 ^ n13112 ^ 1'b0 ;
  assign n16616 = n1944 & ~n13349 ;
  assign n16617 = n10202 & n16616 ;
  assign n16618 = n1525 & ~n9474 ;
  assign n16619 = n16618 ^ n2980 ^ 1'b0 ;
  assign n16620 = n16619 ^ n4916 ^ n4347 ;
  assign n16621 = n3513 ^ n707 ^ 1'b0 ;
  assign n16622 = n15164 | n16621 ;
  assign n16623 = n132 & ~n16622 ;
  assign n16624 = n5314 ^ n2206 ^ 1'b0 ;
  assign n16627 = n9868 & n10619 ;
  assign n16625 = n7839 ^ n5123 ^ 1'b0 ;
  assign n16626 = n11600 & ~n16625 ;
  assign n16628 = n16627 ^ n16626 ^ 1'b0 ;
  assign n16629 = n16628 ^ n12344 ^ 1'b0 ;
  assign n16630 = ( n1636 & ~n10293 ) | ( n1636 & n12179 ) | ( ~n10293 & n12179 ) ;
  assign n16631 = n14600 | n16630 ;
  assign n16632 = n7709 | n16631 ;
  assign n16633 = n4104 & ~n4207 ;
  assign n16634 = n11227 ^ n6482 ^ n5487 ;
  assign n16635 = n11704 ^ n9923 ^ 1'b0 ;
  assign n16636 = n16634 & ~n16635 ;
  assign n16637 = n4419 ^ n3835 ^ 1'b0 ;
  assign n16638 = n16636 & ~n16637 ;
  assign n16639 = ( n1530 & n3758 ) | ( n1530 & ~n6117 ) | ( n3758 & ~n6117 ) ;
  assign n16640 = n8624 | n9008 ;
  assign n16641 = n307 & n7705 ;
  assign n16642 = ~n1017 & n8684 ;
  assign n16643 = n16642 ^ n899 ^ 1'b0 ;
  assign n16644 = n16641 & ~n16643 ;
  assign n16645 = n12021 & n16644 ;
  assign n16646 = ~n13203 & n13765 ;
  assign n16647 = n10306 | n16646 ;
  assign n16650 = ~n3169 & n7899 ;
  assign n16648 = n16329 ^ n1362 ^ 1'b0 ;
  assign n16649 = n12496 | n16648 ;
  assign n16651 = n16650 ^ n16649 ^ 1'b0 ;
  assign n16652 = n1029 & ~n1955 ;
  assign n16653 = n16652 ^ n1451 ^ 1'b0 ;
  assign n16654 = n788 & n8140 ;
  assign n16655 = ~n2028 & n16654 ;
  assign n16656 = n5906 ^ n4481 ^ 1'b0 ;
  assign n16658 = n4039 ^ n1677 ^ 1'b0 ;
  assign n16657 = ~n5752 & n15561 ;
  assign n16659 = n16658 ^ n16657 ^ 1'b0 ;
  assign n16660 = n11549 ^ n1154 ^ 1'b0 ;
  assign n16662 = n5297 & ~n12407 ;
  assign n16663 = n10089 | n16662 ;
  assign n16664 = n1614 | n16663 ;
  assign n16661 = n12205 ^ n8354 ^ n8252 ;
  assign n16665 = n16664 ^ n16661 ^ 1'b0 ;
  assign n16666 = n12665 ^ n1933 ^ 1'b0 ;
  assign n16667 = ~n4855 & n11320 ;
  assign n16668 = n691 & ~n16667 ;
  assign n16669 = n16666 & n16668 ;
  assign n16670 = n5911 & n6330 ;
  assign n16671 = n15182 & n16670 ;
  assign n16672 = n2079 & n4847 ;
  assign n16673 = n422 & ~n8187 ;
  assign n16674 = n8676 & n16673 ;
  assign n16675 = n14861 | n16674 ;
  assign n16676 = n16675 ^ n1420 ^ 1'b0 ;
  assign n16677 = n16672 & ~n16676 ;
  assign n16678 = n7502 | n16677 ;
  assign n16679 = n16678 ^ n14008 ^ 1'b0 ;
  assign n16680 = n7663 & n12474 ;
  assign n16681 = n16680 ^ n4839 ^ 1'b0 ;
  assign n16682 = n15378 ^ n937 ^ 1'b0 ;
  assign n16683 = n14244 & n16682 ;
  assign n16684 = n745 | n5682 ;
  assign n16685 = n16684 ^ n3953 ^ 1'b0 ;
  assign n16686 = ( ~n867 & n1175 ) | ( ~n867 & n3167 ) | ( n1175 & n3167 ) ;
  assign n16687 = n3340 & ~n16686 ;
  assign n16688 = ~n5767 & n16687 ;
  assign n16689 = n6135 ^ n1286 ^ 1'b0 ;
  assign n16690 = n323 & n16689 ;
  assign n16691 = n9015 & n16690 ;
  assign n16694 = ~x6 & n2041 ;
  assign n16692 = n2951 & n4000 ;
  assign n16693 = n6393 & n16692 ;
  assign n16695 = n16694 ^ n16693 ^ n10293 ;
  assign n16696 = n1212 & n13554 ;
  assign n16697 = ~n10990 & n16696 ;
  assign n16698 = ( ~n4297 & n16695 ) | ( ~n4297 & n16697 ) | ( n16695 & n16697 ) ;
  assign n16699 = n9247 ^ n6436 ^ 1'b0 ;
  assign n16700 = n4443 | n15737 ;
  assign n16701 = n16700 ^ n3829 ^ 1'b0 ;
  assign n16702 = n4957 | n13520 ;
  assign n16703 = n16702 ^ n3703 ^ 1'b0 ;
  assign n16704 = n1106 & ~n3169 ;
  assign n16705 = n4964 | n16704 ;
  assign n16706 = n16003 ^ n10597 ^ 1'b0 ;
  assign n16707 = n16706 ^ n2519 ^ n1368 ;
  assign n16708 = n4653 & ~n16707 ;
  assign n16709 = n8526 ^ n8206 ^ 1'b0 ;
  assign n16710 = n11475 ^ n367 ^ 1'b0 ;
  assign n16711 = n16709 & n16710 ;
  assign n16712 = n16711 ^ n9574 ^ 1'b0 ;
  assign n16713 = ~n1452 & n5183 ;
  assign n16714 = n16713 ^ n6631 ^ 1'b0 ;
  assign n16715 = n16714 ^ n7081 ^ 1'b0 ;
  assign n16716 = n5444 ^ n1856 ^ 1'b0 ;
  assign n16717 = n145 & n16716 ;
  assign n16718 = n8160 ^ n1654 ^ 1'b0 ;
  assign n16719 = ~n5747 & n16718 ;
  assign n16720 = n13247 & n16719 ;
  assign n16721 = n16062 & n16720 ;
  assign n16722 = n9776 | n16721 ;
  assign n16723 = n11308 ^ n4962 ^ n547 ;
  assign n16724 = ~n881 & n4925 ;
  assign n16725 = n16724 ^ n4610 ^ 1'b0 ;
  assign n16726 = x35 & ~n6570 ;
  assign n16727 = n16725 & n16726 ;
  assign n16728 = n5410 ^ n2209 ^ 1'b0 ;
  assign n16729 = n9137 ^ n2693 ^ 1'b0 ;
  assign n16730 = n16728 & n16729 ;
  assign n16731 = n4780 ^ n4671 ^ 1'b0 ;
  assign n16732 = n4156 & ~n16731 ;
  assign n16733 = n16732 ^ n2839 ^ n1479 ;
  assign n16734 = n10700 ^ n7488 ^ 1'b0 ;
  assign n16735 = n16734 ^ n5680 ^ 1'b0 ;
  assign n16736 = n16733 | n16735 ;
  assign n16737 = n8075 & ~n16736 ;
  assign n16738 = n2638 ^ n236 ^ 1'b0 ;
  assign n16739 = n16738 ^ n8331 ^ 1'b0 ;
  assign n16740 = n4698 & ~n16739 ;
  assign n16741 = n5808 & ~n8341 ;
  assign n16742 = n7984 & n16741 ;
  assign n16743 = ~n1638 & n16742 ;
  assign n16744 = n16743 ^ n7701 ^ x70 ;
  assign n16748 = n1120 | n3152 ;
  assign n16745 = n1205 | n1677 ;
  assign n16746 = n1103 & ~n6337 ;
  assign n16747 = ~n16745 & n16746 ;
  assign n16749 = n16748 ^ n16747 ^ n9305 ;
  assign n16750 = ( n10704 & ~n15477 ) | ( n10704 & n16100 ) | ( ~n15477 & n16100 ) ;
  assign n16751 = n4545 ^ n1758 ^ 1'b0 ;
  assign n16752 = n8401 | n13323 ;
  assign n16753 = n2266 & ~n16752 ;
  assign n16754 = n10478 ^ n3738 ^ 1'b0 ;
  assign n16755 = ( n4581 & n6464 ) | ( n4581 & n7789 ) | ( n6464 & n7789 ) ;
  assign n16756 = n16755 ^ n2345 ^ 1'b0 ;
  assign n16757 = ~n16754 & n16756 ;
  assign n16758 = n16757 ^ n4342 ^ 1'b0 ;
  assign n16759 = n11799 & n16758 ;
  assign n16760 = n3989 & n16759 ;
  assign n16761 = n7127 & n16760 ;
  assign n16762 = ~n1157 & n7801 ;
  assign n16763 = ~n188 & n16762 ;
  assign n16764 = n7421 & ~n16763 ;
  assign n16765 = n16764 ^ n373 ^ 1'b0 ;
  assign n16766 = n3408 & ~n16765 ;
  assign n16767 = n6830 & n16766 ;
  assign n16768 = n16767 ^ n15629 ^ n13660 ;
  assign n16769 = ( n1452 & ~n1674 ) | ( n1452 & n2492 ) | ( ~n1674 & n2492 ) ;
  assign n16770 = n12897 ^ n7514 ^ 1'b0 ;
  assign n16771 = n16769 | n16770 ;
  assign n16772 = n12827 ^ n3426 ^ 1'b0 ;
  assign n16773 = ~n5747 & n16772 ;
  assign n16774 = n5013 ^ n1489 ^ n463 ;
  assign n16775 = n16774 ^ n1734 ^ 1'b0 ;
  assign n16776 = n16773 | n16775 ;
  assign n16777 = n1197 | n12494 ;
  assign n16778 = n3786 & ~n16777 ;
  assign n16779 = n7787 | n16778 ;
  assign n16780 = n9223 | n16779 ;
  assign n16781 = n6459 & n16780 ;
  assign n16782 = ~n16776 & n16781 ;
  assign n16783 = n12298 ^ n8500 ^ 1'b0 ;
  assign n16784 = n590 | n11761 ;
  assign n16785 = ~n601 & n6333 ;
  assign n16786 = ~n12472 & n16785 ;
  assign n16787 = n15284 & ~n16786 ;
  assign n16788 = n16787 ^ n11384 ^ 1'b0 ;
  assign n16789 = n15033 ^ n1036 ^ 1'b0 ;
  assign n16790 = ( n6532 & n13124 ) | ( n6532 & ~n16789 ) | ( n13124 & ~n16789 ) ;
  assign n16791 = n16790 ^ n11786 ^ n3644 ;
  assign n16793 = ~n5633 & n14083 ;
  assign n16792 = ~n2864 & n3755 ;
  assign n16794 = n16793 ^ n16792 ^ 1'b0 ;
  assign n16803 = n6161 & n9014 ;
  assign n16804 = n16601 & n16803 ;
  assign n16805 = n16804 ^ n6866 ^ 1'b0 ;
  assign n16806 = ~n12157 & n16805 ;
  assign n16799 = n3567 | n12895 ;
  assign n16800 = n13827 & ~n16799 ;
  assign n16795 = n4466 & n13172 ;
  assign n16796 = n6087 & ~n13197 ;
  assign n16797 = ~n11790 & n16796 ;
  assign n16798 = n16795 | n16797 ;
  assign n16801 = n16800 ^ n16798 ^ 1'b0 ;
  assign n16802 = n1054 | n16801 ;
  assign n16807 = n16806 ^ n16802 ^ 1'b0 ;
  assign n16808 = n2069 & n6790 ;
  assign n16809 = n1694 ^ n1484 ^ 1'b0 ;
  assign n16810 = n16808 & n16809 ;
  assign n16811 = n15538 ^ n4622 ^ 1'b0 ;
  assign n16812 = n16810 & ~n16811 ;
  assign n16813 = n9738 ^ n2654 ^ 1'b0 ;
  assign n16814 = n1971 & n16813 ;
  assign n16815 = n16426 ^ n6649 ^ 1'b0 ;
  assign n16816 = n16814 & n16815 ;
  assign n16817 = ~n12819 & n16816 ;
  assign n16818 = n1484 ^ n1103 ^ n592 ;
  assign n16819 = n1639 | n4000 ;
  assign n16820 = n16818 | n16819 ;
  assign n16821 = ( n706 & n16817 ) | ( n706 & ~n16820 ) | ( n16817 & ~n16820 ) ;
  assign n16822 = n3479 & n10340 ;
  assign n16823 = n3083 & ~n6866 ;
  assign n16824 = n16823 ^ n7383 ^ 1'b0 ;
  assign n16825 = ~x27 & n4916 ;
  assign n16826 = n2657 | n16825 ;
  assign n16827 = n16826 ^ n2979 ^ 1'b0 ;
  assign n16828 = ~n4964 & n10095 ;
  assign n16829 = n11167 & n16828 ;
  assign n16830 = ~n2142 & n5503 ;
  assign n16831 = ~x73 & n5356 ;
  assign n16832 = n16831 ^ n3916 ^ 1'b0 ;
  assign n16833 = n8178 ^ n5641 ^ n5207 ;
  assign n16834 = n1484 | n7613 ;
  assign n16835 = n418 & ~n16834 ;
  assign n16836 = n16835 ^ n12702 ^ 1'b0 ;
  assign n16837 = n16433 & ~n16836 ;
  assign n16838 = n12964 ^ n4895 ^ 1'b0 ;
  assign n16839 = n567 & ~n16838 ;
  assign n16840 = ~n3816 & n3994 ;
  assign n16841 = n750 & n16840 ;
  assign n16842 = n11444 ^ n7555 ^ n7415 ;
  assign n16843 = n13700 & n16842 ;
  assign n16849 = n8627 ^ n7920 ^ 1'b0 ;
  assign n16844 = n8790 ^ n6248 ^ n1319 ;
  assign n16845 = n3529 & n16844 ;
  assign n16846 = n16845 ^ n4632 ^ 1'b0 ;
  assign n16847 = n5369 & n16846 ;
  assign n16848 = n16847 ^ n10202 ^ 1'b0 ;
  assign n16850 = n16849 ^ n16848 ^ 1'b0 ;
  assign n16851 = n7496 | n16850 ;
  assign n16852 = n12779 ^ x92 ^ 1'b0 ;
  assign n16853 = n6719 | n16852 ;
  assign n16854 = n14385 | n15798 ;
  assign n16855 = n16853 & ~n16854 ;
  assign n16856 = n582 ^ n418 ^ 1'b0 ;
  assign n16857 = n5749 | n16856 ;
  assign n16858 = n16857 ^ n220 ^ 1'b0 ;
  assign n16860 = n9591 ^ n8854 ^ n6522 ;
  assign n16861 = n5511 | n16860 ;
  assign n16859 = ~n1753 & n12485 ;
  assign n16862 = n16861 ^ n16859 ^ 1'b0 ;
  assign n16863 = n12024 ^ n8691 ^ 1'b0 ;
  assign n16864 = ( n2973 & ~n16862 ) | ( n2973 & n16863 ) | ( ~n16862 & n16863 ) ;
  assign n16865 = n12521 & n13695 ;
  assign n16866 = n16865 ^ x3 ^ 1'b0 ;
  assign n16867 = n909 | n3249 ;
  assign n16868 = n1422 & n3710 ;
  assign n16869 = n3148 & ~n16868 ;
  assign n16873 = n681 & ~n1860 ;
  assign n16874 = n16873 ^ n987 ^ 1'b0 ;
  assign n16875 = n11233 | n16874 ;
  assign n16876 = n16875 ^ n2087 ^ 1'b0 ;
  assign n16870 = ( n433 & ~n6739 ) | ( n433 & n7966 ) | ( ~n6739 & n7966 ) ;
  assign n16871 = n16870 ^ n5036 ^ 1'b0 ;
  assign n16872 = n245 & n16871 ;
  assign n16877 = n16876 ^ n16872 ^ n15801 ;
  assign n16880 = x66 & ~n4653 ;
  assign n16881 = n1573 & n16880 ;
  assign n16878 = n16689 ^ n3304 ^ 1'b0 ;
  assign n16879 = n11930 & n16878 ;
  assign n16882 = n16881 ^ n16879 ^ n10324 ;
  assign n16883 = n14201 ^ n8621 ^ n1929 ;
  assign n16884 = n7887 ^ n2229 ^ x94 ;
  assign n16885 = n984 | n16884 ;
  assign n16886 = n16885 ^ n7453 ^ 1'b0 ;
  assign n16887 = ~n11238 & n14976 ;
  assign n16888 = ~n16886 & n16887 ;
  assign n16889 = ~n6872 & n14788 ;
  assign n16890 = n16889 ^ n3450 ^ 1'b0 ;
  assign n16891 = n3648 | n13793 ;
  assign n16892 = n1412 | n12399 ;
  assign n16893 = n678 | n4195 ;
  assign n16894 = n16893 ^ n7665 ^ n5452 ;
  assign n16895 = n9296 & ~n15693 ;
  assign n16896 = n4713 & n16895 ;
  assign n16897 = n1036 & n16896 ;
  assign n16898 = n5376 & ~n9621 ;
  assign n16899 = n16898 ^ n4065 ^ 1'b0 ;
  assign n16900 = ( x10 & ~n2495 ) | ( x10 & n6808 ) | ( ~n2495 & n6808 ) ;
  assign n16901 = ( n2994 & ~n7116 ) | ( n2994 & n16709 ) | ( ~n7116 & n16709 ) ;
  assign n16902 = n12469 ^ n7589 ^ 1'b0 ;
  assign n16903 = n3393 | n5212 ;
  assign n16904 = n16903 ^ n16672 ^ 1'b0 ;
  assign n16905 = n10563 & n16904 ;
  assign n16906 = n12246 & n16905 ;
  assign n16907 = n1220 & n16906 ;
  assign n16908 = n190 | n7475 ;
  assign n16909 = n16908 ^ n2166 ^ 1'b0 ;
  assign n16910 = n1652 & n16909 ;
  assign n16911 = ~n16907 & n16910 ;
  assign n16912 = n3325 & ~n16911 ;
  assign n16914 = n13668 ^ n9666 ^ 1'b0 ;
  assign n16913 = n12499 | n14170 ;
  assign n16915 = n16914 ^ n16913 ^ 1'b0 ;
  assign n16916 = n16687 ^ n4374 ^ 1'b0 ;
  assign n16917 = n12428 ^ n10738 ^ 1'b0 ;
  assign n16918 = n8826 & ~n16917 ;
  assign n16919 = n9823 & n16918 ;
  assign n16920 = ~n15964 & n16919 ;
  assign n16921 = ~n1611 & n2888 ;
  assign n16922 = ~n1406 & n16921 ;
  assign n16923 = n16922 ^ n2329 ^ 1'b0 ;
  assign n16924 = n3625 | n13626 ;
  assign n16925 = n13959 ^ n3216 ^ 1'b0 ;
  assign n16926 = n4221 | n16925 ;
  assign n16927 = n16926 ^ n10439 ^ 1'b0 ;
  assign n16928 = ( n1008 & ~n1909 ) | ( n1008 & n16927 ) | ( ~n1909 & n16927 ) ;
  assign n16930 = ~n1017 & n1034 ;
  assign n16931 = n1784 & n16930 ;
  assign n16932 = n15742 ^ n8357 ^ 1'b0 ;
  assign n16933 = ~n16931 & n16932 ;
  assign n16929 = ~n4133 & n8915 ;
  assign n16934 = n16933 ^ n16929 ^ 1'b0 ;
  assign n16935 = n11813 | n14170 ;
  assign n16936 = n14639 ^ n9364 ^ 1'b0 ;
  assign n16937 = n6007 ^ n3429 ^ 1'b0 ;
  assign n16938 = n7727 & ~n16937 ;
  assign n16939 = n16938 ^ n7707 ^ 1'b0 ;
  assign n16940 = ( n2510 & n9484 ) | ( n2510 & ~n9647 ) | ( n9484 & ~n9647 ) ;
  assign n16941 = ( n2706 & n14415 ) | ( n2706 & n16940 ) | ( n14415 & n16940 ) ;
  assign n16942 = n16941 ^ n4927 ^ 1'b0 ;
  assign n16943 = n3037 | n7774 ;
  assign n16944 = n16943 ^ n3282 ^ 1'b0 ;
  assign n16945 = n12185 ^ n1528 ^ 1'b0 ;
  assign n16946 = n16944 & n16945 ;
  assign n16947 = n12339 ^ n876 ^ 1'b0 ;
  assign n16948 = x64 & ~n16947 ;
  assign n16949 = n5221 ^ n1711 ^ 1'b0 ;
  assign n16950 = n10542 ^ n5421 ^ 1'b0 ;
  assign n16951 = ~n337 & n13297 ;
  assign n16952 = n16951 ^ n9564 ^ 1'b0 ;
  assign n16953 = n16679 & ~n16952 ;
  assign n16954 = n10990 ^ n7032 ^ 1'b0 ;
  assign n16955 = ~n16671 & n16954 ;
  assign n16956 = n190 & n3767 ;
  assign n16957 = n7040 ^ n4683 ^ 1'b0 ;
  assign n16958 = n7113 & n16957 ;
  assign n16959 = n16958 ^ n10502 ^ n3982 ;
  assign n16960 = n16959 ^ n2155 ^ 1'b0 ;
  assign n16961 = ( n4204 & ~n6614 ) | ( n4204 & n16960 ) | ( ~n6614 & n16960 ) ;
  assign n16962 = ~n7165 & n9156 ;
  assign n16963 = n16962 ^ n4187 ^ 1'b0 ;
  assign n16964 = ( n3826 & n7075 ) | ( n3826 & ~n7575 ) | ( n7075 & ~n7575 ) ;
  assign n16965 = n10464 & n16964 ;
  assign n16966 = n12835 | n16235 ;
  assign n16967 = n16966 ^ n678 ^ 1'b0 ;
  assign n16968 = n3066 | n14544 ;
  assign n16969 = x74 | n16968 ;
  assign n16970 = n4767 ^ n4656 ^ x74 ;
  assign n16971 = n6633 | n8844 ;
  assign n16972 = n16971 ^ n12205 ^ 1'b0 ;
  assign n16973 = n15835 ^ n967 ^ 1'b0 ;
  assign n16974 = ~n5014 & n8611 ;
  assign n16975 = n16974 ^ n11014 ^ 1'b0 ;
  assign n16976 = n3574 & ~n12006 ;
  assign n16977 = n16976 ^ n5682 ^ 1'b0 ;
  assign n16978 = n16977 ^ n12022 ^ n2929 ;
  assign n16979 = n9966 ^ n3223 ^ 1'b0 ;
  assign n16980 = n16979 ^ n5531 ^ 1'b0 ;
  assign n16981 = n16980 ^ n11329 ^ n8259 ;
  assign n16982 = n2607 & n11421 ;
  assign n16983 = ~n399 & n10675 ;
  assign n16984 = n16983 ^ n6304 ^ n4946 ;
  assign n16985 = ~n11710 & n16984 ;
  assign n16986 = n7729 ^ n2309 ^ 1'b0 ;
  assign n16987 = n16360 ^ n4490 ^ 1'b0 ;
  assign n16988 = n2517 & n16987 ;
  assign n16989 = ( n1876 & n6700 ) | ( n1876 & ~n11270 ) | ( n6700 & ~n11270 ) ;
  assign n16990 = ~n5040 & n10738 ;
  assign n16991 = n16990 ^ n4037 ^ 1'b0 ;
  assign n16992 = n16991 ^ n2432 ^ n2260 ;
  assign n16993 = n2859 | n15808 ;
  assign n16994 = ( n13915 & n16992 ) | ( n13915 & ~n16993 ) | ( n16992 & ~n16993 ) ;
  assign n16995 = n8729 & n10134 ;
  assign n16996 = n6876 ^ n2768 ^ 1'b0 ;
  assign n16997 = n3376 & ~n16996 ;
  assign n16998 = ~n3055 & n16997 ;
  assign n16999 = n16998 ^ n7305 ^ 1'b0 ;
  assign n17000 = n5808 & n9322 ;
  assign n17001 = ~n9373 & n17000 ;
  assign n17002 = n2921 & n9134 ;
  assign n17003 = n12177 ^ n11382 ^ 1'b0 ;
  assign n17004 = n14953 ^ n13559 ^ 1'b0 ;
  assign n17005 = n3114 & n17004 ;
  assign n17006 = n11690 & n17005 ;
  assign n17007 = n17006 ^ n425 ^ 1'b0 ;
  assign n17008 = n7533 & n9209 ;
  assign n17009 = n8588 ^ n6771 ^ 1'b0 ;
  assign n17010 = n11745 ^ n4795 ^ n3838 ;
  assign n17011 = n11210 & ~n17010 ;
  assign n17012 = n13233 ^ n7002 ^ n6381 ;
  assign n17013 = n13733 ^ n8834 ^ n4297 ;
  assign n17014 = n11962 ^ n5101 ^ 1'b0 ;
  assign n17015 = n1293 & ~n17014 ;
  assign n17016 = n9189 ^ n282 ^ 1'b0 ;
  assign n17017 = n3353 & n17016 ;
  assign n17018 = n2651 & n17017 ;
  assign n17020 = n4025 & ~n4456 ;
  assign n17019 = n475 | n2133 ;
  assign n17021 = n17020 ^ n17019 ^ 1'b0 ;
  assign n17022 = ~n17018 & n17021 ;
  assign n17023 = n17022 ^ n3396 ^ 1'b0 ;
  assign n17024 = n651 | n3591 ;
  assign n17025 = n17024 ^ n14910 ^ 1'b0 ;
  assign n17026 = ~n3533 & n7090 ;
  assign n17027 = n9873 ^ n8361 ^ 1'b0 ;
  assign n17028 = n4033 & ~n17027 ;
  assign n17029 = n7284 ^ n1633 ^ 1'b0 ;
  assign n17030 = n2423 ^ n601 ^ 1'b0 ;
  assign n17031 = n3324 & n17030 ;
  assign n17032 = n17029 & n17031 ;
  assign n17033 = n8959 ^ n6068 ^ 1'b0 ;
  assign n17034 = n6428 ^ n3439 ^ 1'b0 ;
  assign n17035 = ~n6771 & n17034 ;
  assign n17036 = n17035 ^ n7089 ^ 1'b0 ;
  assign n17037 = n4553 & ~n17036 ;
  assign n17038 = n4451 & n17037 ;
  assign n17039 = n17038 ^ n3924 ^ 1'b0 ;
  assign n17040 = n12474 & ~n17039 ;
  assign n17041 = n11882 ^ n750 ^ 1'b0 ;
  assign n17042 = n6349 & n17041 ;
  assign n17043 = n17042 ^ n712 ^ 1'b0 ;
  assign n17044 = ~n6746 & n7842 ;
  assign n17045 = n3728 & ~n5997 ;
  assign n17046 = ~n17044 & n17045 ;
  assign n17047 = n1519 ^ n1473 ^ 1'b0 ;
  assign n17048 = n10660 & n17047 ;
  assign n17049 = n6279 ^ n4364 ^ 1'b0 ;
  assign n17050 = n479 & ~n4645 ;
  assign n17051 = ~n10376 & n17050 ;
  assign n17052 = n16704 & n17051 ;
  assign n17053 = n8336 ^ n2958 ^ 1'b0 ;
  assign n17054 = n1450 & ~n6850 ;
  assign n17055 = n17054 ^ n10437 ^ 1'b0 ;
  assign n17056 = n3216 & n10686 ;
  assign n17057 = n1813 & n17056 ;
  assign n17058 = n2222 | n17057 ;
  assign n17059 = ~n6211 & n17058 ;
  assign n17060 = n7191 & n17059 ;
  assign n17061 = n7666 & ~n17060 ;
  assign n17062 = n17061 ^ n9257 ^ 1'b0 ;
  assign n17063 = ( ~n3061 & n5600 ) | ( ~n3061 & n8382 ) | ( n5600 & n8382 ) ;
  assign n17074 = n210 | n700 ;
  assign n17076 = n17074 ^ n1675 ^ 1'b0 ;
  assign n17072 = n6681 ^ n840 ^ 1'b0 ;
  assign n17073 = n7124 | n17072 ;
  assign n17075 = n17074 ^ n17073 ^ n3979 ;
  assign n17077 = n17076 ^ n17075 ^ n15524 ;
  assign n17078 = n8534 & ~n17077 ;
  assign n17064 = n16216 ^ n7031 ^ 1'b0 ;
  assign n17065 = x37 & ~n17064 ;
  assign n17066 = ~n225 & n516 ;
  assign n17067 = ~n620 & n17066 ;
  assign n17068 = n17067 ^ n9752 ^ 1'b0 ;
  assign n17069 = n17065 & n17068 ;
  assign n17070 = n11882 | n12490 ;
  assign n17071 = n17069 | n17070 ;
  assign n17079 = n17078 ^ n17071 ^ n5697 ;
  assign n17080 = n3728 ^ n823 ^ 1'b0 ;
  assign n17081 = n17080 ^ n10692 ^ x96 ;
  assign n17083 = ( x97 & ~n8310 ) | ( x97 & n10716 ) | ( ~n8310 & n10716 ) ;
  assign n17082 = n11530 | n15609 ;
  assign n17084 = n17083 ^ n17082 ^ 1'b0 ;
  assign n17085 = n9503 & n17084 ;
  assign n17086 = n7064 & n17085 ;
  assign n17087 = n3148 | n7434 ;
  assign n17088 = n17087 ^ n452 ^ 1'b0 ;
  assign n17089 = ~n3638 & n9466 ;
  assign n17090 = n17088 & ~n17089 ;
  assign n17091 = n17090 ^ n10279 ^ 1'b0 ;
  assign n17092 = n7357 ^ n3158 ^ 1'b0 ;
  assign n17093 = n16277 ^ n11179 ^ 1'b0 ;
  assign n17094 = ( n1743 & n7585 ) | ( n1743 & ~n12210 ) | ( n7585 & ~n12210 ) ;
  assign n17095 = n4186 ^ x108 ^ 1'b0 ;
  assign n17096 = n8929 & ~n17095 ;
  assign n17097 = ( ~n1584 & n14089 ) | ( ~n1584 & n17096 ) | ( n14089 & n17096 ) ;
  assign n17098 = n3768 & ~n4660 ;
  assign n17099 = n15787 ^ n2694 ^ 1'b0 ;
  assign n17100 = n9674 ^ n6266 ^ 1'b0 ;
  assign n17101 = n17099 & ~n17100 ;
  assign n17102 = n2162 | n4087 ;
  assign n17103 = n6148 & n16914 ;
  assign n17104 = n6420 ^ n3662 ^ 1'b0 ;
  assign n17105 = n17104 ^ n5342 ^ 1'b0 ;
  assign n17106 = n17103 | n17105 ;
  assign n17107 = n17106 ^ n9459 ^ 1'b0 ;
  assign n17108 = n12318 ^ n3418 ^ 1'b0 ;
  assign n17109 = n10071 ^ x37 ^ 1'b0 ;
  assign n17110 = n5598 ^ n239 ^ 1'b0 ;
  assign n17111 = ( n4230 & ~n4714 ) | ( n4230 & n5084 ) | ( ~n4714 & n5084 ) ;
  assign n17112 = ( n9934 & ~n17110 ) | ( n9934 & n17111 ) | ( ~n17110 & n17111 ) ;
  assign n17113 = ( n5642 & n17109 ) | ( n5642 & ~n17112 ) | ( n17109 & ~n17112 ) ;
  assign n17114 = n15016 & n17113 ;
  assign n17115 = n11157 ^ n6905 ^ 1'b0 ;
  assign n17116 = n2383 | n17115 ;
  assign n17117 = n8443 & n14075 ;
  assign n17118 = n17117 ^ n3350 ^ 1'b0 ;
  assign n17119 = n10356 ^ n1143 ^ 1'b0 ;
  assign n17120 = n138 & n17119 ;
  assign n17121 = n16326 ^ n5897 ^ 1'b0 ;
  assign n17122 = n8994 ^ n8132 ^ 1'b0 ;
  assign n17123 = n1150 & n17122 ;
  assign n17124 = n3673 & n17123 ;
  assign n17125 = n17124 ^ n4233 ^ 1'b0 ;
  assign n17126 = n5960 & n9339 ;
  assign n17127 = n6301 & n17126 ;
  assign n17128 = ~n9823 & n10932 ;
  assign n17129 = n17127 & ~n17128 ;
  assign n17130 = n14826 ^ n11095 ^ 1'b0 ;
  assign n17131 = ~n17129 & n17130 ;
  assign n17132 = n6845 ^ n3563 ^ 1'b0 ;
  assign n17134 = n13021 ^ n6148 ^ 1'b0 ;
  assign n17135 = n2175 & n17134 ;
  assign n17136 = n5281 ^ n2451 ^ 1'b0 ;
  assign n17137 = n1387 | n17136 ;
  assign n17138 = n17135 | n17137 ;
  assign n17133 = n1981 & ~n3037 ;
  assign n17139 = n17138 ^ n17133 ^ 1'b0 ;
  assign n17140 = n980 & n9662 ;
  assign n17141 = n17140 ^ n9630 ^ 1'b0 ;
  assign n17142 = n10186 & ~n13483 ;
  assign n17143 = n15457 & n17142 ;
  assign n17144 = n7787 ^ n494 ^ 1'b0 ;
  assign n17145 = n2278 & ~n8582 ;
  assign n17146 = n3217 & n17145 ;
  assign n17147 = n17146 ^ n5434 ^ 1'b0 ;
  assign n17148 = n8492 ^ n4565 ^ 1'b0 ;
  assign n17149 = ( ~n141 & n725 ) | ( ~n141 & n17148 ) | ( n725 & n17148 ) ;
  assign n17150 = n3457 ^ n1403 ^ 1'b0 ;
  assign n17151 = n7960 | n17150 ;
  assign n17152 = n17151 ^ n16780 ^ n8153 ;
  assign n17153 = n14603 ^ n9866 ^ 1'b0 ;
  assign n17154 = n3727 | n17153 ;
  assign n17155 = n10742 ^ n10720 ^ n3785 ;
  assign n17156 = n14413 | n17155 ;
  assign n17157 = n16338 & ~n17156 ;
  assign n17158 = n10186 ^ n6866 ^ 1'b0 ;
  assign n17159 = n2947 & ~n17158 ;
  assign n17160 = ( n4734 & n14274 ) | ( n4734 & n17159 ) | ( n14274 & n17159 ) ;
  assign n17161 = n17160 ^ n14626 ^ 1'b0 ;
  assign n17162 = n6022 & ~n13914 ;
  assign n17163 = ~n4600 & n9840 ;
  assign n17164 = n17163 ^ n4667 ^ 1'b0 ;
  assign n17165 = ~n17162 & n17164 ;
  assign n17166 = n1103 & n5314 ;
  assign n17167 = n17166 ^ n12493 ^ 1'b0 ;
  assign n17168 = n17167 ^ n7844 ^ 1'b0 ;
  assign n17169 = ~n7075 & n9778 ;
  assign n17171 = ~n2692 & n2727 ;
  assign n17170 = n1506 & ~n1526 ;
  assign n17172 = n17171 ^ n17170 ^ 1'b0 ;
  assign n17173 = n9659 & n17172 ;
  assign n17174 = n17173 ^ n2588 ^ 1'b0 ;
  assign n17175 = n17174 ^ n7893 ^ n2198 ;
  assign n17176 = n403 & n2443 ;
  assign n17177 = ~n7214 & n17176 ;
  assign n17179 = n10592 ^ n3709 ^ 1'b0 ;
  assign n17178 = n10104 & n14215 ;
  assign n17180 = n17179 ^ n17178 ^ 1'b0 ;
  assign n17187 = n12853 ^ n4199 ^ 1'b0 ;
  assign n17188 = n5216 & n17187 ;
  assign n17185 = n3282 ^ n2069 ^ 1'b0 ;
  assign n17186 = n8437 & ~n17185 ;
  assign n17189 = n17188 ^ n17186 ^ 1'b0 ;
  assign n17181 = n9647 ^ n3036 ^ 1'b0 ;
  assign n17182 = n17181 ^ n12090 ^ 1'b0 ;
  assign n17183 = n2117 | n17182 ;
  assign n17184 = n4076 & ~n17183 ;
  assign n17190 = n17189 ^ n17184 ^ 1'b0 ;
  assign n17191 = n6905 ^ n3627 ^ n3076 ;
  assign n17192 = n6548 & ~n17191 ;
  assign n17193 = n4531 & ~n6333 ;
  assign n17194 = n1165 & ~n17055 ;
  assign n17195 = ~n5517 & n12943 ;
  assign n17196 = n14525 ^ n9096 ^ 1'b0 ;
  assign n17197 = n16096 ^ n14440 ^ 1'b0 ;
  assign n17198 = n5183 & n9634 ;
  assign n17199 = n9396 | n12081 ;
  assign n17200 = n10902 | n11811 ;
  assign n17201 = n15019 ^ n12157 ^ 1'b0 ;
  assign n17202 = ( n2607 & n2800 ) | ( n2607 & ~n4285 ) | ( n2800 & ~n4285 ) ;
  assign n17203 = ( n420 & ~n11423 ) | ( n420 & n17202 ) | ( ~n11423 & n17202 ) ;
  assign n17204 = n9681 & ~n10281 ;
  assign n17205 = ~n245 & n13135 ;
  assign n17206 = n706 & n6798 ;
  assign n17207 = n17206 ^ n10161 ^ 1'b0 ;
  assign n17208 = ~n15538 & n17207 ;
  assign n17209 = n4716 & n17208 ;
  assign n17210 = n6629 ^ n2077 ^ 1'b0 ;
  assign n17211 = n14641 ^ n6494 ^ 1'b0 ;
  assign n17212 = n5342 | n17211 ;
  assign n17213 = n16238 ^ n11577 ^ 1'b0 ;
  assign n17214 = n4939 & ~n17213 ;
  assign n17215 = n7225 & ~n9206 ;
  assign n17216 = ~n6571 & n17215 ;
  assign n17217 = n17216 ^ n11241 ^ 1'b0 ;
  assign n17218 = n11174 & n17217 ;
  assign n17219 = n8976 & ~n10204 ;
  assign n17220 = n6550 ^ n4820 ^ 1'b0 ;
  assign n17221 = n17219 & ~n17220 ;
  assign n17222 = n16666 ^ n8723 ^ 1'b0 ;
  assign n17223 = n3746 & ~n17222 ;
  assign n17228 = n451 & ~n2034 ;
  assign n17229 = n17228 ^ n11945 ^ 1'b0 ;
  assign n17230 = n5885 & ~n17229 ;
  assign n17224 = n1161 & n3828 ;
  assign n17225 = n2028 | n17224 ;
  assign n17226 = n13795 & ~n17225 ;
  assign n17227 = n12214 & n17226 ;
  assign n17231 = n17230 ^ n17227 ^ 1'b0 ;
  assign n17232 = n11391 ^ n3571 ^ 1'b0 ;
  assign n17233 = n5447 & n17232 ;
  assign n17234 = n9703 ^ n8792 ^ 1'b0 ;
  assign n17235 = n13367 | n17234 ;
  assign n17236 = n17235 ^ n2585 ^ 1'b0 ;
  assign n17237 = n15506 ^ n5314 ^ 1'b0 ;
  assign n17238 = n279 & ~n17237 ;
  assign n17239 = n12506 ^ n11609 ^ n9287 ;
  assign n17240 = ( n5190 & ~n10567 ) | ( n5190 & n17239 ) | ( ~n10567 & n17239 ) ;
  assign n17241 = n13666 ^ n10476 ^ n6791 ;
  assign n17242 = n8544 ^ n2440 ^ 1'b0 ;
  assign n17243 = n11794 ^ n4460 ^ 1'b0 ;
  assign n17244 = n6864 ^ n2440 ^ 1'b0 ;
  assign n17245 = n371 & ~n4913 ;
  assign n17246 = n4511 & n17245 ;
  assign n17247 = ( n5638 & ~n9216 ) | ( n5638 & n17246 ) | ( ~n9216 & n17246 ) ;
  assign n17248 = n17244 & n17247 ;
  assign n17249 = n4504 ^ n619 ^ 1'b0 ;
  assign n17250 = n8811 & n17249 ;
  assign n17251 = n6381 ^ n3785 ^ 1'b0 ;
  assign n17252 = n9470 ^ n6972 ^ 1'b0 ;
  assign n17253 = ( x51 & ~x80 ) | ( x51 & n17252 ) | ( ~x80 & n17252 ) ;
  assign n17254 = n14075 ^ n6684 ^ 1'b0 ;
  assign n17255 = n1046 & ~n17254 ;
  assign n17256 = ( ~n1396 & n9498 ) | ( ~n1396 & n17255 ) | ( n9498 & n17255 ) ;
  assign n17257 = ~n6990 & n17256 ;
  assign n17258 = ~n17035 & n17257 ;
  assign n17259 = n1781 & ~n3815 ;
  assign n17260 = n6575 & n7518 ;
  assign n17261 = n17260 ^ n2490 ^ 1'b0 ;
  assign n17262 = ( n11936 & n12881 ) | ( n11936 & ~n17261 ) | ( n12881 & ~n17261 ) ;
  assign n17263 = n11035 & n17262 ;
  assign n17264 = n17259 & n17263 ;
  assign n17266 = ( n4025 & n6010 ) | ( n4025 & ~n9339 ) | ( n6010 & ~n9339 ) ;
  assign n17265 = n5453 & n8287 ;
  assign n17267 = n17266 ^ n17265 ^ n16003 ;
  assign n17268 = n10853 & ~n13037 ;
  assign n17269 = ( n5695 & n7824 ) | ( n5695 & ~n13454 ) | ( n7824 & ~n13454 ) ;
  assign n17270 = n8248 & n17269 ;
  assign n17271 = n17270 ^ n2514 ^ n2249 ;
  assign n17272 = n6215 | n8587 ;
  assign n17273 = n2638 & n9574 ;
  assign n17274 = n10776 | n13805 ;
  assign n17275 = n4833 & ~n17274 ;
  assign n17276 = n676 & ~n1413 ;
  assign n17277 = n345 & ~n6097 ;
  assign n17278 = n3138 ^ x20 ^ 1'b0 ;
  assign n17279 = ~n8624 & n17278 ;
  assign n17280 = n10484 & n17279 ;
  assign n17281 = ~n4154 & n17280 ;
  assign n17284 = x113 & n673 ;
  assign n17285 = ~n2738 & n17284 ;
  assign n17282 = n12529 ^ n2863 ^ 1'b0 ;
  assign n17283 = n13336 | n17282 ;
  assign n17286 = n17285 ^ n17283 ^ 1'b0 ;
  assign n17287 = n1372 ^ n1319 ^ 1'b0 ;
  assign n17288 = n6295 & ~n14391 ;
  assign n17289 = n1721 & ~n10100 ;
  assign n17290 = n2259 | n17289 ;
  assign n17291 = n9649 | n17290 ;
  assign n17292 = n2391 & n14303 ;
  assign n17293 = ( ~n6201 & n10368 ) | ( ~n6201 & n17292 ) | ( n10368 & n17292 ) ;
  assign n17294 = n10234 ^ n1800 ^ 1'b0 ;
  assign n17295 = ~n13429 & n17294 ;
  assign n17297 = n5547 & n8040 ;
  assign n17296 = n2302 & n11781 ;
  assign n17298 = n17297 ^ n17296 ^ 1'b0 ;
  assign n17299 = ~n8548 & n9862 ;
  assign n17300 = n17299 ^ n2331 ^ 1'b0 ;
  assign n17301 = n7421 & ~n16664 ;
  assign n17302 = n2934 & ~n4907 ;
  assign n17303 = n5973 & n17302 ;
  assign n17304 = n387 & n594 ;
  assign n17305 = n7669 & n17304 ;
  assign n17306 = n9634 & ~n17305 ;
  assign n17307 = n6674 & n17306 ;
  assign n17308 = ( n2807 & ~n17303 ) | ( n2807 & n17307 ) | ( ~n17303 & n17307 ) ;
  assign n17309 = n2846 ^ n326 ^ 1'b0 ;
  assign n17310 = ( n571 & n4550 ) | ( n571 & n4839 ) | ( n4550 & n4839 ) ;
  assign n17311 = n15552 ^ n5097 ^ 1'b0 ;
  assign n17312 = ~n11474 & n14828 ;
  assign n17313 = ~n3028 & n17312 ;
  assign n17314 = n17313 ^ n9092 ^ n6311 ;
  assign n17315 = ( ~n2341 & n5495 ) | ( ~n2341 & n6200 ) | ( n5495 & n6200 ) ;
  assign n17316 = ~n17314 & n17315 ;
  assign n17317 = n15634 ^ n11251 ^ 1'b0 ;
  assign n17318 = ~n4485 & n12249 ;
  assign n17319 = n17318 ^ n4872 ^ 1'b0 ;
  assign n17320 = ~n13858 & n17319 ;
  assign n17321 = n2924 ^ n2878 ^ 1'b0 ;
  assign n17322 = n4470 & n9144 ;
  assign n17323 = ~n1724 & n17322 ;
  assign n17324 = ~n17321 & n17323 ;
  assign n17325 = n17324 ^ n11764 ^ n8132 ;
  assign n17326 = n7547 ^ n6778 ^ n4503 ;
  assign n17327 = n17326 ^ n13149 ^ x120 ;
  assign n17328 = n14088 ^ n1236 ^ 1'b0 ;
  assign n17329 = n2017 & n7247 ;
  assign n17330 = n632 & ~n10895 ;
  assign n17331 = n9489 & n17330 ;
  assign n17332 = n17329 | n17331 ;
  assign n17333 = n17332 ^ n3931 ^ 1'b0 ;
  assign n17334 = n210 | n13435 ;
  assign n17335 = n937 | n4369 ;
  assign n17336 = n10095 & n10662 ;
  assign n17337 = n17336 ^ n1688 ^ 1'b0 ;
  assign n17338 = n770 ^ n153 ^ 1'b0 ;
  assign n17339 = x13 | n17338 ;
  assign n17340 = ( ~n7238 & n12813 ) | ( ~n7238 & n17339 ) | ( n12813 & n17339 ) ;
  assign n17341 = n17340 ^ n12813 ^ 1'b0 ;
  assign n17342 = n6927 & n17341 ;
  assign n17343 = ~n17337 & n17342 ;
  assign n17344 = n17343 ^ n9475 ^ n9395 ;
  assign n17345 = n8378 & ~n16992 ;
  assign n17346 = n13948 ^ n6888 ^ n2770 ;
  assign n17347 = ( n9043 & n16280 ) | ( n9043 & ~n17346 ) | ( n16280 & ~n17346 ) ;
  assign n17348 = ~n16894 & n17347 ;
  assign n17349 = n17348 ^ n15306 ^ 1'b0 ;
  assign n17351 = ( n1594 & n5855 ) | ( n1594 & n5981 ) | ( n5855 & n5981 ) ;
  assign n17350 = n3343 & n14294 ;
  assign n17352 = n17351 ^ n17350 ^ 1'b0 ;
  assign n17353 = ( ~n978 & n2829 ) | ( ~n978 & n5009 ) | ( n2829 & n5009 ) ;
  assign n17354 = n17353 ^ n14214 ^ 1'b0 ;
  assign n17355 = n17352 & ~n17354 ;
  assign n17356 = n15592 ^ n14410 ^ 1'b0 ;
  assign n17357 = n17313 & n17356 ;
  assign n17358 = n13644 ^ n11523 ^ n11243 ;
  assign n17359 = n17358 ^ n12490 ^ n1080 ;
  assign n17360 = n11505 & ~n17359 ;
  assign n17361 = n17360 ^ n10799 ^ 1'b0 ;
  assign n17362 = n17361 ^ n11718 ^ n7109 ;
  assign n17363 = n15437 ^ n1217 ^ 1'b0 ;
  assign n17364 = n14032 & n17363 ;
  assign n17367 = n1899 ^ n175 ^ 1'b0 ;
  assign n17368 = n17367 ^ n1231 ^ n892 ;
  assign n17365 = n4404 ^ n280 ^ 1'b0 ;
  assign n17366 = n1276 & ~n17365 ;
  assign n17369 = n17368 ^ n17366 ^ 1'b0 ;
  assign n17370 = n6823 ^ n703 ^ 1'b0 ;
  assign n17371 = n17370 ^ n7479 ^ 1'b0 ;
  assign n17372 = ~n852 & n17371 ;
  assign n17373 = n2207 & n4810 ;
  assign n17374 = ~n1075 & n17373 ;
  assign n17375 = n17374 ^ n4271 ^ n1479 ;
  assign n17376 = ~n6204 & n9619 ;
  assign n17377 = ~n17375 & n17376 ;
  assign n17378 = n11380 ^ n1115 ^ 1'b0 ;
  assign n17379 = n17377 & ~n17378 ;
  assign n17380 = n11737 ^ n6959 ^ 1'b0 ;
  assign n17381 = n8939 & ~n17380 ;
  assign n17382 = n4405 & ~n13001 ;
  assign n17383 = n11859 ^ n3562 ^ 1'b0 ;
  assign n17384 = n17382 & ~n17383 ;
  assign n17385 = n17384 ^ n13432 ^ 1'b0 ;
  assign n17386 = n4364 ^ n2331 ^ 1'b0 ;
  assign n17387 = n218 & n6004 ;
  assign n17388 = n5328 & ~n13424 ;
  assign n17389 = n7090 | n17388 ;
  assign n17391 = n998 | n16979 ;
  assign n17392 = n17391 ^ n7919 ^ 1'b0 ;
  assign n17390 = n10446 ^ n9324 ^ n3562 ;
  assign n17393 = n17392 ^ n17390 ^ n16354 ;
  assign n17394 = n5314 & ~n6448 ;
  assign n17395 = n6410 & ~n9950 ;
  assign n17396 = n17395 ^ n5717 ^ 1'b0 ;
  assign n17397 = n11260 ^ n5874 ^ 1'b0 ;
  assign n17398 = n812 & ~n1412 ;
  assign n17399 = ~n6961 & n17398 ;
  assign n17400 = n8123 | n17399 ;
  assign n17401 = n17397 | n17400 ;
  assign n17402 = n1867 & ~n5882 ;
  assign n17403 = n17402 ^ n10790 ^ 1'b0 ;
  assign n17404 = n4770 | n5380 ;
  assign n17405 = n17404 ^ n3398 ^ 1'b0 ;
  assign n17406 = n461 | n1379 ;
  assign n17407 = n17406 ^ n14398 ^ n4806 ;
  assign n17408 = n3617 ^ n2108 ^ 1'b0 ;
  assign n17409 = n4783 ^ n2631 ^ 1'b0 ;
  assign n17410 = n15144 ^ n10265 ^ 1'b0 ;
  assign n17411 = ~n3014 & n8976 ;
  assign n17412 = n17411 ^ n4827 ^ 1'b0 ;
  assign n17413 = ~n4261 & n17412 ;
  assign n17417 = ~n2529 & n9703 ;
  assign n17418 = ~n9703 & n17417 ;
  assign n17414 = n2682 | n14704 ;
  assign n17415 = n14704 & ~n17414 ;
  assign n17416 = n5717 | n17415 ;
  assign n17419 = n17418 ^ n17416 ^ 1'b0 ;
  assign n17420 = n2351 & n8956 ;
  assign n17421 = n7434 & n17420 ;
  assign n17422 = ~n8226 & n17421 ;
  assign n17423 = n2723 ^ n2469 ^ 1'b0 ;
  assign n17425 = n17074 ^ n6760 ^ n3321 ;
  assign n17426 = ( ~n1198 & n8252 ) | ( ~n1198 & n17425 ) | ( n8252 & n17425 ) ;
  assign n17424 = n2875 & n12298 ;
  assign n17427 = n17426 ^ n17424 ^ 1'b0 ;
  assign n17428 = ( n5746 & n6199 ) | ( n5746 & n17427 ) | ( n6199 & n17427 ) ;
  assign n17429 = n6271 ^ n5419 ^ 1'b0 ;
  assign n17430 = n17429 ^ n4916 ^ 1'b0 ;
  assign n17431 = n14391 ^ n9094 ^ n8523 ;
  assign n17432 = n11581 & n12575 ;
  assign n17433 = n919 & n10597 ;
  assign n17434 = n2368 & ~n2705 ;
  assign n17435 = n17434 ^ n3380 ^ 1'b0 ;
  assign n17436 = n2341 | n5535 ;
  assign n17437 = n1503 | n17436 ;
  assign n17438 = n17437 ^ n5603 ^ 1'b0 ;
  assign n17439 = ~n17435 & n17438 ;
  assign n17443 = n2462 & n8099 ;
  assign n17444 = n13796 & ~n17443 ;
  assign n17445 = n17444 ^ x93 ^ 1'b0 ;
  assign n17440 = n10418 & ~n13765 ;
  assign n17441 = n17440 ^ n7989 ^ 1'b0 ;
  assign n17442 = ~n2259 & n17441 ;
  assign n17446 = n17445 ^ n17442 ^ 1'b0 ;
  assign n17447 = ( n145 & n10073 ) | ( n145 & n17446 ) | ( n10073 & n17446 ) ;
  assign n17448 = n2619 & ~n12683 ;
  assign n17449 = n17448 ^ n859 ^ 1'b0 ;
  assign n17450 = n17449 ^ n10138 ^ n6090 ;
  assign n17451 = n2569 | n17282 ;
  assign n17452 = ~n2098 & n11273 ;
  assign n17453 = n1520 & n17110 ;
  assign n17454 = n4697 & ~n17453 ;
  assign n17455 = n2331 | n17454 ;
  assign n17456 = n10394 & n17455 ;
  assign n17457 = n17452 & n17456 ;
  assign n17458 = n5892 & n7372 ;
  assign n17459 = x50 & ~n17458 ;
  assign n17460 = n3638 ^ n1920 ^ 1'b0 ;
  assign n17461 = ~n6201 & n17460 ;
  assign n17462 = n17461 ^ n8253 ^ n4605 ;
  assign n17463 = n17462 ^ n6436 ^ 1'b0 ;
  assign n17464 = n8212 | n17463 ;
  assign n17465 = n17459 | n17464 ;
  assign n17466 = n5347 | n9327 ;
  assign n17467 = x56 | n17466 ;
  assign n17468 = n6742 ^ n5971 ^ 1'b0 ;
  assign n17469 = n17467 & n17468 ;
  assign n17470 = n6041 | n7657 ;
  assign n17471 = n644 & ~n17470 ;
  assign n17472 = n17471 ^ n16630 ^ 1'b0 ;
  assign n17473 = n8349 ^ n8039 ^ n4865 ;
  assign n17474 = n17473 ^ n12917 ^ n6534 ;
  assign n17481 = n14639 ^ n1597 ^ 1'b0 ;
  assign n17475 = n8939 & n14915 ;
  assign n17476 = n17475 ^ n3329 ^ 1'b0 ;
  assign n17477 = n17476 ^ n2304 ^ 1'b0 ;
  assign n17478 = n10837 | n17477 ;
  assign n17479 = n17478 ^ n9013 ^ 1'b0 ;
  assign n17480 = n9251 & n17479 ;
  assign n17482 = n17481 ^ n17480 ^ n2594 ;
  assign n17483 = ~n11096 & n15869 ;
  assign n17484 = ~n13712 & n17483 ;
  assign n17486 = n3023 | n5952 ;
  assign n17487 = n17486 ^ n12964 ^ 1'b0 ;
  assign n17485 = n2953 & n4400 ;
  assign n17488 = n17487 ^ n17485 ^ 1'b0 ;
  assign n17489 = ~n5059 & n5507 ;
  assign n17490 = ( n8692 & n9327 ) | ( n8692 & ~n17489 ) | ( n9327 & ~n17489 ) ;
  assign n17491 = ( n2194 & n12301 ) | ( n2194 & ~n17490 ) | ( n12301 & ~n17490 ) ;
  assign n17492 = n2671 ^ n512 ^ 1'b0 ;
  assign n17493 = n7739 & n17492 ;
  assign n17494 = x1 | n4820 ;
  assign n17495 = n3435 | n4932 ;
  assign n17496 = n3435 & ~n17495 ;
  assign n17497 = n7160 & ~n17496 ;
  assign n17498 = ~n7160 & n17497 ;
  assign n17499 = n17494 | n17498 ;
  assign n17500 = n6135 & ~n17499 ;
  assign n17501 = ~n2666 & n3569 ;
  assign n17502 = n11676 | n17501 ;
  assign n17503 = ( n5655 & n12068 ) | ( n5655 & n14866 ) | ( n12068 & n14866 ) ;
  assign n17504 = n6450 ^ x3 ^ 1'b0 ;
  assign n17505 = n7420 | n9268 ;
  assign n17506 = n2688 | n17505 ;
  assign n17507 = n12893 | n17506 ;
  assign n17508 = n3919 ^ n497 ^ 1'b0 ;
  assign n17509 = n3966 & n17508 ;
  assign n17510 = n10993 ^ n5719 ^ n191 ;
  assign n17511 = ~n12379 & n17510 ;
  assign n17512 = ~n3137 & n12172 ;
  assign n17513 = ~n1924 & n3471 ;
  assign n17514 = ~n3639 & n17513 ;
  assign n17515 = n7206 & ~n17514 ;
  assign n17518 = n1915 & n2640 ;
  assign n17519 = ~n1919 & n17518 ;
  assign n17520 = ( n2670 & ~n7254 ) | ( n2670 & n17519 ) | ( ~n7254 & n17519 ) ;
  assign n17516 = ~n1781 & n7925 ;
  assign n17517 = ~n9900 & n17516 ;
  assign n17521 = n17520 ^ n17517 ^ 1'b0 ;
  assign n17522 = n3158 & n13713 ;
  assign n17523 = ~n14432 & n17522 ;
  assign n17524 = n12631 ^ n9229 ^ 1'b0 ;
  assign n17525 = n1392 ^ n903 ^ 1'b0 ;
  assign n17526 = n17525 ^ n7689 ^ 1'b0 ;
  assign n17527 = n2107 | n17526 ;
  assign n17528 = n3565 & n6557 ;
  assign n17529 = n17528 ^ n3216 ^ 1'b0 ;
  assign n17530 = x37 & n2750 ;
  assign n17531 = n9341 | n11079 ;
  assign n17532 = n17531 ^ n8576 ^ 1'b0 ;
  assign n17533 = n9950 ^ n7114 ^ 1'b0 ;
  assign n17534 = n10125 ^ n6227 ^ 1'b0 ;
  assign n17535 = n17533 | n17534 ;
  assign n17536 = n323 & n11799 ;
  assign n17537 = ~n6781 & n17536 ;
  assign n17538 = n2710 & ~n17537 ;
  assign n17539 = n13465 | n16360 ;
  assign n17540 = n16274 ^ n11412 ^ 1'b0 ;
  assign n17541 = ~n14231 & n17540 ;
  assign n17542 = n15488 ^ n13476 ^ n11696 ;
  assign n17543 = ( n5824 & n13291 ) | ( n5824 & ~n14052 ) | ( n13291 & ~n14052 ) ;
  assign n17544 = n6393 ^ n3503 ^ 1'b0 ;
  assign n17545 = n2634 | n17544 ;
  assign n17546 = n6450 | n17545 ;
  assign n17547 = n17546 ^ n11552 ^ n6187 ;
  assign n17548 = ( n2845 & n5879 ) | ( n2845 & n17547 ) | ( n5879 & n17547 ) ;
  assign n17549 = n6564 ^ n1803 ^ 1'b0 ;
  assign n17550 = n11432 & n17549 ;
  assign n17551 = n17550 ^ n6778 ^ 1'b0 ;
  assign n17552 = ~n7715 & n17551 ;
  assign n17553 = ~n17548 & n17552 ;
  assign n17554 = ~n3344 & n11750 ;
  assign n17555 = n1012 & ~n17554 ;
  assign n17556 = n9619 & n9953 ;
  assign n17557 = n17555 & n17556 ;
  assign n17558 = n5928 ^ n3694 ^ x124 ;
  assign n17559 = n17558 ^ n1599 ^ 1'b0 ;
  assign n17560 = n6094 & n17559 ;
  assign n17561 = ~n245 & n17560 ;
  assign n17562 = n17561 ^ n10551 ^ n4445 ;
  assign n17566 = n5267 ^ n3952 ^ n1815 ;
  assign n17563 = ~n7681 & n17188 ;
  assign n17564 = n17563 ^ n781 ^ 1'b0 ;
  assign n17565 = n17564 ^ n14486 ^ n11287 ;
  assign n17567 = n17566 ^ n17565 ^ 1'b0 ;
  assign n17568 = n17567 ^ n9786 ^ n4880 ;
  assign n17569 = n14884 ^ n10002 ^ 1'b0 ;
  assign n17570 = n3919 ^ n2254 ^ 1'b0 ;
  assign n17571 = n17570 ^ n7716 ^ 1'b0 ;
  assign n17573 = n1141 & n17074 ;
  assign n17572 = n2897 | n12536 ;
  assign n17574 = n17573 ^ n17572 ^ 1'b0 ;
  assign n17579 = n10980 ^ n320 ^ 1'b0 ;
  assign n17575 = n9703 ^ n5466 ^ n4008 ;
  assign n17576 = n7609 & ~n17575 ;
  assign n17577 = ~n6638 & n17576 ;
  assign n17578 = n12179 | n17577 ;
  assign n17580 = n17579 ^ n17578 ^ 1'b0 ;
  assign n17581 = n889 | n17580 ;
  assign n17582 = n17581 ^ n2860 ^ 1'b0 ;
  assign n17583 = n17574 & n17582 ;
  assign n17584 = ~n8353 & n17080 ;
  assign n17585 = n10440 & n17584 ;
  assign n17586 = n17585 ^ n10625 ^ 1'b0 ;
  assign n17587 = n2721 ^ n1587 ^ 1'b0 ;
  assign n17588 = n17587 ^ n2568 ^ 1'b0 ;
  assign n17589 = n927 & n7192 ;
  assign n17590 = n17589 ^ n8337 ^ 1'b0 ;
  assign n17591 = n17590 ^ n14459 ^ 1'b0 ;
  assign n17592 = n17588 | n17591 ;
  assign n17593 = n5203 | n6676 ;
  assign n17594 = ( n12132 & ~n15968 ) | ( n12132 & n17593 ) | ( ~n15968 & n17593 ) ;
  assign n17595 = n9656 ^ n7478 ^ 1'b0 ;
  assign n17596 = ~n6934 & n12771 ;
  assign n17597 = n5906 & n17596 ;
  assign n17598 = n1208 & ~n11877 ;
  assign n17599 = n17597 & n17598 ;
  assign n17600 = n3075 & n4450 ;
  assign n17601 = n17600 ^ n5618 ^ 1'b0 ;
  assign n17602 = n12328 & n17601 ;
  assign n17603 = n17602 ^ n10919 ^ 1'b0 ;
  assign n17604 = n3252 ^ n2453 ^ 1'b0 ;
  assign n17605 = n10357 ^ n9417 ^ n6428 ;
  assign n17606 = ~x22 & n17605 ;
  assign n17607 = n8230 ^ n3016 ^ 1'b0 ;
  assign n17608 = n17607 ^ n3547 ^ 1'b0 ;
  assign n17609 = n14422 & ~n17608 ;
  assign n17610 = ( n8865 & n11287 ) | ( n8865 & ~n17609 ) | ( n11287 & ~n17609 ) ;
  assign n17611 = n1396 & ~n4348 ;
  assign n17612 = n17611 ^ n6808 ^ 1'b0 ;
  assign n17618 = n10809 ^ n1754 ^ 1'b0 ;
  assign n17616 = ~n466 & n4047 ;
  assign n17613 = n1840 ^ n1089 ^ 1'b0 ;
  assign n17614 = n3163 | n17613 ;
  assign n17615 = n4059 & n17614 ;
  assign n17617 = n17616 ^ n17615 ^ 1'b0 ;
  assign n17619 = n17618 ^ n17617 ^ 1'b0 ;
  assign n17620 = n6384 & n17619 ;
  assign n17621 = n2209 & n5866 ;
  assign n17622 = ~n17326 & n17621 ;
  assign n17623 = n6148 ^ n2234 ^ 1'b0 ;
  assign n17624 = n8611 & n9457 ;
  assign n17625 = ~n10563 & n17624 ;
  assign n17626 = n17623 & ~n17625 ;
  assign n17627 = ( ~n2184 & n6124 ) | ( ~n2184 & n17626 ) | ( n6124 & n17626 ) ;
  assign n17628 = n7876 ^ n2053 ^ 1'b0 ;
  assign n17629 = n8367 | n17628 ;
  assign n17630 = n5944 | n17629 ;
  assign n17631 = ~n1877 & n3946 ;
  assign n17632 = n17631 ^ n9703 ^ 1'b0 ;
  assign n17633 = n12846 ^ n523 ^ 1'b0 ;
  assign n17634 = ~n17089 & n17633 ;
  assign n17635 = n17634 ^ n6506 ^ 1'b0 ;
  assign n17636 = n388 & n13293 ;
  assign n17637 = n11426 ^ x23 ^ 1'b0 ;
  assign n17638 = ( n3860 & n5098 ) | ( n3860 & ~n7210 ) | ( n5098 & ~n7210 ) ;
  assign n17639 = n17638 ^ n910 ^ 1'b0 ;
  assign n17640 = ~n2553 & n10604 ;
  assign n17641 = ( n753 & n3342 ) | ( n753 & n10740 ) | ( n3342 & n10740 ) ;
  assign n17642 = ( n4407 & ~n17640 ) | ( n4407 & n17641 ) | ( ~n17640 & n17641 ) ;
  assign n17643 = n4084 & ~n12897 ;
  assign n17644 = ~n676 & n17643 ;
  assign n17645 = n1362 | n17644 ;
  assign n17646 = n10495 | n17645 ;
  assign n17647 = n13697 & ~n17646 ;
  assign n17648 = n2853 ^ n614 ^ 1'b0 ;
  assign n17649 = n17648 ^ n8617 ^ 1'b0 ;
  assign n17650 = ~n6040 & n6206 ;
  assign n17651 = n17649 & n17650 ;
  assign n17652 = n15285 ^ n4574 ^ n1077 ;
  assign n17653 = ( ~n502 & n5798 ) | ( ~n502 & n8549 ) | ( n5798 & n8549 ) ;
  assign n17654 = n17653 ^ n7415 ^ n2590 ;
  assign n17655 = n10064 | n17654 ;
  assign n17656 = n6643 ^ n2652 ^ 1'b0 ;
  assign n17657 = n809 & ~n2637 ;
  assign n17658 = n17656 & ~n17657 ;
  assign n17659 = ~n3552 & n17658 ;
  assign n17660 = n1811 | n8722 ;
  assign n17661 = n17660 ^ x11 ^ 1'b0 ;
  assign n17662 = n17661 ^ n5353 ^ 1'b0 ;
  assign n17663 = n11629 | n17662 ;
  assign n17664 = n17663 ^ n403 ^ 1'b0 ;
  assign n17665 = n1347 | n5291 ;
  assign n17666 = n17665 ^ n5328 ^ 1'b0 ;
  assign n17667 = n17666 ^ n4047 ^ 1'b0 ;
  assign n17672 = n3615 ^ n2268 ^ 1'b0 ;
  assign n17673 = ~n163 & n17672 ;
  assign n17671 = n6876 ^ n5258 ^ 1'b0 ;
  assign n17669 = n3947 & n12548 ;
  assign n17668 = n4181 & n8024 ;
  assign n17670 = n17669 ^ n17668 ^ 1'b0 ;
  assign n17674 = n17673 ^ n17671 ^ n17670 ;
  assign n17675 = n12835 & n15928 ;
  assign n17679 = ~n1230 & n3061 ;
  assign n17680 = ~n3966 & n17679 ;
  assign n17681 = n2432 & n17680 ;
  assign n17682 = n13959 | n17681 ;
  assign n17683 = n9193 | n17682 ;
  assign n17676 = n3149 & n3560 ;
  assign n17677 = n5225 & n17676 ;
  assign n17678 = n13022 & ~n17677 ;
  assign n17684 = n17683 ^ n17678 ^ 1'b0 ;
  assign n17685 = n2661 | n7577 ;
  assign n17686 = n17685 ^ n12535 ^ 1'b0 ;
  assign n17687 = n17686 ^ n307 ^ 1'b0 ;
  assign n17688 = n746 & n3994 ;
  assign n17689 = n17687 & n17688 ;
  assign n17690 = ~n3151 & n17111 ;
  assign n17691 = n9896 & n17690 ;
  assign n17692 = n17691 ^ n17489 ^ n544 ;
  assign n17693 = n863 & ~n17692 ;
  assign n17694 = ~n3717 & n8753 ;
  assign n17697 = n577 & n7328 ;
  assign n17695 = n9158 & n17370 ;
  assign n17696 = ~n9158 & n17695 ;
  assign n17698 = n17697 ^ n17696 ^ 1'b0 ;
  assign n17699 = n2104 ^ n856 ^ 1'b0 ;
  assign n17700 = n173 & ~n6876 ;
  assign n17701 = ~n12074 & n17700 ;
  assign n17702 = ~n786 & n17701 ;
  assign n17703 = n17702 ^ n3456 ^ 1'b0 ;
  assign n17704 = n193 ^ x110 ^ 1'b0 ;
  assign n17705 = n17703 & ~n17704 ;
  assign n17706 = ( ~n355 & n17699 ) | ( ~n355 & n17705 ) | ( n17699 & n17705 ) ;
  assign n17707 = n8328 ^ n398 ^ 1'b0 ;
  assign n17708 = n14744 ^ n10134 ^ 1'b0 ;
  assign n17709 = n7111 & ~n17708 ;
  assign n17710 = n8981 ^ n6909 ^ 1'b0 ;
  assign n17711 = ~n171 & n17710 ;
  assign n17712 = ~n17709 & n17711 ;
  assign n17713 = n17712 ^ n4806 ^ 1'b0 ;
  assign n17714 = n17707 & ~n17713 ;
  assign n17715 = n1627 & ~n6893 ;
  assign n17716 = n2944 & n17715 ;
  assign n17717 = ( n15025 & n16145 ) | ( n15025 & ~n17687 ) | ( n16145 & ~n17687 ) ;
  assign n17718 = n2713 & ~n15822 ;
  assign n17719 = n15872 ^ n1286 ^ 1'b0 ;
  assign n17720 = ~n379 & n9894 ;
  assign n17721 = ( n6939 & ~n10480 ) | ( n6939 & n17616 ) | ( ~n10480 & n17616 ) ;
  assign n17722 = n11275 ^ n5826 ^ n3282 ;
  assign n17723 = n3396 | n4065 ;
  assign n17724 = n17723 ^ n9265 ^ 1'b0 ;
  assign n17725 = n17724 ^ n6532 ^ 1'b0 ;
  assign n17726 = n8160 & n17725 ;
  assign n17727 = n8249 & n17726 ;
  assign n17728 = ~n1462 & n6278 ;
  assign n17729 = n17728 ^ x86 ^ 1'b0 ;
  assign n17730 = ~n1113 & n1390 ;
  assign n17731 = n17730 ^ n4266 ^ n646 ;
  assign n17732 = n10522 | n17731 ;
  assign n17733 = n9158 ^ n886 ^ n332 ;
  assign n17734 = n3551 | n17733 ;
  assign n17735 = n1603 & ~n17734 ;
  assign n17736 = n17732 | n17735 ;
  assign n17737 = n17729 & ~n17736 ;
  assign n17738 = n3184 | n17737 ;
  assign n17739 = n5285 ^ n5283 ^ n2102 ;
  assign n17740 = ~n1713 & n17441 ;
  assign n17741 = ~n15624 & n17740 ;
  assign n17742 = n17741 ^ n8563 ^ 1'b0 ;
  assign n17743 = n2304 | n7207 ;
  assign n17744 = n8279 ^ n2143 ^ n1605 ;
  assign n17745 = n17744 ^ n9339 ^ 1'b0 ;
  assign n17746 = ~n1784 & n17745 ;
  assign n17747 = ~n1879 & n15634 ;
  assign n17748 = ~n4560 & n17747 ;
  assign n17749 = n10901 ^ n5480 ^ 1'b0 ;
  assign n17750 = ( n2266 & n9216 ) | ( n2266 & ~n17749 ) | ( n9216 & ~n17749 ) ;
  assign n17751 = n5521 ^ n177 ^ 1'b0 ;
  assign n17752 = ( n881 & n8763 ) | ( n881 & n13910 ) | ( n8763 & n13910 ) ;
  assign n17753 = n9092 ^ n1079 ^ 1'b0 ;
  assign n17754 = n16903 & ~n17753 ;
  assign n17755 = ~n4932 & n17754 ;
  assign n17756 = n917 & n17755 ;
  assign n17757 = ( n6003 & n8667 ) | ( n6003 & n17756 ) | ( n8667 & n17756 ) ;
  assign n17758 = n1930 | n7576 ;
  assign n17759 = n8100 | n17758 ;
  assign n17760 = n17759 ^ n11404 ^ 1'b0 ;
  assign n17761 = n7143 ^ n5152 ^ 1'b0 ;
  assign n17762 = n16336 | n17761 ;
  assign n17763 = n15722 & ~n17762 ;
  assign n17764 = n14970 ^ n1578 ^ 1'b0 ;
  assign n17765 = n9966 & n14367 ;
  assign n17766 = n17765 ^ n16046 ^ 1'b0 ;
  assign n17767 = n1504 & ~n14672 ;
  assign n17768 = n17767 ^ n975 ^ 1'b0 ;
  assign n17769 = n17768 ^ n9171 ^ n6522 ;
  assign n17770 = n2608 & ~n2957 ;
  assign n17771 = n7108 ^ n5951 ^ 1'b0 ;
  assign n17772 = n17771 ^ n4149 ^ 1'b0 ;
  assign n17773 = n17236 & ~n17772 ;
  assign n17774 = n5791 | n9737 ;
  assign n17775 = ( n362 & n1692 ) | ( n362 & ~n3608 ) | ( n1692 & ~n3608 ) ;
  assign n17776 = n12900 ^ n8327 ^ 1'b0 ;
  assign n17777 = n11668 ^ n2804 ^ x117 ;
  assign n17778 = n17777 ^ n1765 ^ 1'b0 ;
  assign n17786 = n14266 ^ n3854 ^ 1'b0 ;
  assign n17787 = n9164 ^ n466 ^ 1'b0 ;
  assign n17788 = n9554 & n17787 ;
  assign n17789 = ( n7514 & n9759 ) | ( n7514 & n17788 ) | ( n9759 & n17788 ) ;
  assign n17790 = ( ~n1459 & n5641 ) | ( ~n1459 & n17789 ) | ( n5641 & n17789 ) ;
  assign n17791 = ( n5265 & n17786 ) | ( n5265 & ~n17790 ) | ( n17786 & ~n17790 ) ;
  assign n17780 = n5871 & n6675 ;
  assign n17781 = n6003 & n17780 ;
  assign n17779 = n819 & n2672 ;
  assign n17782 = n17781 ^ n17779 ^ 1'b0 ;
  assign n17783 = n1552 & n17782 ;
  assign n17784 = n17783 ^ n2162 ^ 1'b0 ;
  assign n17785 = n2855 | n17784 ;
  assign n17792 = n17791 ^ n17785 ^ 1'b0 ;
  assign n17793 = n309 & ~n6617 ;
  assign n17794 = n17793 ^ n6092 ^ 1'b0 ;
  assign n17795 = n5920 ^ n1284 ^ 1'b0 ;
  assign n17796 = ~n237 & n17795 ;
  assign n17797 = n17796 ^ n3044 ^ 1'b0 ;
  assign n17798 = n6382 ^ n3755 ^ 1'b0 ;
  assign n17799 = n6680 ^ n6440 ^ 1'b0 ;
  assign n17800 = n6963 | n17799 ;
  assign n17801 = n12549 & ~n17800 ;
  assign n17802 = n370 & n6936 ;
  assign n17803 = n14355 & n17802 ;
  assign n17804 = n7090 ^ n5379 ^ n3708 ;
  assign n17805 = n8257 & n17804 ;
  assign n17806 = ( n601 & ~n6482 ) | ( n601 & n17805 ) | ( ~n6482 & n17805 ) ;
  assign n17807 = n17806 ^ n1434 ^ 1'b0 ;
  assign n17808 = n10161 | n17807 ;
  assign n17809 = n1053 | n17808 ;
  assign n17810 = n11360 ^ n8640 ^ 1'b0 ;
  assign n17811 = n569 | n17810 ;
  assign n17812 = n6514 & n14631 ;
  assign n17813 = ~n10467 & n13034 ;
  assign n17814 = n17813 ^ n4634 ^ 1'b0 ;
  assign n17815 = n2094 & n17814 ;
  assign n17816 = n17815 ^ n14241 ^ n12809 ;
  assign n17820 = n3984 & n5472 ;
  assign n17821 = ~n4933 & n17820 ;
  assign n17822 = ( n2694 & n5493 ) | ( n2694 & ~n17821 ) | ( n5493 & ~n17821 ) ;
  assign n17823 = n1627 & ~n2652 ;
  assign n17824 = ~n17822 & n17823 ;
  assign n17817 = n2456 & n8153 ;
  assign n17818 = n14241 & n17817 ;
  assign n17819 = n778 & ~n17818 ;
  assign n17825 = n17824 ^ n17819 ^ 1'b0 ;
  assign n17826 = ( x89 & n396 ) | ( x89 & n706 ) | ( n396 & n706 ) ;
  assign n17827 = n2907 & n17826 ;
  assign n17828 = n17827 ^ n13454 ^ 1'b0 ;
  assign n17829 = n4454 ^ n427 ^ 1'b0 ;
  assign n17830 = ~n956 & n6466 ;
  assign n17831 = ~n469 & n17830 ;
  assign n17832 = n5628 | n17831 ;
  assign n17833 = n17832 ^ n16049 ^ 1'b0 ;
  assign n17834 = n12485 ^ n3240 ^ 1'b0 ;
  assign n17835 = n4884 | n8530 ;
  assign n17836 = n17834 | n17835 ;
  assign n17837 = ~n6130 & n17836 ;
  assign n17838 = ~n6672 & n17837 ;
  assign n17839 = n8479 & ~n9228 ;
  assign n17840 = n12535 ^ n996 ^ 1'b0 ;
  assign n17843 = n6685 | n6899 ;
  assign n17844 = n17843 ^ n5225 ^ 1'b0 ;
  assign n17842 = n12867 ^ n7623 ^ 1'b0 ;
  assign n17841 = n5255 & n11651 ;
  assign n17845 = n17844 ^ n17842 ^ n17841 ;
  assign n17846 = n9791 ^ n250 ^ 1'b0 ;
  assign n17847 = ~n3979 & n17846 ;
  assign n17848 = n3743 & ~n16201 ;
  assign n17849 = n17848 ^ n1600 ^ 1'b0 ;
  assign n17850 = n17216 ^ n1776 ^ 1'b0 ;
  assign n17851 = n13021 | n17850 ;
  assign n17852 = n11079 ^ n9763 ^ n3845 ;
  assign n17853 = n5017 ^ n2043 ^ 1'b0 ;
  assign n17854 = ~n15966 & n17853 ;
  assign n17855 = n3494 ^ n2752 ^ 1'b0 ;
  assign n17856 = n12502 | n17855 ;
  assign n17857 = n4999 ^ n2535 ^ n2187 ;
  assign n17858 = n14507 ^ n12908 ^ n975 ;
  assign n17859 = n17858 ^ n16876 ^ n311 ;
  assign n17860 = ( n5904 & ~n8169 ) | ( n5904 & n8900 ) | ( ~n8169 & n8900 ) ;
  assign n17861 = ( n17857 & n17859 ) | ( n17857 & n17860 ) | ( n17859 & n17860 ) ;
  assign n17862 = n7008 ^ n372 ^ 1'b0 ;
  assign n17863 = ( n5632 & ~n6523 ) | ( n5632 & n8984 ) | ( ~n6523 & n8984 ) ;
  assign n17864 = n15453 ^ n8404 ^ 1'b0 ;
  assign n17865 = n5797 & n17864 ;
  assign n17866 = n6584 & ~n8996 ;
  assign n17867 = n14968 & ~n17866 ;
  assign n17868 = n2038 ^ n1722 ^ 1'b0 ;
  assign n17869 = n17868 ^ n14323 ^ 1'b0 ;
  assign n17870 = n2987 & ~n17869 ;
  assign n17871 = n6695 & n14595 ;
  assign n17872 = ~n15877 & n17871 ;
  assign n17873 = n3810 ^ n173 ^ 1'b0 ;
  assign n17874 = n3699 | n17873 ;
  assign n17875 = n17874 ^ n4932 ^ 1'b0 ;
  assign n17876 = ~n877 & n10788 ;
  assign n17877 = n17876 ^ n10753 ^ 1'b0 ;
  assign n17880 = n8523 ^ n1118 ^ 1'b0 ;
  assign n17881 = n8914 | n17880 ;
  assign n17878 = n8814 ^ n5402 ^ n4641 ;
  assign n17879 = ~n2845 & n17878 ;
  assign n17882 = n17881 ^ n17879 ^ 1'b0 ;
  assign n17883 = ~n1973 & n10703 ;
  assign n17884 = n17883 ^ n9458 ^ 1'b0 ;
  assign n17885 = n1990 | n9247 ;
  assign n17886 = n17885 ^ n7001 ^ 1'b0 ;
  assign n17887 = n14685 ^ n11311 ^ 1'b0 ;
  assign n17888 = ~n17886 & n17887 ;
  assign n17889 = ~n4492 & n17888 ;
  assign n17890 = ~n6781 & n17889 ;
  assign n17891 = n17890 ^ n1946 ^ 1'b0 ;
  assign n17892 = n17884 & ~n17891 ;
  assign n17893 = n17892 ^ n17593 ^ 1'b0 ;
  assign n17894 = n4664 | n6651 ;
  assign n17895 = n4325 | n14597 ;
  assign n17896 = n2237 & ~n2657 ;
  assign n17900 = n530 & ~n15273 ;
  assign n17901 = n17900 ^ n14900 ^ 1'b0 ;
  assign n17897 = n2637 ^ x12 ^ 1'b0 ;
  assign n17898 = n13849 & ~n17897 ;
  assign n17899 = n17898 ^ n4732 ^ n4608 ;
  assign n17902 = n17901 ^ n17899 ^ n3315 ;
  assign n17903 = n3487 ^ n383 ^ 1'b0 ;
  assign n17904 = ~n11709 & n17903 ;
  assign n17905 = n13811 ^ n4124 ^ 1'b0 ;
  assign n17906 = ~n3344 & n14611 ;
  assign n17907 = n9002 & ~n12085 ;
  assign n17908 = ~n683 & n17907 ;
  assign n17909 = n9667 & ~n17908 ;
  assign n17911 = n14331 ^ n1025 ^ 1'b0 ;
  assign n17912 = n8478 | n17911 ;
  assign n17913 = ( n7314 & n8303 ) | ( n7314 & ~n17912 ) | ( n8303 & ~n17912 ) ;
  assign n17910 = n2359 & n16820 ;
  assign n17914 = n17913 ^ n17910 ^ 1'b0 ;
  assign n17915 = ~n2642 & n17914 ;
  assign n17916 = n6947 ^ n2928 ^ n1791 ;
  assign n17917 = ( n9069 & ~n9545 ) | ( n9069 & n17916 ) | ( ~n9545 & n17916 ) ;
  assign n17918 = n8371 & n16647 ;
  assign n17919 = n17917 & n17918 ;
  assign n17920 = n15570 ^ n4343 ^ 1'b0 ;
  assign n17921 = n17920 ^ n15344 ^ n1000 ;
  assign n17923 = n4839 ^ x75 ^ 1'b0 ;
  assign n17922 = n6346 & ~n10794 ;
  assign n17924 = n17923 ^ n17922 ^ 1'b0 ;
  assign n17925 = n15266 ^ n8481 ^ 1'b0 ;
  assign n17926 = n8328 | n17925 ;
  assign n17927 = n7010 ^ n6937 ^ n975 ;
  assign n17928 = ~n11935 & n13172 ;
  assign n17929 = ~n17927 & n17928 ;
  assign n17930 = n16548 & n17929 ;
  assign n17931 = n12296 ^ n2369 ^ n247 ;
  assign n17932 = n17931 ^ n2316 ^ 1'b0 ;
  assign n17933 = ~n3258 & n17279 ;
  assign n17934 = n17932 & n17933 ;
  assign n17935 = n3623 | n6190 ;
  assign n17936 = n17935 ^ n4854 ^ 1'b0 ;
  assign n17937 = n588 & ~n17936 ;
  assign n17938 = ~n3316 & n17937 ;
  assign n17939 = n642 | n17216 ;
  assign n17940 = n1501 & n6937 ;
  assign n17941 = n17940 ^ n5504 ^ 1'b0 ;
  assign n17942 = n17941 ^ n17375 ^ n2929 ;
  assign n17943 = ( ~n4180 & n7411 ) | ( ~n4180 & n15620 ) | ( n7411 & n15620 ) ;
  assign n17944 = ~n17942 & n17943 ;
  assign n17945 = ~n8331 & n17944 ;
  assign n17946 = ( n8273 & n15748 ) | ( n8273 & ~n17841 ) | ( n15748 & ~n17841 ) ;
  assign n17947 = n8977 ^ n651 ^ 1'b0 ;
  assign n17948 = n3435 ^ n1420 ^ 1'b0 ;
  assign n17949 = n6763 & n17948 ;
  assign n17950 = ~n7960 & n10626 ;
  assign n17951 = n2482 & n17950 ;
  assign n17952 = n9437 & ~n17951 ;
  assign n17953 = n12923 ^ n11718 ^ 1'b0 ;
  assign n17954 = n17411 ^ n2355 ^ 1'b0 ;
  assign n17955 = ( n686 & ~n2720 ) | ( n686 & n17954 ) | ( ~n2720 & n17954 ) ;
  assign n17956 = n2328 | n15801 ;
  assign n17957 = n7718 ^ n4469 ^ 1'b0 ;
  assign n17958 = ( n5710 & ~n17956 ) | ( n5710 & n17957 ) | ( ~n17956 & n17957 ) ;
  assign n17959 = n449 & ~n558 ;
  assign n17960 = n17959 ^ n7085 ^ n4647 ;
  assign n17961 = n16390 ^ n4654 ^ n3031 ;
  assign n17962 = ~n7064 & n17961 ;
  assign n17963 = n2388 & n7222 ;
  assign n17964 = n6257 & n17963 ;
  assign n17965 = n9664 ^ n2362 ^ 1'b0 ;
  assign n17966 = ~n2471 & n17965 ;
  assign n17967 = n16626 ^ n11607 ^ 1'b0 ;
  assign n17968 = n17967 ^ n16100 ^ n11656 ;
  assign n17970 = n14417 | n16862 ;
  assign n17969 = n4827 ^ n2411 ^ n1782 ;
  assign n17971 = n17970 ^ n17969 ^ 1'b0 ;
  assign n17977 = n15796 ^ n863 ^ 1'b0 ;
  assign n17974 = n1971 | n2035 ;
  assign n17972 = n6248 ^ n5824 ^ n2040 ;
  assign n17973 = n3854 & n17972 ;
  assign n17975 = n17974 ^ n17973 ^ 1'b0 ;
  assign n17976 = n17975 ^ n9184 ^ 1'b0 ;
  assign n17978 = n17977 ^ n17976 ^ n651 ;
  assign n17979 = n17978 ^ n5034 ^ 1'b0 ;
  assign n17980 = n758 | n3576 ;
  assign n17981 = n1314 & ~n13536 ;
  assign n17982 = ~n17980 & n17981 ;
  assign n17985 = n4331 & ~n9434 ;
  assign n17986 = ~n1197 & n17985 ;
  assign n17987 = n15216 & n17986 ;
  assign n17983 = n6300 ^ n2164 ^ 1'b0 ;
  assign n17984 = n14170 | n17983 ;
  assign n17988 = n17987 ^ n17984 ^ 1'b0 ;
  assign n17989 = n12885 ^ n5983 ^ 1'b0 ;
  assign n17990 = n9060 ^ n667 ^ 1'b0 ;
  assign n17991 = n8225 & n17990 ;
  assign n17992 = n1206 & n11007 ;
  assign n17993 = n17992 ^ n8915 ^ 1'b0 ;
  assign n17994 = ~n635 & n17993 ;
  assign n17995 = n17987 ^ n9821 ^ 1'b0 ;
  assign n17996 = n11997 & n17995 ;
  assign n17997 = n4654 ^ n3452 ^ n3037 ;
  assign n17998 = n3494 & n10595 ;
  assign n17999 = ~n3658 & n17998 ;
  assign n18000 = n9274 & n13710 ;
  assign n18001 = ~n1585 & n18000 ;
  assign n18002 = n12233 ^ n671 ^ 1'b0 ;
  assign n18003 = n12902 ^ n4471 ^ 1'b0 ;
  assign n18004 = n6133 & ~n18003 ;
  assign n18005 = n12007 ^ n4432 ^ n2917 ;
  assign n18006 = n2019 ^ n619 ^ 1'b0 ;
  assign n18007 = n15768 | n18006 ;
  assign n18008 = n6548 & n7269 ;
  assign n18009 = ~n2589 & n18008 ;
  assign n18010 = n10374 ^ n6201 ^ n6002 ;
  assign n18011 = n18010 ^ n174 ^ 1'b0 ;
  assign n18012 = n10204 & n13216 ;
  assign n18013 = n7471 & n18012 ;
  assign n18014 = x31 | n1853 ;
  assign n18015 = n18014 ^ n5274 ^ 1'b0 ;
  assign n18016 = n18015 ^ n10167 ^ 1'b0 ;
  assign n18017 = n218 & n875 ;
  assign n18018 = ~n218 & n18017 ;
  assign n18019 = ~n4791 & n18018 ;
  assign n18020 = ~n3055 & n8482 ;
  assign n18021 = ~n18019 & n18020 ;
  assign n18022 = ~n12784 & n13793 ;
  assign n18023 = n5185 & n11000 ;
  assign n18024 = n18023 ^ n1476 ^ 1'b0 ;
  assign n18025 = ~n3900 & n16817 ;
  assign n18026 = n1168 & ~n3607 ;
  assign n18027 = n9468 & n18026 ;
  assign n18028 = n18027 ^ n740 ^ 1'b0 ;
  assign n18029 = ~n15426 & n18028 ;
  assign n18030 = n18029 ^ n6434 ^ 1'b0 ;
  assign n18031 = ~n828 & n16370 ;
  assign n18032 = n18031 ^ n8397 ^ 1'b0 ;
  assign n18033 = ( n879 & n4376 ) | ( n879 & ~n18032 ) | ( n4376 & ~n18032 ) ;
  assign n18034 = n14486 & n17873 ;
  assign n18035 = n18034 ^ n13375 ^ 1'b0 ;
  assign n18036 = ~n16126 & n18035 ;
  assign n18037 = n8064 & n18036 ;
  assign n18038 = n18033 & n18037 ;
  assign n18039 = n1012 & ~n11790 ;
  assign n18040 = n18039 ^ n13052 ^ 1'b0 ;
  assign n18041 = n375 | n959 ;
  assign n18042 = n7161 & ~n18041 ;
  assign n18043 = ~n3147 & n8649 ;
  assign n18044 = n18042 & n18043 ;
  assign n18045 = n12991 ^ n6998 ^ 1'b0 ;
  assign n18046 = n18044 | n18045 ;
  assign n18047 = ~n7771 & n18046 ;
  assign n18048 = ( n3597 & n4419 ) | ( n3597 & n17087 ) | ( n4419 & n17087 ) ;
  assign n18049 = ~n4675 & n8425 ;
  assign n18050 = n18049 ^ n2751 ^ 1'b0 ;
  assign n18051 = n14595 & n18050 ;
  assign n18052 = ~n18048 & n18051 ;
  assign n18053 = n6517 ^ n998 ^ 1'b0 ;
  assign n18054 = n8733 & ~n18053 ;
  assign n18055 = n1379 | n7814 ;
  assign n18056 = n9356 ^ n9214 ^ n6900 ;
  assign n18057 = n2313 ^ n342 ^ 1'b0 ;
  assign n18058 = n4538 & n18057 ;
  assign n18059 = n12188 & n18058 ;
  assign n18060 = n14640 ^ n2221 ^ 1'b0 ;
  assign n18061 = n5312 & ~n18060 ;
  assign n18062 = n1938 & ~n18061 ;
  assign n18063 = n176 & ~n18062 ;
  assign n18064 = n5203 | n8281 ;
  assign n18065 = n18064 ^ n2328 ^ 1'b0 ;
  assign n18066 = n14993 ^ n12129 ^ 1'b0 ;
  assign n18067 = n16207 & ~n18066 ;
  assign n18068 = n10448 & n12485 ;
  assign n18069 = n8437 ^ n1379 ^ n857 ;
  assign n18070 = ~x118 & n7729 ;
  assign n18071 = x17 & ~n17971 ;
  assign n18072 = ~n3562 & n18071 ;
  assign n18074 = n9265 ^ n4647 ^ 1'b0 ;
  assign n18075 = n3519 | n18074 ;
  assign n18073 = n4068 & ~n6255 ;
  assign n18076 = n18075 ^ n18073 ^ 1'b0 ;
  assign n18077 = n8069 & n17551 ;
  assign n18078 = n18077 ^ n6378 ^ 1'b0 ;
  assign n18079 = n2404 ^ n2233 ^ n1832 ;
  assign n18080 = ~n9979 & n18079 ;
  assign n18081 = n2147 & ~n7103 ;
  assign n18082 = n6906 & ~n7922 ;
  assign n18083 = n18081 & n18082 ;
  assign n18084 = ~n5043 & n9381 ;
  assign n18085 = n18083 | n18084 ;
  assign n18086 = n18085 ^ n4078 ^ 1'b0 ;
  assign n18087 = n6094 ^ n4012 ^ 1'b0 ;
  assign n18088 = n17667 ^ n10627 ^ 1'b0 ;
  assign n18089 = n15858 ^ n2317 ^ 1'b0 ;
  assign n18091 = n6380 & ~n7357 ;
  assign n18090 = n9271 ^ n1710 ^ 1'b0 ;
  assign n18092 = n18091 ^ n18090 ^ n4097 ;
  assign n18093 = n13293 ^ n4222 ^ 1'b0 ;
  assign n18094 = ~n2419 & n9178 ;
  assign n18095 = n2973 & ~n8628 ;
  assign n18096 = ~n2554 & n18095 ;
  assign n18097 = n4848 ^ n3660 ^ 1'b0 ;
  assign n18098 = ~n10239 & n18097 ;
  assign n18099 = n18098 ^ n14075 ^ 1'b0 ;
  assign n18100 = n6344 ^ n4053 ^ 1'b0 ;
  assign n18101 = ~n9713 & n18100 ;
  assign n18102 = n18101 ^ n17667 ^ 1'b0 ;
  assign n18103 = ~n4557 & n18102 ;
  assign n18104 = n13386 ^ n3256 ^ 1'b0 ;
  assign n18105 = ~n2850 & n18104 ;
  assign n18106 = n2859 & n10893 ;
  assign n18107 = n18105 & n18106 ;
  assign n18108 = n389 & n3223 ;
  assign n18109 = n18108 ^ n4394 ^ 1'b0 ;
  assign n18110 = n13667 & ~n18109 ;
  assign n18111 = n5039 ^ n3608 ^ 1'b0 ;
  assign n18112 = n18111 ^ n15769 ^ n9323 ;
  assign n18113 = n18112 ^ n6453 ^ 1'b0 ;
  assign n18114 = n18110 & ~n18113 ;
  assign n18115 = n5916 ^ n4373 ^ 1'b0 ;
  assign n18116 = ( n7781 & ~n9268 ) | ( n7781 & n18115 ) | ( ~n9268 & n18115 ) ;
  assign n18117 = n7550 & ~n10600 ;
  assign n18118 = n18116 & ~n18117 ;
  assign n18119 = n557 & ~n12999 ;
  assign n18120 = n18119 ^ n9474 ^ 1'b0 ;
  assign n18121 = ~n1632 & n13363 ;
  assign n18122 = ~n1248 & n18121 ;
  assign n18123 = n18122 ^ n4730 ^ 1'b0 ;
  assign n18124 = ~n2451 & n4990 ;
  assign n18125 = n4285 & n6109 ;
  assign n18126 = ~n3191 & n10396 ;
  assign n18127 = n6478 ^ n1160 ^ 1'b0 ;
  assign n18128 = n18127 ^ n3786 ^ 1'b0 ;
  assign n18129 = n7880 & n18128 ;
  assign n18130 = n11570 ^ n243 ^ 1'b0 ;
  assign n18131 = n18129 & ~n18130 ;
  assign n18136 = n8790 ^ n337 ^ 1'b0 ;
  assign n18132 = n4038 & n4239 ;
  assign n18133 = n3401 & n18132 ;
  assign n18134 = n12339 ^ n6506 ^ 1'b0 ;
  assign n18135 = ~n18133 & n18134 ;
  assign n18137 = n18136 ^ n18135 ^ n1230 ;
  assign n18138 = n1338 & n17607 ;
  assign n18139 = n14189 & n18138 ;
  assign n18140 = n1345 & ~n18139 ;
  assign n18141 = ~n18137 & n18140 ;
  assign n18142 = n4812 & ~n9574 ;
  assign n18146 = n1452 ^ n438 ^ 1'b0 ;
  assign n18143 = n8606 ^ n5820 ^ 1'b0 ;
  assign n18144 = x51 & n18143 ;
  assign n18145 = n18144 ^ n5191 ^ n4462 ;
  assign n18147 = n18146 ^ n18145 ^ 1'b0 ;
  assign n18148 = n15581 ^ n13655 ^ n10682 ;
  assign n18149 = n17446 ^ n3389 ^ x51 ;
  assign n18150 = n1745 & n3649 ;
  assign n18151 = n4456 & n18150 ;
  assign n18152 = ~n2112 & n17519 ;
  assign n18153 = n4541 | n18152 ;
  assign n18154 = ( n2730 & n3147 ) | ( n2730 & n13598 ) | ( n3147 & n13598 ) ;
  assign n18155 = n2091 & ~n18154 ;
  assign n18156 = n7890 & n18155 ;
  assign n18157 = n3055 & ~n13975 ;
  assign n18158 = n18157 ^ n2425 ^ 1'b0 ;
  assign n18159 = ~n7206 & n18158 ;
  assign n18160 = n18159 ^ n12877 ^ 1'b0 ;
  assign n18161 = n3192 & n8826 ;
  assign n18162 = n18161 ^ n1034 ^ 1'b0 ;
  assign n18163 = ~n2062 & n3876 ;
  assign n18164 = ( n718 & n18162 ) | ( n718 & ~n18163 ) | ( n18162 & ~n18163 ) ;
  assign n18165 = n6522 & n9904 ;
  assign n18168 = n15201 ^ n4187 ^ 1'b0 ;
  assign n18169 = n18168 ^ n13955 ^ n5584 ;
  assign n18166 = ~n918 & n2010 ;
  assign n18167 = n18166 ^ n3472 ^ 1'b0 ;
  assign n18170 = n18169 ^ n18167 ^ 1'b0 ;
  assign n18171 = n17069 ^ n14105 ^ n11128 ;
  assign n18172 = n3861 & ~n10312 ;
  assign n18173 = n18172 ^ n10363 ^ 1'b0 ;
  assign n18174 = n3188 ^ x62 ^ 1'b0 ;
  assign n18175 = n18173 & n18174 ;
  assign n18176 = n16860 ^ n8905 ^ n3173 ;
  assign n18177 = ~n3959 & n18176 ;
  assign n18178 = n3446 | n11614 ;
  assign n18179 = n18177 | n18178 ;
  assign n18180 = ~n1374 & n15723 ;
  assign n18181 = n1374 & ~n10114 ;
  assign n18182 = n18181 ^ n15739 ^ 1'b0 ;
  assign n18184 = n12531 & ~n12667 ;
  assign n18183 = n6473 & n16734 ;
  assign n18185 = n18184 ^ n18183 ^ 1'b0 ;
  assign n18186 = n6895 ^ n4283 ^ 1'b0 ;
  assign n18187 = n7268 | n18186 ;
  assign n18188 = n18187 ^ n3380 ^ 1'b0 ;
  assign n18189 = ( n527 & n7793 ) | ( n527 & n18188 ) | ( n7793 & n18188 ) ;
  assign n18190 = n18189 ^ n5458 ^ 1'b0 ;
  assign n18191 = ~n2921 & n5124 ;
  assign n18192 = n791 | n11325 ;
  assign n18193 = ( n8717 & n18191 ) | ( n8717 & ~n18192 ) | ( n18191 & ~n18192 ) ;
  assign n18194 = n15140 & ~n16099 ;
  assign n18195 = n12917 ^ n2912 ^ 1'b0 ;
  assign n18196 = n250 & ~n18195 ;
  assign n18197 = n2024 & ~n10872 ;
  assign n18198 = n918 & n18197 ;
  assign n18201 = n9963 ^ n7314 ^ n4181 ;
  assign n18199 = n4617 & n15451 ;
  assign n18200 = ~n4617 & n18199 ;
  assign n18202 = n18201 ^ n18200 ^ n10275 ;
  assign n18203 = ( ~x50 & n1775 ) | ( ~x50 & n5097 ) | ( n1775 & n5097 ) ;
  assign n18204 = ~n9195 & n9303 ;
  assign n18205 = ~n18203 & n18204 ;
  assign n18206 = n18205 ^ n10619 ^ n2602 ;
  assign n18208 = n6135 ^ n2703 ^ 1'b0 ;
  assign n18209 = n11178 | n18208 ;
  assign n18207 = n7831 | n13853 ;
  assign n18210 = n18209 ^ n18207 ^ 1'b0 ;
  assign n18211 = n16499 ^ n13039 ^ 1'b0 ;
  assign n18212 = n13579 ^ n5745 ^ n4841 ;
  assign n18213 = n13109 ^ n6670 ^ 1'b0 ;
  assign n18214 = n7111 & n18213 ;
  assign n18215 = n16927 ^ n10416 ^ n7111 ;
  assign n18216 = n6145 | n6667 ;
  assign n18217 = n18216 ^ n310 ^ 1'b0 ;
  assign n18218 = n18217 ^ n387 ^ 1'b0 ;
  assign n18219 = n16174 ^ n5205 ^ 1'b0 ;
  assign n18220 = n16963 ^ n10221 ^ 1'b0 ;
  assign n18221 = n17677 ^ n9158 ^ 1'b0 ;
  assign n18222 = n5458 & ~n18221 ;
  assign n18223 = n16648 ^ n11095 ^ n9554 ;
  assign n18224 = n4283 | n14410 ;
  assign n18225 = ( x16 & n8692 ) | ( x16 & n11364 ) | ( n8692 & n11364 ) ;
  assign n18226 = n7962 ^ n189 ^ 1'b0 ;
  assign n18227 = n18226 ^ n1124 ^ 1'b0 ;
  assign n18228 = n13449 ^ n5231 ^ 1'b0 ;
  assign n18229 = n3424 & n5152 ;
  assign n18230 = n18228 & n18229 ;
  assign n18231 = n5892 | n18230 ;
  assign n18232 = n11396 & ~n18231 ;
  assign n18233 = n5158 & n6354 ;
  assign n18234 = n18233 ^ n7507 ^ n5032 ;
  assign n18235 = n1044 | n13731 ;
  assign n18237 = ~n3108 & n4610 ;
  assign n18236 = ~n5584 & n14124 ;
  assign n18238 = n18237 ^ n18236 ^ 1'b0 ;
  assign n18239 = n18238 ^ n9214 ^ 1'b0 ;
  assign n18240 = ~n969 & n18239 ;
  assign n18241 = n18240 ^ n4252 ^ 1'b0 ;
  assign n18242 = n8537 & ~n17383 ;
  assign n18243 = n12579 & n18242 ;
  assign n18244 = n18243 ^ n1791 ^ 1'b0 ;
  assign n18245 = n962 & ~n18244 ;
  assign n18246 = n9374 ^ n6204 ^ n5530 ;
  assign n18247 = ~n2788 & n9591 ;
  assign n18248 = n3995 & n5781 ;
  assign n18249 = n18248 ^ n1143 ^ 1'b0 ;
  assign n18250 = n18249 ^ n4070 ^ n3014 ;
  assign n18251 = n13926 & ~n18250 ;
  assign n18252 = ( n2375 & ~n10173 ) | ( n2375 & n18251 ) | ( ~n10173 & n18251 ) ;
  assign n18254 = n9422 ^ n2865 ^ 1'b0 ;
  assign n18253 = n454 & n8385 ;
  assign n18255 = n18254 ^ n18253 ^ 1'b0 ;
  assign n18259 = n1693 ^ n1106 ^ 1'b0 ;
  assign n18256 = ~n6711 & n14915 ;
  assign n18257 = n9366 & ~n18256 ;
  assign n18258 = n13977 | n18257 ;
  assign n18260 = n18259 ^ n18258 ^ 1'b0 ;
  assign n18261 = ~n7792 & n9728 ;
  assign n18262 = ( n4281 & n6218 ) | ( n4281 & n18261 ) | ( n6218 & n18261 ) ;
  assign n18263 = n13764 ^ n9092 ^ 1'b0 ;
  assign n18264 = n14032 ^ n7347 ^ 1'b0 ;
  assign n18268 = n11562 ^ n2796 ^ 1'b0 ;
  assign n18269 = n12411 & ~n18268 ;
  assign n18265 = n2484 ^ n1547 ^ 1'b0 ;
  assign n18266 = n1771 & n18265 ;
  assign n18267 = ( n1286 & n3208 ) | ( n1286 & n18266 ) | ( n3208 & n18266 ) ;
  assign n18270 = n18269 ^ n18267 ^ 1'b0 ;
  assign n18271 = n10981 | n18270 ;
  assign n18272 = n14869 | n18271 ;
  assign n18273 = n18272 ^ n11235 ^ 1'b0 ;
  assign n18274 = n901 | n7743 ;
  assign n18275 = n18274 ^ n12596 ^ 1'b0 ;
  assign n18276 = n14716 ^ n4752 ^ 1'b0 ;
  assign n18277 = n18276 ^ n14251 ^ 1'b0 ;
  assign n18278 = n7012 & ~n18277 ;
  assign n18279 = ( n7028 & n8084 ) | ( n7028 & n13548 ) | ( n8084 & n13548 ) ;
  assign n18280 = ( n3557 & n9276 ) | ( n3557 & ~n10160 ) | ( n9276 & ~n10160 ) ;
  assign n18281 = n10565 ^ n1582 ^ 1'b0 ;
  assign n18282 = n1106 | n18281 ;
  assign n18283 = n5822 & ~n18282 ;
  assign n18284 = n1300 & n18283 ;
  assign n18285 = n17842 ^ n4987 ^ n3791 ;
  assign n18286 = n3652 & ~n18285 ;
  assign n18288 = n13460 ^ n6516 ^ 1'b0 ;
  assign n18287 = n6116 & n17570 ;
  assign n18289 = n18288 ^ n18287 ^ 1'b0 ;
  assign n18290 = n18289 ^ n14357 ^ 1'b0 ;
  assign n18291 = n7972 & n12127 ;
  assign n18292 = n18291 ^ n6623 ^ 1'b0 ;
  assign n18293 = n3189 & ~n7402 ;
  assign n18294 = n18293 ^ n1918 ^ 1'b0 ;
  assign n18295 = n18292 & ~n18294 ;
  assign n18296 = n1238 & ~n3684 ;
  assign n18297 = n12971 ^ n8645 ^ 1'b0 ;
  assign n18298 = n14510 & ~n18297 ;
  assign n18299 = n18298 ^ n13839 ^ 1'b0 ;
  assign n18300 = ( n7768 & ~n18296 ) | ( n7768 & n18299 ) | ( ~n18296 & n18299 ) ;
  assign n18301 = ( n2654 & n2673 ) | ( n2654 & n3959 ) | ( n2673 & n3959 ) ;
  assign n18304 = n4186 | n7370 ;
  assign n18302 = n12350 ^ n4927 ^ 1'b0 ;
  assign n18303 = n17202 & ~n18302 ;
  assign n18305 = n18304 ^ n18303 ^ n17065 ;
  assign n18306 = n16181 ^ n10767 ^ 1'b0 ;
  assign n18307 = n2806 & ~n4996 ;
  assign n18308 = n6705 & n18307 ;
  assign n18309 = n4167 & ~n5918 ;
  assign n18310 = n18309 ^ n9065 ^ n1197 ;
  assign n18311 = n6939 ^ n551 ^ 1'b0 ;
  assign n18312 = n7559 | n18311 ;
  assign n18313 = n18312 ^ n8936 ^ 1'b0 ;
  assign n18314 = n7330 | n7384 ;
  assign n18315 = n16857 ^ n11702 ^ n616 ;
  assign n18316 = ~n16101 & n18315 ;
  assign n18317 = n18314 & n18316 ;
  assign n18318 = n3415 & ~n3638 ;
  assign n18319 = n18318 ^ n8453 ^ 1'b0 ;
  assign n18320 = n2041 & ~n4161 ;
  assign n18321 = ~n7518 & n18320 ;
  assign n18322 = n13478 | n18321 ;
  assign n18323 = ~n740 & n16958 ;
  assign n18324 = ~n3321 & n5504 ;
  assign n18325 = n7701 & n9540 ;
  assign n18326 = n8498 & n18325 ;
  assign n18327 = n4471 | n18326 ;
  assign n18328 = ( n7966 & n8137 ) | ( n7966 & ~n11692 ) | ( n8137 & ~n11692 ) ;
  assign n18329 = n1681 & ~n11180 ;
  assign n18330 = ( n10668 & ~n18328 ) | ( n10668 & n18329 ) | ( ~n18328 & n18329 ) ;
  assign n18331 = n3590 & n6392 ;
  assign n18332 = ~n215 & n6658 ;
  assign n18333 = n18331 & n18332 ;
  assign n18334 = n13064 & ~n18333 ;
  assign n18335 = n18330 & n18334 ;
  assign n18336 = ~n7219 & n9584 ;
  assign n18337 = n3411 & ~n13406 ;
  assign n18338 = ~n7346 & n7750 ;
  assign n18339 = ~n5967 & n6607 ;
  assign n18340 = ~n3167 & n18339 ;
  assign n18341 = n16313 ^ n869 ^ 1'b0 ;
  assign n18342 = n17421 ^ n2508 ^ 1'b0 ;
  assign n18343 = n2543 & n3528 ;
  assign n18344 = ( ~n8834 & n11442 ) | ( ~n8834 & n13814 ) | ( n11442 & n13814 ) ;
  assign n18345 = n18343 & n18344 ;
  assign n18346 = n14340 ^ n13529 ^ 1'b0 ;
  assign n18347 = ~n3999 & n18346 ;
  assign n18348 = n395 & ~n8190 ;
  assign n18350 = n2945 ^ n2892 ^ 1'b0 ;
  assign n18351 = n5503 & n18350 ;
  assign n18349 = n3976 | n11859 ;
  assign n18352 = n18351 ^ n18349 ^ 1'b0 ;
  assign n18353 = n4076 & ~n5361 ;
  assign n18354 = n18353 ^ n8516 ^ 1'b0 ;
  assign n18355 = ~n8075 & n18354 ;
  assign n18356 = n18352 & n18355 ;
  assign n18357 = n17584 & n18356 ;
  assign n18358 = n8530 & n18357 ;
  assign n18359 = ~n1462 & n13299 ;
  assign n18360 = n8761 ^ n1212 ^ 1'b0 ;
  assign n18361 = n2113 | n18360 ;
  assign n18362 = n1046 & ~n4651 ;
  assign n18363 = ~n18361 & n18362 ;
  assign n18364 = n7949 ^ n4466 ^ n945 ;
  assign n18365 = n7719 ^ n1826 ^ 1'b0 ;
  assign n18366 = n3701 | n14976 ;
  assign n18367 = n910 & n1584 ;
  assign n18368 = n11930 & ~n18367 ;
  assign n18369 = n15864 ^ n11294 ^ n5218 ;
  assign n18370 = n18368 | n18369 ;
  assign n18371 = ( n1630 & n9655 ) | ( n1630 & ~n10029 ) | ( n9655 & ~n10029 ) ;
  assign n18372 = n18014 ^ n9977 ^ 1'b0 ;
  assign n18373 = n1499 & n7939 ;
  assign n18374 = n15131 | n18373 ;
  assign n18375 = x123 & n18374 ;
  assign n18376 = n11614 & n16489 ;
  assign n18377 = n11603 ^ n11447 ^ n1743 ;
  assign n18382 = n5490 ^ n4897 ^ 1'b0 ;
  assign n18383 = n1057 & n18382 ;
  assign n18379 = x88 & n1173 ;
  assign n18380 = n4309 & n18379 ;
  assign n18381 = n18380 ^ n452 ^ x36 ;
  assign n18378 = n14152 ^ n10621 ^ 1'b0 ;
  assign n18384 = n18383 ^ n18381 ^ n18378 ;
  assign n18385 = x106 | n7158 ;
  assign n18386 = n6815 ^ n143 ^ 1'b0 ;
  assign n18387 = ~n10631 & n18386 ;
  assign n18388 = ~n10366 & n14601 ;
  assign n18389 = n14932 & ~n18388 ;
  assign n18390 = n6627 ^ n5127 ^ 1'b0 ;
  assign n18391 = n11179 ^ n9018 ^ n2958 ;
  assign n18393 = n2030 & ~n4017 ;
  assign n18394 = n2264 & n18393 ;
  assign n18395 = n18394 ^ n8555 ^ 1'b0 ;
  assign n18392 = n9349 | n13360 ;
  assign n18396 = n18395 ^ n18392 ^ 1'b0 ;
  assign n18397 = n7707 ^ n616 ^ 1'b0 ;
  assign n18398 = n14907 & n18397 ;
  assign n18399 = n5043 & n13882 ;
  assign n18400 = n17934 ^ n8807 ^ 1'b0 ;
  assign n18401 = n5785 & ~n18400 ;
  assign n18402 = ( n13668 & ~n18399 ) | ( n13668 & n18401 ) | ( ~n18399 & n18401 ) ;
  assign n18403 = n5456 ^ n4992 ^ 1'b0 ;
  assign n18404 = n6337 | n16703 ;
  assign n18405 = n5304 | n12221 ;
  assign n18406 = n18405 ^ n1918 ^ 1'b0 ;
  assign n18407 = n6784 | n18406 ;
  assign n18408 = n18407 ^ n6240 ^ 1'b0 ;
  assign n18409 = n15099 ^ n3775 ^ n2725 ;
  assign n18410 = n2493 ^ n817 ^ 1'b0 ;
  assign n18411 = n3108 & ~n18410 ;
  assign n18412 = n16548 ^ n6194 ^ 1'b0 ;
  assign n18413 = ( n14412 & n18411 ) | ( n14412 & ~n18412 ) | ( n18411 & ~n18412 ) ;
  assign n18414 = ~n2062 & n2295 ;
  assign n18415 = ~n5888 & n18414 ;
  assign n18416 = n18415 ^ n11940 ^ 1'b0 ;
  assign n18417 = ~n3199 & n18416 ;
  assign n18418 = n18417 ^ n16347 ^ n2839 ;
  assign n18419 = ~n6756 & n11406 ;
  assign n18420 = n842 & n12531 ;
  assign n18421 = n1648 & n18420 ;
  assign n18422 = n4107 | n18421 ;
  assign n18423 = n7962 ^ n1684 ^ 1'b0 ;
  assign n18424 = ~n16479 & n18423 ;
  assign n18425 = n11688 ^ n683 ^ 1'b0 ;
  assign n18426 = n9417 & ~n18425 ;
  assign n18429 = ~n5089 & n6231 ;
  assign n18427 = n11311 ^ n4361 ^ n2285 ;
  assign n18428 = n18427 ^ n13264 ^ 1'b0 ;
  assign n18430 = n18429 ^ n18428 ^ n9158 ;
  assign n18431 = n11061 ^ n7989 ^ n884 ;
  assign n18432 = n7501 ^ n7321 ^ 1'b0 ;
  assign n18433 = ( n1512 & n14841 ) | ( n1512 & n18432 ) | ( n14841 & n18432 ) ;
  assign n18434 = n3638 ^ n3399 ^ 1'b0 ;
  assign n18435 = ~n13497 & n18434 ;
  assign n18436 = n5606 & n14439 ;
  assign n18437 = ~n1800 & n17437 ;
  assign n18438 = ( n2958 & n14178 ) | ( n2958 & ~n18331 ) | ( n14178 & ~n18331 ) ;
  assign n18439 = n12809 ^ n3930 ^ 1'b0 ;
  assign n18440 = n5262 | n18439 ;
  assign n18441 = n6761 ^ n3703 ^ 1'b0 ;
  assign n18442 = n18440 | n18441 ;
  assign n18443 = n18442 ^ n13105 ^ 1'b0 ;
  assign n18444 = ( n3785 & ~n6283 ) | ( n3785 & n18443 ) | ( ~n6283 & n18443 ) ;
  assign n18445 = ~n1059 & n3835 ;
  assign n18446 = n3169 & n18445 ;
  assign n18447 = n18446 ^ n1627 ^ n1033 ;
  assign n18448 = n1575 & ~n2083 ;
  assign n18449 = n4351 & n18448 ;
  assign n18450 = n18447 | n18449 ;
  assign n18451 = n18450 ^ n17264 ^ 1'b0 ;
  assign n18454 = x3 | n2306 ;
  assign n18455 = n18454 ^ n16842 ^ 1'b0 ;
  assign n18456 = n1481 & ~n18455 ;
  assign n18452 = ~n707 & n8922 ;
  assign n18453 = n1403 | n18452 ;
  assign n18457 = n18456 ^ n18453 ^ 1'b0 ;
  assign n18458 = ~n2049 & n14512 ;
  assign n18459 = ~n875 & n18458 ;
  assign n18460 = n17055 ^ n4745 ^ 1'b0 ;
  assign n18461 = n7567 ^ n6208 ^ 1'b0 ;
  assign n18462 = n18461 ^ n9862 ^ n7742 ;
  assign n18463 = n12177 ^ n11416 ^ n5290 ;
  assign n18464 = n15227 ^ n3363 ^ 1'b0 ;
  assign n18465 = n8287 | n18464 ;
  assign n18466 = n11031 | n18465 ;
  assign n18467 = n18463 & ~n18466 ;
  assign n18468 = n12149 ^ n2654 ^ 1'b0 ;
  assign n18469 = n5001 | n18468 ;
  assign n18470 = n831 & ~n18469 ;
  assign n18471 = n18470 ^ n8132 ^ 1'b0 ;
  assign n18472 = n13195 ^ n9398 ^ 1'b0 ;
  assign n18473 = n7920 & n18472 ;
  assign n18474 = n13414 ^ n9830 ^ 1'b0 ;
  assign n18476 = n6452 & ~n7473 ;
  assign n18477 = n4402 & n18476 ;
  assign n18478 = ~n17351 & n18477 ;
  assign n18475 = ( n6367 & n7605 ) | ( n6367 & n8737 ) | ( n7605 & n8737 ) ;
  assign n18479 = n18478 ^ n18475 ^ 1'b0 ;
  assign n18480 = ( x51 & ~n8144 ) | ( x51 & n12239 ) | ( ~n8144 & n12239 ) ;
  assign n18481 = ( n176 & n13796 ) | ( n176 & ~n18480 ) | ( n13796 & ~n18480 ) ;
  assign n18482 = ~n16642 & n18481 ;
  assign n18483 = ~n372 & n2222 ;
  assign n18484 = n2436 & n18483 ;
  assign n18485 = n7754 & ~n13950 ;
  assign n18486 = n7258 ^ n2219 ^ 1'b0 ;
  assign n18487 = n13454 ^ n4121 ^ 1'b0 ;
  assign n18488 = n15253 | n18487 ;
  assign n18489 = n7217 | n10722 ;
  assign n18490 = n8862 ^ n1935 ^ 1'b0 ;
  assign n18491 = n681 & ~n11899 ;
  assign n18492 = ~n12995 & n18491 ;
  assign n18493 = n18490 & n18492 ;
  assign n18494 = n11971 ^ n4472 ^ 1'b0 ;
  assign n18495 = n10104 ^ n9661 ^ 1'b0 ;
  assign n18496 = n4691 ^ n3908 ^ n3831 ;
  assign n18497 = n10198 & ~n12994 ;
  assign n18498 = n6651 & n18497 ;
  assign n18499 = n18496 & ~n18498 ;
  assign n18500 = ~n18495 & n18499 ;
  assign n18501 = n11618 & n17111 ;
  assign n18502 = n18501 ^ n15747 ^ 1'b0 ;
  assign n18503 = n8797 ^ n7758 ^ n4494 ;
  assign n18504 = n18503 ^ n599 ^ 1'b0 ;
  assign n18505 = n18502 | n18504 ;
  assign n18508 = n4783 ^ x115 ^ 1'b0 ;
  assign n18509 = n4010 & n18508 ;
  assign n18506 = n1499 | n4981 ;
  assign n18507 = n1476 & n18506 ;
  assign n18510 = n18509 ^ n18507 ^ 1'b0 ;
  assign n18511 = n1892 & ~n13043 ;
  assign n18512 = n8404 & n18511 ;
  assign n18513 = n5373 & n18512 ;
  assign n18514 = ~n1880 & n18513 ;
  assign n18515 = n8256 & ~n14940 ;
  assign n18516 = n11517 | n13374 ;
  assign n18517 = n18516 ^ n13929 ^ 1'b0 ;
  assign n18518 = n3832 ^ n425 ^ 1'b0 ;
  assign n18519 = ~n10910 & n18518 ;
  assign n18520 = n18517 & n18519 ;
  assign n18522 = n2609 & ~n12399 ;
  assign n18521 = ~n220 & n14718 ;
  assign n18523 = n18522 ^ n18521 ^ 1'b0 ;
  assign n18524 = n10733 ^ n1765 ^ 1'b0 ;
  assign n18525 = n323 & ~n4858 ;
  assign n18526 = n18525 ^ n17374 ^ 1'b0 ;
  assign n18527 = n11699 ^ n6362 ^ n1637 ;
  assign n18528 = n18527 ^ n7478 ^ 1'b0 ;
  assign n18529 = ~n14636 & n18528 ;
  assign n18530 = n9577 ^ n6828 ^ n403 ;
  assign n18531 = ~n353 & n18530 ;
  assign n18532 = n6330 & n11432 ;
  assign n18533 = ~n5116 & n18532 ;
  assign n18534 = n18533 ^ n2926 ^ 1'b0 ;
  assign n18535 = ~n11300 & n17558 ;
  assign n18536 = n18535 ^ n5333 ^ 1'b0 ;
  assign n18537 = n2035 & n3786 ;
  assign n18538 = n3348 | n14340 ;
  assign n18539 = n3972 | n18538 ;
  assign n18540 = n18537 & n18539 ;
  assign n18541 = n17537 & n18540 ;
  assign n18542 = n11292 & ~n18541 ;
  assign n18543 = n18542 ^ n2809 ^ 1'b0 ;
  assign n18544 = n18543 ^ n2706 ^ n1095 ;
  assign n18548 = n15730 ^ n9681 ^ n2970 ;
  assign n18545 = n1171 & n5551 ;
  assign n18546 = ~n2532 & n14322 ;
  assign n18547 = ~n18545 & n18546 ;
  assign n18549 = n18548 ^ n18547 ^ n1995 ;
  assign n18550 = ~n6431 & n11525 ;
  assign n18551 = n13536 ^ n3708 ^ n1684 ;
  assign n18552 = ~n3203 & n6391 ;
  assign n18553 = n5567 & ~n17691 ;
  assign n18554 = ~n2826 & n18553 ;
  assign n18555 = n12546 ^ n5259 ^ 1'b0 ;
  assign n18556 = n615 & n18555 ;
  assign n18557 = n935 & n18556 ;
  assign n18558 = n18557 ^ n7025 ^ n3578 ;
  assign n18559 = n1055 ^ n469 ^ 1'b0 ;
  assign n18560 = ( ~n8860 & n10763 ) | ( ~n8860 & n18559 ) | ( n10763 & n18559 ) ;
  assign n18561 = n17661 ^ n4981 ^ n3767 ;
  assign n18562 = n11818 ^ n4078 ^ 1'b0 ;
  assign n18563 = n7056 | n18562 ;
  assign n18564 = n9474 ^ n1085 ^ n1057 ;
  assign n18565 = ( ~n3339 & n11903 ) | ( ~n3339 & n18564 ) | ( n11903 & n18564 ) ;
  assign n18566 = ( n1989 & ~n8976 ) | ( n1989 & n18565 ) | ( ~n8976 & n18565 ) ;
  assign n18567 = n1154 & ~n8090 ;
  assign n18568 = n18566 & n18567 ;
  assign n18569 = n239 & n15569 ;
  assign n18570 = n18569 ^ n11300 ^ 1'b0 ;
  assign n18571 = n11611 ^ n4841 ^ 1'b0 ;
  assign n18572 = n6778 ^ n2914 ^ 1'b0 ;
  assign n18573 = n18571 & ~n18572 ;
  assign n18574 = n1575 & ~n3142 ;
  assign n18575 = n3528 & n18574 ;
  assign n18576 = ( n12496 & n17937 ) | ( n12496 & ~n18575 ) | ( n17937 & ~n18575 ) ;
  assign n18577 = ~n1156 & n3718 ;
  assign n18578 = n4524 | n18577 ;
  assign n18579 = n678 & ~n5029 ;
  assign n18580 = n18579 ^ n11340 ^ 1'b0 ;
  assign n18581 = n17603 ^ n1179 ^ 1'b0 ;
  assign n18582 = n14114 & ~n18581 ;
  assign n18583 = n17686 ^ n17109 ^ n16329 ;
  assign n18584 = ~n2550 & n9092 ;
  assign n18585 = ( n3145 & ~n4627 ) | ( n3145 & n7284 ) | ( ~n4627 & n7284 ) ;
  assign n18586 = n5126 & ~n6056 ;
  assign n18587 = n18585 & n18586 ;
  assign n18588 = n2844 | n7639 ;
  assign n18589 = n3589 & n8695 ;
  assign n18590 = n15872 ^ n15711 ^ 1'b0 ;
  assign n18591 = ~n18589 & n18590 ;
  assign n18592 = n711 & ~n12188 ;
  assign n18593 = n642 | n4749 ;
  assign n18594 = n10459 | n14811 ;
  assign n18595 = n18594 ^ n18469 ^ 1'b0 ;
  assign n18596 = n3861 ^ n2886 ^ 1'b0 ;
  assign n18597 = n8132 & n8341 ;
  assign n18598 = n18597 ^ n17108 ^ 1'b0 ;
  assign n18599 = n18596 | n18598 ;
  assign n18600 = n13713 ^ n2847 ^ n1909 ;
  assign n18601 = ( ~n5352 & n15728 ) | ( ~n5352 & n18600 ) | ( n15728 & n18600 ) ;
  assign n18602 = ~n4857 & n5402 ;
  assign n18603 = ~n5402 & n18602 ;
  assign n18604 = n856 & ~n18603 ;
  assign n18605 = n2892 & ~n18604 ;
  assign n18606 = n18604 & n18605 ;
  assign n18607 = n13989 ^ n8226 ^ 1'b0 ;
  assign n18610 = n5452 & ~n5749 ;
  assign n18611 = n18610 ^ n7566 ^ 1'b0 ;
  assign n18608 = n5711 & ~n14618 ;
  assign n18609 = n5812 | n18608 ;
  assign n18612 = n18611 ^ n18609 ^ 1'b0 ;
  assign n18613 = n4233 ^ n3292 ^ 1'b0 ;
  assign n18614 = ( n1449 & n9554 ) | ( n1449 & n13437 ) | ( n9554 & n13437 ) ;
  assign n18615 = n569 ^ x68 ^ 1'b0 ;
  assign n18616 = n8199 & ~n18615 ;
  assign n18617 = n18616 ^ n3149 ^ 1'b0 ;
  assign n18618 = n4410 ^ n786 ^ 1'b0 ;
  assign n18619 = n3510 & ~n18618 ;
  assign n18620 = n9766 | n13247 ;
  assign n18621 = n18620 ^ n7918 ^ 1'b0 ;
  assign n18622 = n2039 | n16484 ;
  assign n18623 = n18621 | n18622 ;
  assign n18624 = n551 & n18464 ;
  assign n18625 = ( n247 & n1086 ) | ( n247 & n14249 ) | ( n1086 & n14249 ) ;
  assign n18626 = n18625 ^ n12054 ^ n6241 ;
  assign n18627 = ~n4348 & n11184 ;
  assign n18628 = n2883 & n18627 ;
  assign n18629 = n18628 ^ n5057 ^ n1271 ;
  assign n18630 = ( n5569 & n9489 ) | ( n5569 & n18629 ) | ( n9489 & n18629 ) ;
  assign n18631 = n10126 & n18630 ;
  assign n18632 = n18631 ^ n7813 ^ 1'b0 ;
  assign n18633 = n5665 | n18632 ;
  assign n18634 = n6872 | n17313 ;
  assign n18635 = n18634 ^ n10327 ^ 1'b0 ;
  assign n18636 = ( n3797 & n12066 ) | ( n3797 & ~n18635 ) | ( n12066 & ~n18635 ) ;
  assign n18639 = n4189 & n11444 ;
  assign n18637 = n7170 & n10747 ;
  assign n18638 = x80 & ~n18637 ;
  assign n18640 = n18639 ^ n18638 ^ 1'b0 ;
  assign n18641 = n1535 | n18640 ;
  assign n18642 = ( n967 & n1454 ) | ( n967 & n7413 ) | ( n1454 & n7413 ) ;
  assign n18643 = n6219 & n18642 ;
  assign n18644 = n18643 ^ n1288 ^ 1'b0 ;
  assign n18645 = ( n7620 & n9573 ) | ( n7620 & n13577 ) | ( n9573 & n13577 ) ;
  assign n18646 = ~n13595 & n18645 ;
  assign n18647 = ~n18644 & n18646 ;
  assign n18649 = n231 | n7018 ;
  assign n18650 = n18649 ^ n4285 ^ 1'b0 ;
  assign n18648 = n3155 ^ n1779 ^ 1'b0 ;
  assign n18651 = n18650 ^ n18648 ^ 1'b0 ;
  assign n18652 = n3781 | n18651 ;
  assign n18653 = n3557 | n3845 ;
  assign n18654 = n18653 ^ n1730 ^ 1'b0 ;
  assign n18655 = ( x69 & n3220 ) | ( x69 & ~n6519 ) | ( n3220 & ~n6519 ) ;
  assign n18656 = n5594 | n10332 ;
  assign n18657 = n18656 ^ n3847 ^ 1'b0 ;
  assign n18658 = n18657 ^ n285 ^ 1'b0 ;
  assign n18659 = n15852 & ~n18658 ;
  assign n18660 = ~n8617 & n18659 ;
  assign n18661 = ( n7882 & n9840 ) | ( n7882 & n18660 ) | ( n9840 & n18660 ) ;
  assign n18662 = n1627 & n5507 ;
  assign n18665 = n9881 ^ n7150 ^ n6348 ;
  assign n18666 = n18665 ^ n10800 ^ 1'b0 ;
  assign n18663 = n18044 ^ n17564 ^ n11752 ;
  assign n18664 = n6056 | n18663 ;
  assign n18667 = n18666 ^ n18664 ^ 1'b0 ;
  assign n18669 = n17878 ^ n5786 ^ 1'b0 ;
  assign n18670 = ~n3765 & n15748 ;
  assign n18671 = n18670 ^ n12516 ^ 1'b0 ;
  assign n18672 = ~n18669 & n18671 ;
  assign n18668 = n12433 | n14708 ;
  assign n18673 = n18672 ^ n18668 ^ 1'b0 ;
  assign n18674 = n11055 & ~n18673 ;
  assign n18675 = n18674 ^ n11021 ^ 1'b0 ;
  assign n18676 = n1721 | n11340 ;
  assign n18677 = n2843 | n18676 ;
  assign n18678 = n16707 ^ n4562 ^ 1'b0 ;
  assign n18679 = n2956 & ~n7792 ;
  assign n18680 = n18679 ^ n9551 ^ 1'b0 ;
  assign n18681 = n18678 | n18680 ;
  assign n18682 = n2932 | n6561 ;
  assign n18683 = n18682 ^ n4851 ^ n1062 ;
  assign n18684 = n3000 | n10579 ;
  assign n18685 = n8515 & ~n18684 ;
  assign n18686 = ( ~n3228 & n3878 ) | ( ~n3228 & n18685 ) | ( n3878 & n18685 ) ;
  assign n18687 = n977 | n1106 ;
  assign n18688 = n18687 ^ n8089 ^ n6104 ;
  assign n18689 = n4954 | n6034 ;
  assign n18690 = n18689 ^ n6261 ^ 1'b0 ;
  assign n18691 = n4348 & ~n18690 ;
  assign n18692 = ~n15837 & n15930 ;
  assign n18693 = n18692 ^ n14651 ^ 1'b0 ;
  assign n18694 = n3216 ^ n917 ^ 1'b0 ;
  assign n18695 = n18693 | n18694 ;
  assign n18697 = n2234 & ~n8093 ;
  assign n18698 = n18697 ^ n3826 ^ 1'b0 ;
  assign n18696 = n1139 & ~n6876 ;
  assign n18699 = n18698 ^ n18696 ^ 1'b0 ;
  assign n18700 = ( n5446 & ~n16245 ) | ( n5446 & n18699 ) | ( ~n16245 & n18699 ) ;
  assign n18701 = n15284 ^ n4268 ^ 1'b0 ;
  assign n18702 = ~n4567 & n18701 ;
  assign n18703 = n6914 & n18702 ;
  assign n18704 = n18703 ^ n16499 ^ 1'b0 ;
  assign n18705 = n14154 ^ n3557 ^ 1'b0 ;
  assign n18706 = n11396 ^ n5387 ^ n166 ;
  assign n18707 = ( n2755 & n18091 ) | ( n2755 & ~n18706 ) | ( n18091 & ~n18706 ) ;
  assign n18708 = ( n15638 & n18705 ) | ( n15638 & n18707 ) | ( n18705 & n18707 ) ;
  assign n18709 = n496 | n2544 ;
  assign n18710 = ~n5696 & n18709 ;
  assign n18711 = n18710 ^ n6196 ^ 1'b0 ;
  assign n18712 = ( ~n3835 & n11227 ) | ( ~n3835 & n13724 ) | ( n11227 & n13724 ) ;
  assign n18713 = n5069 | n6046 ;
  assign n18714 = n18712 & ~n18713 ;
  assign n18715 = n10420 | n18714 ;
  assign n18716 = n9282 & ~n18715 ;
  assign n18717 = n13901 ^ n4426 ^ 1'b0 ;
  assign n18718 = n5580 ^ n2275 ^ 1'b0 ;
  assign n18719 = n1849 & n18718 ;
  assign n18720 = n12927 ^ n1150 ^ 1'b0 ;
  assign n18721 = n7970 ^ n6479 ^ n5365 ;
  assign n18722 = n18721 ^ n4845 ^ 1'b0 ;
  assign n18723 = n18722 ^ n11115 ^ n791 ;
  assign n18724 = n2166 ^ n1089 ^ 1'b0 ;
  assign n18725 = n3670 & n18724 ;
  assign n18726 = n280 ^ x14 ^ 1'b0 ;
  assign n18727 = n18726 ^ n10126 ^ 1'b0 ;
  assign n18728 = n1257 & n18727 ;
  assign n18729 = ~n7332 & n18728 ;
  assign n18730 = n1521 & n18729 ;
  assign n18731 = n8657 ^ n7238 ^ 1'b0 ;
  assign n18732 = n6701 & ~n18731 ;
  assign n18733 = n18732 ^ n1281 ^ 1'b0 ;
  assign n18734 = ~n13002 & n15324 ;
  assign n18735 = n4562 & n7503 ;
  assign n18736 = n18735 ^ n1017 ^ 1'b0 ;
  assign n18737 = n17851 & ~n18736 ;
  assign n18738 = x68 | n11179 ;
  assign n18739 = n5463 | n6658 ;
  assign n18740 = n18739 ^ n7402 ^ n4664 ;
  assign n18741 = ( ~n2089 & n5389 ) | ( ~n2089 & n5971 ) | ( n5389 & n5971 ) ;
  assign n18742 = ~n6632 & n18741 ;
  assign n18743 = ( ~n1263 & n12412 ) | ( ~n1263 & n15629 ) | ( n12412 & n15629 ) ;
  assign n18744 = ~n5631 & n18743 ;
  assign n18745 = n12717 & n18744 ;
  assign n18746 = n12676 ^ n3414 ^ 1'b0 ;
  assign n18747 = n18746 ^ n18548 ^ n1795 ;
  assign n18748 = n12779 | n18747 ;
  assign n18749 = n18745 & ~n18748 ;
  assign n18750 = n9496 | n13675 ;
  assign n18751 = ( n2552 & ~n4388 ) | ( n2552 & n17390 ) | ( ~n4388 & n17390 ) ;
  assign n18752 = n6633 & n11225 ;
  assign n18753 = ( n6388 & n15544 ) | ( n6388 & ~n18752 ) | ( n15544 & ~n18752 ) ;
  assign n18754 = n8609 & ~n18753 ;
  assign n18755 = ~n11206 & n18754 ;
  assign n18756 = n188 & n6171 ;
  assign n18757 = n8360 ^ n3585 ^ 1'b0 ;
  assign n18761 = n18383 ^ n6072 ^ 1'b0 ;
  assign n18762 = n14186 | n18761 ;
  assign n18763 = ( ~n469 & n10168 ) | ( ~n469 & n18762 ) | ( n10168 & n18762 ) ;
  assign n18760 = n12308 & ~n15950 ;
  assign n18758 = n521 ^ x50 ^ 1'b0 ;
  assign n18759 = n1327 & n18758 ;
  assign n18764 = n18763 ^ n18760 ^ n18759 ;
  assign n18765 = n7160 ^ n2117 ^ n1761 ;
  assign n18766 = n2824 & ~n18765 ;
  assign n18767 = ~n6741 & n18766 ;
  assign n18768 = n1588 ^ n1117 ^ 1'b0 ;
  assign n18769 = n18768 ^ n7851 ^ n507 ;
  assign n18770 = n3044 ^ n3016 ^ 1'b0 ;
  assign n18771 = n18770 ^ n12676 ^ 1'b0 ;
  assign n18772 = n18771 ^ n730 ^ 1'b0 ;
  assign n18773 = n2006 | n3172 ;
  assign n18774 = n2637 | n7701 ;
  assign n18775 = n18773 & n18774 ;
  assign n18776 = ~n18772 & n18775 ;
  assign n18777 = n8779 ^ n4407 ^ 1'b0 ;
  assign n18778 = n3265 ^ n2016 ^ 1'b0 ;
  assign n18779 = n6738 ^ n5861 ^ 1'b0 ;
  assign n18780 = n3901 | n10257 ;
  assign n18781 = n3696 & ~n18780 ;
  assign n18782 = n7305 & n18781 ;
  assign n18783 = ( n2912 & n12012 ) | ( n2912 & ~n18782 ) | ( n12012 & ~n18782 ) ;
  assign n18784 = n18779 | n18783 ;
  assign n18785 = n3357 ^ n1293 ^ 1'b0 ;
  assign n18786 = n18784 | n18785 ;
  assign n18787 = ~n12495 & n15298 ;
  assign n18788 = ~n4194 & n6877 ;
  assign n18789 = ~n4898 & n13432 ;
  assign n18790 = n18789 ^ n16996 ^ n1123 ;
  assign n18791 = n15443 | n15892 ;
  assign n18792 = n3103 & ~n5829 ;
  assign n18793 = n18792 ^ n14145 ^ 1'b0 ;
  assign n18797 = n17982 ^ n8341 ^ n5453 ;
  assign n18794 = n17365 ^ n1222 ^ 1'b0 ;
  assign n18795 = n18794 ^ n2117 ^ 1'b0 ;
  assign n18796 = n7787 | n18795 ;
  assign n18798 = n18797 ^ n18796 ^ 1'b0 ;
  assign n18799 = n5899 | n7850 ;
  assign n18800 = n18673 | n18799 ;
  assign n18801 = n336 & ~n4440 ;
  assign n18802 = n14265 & ~n18801 ;
  assign n18803 = n5069 & ~n12084 ;
  assign n18804 = ~n1485 & n10941 ;
  assign n18805 = n18804 ^ n11962 ^ 1'b0 ;
  assign n18806 = n13425 & n18805 ;
  assign n18807 = ~n7920 & n14407 ;
  assign n18809 = n4574 | n6504 ;
  assign n18810 = n18809 ^ n10622 ^ 1'b0 ;
  assign n18811 = ( ~n11768 & n14166 ) | ( ~n11768 & n18810 ) | ( n14166 & n18810 ) ;
  assign n18808 = n3179 & ~n7099 ;
  assign n18812 = n18811 ^ n18808 ^ 1'b0 ;
  assign n18813 = n1177 | n7393 ;
  assign n18814 = n18813 ^ n3182 ^ 1'b0 ;
  assign n18815 = n982 | n18814 ;
  assign n18816 = n13708 | n18815 ;
  assign n18817 = n4722 ^ n2304 ^ 1'b0 ;
  assign n18818 = ~n6760 & n18817 ;
  assign n18819 = n4563 & ~n12379 ;
  assign n18820 = ~n18818 & n18819 ;
  assign n18821 = n13090 | n18820 ;
  assign n18823 = ~n227 & n1713 ;
  assign n18822 = ~n5378 & n11421 ;
  assign n18824 = n18823 ^ n18822 ^ 1'b0 ;
  assign n18825 = n2922 & n5318 ;
  assign n18826 = ( ~n7619 & n9743 ) | ( ~n7619 & n18825 ) | ( n9743 & n18825 ) ;
  assign n18827 = n18191 ^ n10028 ^ 1'b0 ;
  assign n18828 = n17735 ^ n16528 ^ 1'b0 ;
  assign n18829 = ~n10437 & n18828 ;
  assign n18830 = n18314 ^ n4032 ^ 1'b0 ;
  assign n18831 = n3710 | n18830 ;
  assign n18832 = n5178 & n18831 ;
  assign n18833 = ~n295 & n6286 ;
  assign n18834 = n18833 ^ n5562 ^ 1'b0 ;
  assign n18835 = n11323 & n18834 ;
  assign n18836 = n18835 ^ n6456 ^ 1'b0 ;
  assign n18837 = n4221 ^ n590 ^ 1'b0 ;
  assign n18838 = ~n18836 & n18837 ;
  assign n18839 = ( n404 & n1436 ) | ( n404 & ~n18838 ) | ( n1436 & ~n18838 ) ;
  assign n18840 = ( n3412 & ~n13154 ) | ( n3412 & n13219 ) | ( ~n13154 & n13219 ) ;
  assign n18841 = n8212 & ~n18840 ;
  assign n18842 = ( n508 & ~n9086 ) | ( n508 & n18841 ) | ( ~n9086 & n18841 ) ;
  assign n18843 = n12312 ^ n150 ^ 1'b0 ;
  assign n18844 = n5076 & ~n18843 ;
  assign n18845 = n18844 ^ n18635 ^ 1'b0 ;
  assign n18846 = n9261 & n18845 ;
  assign n18847 = n18846 ^ n3195 ^ 1'b0 ;
  assign n18848 = n4499 & n18847 ;
  assign n18849 = n18848 ^ n10281 ^ n3513 ;
  assign n18850 = n359 & ~n6676 ;
  assign n18851 = n15504 ^ n3927 ^ 1'b0 ;
  assign n18852 = n4384 | n18851 ;
  assign n18853 = ~n404 & n2741 ;
  assign n18854 = ( x42 & n16114 ) | ( x42 & n18853 ) | ( n16114 & n18853 ) ;
  assign n18855 = n18854 ^ n12741 ^ x69 ;
  assign n18856 = ( ~n8900 & n14585 ) | ( ~n8900 & n15222 ) | ( n14585 & n15222 ) ;
  assign n18857 = n18856 ^ n2326 ^ 1'b0 ;
  assign n18858 = n3540 ^ n793 ^ 1'b0 ;
  assign n18859 = ( n13158 & n14680 ) | ( n13158 & ~n18858 ) | ( n14680 & ~n18858 ) ;
  assign n18860 = n11087 ^ n7604 ^ 1'b0 ;
  assign n18861 = ~n2562 & n18860 ;
  assign n18862 = n16063 ^ n7547 ^ 1'b0 ;
  assign n18863 = n6003 | n18862 ;
  assign n18864 = n2034 & ~n18863 ;
  assign n18865 = n9335 & n18864 ;
  assign n18866 = n11297 ^ n8956 ^ 1'b0 ;
  assign n18867 = n17352 ^ n13743 ^ 1'b0 ;
  assign n18868 = n6899 ^ n791 ^ 1'b0 ;
  assign n18869 = n16650 ^ n3130 ^ 1'b0 ;
  assign n18870 = n9413 | n18869 ;
  assign n18871 = n10414 ^ n6607 ^ n1271 ;
  assign n18872 = n18871 ^ n1235 ^ 1'b0 ;
  assign n18873 = n18870 | n18872 ;
  assign n18874 = ~n9923 & n18526 ;
  assign n18875 = n18874 ^ n1286 ^ 1'b0 ;
  assign n18876 = n15654 ^ n8549 ^ 1'b0 ;
  assign n18877 = n3662 & ~n18876 ;
  assign n18878 = n18877 ^ n10796 ^ 1'b0 ;
  assign n18879 = n3313 & n18878 ;
  assign n18880 = n1422 & n2570 ;
  assign n18881 = ~n2570 & n18880 ;
  assign n18882 = n10931 & ~n18881 ;
  assign n18883 = n5123 & n18882 ;
  assign n18884 = n824 & n11518 ;
  assign n18885 = n18883 | n18884 ;
  assign n18887 = n5579 ^ n2236 ^ 1'b0 ;
  assign n18888 = ( ~n3808 & n6599 ) | ( ~n3808 & n18887 ) | ( n6599 & n18887 ) ;
  assign n18886 = n387 & ~n8835 ;
  assign n18889 = n18888 ^ n18886 ^ 1'b0 ;
  assign n18890 = n13733 ^ n10221 ^ 1'b0 ;
  assign n18891 = n1519 | n18890 ;
  assign n18892 = n18891 ^ n12456 ^ 1'b0 ;
  assign n18893 = n18889 & n18892 ;
  assign n18894 = n15019 ^ n11343 ^ 1'b0 ;
  assign n18895 = n12632 ^ n920 ^ 1'b0 ;
  assign n18896 = n165 | n5046 ;
  assign n18897 = n2325 & n18896 ;
  assign n18898 = n18897 ^ n7174 ^ 1'b0 ;
  assign n18899 = ~n2521 & n13774 ;
  assign n18900 = n2521 & n18899 ;
  assign n18901 = n231 & n18900 ;
  assign n18902 = n1644 & n18901 ;
  assign n18903 = n18902 ^ n2740 ^ 1'b0 ;
  assign n18904 = ~n4874 & n15928 ;
  assign n18905 = n18904 ^ n8992 ^ 1'b0 ;
  assign n18906 = ( n13428 & ~n13903 ) | ( n13428 & n15340 ) | ( ~n13903 & n15340 ) ;
  assign n18907 = n5078 | n11008 ;
  assign n18908 = ~n2642 & n5216 ;
  assign n18909 = ~n2839 & n18908 ;
  assign n18910 = n18909 ^ n5822 ^ n5285 ;
  assign n18911 = n18910 ^ n2450 ^ 1'b0 ;
  assign n18912 = n1561 & n3059 ;
  assign n18913 = n18911 & n18912 ;
  assign n18914 = n6742 ^ n6367 ^ 1'b0 ;
  assign n18915 = n11454 & ~n18914 ;
  assign n18916 = ~n8120 & n18915 ;
  assign n18917 = n11043 & n18916 ;
  assign n18918 = ~n4297 & n4984 ;
  assign n18919 = ~n12411 & n18918 ;
  assign n18920 = n1765 & ~n18919 ;
  assign n18921 = n2197 & ~n14889 ;
  assign n18922 = n3265 | n11829 ;
  assign n18924 = n6330 ^ n431 ^ 1'b0 ;
  assign n18925 = n18924 ^ n12541 ^ 1'b0 ;
  assign n18926 = n11423 & ~n18925 ;
  assign n18923 = n2750 | n5001 ;
  assign n18927 = n18926 ^ n18923 ^ 1'b0 ;
  assign n18928 = n3127 & n5517 ;
  assign n18929 = n2515 & n18928 ;
  assign n18930 = n7578 & n14015 ;
  assign n18931 = n10170 & n18930 ;
  assign n18932 = n18929 | n18931 ;
  assign n18935 = n1644 & n7899 ;
  assign n18936 = n1658 | n18935 ;
  assign n18937 = n18936 ^ n12814 ^ 1'b0 ;
  assign n18933 = n6911 & n8371 ;
  assign n18934 = n18933 ^ n5613 ^ 1'b0 ;
  assign n18938 = n18937 ^ n18934 ^ n10997 ;
  assign n18939 = n4042 & ~n12351 ;
  assign n18940 = n18938 & n18939 ;
  assign n18941 = n5340 & n14756 ;
  assign n18942 = n15156 & n16332 ;
  assign n18943 = n17269 ^ n4281 ^ 1'b0 ;
  assign n18946 = ~n4344 & n11708 ;
  assign n18947 = n18946 ^ n3065 ^ 1'b0 ;
  assign n18944 = n8073 & ~n9935 ;
  assign n18945 = ( n1860 & n3200 ) | ( n1860 & ~n18944 ) | ( n3200 & ~n18944 ) ;
  assign n18948 = n18947 ^ n18945 ^ 1'b0 ;
  assign n18949 = n5429 | n15433 ;
  assign n18950 = n18949 ^ n636 ^ 1'b0 ;
  assign n18951 = n7626 ^ n7411 ^ 1'b0 ;
  assign n18952 = n2596 | n18951 ;
  assign n18953 = n18950 | n18952 ;
  assign n18954 = n18953 ^ n15223 ^ n1021 ;
  assign n18955 = n8661 | n12853 ;
  assign n18956 = n18955 ^ n1240 ^ 1'b0 ;
  assign n18957 = n18956 ^ n8771 ^ x67 ;
  assign n18958 = n9255 ^ n5546 ^ n2841 ;
  assign n18959 = x30 & n3417 ;
  assign n18960 = ~n18958 & n18959 ;
  assign n18961 = n8530 | n14647 ;
  assign n18962 = n7455 & ~n18961 ;
  assign n18963 = n18960 & n18962 ;
  assign n18964 = n5316 | n18963 ;
  assign n18965 = n18964 ^ n9396 ^ 1'b0 ;
  assign n18966 = n1655 & ~n5338 ;
  assign n18967 = n18966 ^ n17146 ^ 1'b0 ;
  assign n18970 = n2033 ^ n799 ^ 1'b0 ;
  assign n18971 = n8854 & n18970 ;
  assign n18972 = n2713 & ~n12127 ;
  assign n18973 = ~n18971 & n18972 ;
  assign n18968 = n16857 ^ n1996 ^ 1'b0 ;
  assign n18969 = n17003 & ~n18968 ;
  assign n18974 = n18973 ^ n18969 ^ 1'b0 ;
  assign n18975 = ~n9583 & n15229 ;
  assign n18976 = n10381 & n18975 ;
  assign n18977 = n377 & n5930 ;
  assign n18978 = n8046 ^ n6319 ^ 1'b0 ;
  assign n18979 = n5149 | n18978 ;
  assign n18980 = n716 | n18979 ;
  assign n18981 = ~n277 & n3055 ;
  assign n18982 = n18981 ^ n14869 ^ n2551 ;
  assign n18983 = n395 | n5691 ;
  assign n18984 = n2850 & ~n18983 ;
  assign n18985 = n8667 & ~n17733 ;
  assign n18986 = n17733 & n18985 ;
  assign n18987 = ( n18982 & ~n18984 ) | ( n18982 & n18986 ) | ( ~n18984 & n18986 ) ;
  assign n18988 = n12817 ^ n11620 ^ 1'b0 ;
  assign n18989 = n707 & ~n15223 ;
  assign n18990 = n11280 ^ n10267 ^ 1'b0 ;
  assign n18991 = n6138 & n13575 ;
  assign n18992 = n3876 & n18991 ;
  assign n18993 = n18992 ^ n8835 ^ n8035 ;
  assign n18995 = n11062 ^ n4508 ^ 1'b0 ;
  assign n18996 = n18133 | n18995 ;
  assign n18994 = n510 | n5910 ;
  assign n18997 = n18996 ^ n18994 ^ n7717 ;
  assign n18998 = n12893 | n15022 ;
  assign n18999 = n18896 ^ n5808 ^ 1'b0 ;
  assign n19000 = n336 & n502 ;
  assign n19001 = n9341 & n19000 ;
  assign n19002 = n1561 ^ n261 ^ 1'b0 ;
  assign n19003 = n1958 ^ n744 ^ 1'b0 ;
  assign n19004 = n19002 & ~n19003 ;
  assign n19005 = n17084 ^ n4491 ^ 1'b0 ;
  assign n19006 = n19005 ^ n16480 ^ 1'b0 ;
  assign n19007 = ( ~n696 & n3518 ) | ( ~n696 & n4188 ) | ( n3518 & n4188 ) ;
  assign n19008 = n7072 & n10308 ;
  assign n19009 = ~n19007 & n19008 ;
  assign n19010 = n13942 | n18994 ;
  assign n19011 = n11298 ^ n10127 ^ 1'b0 ;
  assign n19012 = n409 & ~n1044 ;
  assign n19013 = n19012 ^ n10916 ^ n10649 ;
  assign n19014 = n1710 & n5330 ;
  assign n19015 = n2377 & n19014 ;
  assign n19016 = n19015 ^ n10586 ^ n5084 ;
  assign n19017 = n11118 ^ n3200 ^ 1'b0 ;
  assign n19018 = n19016 | n19017 ;
  assign n19019 = n129 & n10521 ;
  assign n19020 = n17794 | n19019 ;
  assign n19021 = n19020 ^ n14101 ^ 1'b0 ;
  assign n19022 = n11690 & ~n19021 ;
  assign n19023 = ~n2726 & n6166 ;
  assign n19024 = n19023 ^ x23 ^ 1'b0 ;
  assign n19025 = n17951 & ~n19024 ;
  assign n19026 = n7379 | n11653 ;
  assign n19027 = ( n7967 & n10111 ) | ( n7967 & ~n19026 ) | ( n10111 & ~n19026 ) ;
  assign n19033 = n8361 ^ n6846 ^ n5463 ;
  assign n19029 = n3111 | n3403 ;
  assign n19030 = n19029 ^ n11055 ^ 1'b0 ;
  assign n19028 = n14338 & ~n17723 ;
  assign n19031 = n19030 ^ n19028 ^ n6543 ;
  assign n19032 = n6372 | n19031 ;
  assign n19034 = n19033 ^ n19032 ^ 1'b0 ;
  assign n19035 = n10605 ^ n9374 ^ n1899 ;
  assign n19036 = n19035 ^ n5091 ^ 1'b0 ;
  assign n19037 = ( ~x100 & n10764 ) | ( ~x100 & n19036 ) | ( n10764 & n19036 ) ;
  assign n19038 = n12457 ^ n5669 ^ 1'b0 ;
  assign n19039 = n19037 & ~n19038 ;
  assign n19040 = n10627 ^ n234 ^ 1'b0 ;
  assign n19041 = ~n9829 & n19040 ;
  assign n19042 = n1520 & n9948 ;
  assign n19043 = ~n1581 & n19042 ;
  assign n19044 = n11993 ^ n2688 ^ 1'b0 ;
  assign n19045 = ~n5565 & n6428 ;
  assign n19046 = n13869 ^ n4397 ^ 1'b0 ;
  assign n19047 = ~n4580 & n19046 ;
  assign n19048 = ( n3803 & n19045 ) | ( n3803 & ~n19047 ) | ( n19045 & ~n19047 ) ;
  assign n19049 = n8169 | n15822 ;
  assign n19050 = n12127 | n19049 ;
  assign n19051 = n1553 | n5664 ;
  assign n19052 = n12428 ^ n6400 ^ n6071 ;
  assign n19058 = n10855 ^ n10481 ^ 1'b0 ;
  assign n19053 = n8818 ^ n4100 ^ n3142 ;
  assign n19054 = n678 & n11067 ;
  assign n19055 = n19054 ^ n2850 ^ 1'b0 ;
  assign n19056 = ~n19053 & n19055 ;
  assign n19057 = n19056 ^ n18773 ^ 1'b0 ;
  assign n19059 = n19058 ^ n19057 ^ n9456 ;
  assign n19060 = n18322 ^ n17236 ^ 1'b0 ;
  assign n19061 = ~n3967 & n19060 ;
  assign n19062 = n19061 ^ n12759 ^ 1'b0 ;
  assign n19064 = ~n7934 & n17174 ;
  assign n19063 = n7726 | n7876 ;
  assign n19065 = n19064 ^ n19063 ^ 1'b0 ;
  assign n19066 = n3738 & ~n4303 ;
  assign n19067 = n9968 ^ n5945 ^ 1'b0 ;
  assign n19068 = n3426 & n19067 ;
  assign n19069 = ( n2032 & n13743 ) | ( n2032 & n15271 ) | ( n13743 & n15271 ) ;
  assign n19070 = ~n1511 & n2464 ;
  assign n19071 = ~n19069 & n19070 ;
  assign n19072 = n16876 ^ n1151 ^ n243 ;
  assign n19073 = ( n707 & ~n10693 ) | ( n707 & n19072 ) | ( ~n10693 & n19072 ) ;
  assign n19074 = n7218 ^ n4950 ^ 1'b0 ;
  assign n19075 = n6884 ^ n3634 ^ n2437 ;
  assign n19076 = ( n4368 & ~n6657 ) | ( n4368 & n19075 ) | ( ~n6657 & n19075 ) ;
  assign n19077 = ( n9210 & n12490 ) | ( n9210 & n19076 ) | ( n12490 & n19076 ) ;
  assign n19078 = x41 & n9949 ;
  assign n19079 = n11326 ^ n7025 ^ 1'b0 ;
  assign n19080 = n7305 & n19079 ;
  assign n19081 = n3176 & ~n6020 ;
  assign n19082 = n6209 & n19081 ;
  assign n19083 = n17961 ^ n16944 ^ 1'b0 ;
  assign n19084 = n2945 | n17794 ;
  assign n19085 = n19084 ^ n17281 ^ n16124 ;
  assign n19086 = n3614 ^ n1409 ^ 1'b0 ;
  assign n19087 = ~n2223 & n19086 ;
  assign n19088 = n4639 ^ x25 ^ 1'b0 ;
  assign n19089 = n19087 & ~n19088 ;
  assign n19090 = ~n10622 & n19089 ;
  assign n19091 = n1412 & n19090 ;
  assign n19092 = n6713 ^ n3316 ^ 1'b0 ;
  assign n19093 = n8206 & ~n19092 ;
  assign n19094 = n19093 ^ n7123 ^ n618 ;
  assign n19095 = ( ~n956 & n6430 ) | ( ~n956 & n19094 ) | ( n6430 & n19094 ) ;
  assign n19096 = ( n872 & n7328 ) | ( n872 & ~n19095 ) | ( n7328 & ~n19095 ) ;
  assign n19097 = n8502 | n8765 ;
  assign n19098 = n13066 | n19097 ;
  assign n19099 = n19098 ^ n7124 ^ 1'b0 ;
  assign n19100 = n1718 & n8849 ;
  assign n19101 = n19100 ^ n16847 ^ 1'b0 ;
  assign n19102 = ~n5278 & n16014 ;
  assign n19106 = ( n1833 & n2860 ) | ( n1833 & n9890 ) | ( n2860 & n9890 ) ;
  assign n19104 = n13034 ^ n731 ^ 1'b0 ;
  assign n19105 = n3547 | n19104 ;
  assign n19107 = n19106 ^ n19105 ^ 1'b0 ;
  assign n19108 = ~n6573 & n19107 ;
  assign n19103 = n7047 | n8991 ;
  assign n19109 = n19108 ^ n19103 ^ 1'b0 ;
  assign n19110 = n7812 & ~n18709 ;
  assign n19111 = n7718 ^ n4555 ^ 1'b0 ;
  assign n19112 = n15127 & n19111 ;
  assign n19113 = ~n19110 & n19112 ;
  assign n19114 = n19109 & ~n19113 ;
  assign n19115 = ~n9761 & n19114 ;
  assign n19116 = n8040 ^ n7558 ^ 1'b0 ;
  assign n19117 = n2839 ^ n1046 ^ 1'b0 ;
  assign n19118 = n6250 & ~n19117 ;
  assign n19119 = x27 & n3959 ;
  assign n19120 = ~n19118 & n19119 ;
  assign n19121 = n19120 ^ n6801 ^ 1'b0 ;
  assign n19122 = n18539 & ~n19121 ;
  assign n19123 = n18950 ^ n6876 ^ n3487 ;
  assign n19124 = n19074 ^ n11219 ^ 1'b0 ;
  assign n19125 = n19123 & ~n19124 ;
  assign n19126 = ~n2682 & n3858 ;
  assign n19127 = n19126 ^ n8132 ^ 1'b0 ;
  assign n19128 = n14792 ^ n9913 ^ 1'b0 ;
  assign n19129 = x74 & n16849 ;
  assign n19130 = ( ~n3516 & n12000 ) | ( ~n3516 & n13593 ) | ( n12000 & n13593 ) ;
  assign n19131 = n13533 & n19130 ;
  assign n19132 = n13691 & n19131 ;
  assign n19133 = ~n3113 & n6104 ;
  assign n19134 = n11539 ^ n1418 ^ 1'b0 ;
  assign n19135 = n18858 ^ n5687 ^ 1'b0 ;
  assign n19136 = n19135 ^ n7683 ^ 1'b0 ;
  assign n19137 = ~n2547 & n19136 ;
  assign n19138 = n11398 ^ n5183 ^ 1'b0 ;
  assign n19139 = n403 & ~n19138 ;
  assign n19140 = n10010 ^ n8935 ^ n1258 ;
  assign n19141 = n4624 ^ n2818 ^ 1'b0 ;
  assign n19142 = n10266 ^ n2839 ^ 1'b0 ;
  assign n19143 = n305 ^ n299 ^ 1'b0 ;
  assign n19144 = ~n12494 & n19143 ;
  assign n19145 = n19142 & n19144 ;
  assign n19146 = n9857 ^ n6399 ^ 1'b0 ;
  assign n19147 = n7445 ^ n4504 ^ 1'b0 ;
  assign n19148 = n4195 | n19147 ;
  assign n19149 = n7095 & n19148 ;
  assign n19150 = n4460 ^ n1743 ^ 1'b0 ;
  assign n19151 = n19149 | n19150 ;
  assign n19152 = n5085 & n10348 ;
  assign n19153 = n19152 ^ n12905 ^ 1'b0 ;
  assign n19154 = n13429 ^ n4017 ^ 1'b0 ;
  assign n19155 = n19153 & n19154 ;
  assign n19156 = n15663 & n19155 ;
  assign n19157 = n15582 ^ n7583 ^ n986 ;
  assign n19158 = n7887 ^ n4626 ^ 1'b0 ;
  assign n19159 = n2193 & n11631 ;
  assign n19160 = n19159 ^ n14096 ^ 1'b0 ;
  assign n19161 = n9310 ^ n840 ^ 1'b0 ;
  assign n19162 = n18939 ^ n9233 ^ 1'b0 ;
  assign n19163 = ~n19161 & n19162 ;
  assign n19165 = ( ~n2289 & n3842 ) | ( ~n2289 & n6858 ) | ( n3842 & n6858 ) ;
  assign n19164 = ~n3939 & n5039 ;
  assign n19166 = n19165 ^ n19164 ^ 1'b0 ;
  assign n19167 = ~n1358 & n8869 ;
  assign n19168 = n12195 & n15118 ;
  assign n19169 = n1432 ^ n635 ^ 1'b0 ;
  assign n19170 = ~n6225 & n14637 ;
  assign n19171 = n5144 & n9274 ;
  assign n19172 = n13649 & n19171 ;
  assign n19173 = n10847 & n12205 ;
  assign n19174 = n19173 ^ n7925 ^ 1'b0 ;
  assign n19175 = n1330 & ~n8491 ;
  assign n19176 = ~n770 & n19175 ;
  assign n19177 = x125 & n13244 ;
  assign n19178 = n19177 ^ n9152 ^ 1'b0 ;
  assign n19179 = ~n19176 & n19178 ;
  assign n19180 = ~n8091 & n19179 ;
  assign n19181 = n8778 & n19180 ;
  assign n19182 = n4068 & n19181 ;
  assign n19183 = ~n6948 & n9085 ;
  assign n19184 = n19183 ^ n12544 ^ n5221 ;
  assign n19185 = ( n8606 & n13993 ) | ( n8606 & n19184 ) | ( n13993 & n19184 ) ;
  assign n19186 = n18117 ^ n14808 ^ n13172 ;
  assign n19187 = n12660 ^ n9862 ^ n9251 ;
  assign n19188 = n14166 & n19187 ;
  assign n19189 = n19188 ^ n3016 ^ 1'b0 ;
  assign n19190 = n13908 & n19189 ;
  assign n19191 = n19190 ^ n16357 ^ 1'b0 ;
  assign n19193 = n630 & n16199 ;
  assign n19192 = n2401 & n6251 ;
  assign n19194 = n19193 ^ n19192 ^ 1'b0 ;
  assign n19195 = n16814 ^ n10772 ^ 1'b0 ;
  assign n19196 = n6386 & ~n19195 ;
  assign n19197 = n19196 ^ n3714 ^ 1'b0 ;
  assign n19198 = n19197 ^ n9659 ^ 1'b0 ;
  assign n19199 = ~n2627 & n7124 ;
  assign n19200 = n19199 ^ n9014 ^ 1'b0 ;
  assign n19202 = n2066 | n9018 ;
  assign n19203 = n12546 & ~n19202 ;
  assign n19201 = n2222 | n9728 ;
  assign n19204 = n19203 ^ n19201 ^ 1'b0 ;
  assign n19205 = ~n5092 & n8735 ;
  assign n19206 = n9874 & n19205 ;
  assign n19207 = n5866 & ~n19206 ;
  assign n19208 = ~n12881 & n19207 ;
  assign n19209 = ~n13758 & n19208 ;
  assign n19210 = n19209 ^ n4935 ^ 1'b0 ;
  assign n19211 = ~n19204 & n19210 ;
  assign n19212 = n19211 ^ n10874 ^ 1'b0 ;
  assign n19213 = n5342 ^ n4759 ^ n3625 ;
  assign n19214 = n13910 & ~n17111 ;
  assign n19215 = n2071 ^ n983 ^ 1'b0 ;
  assign n19216 = n1188 | n19215 ;
  assign n19217 = n2199 | n19216 ;
  assign n19218 = n19216 & ~n19217 ;
  assign n19219 = x31 & ~n997 ;
  assign n19220 = ~x31 & n19219 ;
  assign n19221 = n19218 & ~n19220 ;
  assign n19222 = ~n5205 & n19221 ;
  assign n19223 = n2785 & n19222 ;
  assign n19224 = n12853 ^ n1375 ^ 1'b0 ;
  assign n19225 = ~n19223 & n19224 ;
  assign n19227 = n764 & ~n5659 ;
  assign n19228 = ~n764 & n19227 ;
  assign n19229 = n4217 | n19228 ;
  assign n19230 = n4217 & ~n19229 ;
  assign n19231 = n11370 & n19230 ;
  assign n19232 = n6819 & ~n19231 ;
  assign n19226 = ( ~n623 & n6213 ) | ( ~n623 & n9371 ) | ( n6213 & n9371 ) ;
  assign n19233 = n19232 ^ n19226 ^ 1'b0 ;
  assign n19234 = n19225 & n19233 ;
  assign n19235 = n2011 | n2988 ;
  assign n19236 = n19235 ^ n15651 ^ n3444 ;
  assign n19237 = ~n18864 & n19236 ;
  assign n19238 = n3559 ^ n2966 ^ 1'b0 ;
  assign n19239 = n14859 & ~n19238 ;
  assign n19241 = n944 & ~n9887 ;
  assign n19240 = n4921 & ~n12759 ;
  assign n19242 = n19241 ^ n19240 ^ 1'b0 ;
  assign n19243 = n19242 ^ n484 ^ 1'b0 ;
  assign n19244 = n19243 ^ n13872 ^ n8491 ;
  assign n19245 = n14373 ^ n4380 ^ 1'b0 ;
  assign n19246 = ~n5633 & n19245 ;
  assign n19247 = n9830 ^ n8143 ^ 1'b0 ;
  assign n19248 = n19246 & n19247 ;
  assign n19249 = n9274 ^ n1771 ^ 1'b0 ;
  assign n19250 = ~n7012 & n11609 ;
  assign n19251 = n7778 ^ n316 ^ 1'b0 ;
  assign n19252 = n11627 & n19251 ;
  assign n19253 = n14328 ^ n2369 ^ 1'b0 ;
  assign n19254 = n12728 ^ n7959 ^ 1'b0 ;
  assign n19255 = ~n12905 & n19254 ;
  assign n19256 = n7662 | n10968 ;
  assign n19257 = n19256 ^ n16041 ^ 1'b0 ;
  assign n19258 = n8254 ^ n6751 ^ n5731 ;
  assign n19259 = n1617 | n2143 ;
  assign n19260 = n19258 | n19259 ;
  assign n19261 = n3625 & ~n4397 ;
  assign n19262 = ~n14426 & n19261 ;
  assign n19265 = n18825 ^ n6993 ^ 1'b0 ;
  assign n19266 = n3775 | n19265 ;
  assign n19267 = n19266 ^ n14924 ^ 1'b0 ;
  assign n19263 = n13589 ^ n2000 ^ 1'b0 ;
  assign n19264 = ( n12383 & n15734 ) | ( n12383 & ~n19263 ) | ( n15734 & ~n19263 ) ;
  assign n19268 = n19267 ^ n19264 ^ 1'b0 ;
  assign n19269 = n9907 ^ n6489 ^ 1'b0 ;
  assign n19270 = n19269 ^ n9096 ^ 1'b0 ;
  assign n19271 = ( n4087 & n4391 ) | ( n4087 & ~n12412 ) | ( n4391 & ~n12412 ) ;
  assign n19272 = n19271 ^ n18503 ^ 1'b0 ;
  assign n19273 = n17510 & n19272 ;
  assign n19274 = n8013 ^ n636 ^ 1'b0 ;
  assign n19275 = n19273 & ~n19274 ;
  assign n19276 = n2852 ^ n2340 ^ 1'b0 ;
  assign n19277 = n5371 ^ n369 ^ 1'b0 ;
  assign n19278 = n13551 | n19277 ;
  assign n19279 = ( n5001 & ~n11222 ) | ( n5001 & n19278 ) | ( ~n11222 & n19278 ) ;
  assign n19280 = n8034 ^ n6940 ^ n5119 ;
  assign n19281 = n4439 ^ x110 ^ 1'b0 ;
  assign n19282 = n13882 & ~n19281 ;
  assign n19283 = n1245 | n5664 ;
  assign n19284 = n13956 & ~n19283 ;
  assign n19285 = n12061 & n19284 ;
  assign n19286 = ~n14292 & n18693 ;
  assign n19287 = n18648 ^ n1409 ^ 1'b0 ;
  assign n19288 = ~n9775 & n19287 ;
  assign n19289 = n11061 & n19288 ;
  assign n19290 = n4357 & ~n14659 ;
  assign n19291 = n19290 ^ n6279 ^ 1'b0 ;
  assign n19292 = ~n2081 & n8122 ;
  assign n19293 = ~n12761 & n13807 ;
  assign n19294 = ~n19292 & n19293 ;
  assign n19295 = n12094 & n18325 ;
  assign n19296 = ~n11781 & n19295 ;
  assign n19297 = ~n2449 & n5463 ;
  assign n19298 = n7974 ^ n2637 ^ 1'b0 ;
  assign n19299 = n3130 & n5216 ;
  assign n19300 = n19299 ^ n5464 ^ 1'b0 ;
  assign n19301 = n6547 ^ n3551 ^ 1'b0 ;
  assign n19302 = n1275 & n19301 ;
  assign n19303 = n19302 ^ n4183 ^ 1'b0 ;
  assign n19304 = n15179 & ~n19303 ;
  assign n19305 = n4640 & ~n8378 ;
  assign n19306 = ~n8389 & n19305 ;
  assign n19307 = n10871 & n11226 ;
  assign n19308 = n19306 & n19307 ;
  assign n19310 = n10058 ^ n7873 ^ 1'b0 ;
  assign n19309 = n4550 & ~n13529 ;
  assign n19311 = n19310 ^ n19309 ^ 1'b0 ;
  assign n19312 = ( n1694 & n3205 ) | ( n1694 & n18527 ) | ( n3205 & n18527 ) ;
  assign n19313 = n15337 ^ n1893 ^ 1'b0 ;
  assign n19314 = x16 | n12188 ;
  assign n19315 = ~n8820 & n11978 ;
  assign n19316 = n1272 & n19315 ;
  assign n19317 = ( n1827 & n3468 ) | ( n1827 & ~n4246 ) | ( n3468 & ~n4246 ) ;
  assign n19318 = n19317 ^ n8584 ^ n914 ;
  assign n19319 = n19064 & n19318 ;
  assign n19320 = n19316 & n19319 ;
  assign n19321 = n5950 ^ n663 ^ 1'b0 ;
  assign n19322 = n2756 & ~n19321 ;
  assign n19323 = n12785 ^ n6529 ^ 1'b0 ;
  assign n19324 = n1251 & ~n11460 ;
  assign n19325 = ~n8443 & n19324 ;
  assign n19326 = ( n3954 & n6543 ) | ( n3954 & ~n19325 ) | ( n6543 & ~n19325 ) ;
  assign n19327 = n8377 ^ n2622 ^ 1'b0 ;
  assign n19328 = ~n8341 & n19327 ;
  assign n19329 = n5443 & n11092 ;
  assign n19330 = n17653 ^ n1160 ^ 1'b0 ;
  assign n19331 = n8681 ^ n2389 ^ 1'b0 ;
  assign n19332 = ~n380 & n19331 ;
  assign n19333 = n19332 ^ n12106 ^ 1'b0 ;
  assign n19334 = n10481 ^ n8996 ^ 1'b0 ;
  assign n19335 = n19334 ^ n11986 ^ n2489 ;
  assign n19336 = n341 & ~n19335 ;
  assign n19337 = n19336 ^ n7210 ^ 1'b0 ;
  assign n19338 = x37 & n5113 ;
  assign n19339 = ( n5318 & n8657 ) | ( n5318 & n19338 ) | ( n8657 & n19338 ) ;
  assign n19340 = n19339 ^ n13181 ^ 1'b0 ;
  assign n19341 = n10901 ^ n1927 ^ 1'b0 ;
  assign n19342 = n10275 & n17109 ;
  assign n19343 = n19342 ^ n17005 ^ 1'b0 ;
  assign n19344 = n11222 | n13972 ;
  assign n19345 = ~n17256 & n18303 ;
  assign n19346 = n19345 ^ n6322 ^ 1'b0 ;
  assign n19347 = n17520 | n19346 ;
  assign n19348 = n1345 | n9583 ;
  assign n19349 = n13724 ^ n2705 ^ 1'b0 ;
  assign n19350 = ~n1646 & n13195 ;
  assign n19351 = ~n17901 & n19350 ;
  assign n19352 = n19351 ^ n17527 ^ 1'b0 ;
  assign n19353 = n19349 & ~n19352 ;
  assign n19354 = n16485 ^ n13474 ^ 1'b0 ;
  assign n19355 = ( n2207 & ~n7945 ) | ( n2207 & n19354 ) | ( ~n7945 & n19354 ) ;
  assign n19356 = n19355 ^ n2038 ^ 1'b0 ;
  assign n19357 = ( n2618 & n11708 ) | ( n2618 & ~n16686 ) | ( n11708 & ~n16686 ) ;
  assign n19358 = ( n1800 & ~n16350 ) | ( n1800 & n19357 ) | ( ~n16350 & n19357 ) ;
  assign n19359 = n1263 | n16402 ;
  assign n19360 = n3240 & ~n3622 ;
  assign n19361 = n12566 & n19360 ;
  assign n19362 = n6743 | n7922 ;
  assign n19363 = n13565 ^ n2087 ^ 1'b0 ;
  assign n19364 = ( n14817 & n19362 ) | ( n14817 & n19363 ) | ( n19362 & n19363 ) ;
  assign n19365 = n19364 ^ n5572 ^ 1'b0 ;
  assign n19366 = ~n960 & n19365 ;
  assign n19367 = n15490 ^ n4260 ^ 1'b0 ;
  assign n19368 = n10226 ^ n2411 ^ 1'b0 ;
  assign n19369 = n7176 & n19368 ;
  assign n19370 = n19369 ^ x55 ^ 1'b0 ;
  assign n19371 = n6046 ^ n2613 ^ 1'b0 ;
  assign n19372 = ~n4079 & n9968 ;
  assign n19373 = x93 & ~n19372 ;
  assign n19374 = n19373 ^ n4270 ^ 1'b0 ;
  assign n19375 = n19374 ^ n6122 ^ n4946 ;
  assign n19376 = ( ~n770 & n6770 ) | ( ~n770 & n12470 ) | ( n6770 & n12470 ) ;
  assign n19377 = n11403 ^ n399 ^ 1'b0 ;
  assign n19379 = ( n341 & n884 ) | ( n341 & n3127 ) | ( n884 & n3127 ) ;
  assign n19380 = n19379 ^ n18935 ^ 1'b0 ;
  assign n19378 = ~n2423 & n12987 ;
  assign n19381 = n19380 ^ n19378 ^ 1'b0 ;
  assign n19382 = ~n876 & n19381 ;
  assign n19383 = n3270 | n5561 ;
  assign n19384 = n13697 ^ n10218 ^ n8599 ;
  assign n19385 = n831 & n13884 ;
  assign n19386 = ~n11905 & n19385 ;
  assign n19387 = n1467 | n8861 ;
  assign n19388 = n7359 | n12425 ;
  assign n19389 = n12193 | n19388 ;
  assign n19390 = n389 | n19389 ;
  assign n19391 = ~n4025 & n5339 ;
  assign n19392 = n1123 | n19391 ;
  assign n19394 = ~n6387 & n8766 ;
  assign n19393 = n17307 | n17504 ;
  assign n19395 = n19394 ^ n19393 ^ 1'b0 ;
  assign n19396 = n18673 ^ n10890 ^ n345 ;
  assign n19397 = n7529 ^ n6420 ^ n4371 ;
  assign n19398 = ( ~n8738 & n17519 ) | ( ~n8738 & n19397 ) | ( n17519 & n19397 ) ;
  assign n19399 = n7284 ^ n2154 ^ 1'b0 ;
  assign n19400 = n7490 & ~n19399 ;
  assign n19401 = n19400 ^ n4585 ^ 1'b0 ;
  assign n19402 = n2883 ^ n443 ^ 1'b0 ;
  assign n19403 = n11210 | n19402 ;
  assign n19404 = ( n1072 & n1120 ) | ( n1072 & n1949 ) | ( n1120 & n1949 ) ;
  assign n19405 = ( ~n3037 & n16173 ) | ( ~n3037 & n19404 ) | ( n16173 & n19404 ) ;
  assign n19406 = ~n2062 & n19405 ;
  assign n19407 = n254 & n19406 ;
  assign n19408 = n5356 & n5715 ;
  assign n19409 = ~n5356 & n19408 ;
  assign n19410 = n7627 | n19409 ;
  assign n19411 = n5886 & ~n9453 ;
  assign n19412 = n19410 & n19411 ;
  assign n19413 = n7564 & n14533 ;
  assign n19414 = n4786 & n19413 ;
  assign n19415 = n19414 ^ n10153 ^ 1'b0 ;
  assign n19416 = n2672 & n19415 ;
  assign n19417 = n6428 & n18790 ;
  assign n19418 = ~n19416 & n19417 ;
  assign n19419 = n5185 & n15937 ;
  assign n19420 = n19419 ^ n10355 ^ n6947 ;
  assign n19422 = n1237 & ~n7018 ;
  assign n19423 = n19422 ^ n3313 ^ 1'b0 ;
  assign n19421 = n6794 & n15760 ;
  assign n19424 = n19423 ^ n19421 ^ 1'b0 ;
  assign n19425 = n1492 | n3116 ;
  assign n19426 = n19425 ^ n18632 ^ 1'b0 ;
  assign n19427 = ~n7191 & n8247 ;
  assign n19428 = n14730 & ~n19427 ;
  assign n19429 = n4419 & ~n7763 ;
  assign n19430 = n16707 ^ n1901 ^ 1'b0 ;
  assign n19431 = ~n19429 & n19430 ;
  assign n19432 = ( n3371 & n7253 ) | ( n3371 & ~n19339 ) | ( n7253 & ~n19339 ) ;
  assign n19433 = n8685 ^ n7580 ^ 1'b0 ;
  assign n19434 = n13880 & ~n15655 ;
  assign n19435 = n19434 ^ n13575 ^ 1'b0 ;
  assign n19436 = n1835 | n19435 ;
  assign n19437 = n11954 | n19436 ;
  assign n19438 = n2642 | n19224 ;
  assign n19439 = n11179 ^ n6457 ^ 1'b0 ;
  assign n19440 = n5074 & n5516 ;
  assign n19441 = n19440 ^ n10803 ^ 1'b0 ;
  assign n19442 = n10295 | n10640 ;
  assign n19443 = n4531 | n5273 ;
  assign n19444 = ~n10994 & n19443 ;
  assign n19445 = ~n19442 & n19444 ;
  assign n19446 = n19445 ^ n7778 ^ 1'b0 ;
  assign n19447 = n197 & ~n1410 ;
  assign n19448 = ~n4420 & n19447 ;
  assign n19449 = n6476 & ~n19448 ;
  assign n19450 = n19449 ^ n19084 ^ 1'b0 ;
  assign n19451 = n8709 ^ n2541 ^ 1'b0 ;
  assign n19452 = n9091 | n19451 ;
  assign n19453 = n19452 ^ n15290 ^ n912 ;
  assign n19454 = n6669 ^ n6527 ^ 1'b0 ;
  assign n19455 = n7623 | n19454 ;
  assign n19456 = n19455 ^ n10139 ^ 1'b0 ;
  assign n19457 = ~n2726 & n10067 ;
  assign n19458 = ~n12809 & n19457 ;
  assign n19459 = n19458 ^ n15594 ^ n11602 ;
  assign n19460 = n2870 | n8042 ;
  assign n19461 = n9520 & n19460 ;
  assign n19462 = n1283 & ~n18666 ;
  assign n19463 = ~n2451 & n11174 ;
  assign n19464 = n17453 ^ n5553 ^ 1'b0 ;
  assign n19465 = ( n4443 & n19463 ) | ( n4443 & n19464 ) | ( n19463 & n19464 ) ;
  assign n19466 = n681 | n7900 ;
  assign n19467 = ~n9069 & n14137 ;
  assign n19468 = n15729 & n19467 ;
  assign n19469 = ~n5902 & n19468 ;
  assign n19470 = ~n7012 & n8094 ;
  assign n19471 = n19470 ^ n11036 ^ 1'b0 ;
  assign n19472 = ~n10414 & n14673 ;
  assign n19473 = ~n2929 & n7008 ;
  assign n19474 = n16969 & ~n19473 ;
  assign n19475 = ~n2189 & n5381 ;
  assign n19476 = n7808 & n19475 ;
  assign n19477 = n4436 ^ n3897 ^ 1'b0 ;
  assign n19478 = n680 | n11469 ;
  assign n19479 = n7800 & n19478 ;
  assign n19480 = n1455 & ~n19479 ;
  assign n19481 = ~n2652 & n13950 ;
  assign n19482 = ~n2857 & n19481 ;
  assign n19483 = n5434 & ~n19482 ;
  assign n19484 = n19483 ^ n3170 ^ 1'b0 ;
  assign n19485 = n17358 ^ n3249 ^ 1'b0 ;
  assign n19486 = n998 | n19485 ;
  assign n19487 = n13419 & ~n19486 ;
  assign n19488 = n5530 ^ n3808 ^ n1753 ;
  assign n19489 = n4232 & n5356 ;
  assign n19490 = n19488 & n19489 ;
  assign n19491 = n2934 & ~n5901 ;
  assign n19492 = n19491 ^ n5002 ^ 1'b0 ;
  assign n19493 = n16653 & n17080 ;
  assign n19494 = x105 | n15199 ;
  assign n19495 = n9993 ^ n5806 ^ 1'b0 ;
  assign n19496 = ~n6099 & n19495 ;
  assign n19497 = ( n4294 & n7158 ) | ( n4294 & ~n12671 ) | ( n7158 & ~n12671 ) ;
  assign n19498 = n1393 & ~n4050 ;
  assign n19499 = n19498 ^ n4585 ^ 1'b0 ;
  assign n19500 = n19499 ^ n4758 ^ 1'b0 ;
  assign n19501 = n10592 | n19500 ;
  assign n19502 = n19497 & ~n19501 ;
  assign n19503 = n8172 & ~n19502 ;
  assign n19504 = n19503 ^ n1504 ^ 1'b0 ;
  assign n19505 = n5142 ^ n1013 ^ 1'b0 ;
  assign n19506 = n194 & n19505 ;
  assign n19507 = n3011 ^ n254 ^ 1'b0 ;
  assign n19508 = ~n7352 & n8709 ;
  assign n19509 = n17633 ^ n7377 ^ 1'b0 ;
  assign n19510 = ~n19508 & n19509 ;
  assign n19511 = n19507 & n19510 ;
  assign n19512 = n7538 | n8415 ;
  assign n19513 = n2940 & n14530 ;
  assign n19514 = n19513 ^ n10107 ^ 1'b0 ;
  assign n19515 = n19514 ^ n5231 ^ 1'b0 ;
  assign n19516 = n3574 & n10740 ;
  assign n19517 = ~n11207 & n19516 ;
  assign n19518 = n13270 ^ n8994 ^ 1'b0 ;
  assign n19519 = ( n6926 & n11552 ) | ( n6926 & n19518 ) | ( n11552 & n19518 ) ;
  assign n19520 = n19519 ^ n16935 ^ 1'b0 ;
  assign n19521 = n19517 | n19520 ;
  assign n19522 = n2302 & ~n5746 ;
  assign n19523 = n6470 & ~n8587 ;
  assign n19524 = n19523 ^ x48 ^ 1'b0 ;
  assign n19527 = n2023 | n3320 ;
  assign n19525 = n10458 ^ x3 ^ 1'b0 ;
  assign n19526 = ~n12651 & n19525 ;
  assign n19528 = n19527 ^ n19526 ^ n1080 ;
  assign n19529 = n4365 ^ n1258 ^ 1'b0 ;
  assign n19530 = n5603 ^ n1589 ^ 1'b0 ;
  assign n19531 = n19530 ^ n13795 ^ n6706 ;
  assign n19532 = n19531 ^ n12492 ^ 1'b0 ;
  assign n19533 = n3871 | n19532 ;
  assign n19534 = n8531 ^ n7377 ^ 1'b0 ;
  assign n19535 = n4555 & ~n19534 ;
  assign n19536 = n6126 ^ n5631 ^ 1'b0 ;
  assign n19537 = n19535 & ~n19536 ;
  assign n19538 = ~n2483 & n2666 ;
  assign n19539 = n19538 ^ n18027 ^ n10567 ;
  assign n19540 = ( n892 & n1041 ) | ( n892 & ~n17878 ) | ( n1041 & ~n17878 ) ;
  assign n19541 = n1628 & n7796 ;
  assign n19542 = n19541 ^ n290 ^ 1'b0 ;
  assign n19543 = n14165 ^ n3482 ^ 1'b0 ;
  assign n19544 = n869 & ~n19543 ;
  assign n19545 = n15595 | n19544 ;
  assign n19546 = x65 | n13536 ;
  assign n19547 = n11043 & n19546 ;
  assign n19548 = n156 & ~n569 ;
  assign n19549 = n19548 ^ n14304 ^ 1'b0 ;
  assign n19550 = n2388 ^ n1827 ^ 1'b0 ;
  assign n19551 = n19549 | n19550 ;
  assign n19552 = n674 & n16257 ;
  assign n19553 = n16558 ^ n10790 ^ n5034 ;
  assign n19554 = ( n8785 & n15794 ) | ( n8785 & ~n19553 ) | ( n15794 & ~n19553 ) ;
  assign n19555 = n13520 ^ n1089 ^ 1'b0 ;
  assign n19556 = n18309 & ~n19555 ;
  assign n19559 = n8308 | n10754 ;
  assign n19560 = n4270 | n19559 ;
  assign n19558 = n18133 ^ n6399 ^ n1492 ;
  assign n19561 = n19560 ^ n19558 ^ 1'b0 ;
  assign n19557 = n8460 & ~n19187 ;
  assign n19562 = n19561 ^ n19557 ^ 1'b0 ;
  assign n19563 = n19556 & n19562 ;
  assign n19564 = n17781 ^ n4088 ^ 1'b0 ;
  assign n19565 = ~n2917 & n19564 ;
  assign n19566 = n11961 ^ n5897 ^ 1'b0 ;
  assign n19567 = n19566 ^ n6573 ^ n6564 ;
  assign n19568 = n15949 ^ n7185 ^ 1'b0 ;
  assign n19569 = n8341 ^ n4138 ^ 1'b0 ;
  assign n19570 = n2152 & ~n19569 ;
  assign n19571 = ~n2278 & n19570 ;
  assign n19572 = n19568 | n19571 ;
  assign n19573 = n19572 ^ n11058 ^ n7915 ;
  assign n19574 = ~n5585 & n8417 ;
  assign n19575 = ~n2254 & n19574 ;
  assign n19576 = n19575 ^ n15594 ^ 1'b0 ;
  assign n19577 = n17664 ^ n11819 ^ 1'b0 ;
  assign n19578 = n14114 & ~n19577 ;
  assign n19583 = n3740 ^ n562 ^ 1'b0 ;
  assign n19584 = ~n6607 & n19583 ;
  assign n19585 = n14621 & n19584 ;
  assign n19579 = n18166 ^ n6315 ^ 1'b0 ;
  assign n19580 = ~n17917 & n19579 ;
  assign n19581 = n19580 ^ n9781 ^ 1'b0 ;
  assign n19582 = ~n498 & n19581 ;
  assign n19586 = n19585 ^ n19582 ^ 1'b0 ;
  assign n19587 = ~n8496 & n15219 ;
  assign n19588 = n1153 & ~n19587 ;
  assign n19589 = n19588 ^ n3105 ^ 1'b0 ;
  assign n19590 = ~n4981 & n19369 ;
  assign n19591 = n19590 ^ n6729 ^ 1'b0 ;
  assign n19592 = n19130 & ~n19591 ;
  assign n19593 = ~n5114 & n19592 ;
  assign n19594 = n14207 ^ n4697 ^ 1'b0 ;
  assign n19595 = ~n19593 & n19594 ;
  assign n19596 = ( n250 & n2654 ) | ( n250 & n12558 ) | ( n2654 & n12558 ) ;
  assign n19597 = ( n8001 & n18896 ) | ( n8001 & n19596 ) | ( n18896 & n19596 ) ;
  assign n19598 = ~n717 & n1864 ;
  assign n19599 = n19598 ^ n3914 ^ 1'b0 ;
  assign n19600 = n6310 ^ n4860 ^ 1'b0 ;
  assign n19601 = n7804 & ~n19600 ;
  assign n19602 = ~n5743 & n19601 ;
  assign n19603 = n19602 ^ n3574 ^ 1'b0 ;
  assign n19604 = n19599 & n19603 ;
  assign n19605 = n19604 ^ n10234 ^ 1'b0 ;
  assign n19606 = ( ~n10183 & n19597 ) | ( ~n10183 & n19605 ) | ( n19597 & n19605 ) ;
  assign n19607 = x28 & ~n5923 ;
  assign n19608 = n18080 ^ n677 ^ 1'b0 ;
  assign n19609 = n10682 ^ n5530 ^ 1'b0 ;
  assign n19610 = n11328 ^ n4291 ^ n2307 ;
  assign n19611 = n19610 ^ n12089 ^ 1'b0 ;
  assign n19612 = ~n10170 & n14236 ;
  assign n19613 = n3831 ^ n1108 ^ 1'b0 ;
  assign n19614 = n2701 | n19613 ;
  assign n19615 = n4038 | n19614 ;
  assign n19616 = n19615 ^ n10773 ^ n8106 ;
  assign n19617 = n1918 | n17622 ;
  assign n19618 = n19617 ^ n13361 ^ 1'b0 ;
  assign n19619 = n3033 | n5259 ;
  assign n19620 = n10228 | n19619 ;
  assign n19621 = n6657 ^ n3669 ^ 1'b0 ;
  assign n19622 = n13233 & n19621 ;
  assign n19623 = ~n9156 & n16675 ;
  assign n19624 = ~n10738 & n19623 ;
  assign n19625 = n892 & ~n16207 ;
  assign n19626 = n398 & ~n10540 ;
  assign n19627 = ( n335 & n8603 ) | ( n335 & n19626 ) | ( n8603 & n19626 ) ;
  assign n19628 = n2419 & n2467 ;
  assign n19629 = n6031 | n6891 ;
  assign n19630 = n13723 & n19629 ;
  assign n19631 = ~n14347 & n19630 ;
  assign n19632 = n14637 ^ n3107 ^ 1'b0 ;
  assign n19633 = n19631 | n19632 ;
  assign n19634 = n10918 ^ n10504 ^ 1'b0 ;
  assign n19635 = n9240 | n10999 ;
  assign n19636 = n19634 | n19635 ;
  assign n19637 = n16140 & n19636 ;
  assign n19638 = n10682 & n19637 ;
  assign n19639 = n10594 ^ n830 ^ 1'b0 ;
  assign n19640 = n2461 & n19639 ;
  assign n19641 = n1074 & n3312 ;
  assign n19642 = ~n2522 & n19641 ;
  assign n19643 = ~n1051 & n2607 ;
  assign n19644 = n19643 ^ n1765 ^ 1'b0 ;
  assign n19645 = n3152 | n19644 ;
  assign n19646 = ~n19642 & n19645 ;
  assign n19647 = n19646 ^ n7035 ^ 1'b0 ;
  assign n19648 = n7740 ^ n3882 ^ 1'b0 ;
  assign n19649 = n2493 & n4131 ;
  assign n19650 = n19649 ^ n10210 ^ 1'b0 ;
  assign n19651 = n7473 | n18745 ;
  assign n19652 = n19651 ^ n15806 ^ 1'b0 ;
  assign n19653 = n19652 ^ n4469 ^ 1'b0 ;
  assign n19654 = ~n6422 & n19653 ;
  assign n19655 = n1134 & n1430 ;
  assign n19656 = ~n6839 & n19655 ;
  assign n19657 = n11180 ^ n7027 ^ 1'b0 ;
  assign n19658 = n5791 & n19657 ;
  assign n19659 = ( n245 & n14659 ) | ( n245 & ~n19658 ) | ( n14659 & ~n19658 ) ;
  assign n19660 = n2711 & n3276 ;
  assign n19661 = n19660 ^ n576 ^ 1'b0 ;
  assign n19662 = n19036 & n19661 ;
  assign n19663 = n12922 ^ n3868 ^ 1'b0 ;
  assign n19664 = ~n19662 & n19663 ;
  assign n19665 = ~n8640 & n18944 ;
  assign n19666 = n7372 | n9754 ;
  assign n19667 = n8225 ^ n3455 ^ 1'b0 ;
  assign n19668 = n5547 & ~n19667 ;
  assign n19669 = n19666 | n19668 ;
  assign n19670 = n4645 | n19669 ;
  assign n19671 = n16736 ^ n15721 ^ n9424 ;
  assign n19672 = n1387 | n8458 ;
  assign n19673 = n19401 & n19672 ;
  assign n19674 = n17579 ^ n8886 ^ n5428 ;
  assign n19675 = n9763 ^ n1396 ^ 1'b0 ;
  assign n19676 = x49 & n19675 ;
  assign n19677 = n1141 ^ n469 ^ 1'b0 ;
  assign n19678 = n2249 & n19677 ;
  assign n19679 = ( n307 & n12417 ) | ( n307 & ~n19678 ) | ( n12417 & ~n19678 ) ;
  assign n19680 = n14032 ^ n10041 ^ 1'b0 ;
  assign n19681 = n12308 ^ n2112 ^ 1'b0 ;
  assign n19682 = ~n19680 & n19681 ;
  assign n19683 = ~n15443 & n19682 ;
  assign n19684 = n19683 ^ n13722 ^ 1'b0 ;
  assign n19685 = n19679 & n19684 ;
  assign n19686 = n16707 ^ n16420 ^ n5881 ;
  assign n19687 = n9287 ^ n3954 ^ 1'b0 ;
  assign n19688 = n5392 & n10544 ;
  assign n19689 = ~n10250 & n19688 ;
  assign n19690 = n7471 & ~n10767 ;
  assign n19691 = ( n6966 & ~n8959 ) | ( n6966 & n11691 ) | ( ~n8959 & n11691 ) ;
  assign n19692 = n2154 & ~n19691 ;
  assign n19693 = n13395 & n19692 ;
  assign n19694 = n3228 | n9327 ;
  assign n19695 = n19693 | n19694 ;
  assign n19696 = n509 & ~n6179 ;
  assign n19697 = n3630 | n13959 ;
  assign n19698 = n19697 ^ n5077 ^ 1'b0 ;
  assign n19699 = n10476 ^ n4378 ^ n3152 ;
  assign n19700 = n19699 ^ n11638 ^ n1688 ;
  assign n19701 = ( n14098 & n16100 ) | ( n14098 & n19700 ) | ( n16100 & n19700 ) ;
  assign n19702 = n9908 ^ n2431 ^ 1'b0 ;
  assign n19703 = n4723 & n19702 ;
  assign n19704 = n19703 ^ n8776 ^ 1'b0 ;
  assign n19705 = ~n11344 & n12809 ;
  assign n19706 = ~n12809 & n19705 ;
  assign n19707 = ( ~n3684 & n6209 ) | ( ~n3684 & n7299 ) | ( n6209 & n7299 ) ;
  assign n19708 = n19707 ^ n3302 ^ 1'b0 ;
  assign n19709 = n19706 | n19708 ;
  assign n19710 = n10784 & ~n19709 ;
  assign n19711 = n19709 & n19710 ;
  assign n19712 = n19711 ^ n9364 ^ n3554 ;
  assign n19713 = n12078 ^ n9840 ^ 1'b0 ;
  assign n19714 = ~n5487 & n10943 ;
  assign n19715 = n19714 ^ n11985 ^ 1'b0 ;
  assign n19716 = n13264 ^ n3155 ^ 1'b0 ;
  assign n19717 = ~n16786 & n19716 ;
  assign n19718 = n2098 ^ n1311 ^ 1'b0 ;
  assign n19719 = ~n3901 & n19718 ;
  assign n19720 = n19719 ^ n2712 ^ 1'b0 ;
  assign n19721 = n18144 ^ n8108 ^ 1'b0 ;
  assign n19722 = n1552 | n9271 ;
  assign n19723 = n11129 ^ n745 ^ 1'b0 ;
  assign n19724 = n7116 & ~n7567 ;
  assign n19725 = n1380 & n19724 ;
  assign n19726 = ~n1226 & n12205 ;
  assign n19727 = n19725 & n19726 ;
  assign n19728 = n19727 ^ n3226 ^ n681 ;
  assign n19729 = n9216 | n19442 ;
  assign n19730 = n19729 ^ n5969 ^ 1'b0 ;
  assign n19731 = ( ~n1675 & n16748 ) | ( ~n1675 & n19730 ) | ( n16748 & n19730 ) ;
  assign n19732 = n8994 & ~n9744 ;
  assign n19733 = ~n6181 & n19732 ;
  assign n19734 = n19733 ^ n5542 ^ 1'b0 ;
  assign n19735 = ~n8166 & n18535 ;
  assign n19736 = n15632 | n15790 ;
  assign n19737 = n10361 | n15638 ;
  assign n19738 = n19737 ^ n6218 ^ 1'b0 ;
  assign n19739 = n19738 ^ n6463 ^ 1'b0 ;
  assign n19740 = n6799 & ~n10463 ;
  assign n19741 = n11790 & n19740 ;
  assign n19742 = n5868 & n12931 ;
  assign n19743 = n19742 ^ n9726 ^ n7650 ;
  assign n19744 = n10908 ^ n2306 ^ n1944 ;
  assign n19748 = ( n1188 & ~n3857 ) | ( n1188 & n4749 ) | ( ~n3857 & n4749 ) ;
  assign n19749 = n19748 ^ n12872 ^ n9882 ;
  assign n19750 = n3738 & ~n19749 ;
  assign n19751 = n19750 ^ n2198 ^ 1'b0 ;
  assign n19752 = n19751 ^ n5480 ^ 1'b0 ;
  assign n19753 = ~n644 & n19752 ;
  assign n19745 = x51 & ~n425 ;
  assign n19746 = n1238 & n19745 ;
  assign n19747 = n7724 | n19746 ;
  assign n19754 = n19753 ^ n19747 ^ 1'b0 ;
  assign n19755 = n11328 ^ n3446 ^ 1'b0 ;
  assign n19756 = n4330 & ~n19755 ;
  assign n19757 = n18477 ^ n12682 ^ n8919 ;
  assign n19758 = ~n4342 & n19757 ;
  assign n19759 = n7577 & n19758 ;
  assign n19760 = ~n7347 & n9063 ;
  assign n19761 = n16114 & ~n19760 ;
  assign n19762 = n18174 ^ n2611 ^ 1'b0 ;
  assign n19763 = n19761 & n19762 ;
  assign n19764 = n1907 | n18956 ;
  assign n19765 = n19764 ^ n1703 ^ 1'b0 ;
  assign n19766 = n497 & n19765 ;
  assign n19767 = n19766 ^ n6148 ^ 1'b0 ;
  assign n19768 = n1953 & n3805 ;
  assign n19769 = n19768 ^ n1324 ^ 1'b0 ;
  assign n19770 = n19769 ^ n4759 ^ 1'b0 ;
  assign n19771 = ~n2715 & n19770 ;
  assign n19772 = n10959 ^ n8685 ^ 1'b0 ;
  assign n19773 = n19771 & ~n19772 ;
  assign n19774 = n19773 ^ n15630 ^ 1'b0 ;
  assign n19775 = n11995 ^ n4828 ^ 1'b0 ;
  assign n19776 = ( n3210 & ~n5953 ) | ( n3210 & n7444 ) | ( ~n5953 & n7444 ) ;
  assign n19777 = ~n2283 & n19776 ;
  assign n19778 = n19777 ^ n16005 ^ n6018 ;
  assign n19779 = n19775 & n19778 ;
  assign n19780 = n3767 | n9216 ;
  assign n19781 = n14402 & n16496 ;
  assign n19782 = n19781 ^ n7560 ^ 1'b0 ;
  assign n19783 = n869 & ~n7797 ;
  assign n19784 = n19783 ^ n5940 ^ 1'b0 ;
  assign n19785 = n3230 | n11340 ;
  assign n19786 = n15565 ^ n10647 ^ 1'b0 ;
  assign n19787 = n1251 ^ n872 ^ 1'b0 ;
  assign n19788 = n4253 ^ n3307 ^ 1'b0 ;
  assign n19789 = n1353 & n10216 ;
  assign n19790 = ~n1115 & n19789 ;
  assign n19791 = n19788 | n19790 ;
  assign n19792 = n19791 ^ n12564 ^ 1'b0 ;
  assign n19793 = x18 & ~n5043 ;
  assign n19794 = n2339 & n19793 ;
  assign n19795 = n9189 | n19794 ;
  assign n19796 = n6806 | n10424 ;
  assign n19797 = n19795 & ~n19796 ;
  assign n19798 = n19797 ^ n3981 ^ 1'b0 ;
  assign n19799 = n15209 & n19798 ;
  assign n19800 = n3334 ^ n809 ^ 1'b0 ;
  assign n19801 = n5326 ^ n5046 ^ n1695 ;
  assign n19802 = ( n10244 & n14018 ) | ( n10244 & ~n19788 ) | ( n14018 & ~n19788 ) ;
  assign n19803 = n10537 | n18401 ;
  assign n19804 = ( ~n202 & n4165 ) | ( ~n202 & n6458 ) | ( n4165 & n6458 ) ;
  assign n19805 = ( n6131 & n10234 ) | ( n6131 & n19804 ) | ( n10234 & n19804 ) ;
  assign n19806 = n14438 ^ n11272 ^ 1'b0 ;
  assign n19807 = n19806 ^ n134 ^ 1'b0 ;
  assign n19808 = n2271 & n12086 ;
  assign n19809 = n15255 & n17063 ;
  assign n19810 = ~n623 & n17553 ;
  assign n19811 = ( ~n5686 & n15937 ) | ( ~n5686 & n18292 ) | ( n15937 & n18292 ) ;
  assign n19812 = n1064 & ~n11985 ;
  assign n19813 = ( n450 & n4307 ) | ( n450 & ~n19812 ) | ( n4307 & ~n19812 ) ;
  assign n19814 = n4504 & ~n7197 ;
  assign n19815 = n8232 & n19814 ;
  assign n19816 = n19813 & n19815 ;
  assign n19817 = ( n1229 & ~n10808 ) | ( n1229 & n19816 ) | ( ~n10808 & n19816 ) ;
  assign n19818 = n11031 ^ n8198 ^ 1'b0 ;
  assign n19819 = n4398 | n4907 ;
  assign n19820 = n5778 ^ n856 ^ 1'b0 ;
  assign n19821 = n19820 ^ n14968 ^ 1'b0 ;
  assign n19822 = ~n19819 & n19821 ;
  assign n19823 = n13386 ^ n3179 ^ n1062 ;
  assign n19824 = n19822 & ~n19823 ;
  assign n19825 = n15136 ^ n7561 ^ 1'b0 ;
  assign n19826 = ~n5948 & n19122 ;
  assign n19827 = ~n5419 & n19826 ;
  assign n19828 = n1710 | n4018 ;
  assign n19829 = n19828 ^ n6085 ^ 1'b0 ;
  assign n19830 = n8081 | n10364 ;
  assign n19831 = ~n8643 & n19830 ;
  assign n19832 = ~n845 & n19831 ;
  assign n19833 = n19832 ^ n8617 ^ 1'b0 ;
  assign n19834 = n10231 & ~n19833 ;
  assign n19835 = n13189 ^ n6616 ^ 1'b0 ;
  assign n19836 = n13510 & n19835 ;
  assign n19837 = ( ~n6582 & n16884 ) | ( ~n6582 & n19836 ) | ( n16884 & n19836 ) ;
  assign n19838 = n11914 | n12487 ;
  assign n19839 = n1976 | n12603 ;
  assign n19840 = ~n6573 & n14595 ;
  assign n19841 = n19840 ^ n10293 ^ 1'b0 ;
  assign n19842 = n10735 ^ n10332 ^ n9765 ;
  assign n19843 = ~n3446 & n19842 ;
  assign n19844 = n942 | n4267 ;
  assign n19845 = n19844 ^ n4593 ^ 1'b0 ;
  assign n19846 = ~n2466 & n14332 ;
  assign n19847 = n19846 ^ n7957 ^ 1'b0 ;
  assign n19848 = n19847 ^ n3568 ^ n574 ;
  assign n19849 = n11055 ^ n2001 ^ 1'b0 ;
  assign n19850 = n5141 ^ n4647 ^ 1'b0 ;
  assign n19851 = x79 & ~n11085 ;
  assign n19852 = n19850 & n19851 ;
  assign n19853 = n15785 | n19852 ;
  assign n19854 = n19849 & ~n19853 ;
  assign n19855 = n3460 & n12563 ;
  assign n19856 = n10160 | n19855 ;
  assign n19857 = ( n2596 & n5937 ) | ( n2596 & ~n7536 ) | ( n5937 & ~n7536 ) ;
  assign n19858 = n19857 ^ n13928 ^ 1'b0 ;
  assign n19859 = n19858 ^ n2958 ^ 1'b0 ;
  assign n19860 = n13578 ^ n523 ^ 1'b0 ;
  assign n19861 = n18709 & ~n19860 ;
  assign n19862 = ~n753 & n11683 ;
  assign n19863 = ~n7967 & n19862 ;
  assign n19864 = n1186 & n12214 ;
  assign n19865 = n19864 ^ n15266 ^ 1'b0 ;
  assign n19866 = n6647 ^ n2662 ^ 1'b0 ;
  assign n19867 = n19866 ^ n3868 ^ 1'b0 ;
  assign n19868 = n850 | n7761 ;
  assign n19869 = ~n6010 & n10834 ;
  assign n19870 = n19869 ^ n15732 ^ 1'b0 ;
  assign n19872 = n7850 ^ n578 ^ 1'b0 ;
  assign n19873 = n5328 & n19872 ;
  assign n19871 = n1277 | n13578 ;
  assign n19874 = n19873 ^ n19871 ^ 1'b0 ;
  assign n19875 = n15489 ^ n10066 ^ n3135 ;
  assign n19876 = n2972 | n10259 ;
  assign n19877 = n19876 ^ n2691 ^ 1'b0 ;
  assign n19878 = n14595 & n19877 ;
  assign n19879 = ( n10052 & n15237 ) | ( n10052 & n19878 ) | ( n15237 & n19878 ) ;
  assign n19880 = n163 & n18728 ;
  assign n19881 = ( x27 & n11394 ) | ( x27 & ~n13368 ) | ( n11394 & ~n13368 ) ;
  assign n19882 = n2979 & n19881 ;
  assign n19883 = n19882 ^ n13330 ^ 1'b0 ;
  assign n19887 = n13981 ^ n586 ^ 1'b0 ;
  assign n19888 = n677 | n19887 ;
  assign n19885 = n10094 ^ n1952 ^ 1'b0 ;
  assign n19884 = n3456 | n11460 ;
  assign n19886 = n19885 ^ n19884 ^ 1'b0 ;
  assign n19889 = n19888 ^ n19886 ^ n425 ;
  assign n19890 = n10087 ^ n6435 ^ 1'b0 ;
  assign n19891 = ~n1374 & n19890 ;
  assign n19892 = n12050 ^ n11110 ^ 1'b0 ;
  assign n19893 = ~n865 & n19892 ;
  assign n19894 = n18293 ^ n11587 ^ n7761 ;
  assign n19895 = ( n7316 & ~n13085 ) | ( n7316 & n19894 ) | ( ~n13085 & n19894 ) ;
  assign n19896 = n1599 ^ n567 ^ 1'b0 ;
  assign n19897 = ( n2214 & ~n19895 ) | ( n2214 & n19896 ) | ( ~n19895 & n19896 ) ;
  assign n19898 = n4016 | n19402 ;
  assign n19899 = ( n3259 & n6490 ) | ( n3259 & n19898 ) | ( n6490 & n19898 ) ;
  assign n19900 = n9540 ^ n2611 ^ 1'b0 ;
  assign n19901 = n148 & n4164 ;
  assign n19902 = n19901 ^ n12344 ^ 1'b0 ;
  assign n19903 = n19902 ^ n2203 ^ 1'b0 ;
  assign n19904 = n14222 ^ n7432 ^ 1'b0 ;
  assign n19905 = n10183 ^ n2176 ^ 1'b0 ;
  assign n19911 = n745 | n10924 ;
  assign n19912 = n5585 & ~n19911 ;
  assign n19907 = n2551 & ~n9321 ;
  assign n19908 = n15016 & n19005 ;
  assign n19909 = n19907 & n19908 ;
  assign n19910 = n19909 ^ n3802 ^ 1'b0 ;
  assign n19906 = ( n3721 & n8040 ) | ( n3721 & n9395 ) | ( n8040 & n9395 ) ;
  assign n19913 = n19912 ^ n19910 ^ n19906 ;
  assign n19914 = x52 & ~n3167 ;
  assign n19915 = n5366 & n19914 ;
  assign n19916 = n2786 & n15443 ;
  assign n19917 = n19916 ^ n7311 ^ 1'b0 ;
  assign n19918 = n18305 ^ n1882 ^ 1'b0 ;
  assign n19919 = n8319 & n12364 ;
  assign n19920 = n11859 & n19919 ;
  assign n19921 = n9247 ^ n5728 ^ 1'b0 ;
  assign n19922 = ~n1149 & n19921 ;
  assign n19923 = n12989 ^ n12871 ^ n3609 ;
  assign n19924 = n13842 ^ n13403 ^ n7553 ;
  assign n19925 = n15812 ^ n1064 ^ 1'b0 ;
  assign n19926 = n4221 | n14575 ;
  assign n19927 = n19926 ^ n15490 ^ 1'b0 ;
  assign n19928 = n11446 & ~n19927 ;
  assign n19929 = n2256 & ~n8331 ;
  assign n19930 = n17706 & n19929 ;
  assign n19932 = n6079 ^ n4927 ^ 1'b0 ;
  assign n19933 = ( n3053 & ~n7669 ) | ( n3053 & n10895 ) | ( ~n7669 & n10895 ) ;
  assign n19934 = ~n19932 & n19933 ;
  assign n19935 = n19934 ^ n1410 ^ 1'b0 ;
  assign n19931 = ( ~n6483 & n7522 ) | ( ~n6483 & n15150 ) | ( n7522 & n15150 ) ;
  assign n19936 = n19935 ^ n19931 ^ n15374 ;
  assign n19937 = n9787 & n10401 ;
  assign n19938 = n7075 & n19937 ;
  assign n19939 = n372 | n19938 ;
  assign n19940 = n19939 ^ n7230 ^ 1'b0 ;
  assign n19941 = n1350 ^ n431 ^ 1'b0 ;
  assign n19942 = ( ~n3070 & n6261 ) | ( ~n3070 & n12875 ) | ( n6261 & n12875 ) ;
  assign n19946 = ( n4314 & n8504 ) | ( n4314 & ~n18690 ) | ( n8504 & ~n18690 ) ;
  assign n19947 = ~n2092 & n19946 ;
  assign n19948 = n19947 ^ n12541 ^ 1'b0 ;
  assign n19943 = n8885 ^ n535 ^ 1'b0 ;
  assign n19944 = n7173 & n19943 ;
  assign n19945 = ~n6049 & n19944 ;
  assign n19949 = n19948 ^ n19945 ^ 1'b0 ;
  assign n19950 = ~n3976 & n6041 ;
  assign n19951 = n2207 & ~n19950 ;
  assign n19952 = n19951 ^ n10686 ^ 1'b0 ;
  assign n19953 = n2735 ^ n1154 ^ 1'b0 ;
  assign n19954 = n4000 & ~n19953 ;
  assign n19955 = n2824 & n19954 ;
  assign n19956 = n4247 & n19955 ;
  assign n19957 = n19956 ^ n17213 ^ n3243 ;
  assign n19958 = n19957 ^ n19707 ^ n7931 ;
  assign n19959 = n6789 & n8437 ;
  assign n19960 = ~n5730 & n19959 ;
  assign n19961 = n10279 | n19960 ;
  assign n19962 = n19961 ^ n17172 ^ n9672 ;
  assign n19963 = n19962 ^ n15215 ^ 1'b0 ;
  assign n19964 = n4855 | n11087 ;
  assign n19965 = n13784 & ~n19964 ;
  assign n19966 = n5541 & ~n13995 ;
  assign n19967 = ~n9955 & n14559 ;
  assign n19968 = ~n14462 & n15943 ;
  assign n19969 = n7648 & ~n14410 ;
  assign n19970 = ( n4690 & n14704 ) | ( n4690 & n19969 ) | ( n14704 & n19969 ) ;
  assign n19971 = ~n1302 & n9329 ;
  assign n19972 = n19971 ^ n4614 ^ 1'b0 ;
  assign n19973 = n13260 ^ x95 ^ 1'b0 ;
  assign n19974 = n18864 ^ n1799 ^ 1'b0 ;
  assign n19975 = ~n6617 & n13682 ;
  assign n19976 = n11253 & ~n19975 ;
  assign n19977 = ~n884 & n3746 ;
  assign n19978 = ~n4091 & n19977 ;
  assign n19979 = n14852 ^ n4183 ^ 1'b0 ;
  assign n19980 = n3391 & ~n19979 ;
  assign n19981 = ~n19978 & n19980 ;
  assign n19982 = n19981 ^ n4860 ^ 1'b0 ;
  assign n19983 = n19982 ^ n11544 ^ n5689 ;
  assign n19984 = ( n1149 & ~n2940 ) | ( n1149 & n4266 ) | ( ~n2940 & n4266 ) ;
  assign n19985 = n19984 ^ n7395 ^ 1'b0 ;
  assign n19986 = n19985 ^ n12548 ^ n3211 ;
  assign n19987 = ~x55 & n2345 ;
  assign n19988 = n19987 ^ n10763 ^ 1'b0 ;
  assign n19989 = n12172 ^ n3914 ^ n2040 ;
  assign n19990 = ~n6060 & n19989 ;
  assign n19994 = n11825 ^ n5577 ^ 1'b0 ;
  assign n19995 = x65 | n8936 ;
  assign n19996 = n19995 ^ n13085 ^ 1'b0 ;
  assign n19997 = ~n8332 & n19996 ;
  assign n19998 = ( n1323 & n19994 ) | ( n1323 & n19997 ) | ( n19994 & n19997 ) ;
  assign n19991 = n922 | n15665 ;
  assign n19992 = n19991 ^ n6923 ^ 1'b0 ;
  assign n19993 = n19992 ^ n4685 ^ 1'b0 ;
  assign n19999 = n19998 ^ n19993 ^ 1'b0 ;
  assign n20000 = n4162 & ~n11548 ;
  assign n20003 = n3765 ^ n1445 ^ 1'b0 ;
  assign n20001 = n1088 & n3647 ;
  assign n20002 = n20001 ^ n5365 ^ 1'b0 ;
  assign n20004 = n20003 ^ n20002 ^ n12487 ;
  assign n20005 = n20004 ^ n13093 ^ n459 ;
  assign n20006 = n13767 ^ n2549 ^ 1'b0 ;
  assign n20007 = ~n9092 & n20006 ;
  assign n20008 = n20007 ^ n5559 ^ 1'b0 ;
  assign n20009 = n8520 & ~n20008 ;
  assign n20010 = n2321 & n4353 ;
  assign n20011 = n3556 & n16909 ;
  assign n20012 = n9601 & n20011 ;
  assign n20013 = n615 & ~n10522 ;
  assign n20014 = n20013 ^ n12935 ^ 1'b0 ;
  assign n20015 = n2354 & n5359 ;
  assign n20016 = ~n1153 & n20015 ;
  assign n20017 = n175 & ~n1874 ;
  assign n20018 = n17018 ^ n4737 ^ 1'b0 ;
  assign n20019 = n13810 | n19842 ;
  assign n20020 = n9399 & ~n14163 ;
  assign n20021 = ~n8036 & n20020 ;
  assign n20022 = n20021 ^ n5810 ^ 1'b0 ;
  assign n20023 = ~n18285 & n20022 ;
  assign n20024 = n5479 ^ n805 ^ 1'b0 ;
  assign n20025 = n17644 | n18411 ;
  assign n20026 = n2355 | n9811 ;
  assign n20027 = n20025 & ~n20026 ;
  assign n20028 = ( ~n2988 & n5936 ) | ( ~n2988 & n7042 ) | ( n5936 & n7042 ) ;
  assign n20029 = n20028 ^ n1266 ^ 1'b0 ;
  assign n20030 = n2703 | n20029 ;
  assign n20031 = n17710 | n20030 ;
  assign n20032 = n6546 ^ n6520 ^ 1'b0 ;
  assign n20033 = n13167 & n20032 ;
  assign n20034 = ~n259 & n582 ;
  assign n20035 = ~n3838 & n20034 ;
  assign n20036 = n8811 & ~n20035 ;
  assign n20037 = n16372 & n20036 ;
  assign n20038 = ( n3994 & ~n4836 ) | ( n3994 & n8218 ) | ( ~n4836 & n8218 ) ;
  assign n20039 = n20037 | n20038 ;
  assign n20040 = n1268 & n5971 ;
  assign n20041 = n20040 ^ n2106 ^ n1965 ;
  assign n20042 = n5937 ^ n5240 ^ 1'b0 ;
  assign n20043 = n19502 | n20042 ;
  assign n20044 = n1566 | n20043 ;
  assign n20045 = n7867 ^ n6095 ^ 1'b0 ;
  assign n20046 = ( n6939 & ~n10202 ) | ( n6939 & n16693 ) | ( ~n10202 & n16693 ) ;
  assign n20047 = ~n15123 & n20046 ;
  assign n20048 = n196 | n20047 ;
  assign n20049 = ~n9317 & n10654 ;
  assign n20050 = n1567 & n20049 ;
  assign n20051 = n20050 ^ n11412 ^ n4127 ;
  assign n20052 = n19743 & n20051 ;
  assign n20053 = n17494 ^ n15399 ^ n11581 ;
  assign n20054 = n1980 & n3747 ;
  assign n20055 = n17352 ^ n3927 ^ 1'b0 ;
  assign n20056 = n20054 & n20055 ;
  assign n20057 = ~n4497 & n14054 ;
  assign n20058 = n20057 ^ n15033 ^ 1'b0 ;
  assign n20059 = n3647 & ~n20058 ;
  assign n20060 = n20056 & n20059 ;
  assign n20063 = ~n7295 & n9081 ;
  assign n20064 = ~n1424 & n20063 ;
  assign n20065 = n7670 ^ n1186 ^ 1'b0 ;
  assign n20066 = ~n20064 & n20065 ;
  assign n20061 = n10662 ^ n3485 ^ 1'b0 ;
  assign n20062 = n20061 ^ n2921 ^ n1582 ;
  assign n20067 = n20066 ^ n20062 ^ n15544 ;
  assign n20068 = ~n8207 & n15328 ;
  assign n20069 = n20067 & ~n20068 ;
  assign n20070 = ( n2909 & n4858 ) | ( n2909 & ~n5107 ) | ( n4858 & ~n5107 ) ;
  assign n20071 = n20070 ^ n582 ^ 1'b0 ;
  assign n20072 = n6931 & ~n20071 ;
  assign n20073 = x111 & ~n3053 ;
  assign n20074 = ~n13085 & n20073 ;
  assign n20075 = ( n3034 & ~n3344 ) | ( n3034 & n3987 ) | ( ~n3344 & n3987 ) ;
  assign n20076 = n20075 ^ n18564 ^ n7151 ;
  assign n20077 = n3694 ^ n2411 ^ n2074 ;
  assign n20078 = n20077 ^ n1309 ^ 1'b0 ;
  assign n20079 = n20078 ^ n18804 ^ n3138 ;
  assign n20080 = ~n2182 & n19271 ;
  assign n20081 = n20080 ^ n19046 ^ 1'b0 ;
  assign n20082 = n17155 ^ n12153 ^ 1'b0 ;
  assign n20083 = n11147 ^ n1645 ^ 1'b0 ;
  assign n20084 = n3176 & n20083 ;
  assign n20085 = ~n10279 & n19983 ;
  assign n20086 = n19113 & n20085 ;
  assign n20087 = n6494 | n12154 ;
  assign n20088 = n14708 & ~n20087 ;
  assign n20089 = n20088 ^ n5446 ^ 1'b0 ;
  assign n20090 = n14145 & n20089 ;
  assign n20091 = n10152 & ~n19643 ;
  assign n20092 = n14997 & n20091 ;
  assign n20093 = n13888 ^ n12369 ^ 1'b0 ;
  assign n20094 = ~n6012 & n20093 ;
  assign n20095 = n20094 ^ n9607 ^ 1'b0 ;
  assign n20096 = ~n909 & n17903 ;
  assign n20097 = ~n8480 & n20096 ;
  assign n20098 = n654 ^ n305 ^ 1'b0 ;
  assign n20099 = n19858 | n20098 ;
  assign n20100 = n16499 | n20099 ;
  assign n20101 = n1953 & ~n9551 ;
  assign n20102 = ~n1189 & n7873 ;
  assign n20103 = n20102 ^ n15746 ^ 1'b0 ;
  assign n20104 = ~n13930 & n15284 ;
  assign n20105 = x67 & ~n4983 ;
  assign n20106 = ~n257 & n20105 ;
  assign n20107 = n9020 & ~n20106 ;
  assign n20108 = ( ~n3563 & n20104 ) | ( ~n3563 & n20107 ) | ( n20104 & n20107 ) ;
  assign n20109 = n20103 & ~n20108 ;
  assign n20110 = n5778 & ~n8110 ;
  assign n20111 = n8836 & n20110 ;
  assign n20112 = n11568 ^ n7639 ^ n6729 ;
  assign n20113 = n10505 ^ n1318 ^ 1'b0 ;
  assign n20114 = n20112 | n20113 ;
  assign n20115 = ( n6245 & ~n20111 ) | ( n6245 & n20114 ) | ( ~n20111 & n20114 ) ;
  assign n20116 = n4617 ^ n3418 ^ x104 ;
  assign n20117 = n20116 ^ n8288 ^ 1'b0 ;
  assign n20118 = ~n7711 & n11600 ;
  assign n20119 = n5902 & n20118 ;
  assign n20120 = ( n2564 & ~n3604 ) | ( n2564 & n3994 ) | ( ~n3604 & n3994 ) ;
  assign n20121 = ~n1963 & n20120 ;
  assign n20122 = n20121 ^ n10188 ^ 1'b0 ;
  assign n20123 = n3413 & ~n20122 ;
  assign n20124 = ~n1933 & n5328 ;
  assign n20125 = n17455 ^ n2145 ^ 1'b0 ;
  assign n20126 = n145 & n7726 ;
  assign n20127 = ~n4841 & n20126 ;
  assign n20128 = n6049 ^ n3172 ^ 1'b0 ;
  assign n20129 = n3755 & n20128 ;
  assign n20130 = n20129 ^ n14246 ^ 1'b0 ;
  assign n20131 = ~n15713 & n20130 ;
  assign n20132 = n20127 | n20131 ;
  assign n20133 = n20132 ^ n11270 ^ 1'b0 ;
  assign n20134 = n16275 & ~n20133 ;
  assign n20135 = n594 & ~n8558 ;
  assign n20136 = ~n8813 & n20135 ;
  assign n20137 = n20136 ^ n7443 ^ 1'b0 ;
  assign n20138 = n20137 ^ n8488 ^ n7471 ;
  assign n20139 = n10188 ^ n2355 ^ n867 ;
  assign n20141 = n2058 & ~n9035 ;
  assign n20142 = ~n14305 & n20141 ;
  assign n20140 = n279 & ~n2333 ;
  assign n20143 = n20142 ^ n20140 ^ 1'b0 ;
  assign n20144 = n2006 ^ n884 ^ x51 ;
  assign n20145 = ( n3237 & ~n6117 ) | ( n3237 & n20144 ) | ( ~n6117 & n20144 ) ;
  assign n20146 = n11338 ^ n6307 ^ 1'b0 ;
  assign n20147 = n20145 | n20146 ;
  assign n20148 = n20147 ^ n1042 ^ 1'b0 ;
  assign n20149 = n3612 & n11193 ;
  assign n20150 = n14263 ^ n1514 ^ n1106 ;
  assign n20151 = n8914 & ~n9923 ;
  assign n20152 = n7176 ^ n6222 ^ n5389 ;
  assign n20153 = n16753 & n17297 ;
  assign n20154 = ( n20151 & n20152 ) | ( n20151 & ~n20153 ) | ( n20152 & ~n20153 ) ;
  assign n20155 = ~n6317 & n16675 ;
  assign n20156 = n20155 ^ n5773 ^ 1'b0 ;
  assign n20157 = n6201 | n13486 ;
  assign n20158 = n1086 | n16130 ;
  assign n20159 = n962 & ~n20158 ;
  assign n20160 = n20159 ^ n19130 ^ 1'b0 ;
  assign n20161 = n9919 ^ n5531 ^ 1'b0 ;
  assign n20162 = n6156 & ~n20161 ;
  assign n20163 = ~n2827 & n20162 ;
  assign n20164 = n319 | n5003 ;
  assign n20165 = n20164 ^ n802 ^ 1'b0 ;
  assign n20166 = ~n18658 & n20165 ;
  assign n20167 = n20166 ^ n15645 ^ 1'b0 ;
  assign n20168 = n3424 & ~n20167 ;
  assign n20169 = n14326 & n20168 ;
  assign n20170 = n1465 & n12893 ;
  assign n20171 = n1854 & ~n10867 ;
  assign n20172 = n4468 | n14727 ;
  assign n20173 = n9947 & ~n20172 ;
  assign n20174 = n12559 ^ n4802 ^ 1'b0 ;
  assign n20175 = n20173 | n20174 ;
  assign n20176 = n20175 ^ n8523 ^ 1'b0 ;
  assign n20177 = ~n10590 & n16393 ;
  assign n20178 = n2448 & n4390 ;
  assign n20179 = n17472 & n20178 ;
  assign n20180 = n20179 ^ n1581 ^ 1'b0 ;
  assign n20181 = n20177 & ~n20180 ;
  assign n20182 = n3270 ^ n1034 ^ 1'b0 ;
  assign n20183 = n8966 | n20182 ;
  assign n20184 = n20182 & ~n20183 ;
  assign n20185 = n20184 ^ n2457 ^ 1'b0 ;
  assign n20188 = n896 | n10651 ;
  assign n20189 = n896 & ~n20188 ;
  assign n20190 = n4184 & ~n20189 ;
  assign n20191 = n20189 & n20190 ;
  assign n20186 = ~n6363 & n17570 ;
  assign n20187 = ~n17570 & n20186 ;
  assign n20192 = n20191 ^ n20187 ^ 1'b0 ;
  assign n20193 = ~n20185 & n20192 ;
  assign n20194 = n1050 & n13124 ;
  assign n20195 = n20194 ^ n9575 ^ 1'b0 ;
  assign n20196 = n10033 & n15638 ;
  assign n20197 = n18406 ^ n11288 ^ 1'b0 ;
  assign n20203 = ~n1321 & n7092 ;
  assign n20200 = n15722 ^ n12249 ^ 1'b0 ;
  assign n20201 = n8337 & ~n20200 ;
  assign n20198 = n1062 & ~n19860 ;
  assign n20199 = n4739 & n20198 ;
  assign n20202 = n20201 ^ n20199 ^ 1'b0 ;
  assign n20204 = n20203 ^ n20202 ^ n12562 ;
  assign n20206 = ( n700 & n5980 ) | ( n700 & n7471 ) | ( n5980 & n7471 ) ;
  assign n20205 = x1 & n1407 ;
  assign n20207 = n20206 ^ n20205 ^ 1'b0 ;
  assign n20208 = n462 | n13192 ;
  assign n20209 = n5509 & n17836 ;
  assign n20210 = n10952 ^ n1017 ^ 1'b0 ;
  assign n20211 = n9507 & ~n20210 ;
  assign n20212 = n3424 | n7862 ;
  assign n20213 = n20212 ^ n18846 ^ 1'b0 ;
  assign n20214 = n5330 & ~n9745 ;
  assign n20215 = ~n6165 & n20214 ;
  assign n20216 = n425 ^ x57 ^ 1'b0 ;
  assign n20217 = ~n20215 & n20216 ;
  assign n20218 = n10172 ^ n3206 ^ 1'b0 ;
  assign n20219 = n17905 & ~n20218 ;
  assign n20220 = n20219 ^ n16149 ^ 1'b0 ;
  assign n20221 = n4312 ^ n2679 ^ 1'b0 ;
  assign n20222 = n9914 & ~n14222 ;
  assign n20223 = ~n17686 & n20222 ;
  assign n20224 = n6308 ^ n5002 ^ 1'b0 ;
  assign n20225 = n6223 & ~n20224 ;
  assign n20226 = ( ~n3511 & n7256 ) | ( ~n3511 & n11675 ) | ( n7256 & n11675 ) ;
  assign n20227 = n3252 | n20226 ;
  assign n20228 = ~n4526 & n14975 ;
  assign n20229 = n20228 ^ n19776 ^ n17337 ;
  assign n20230 = n5542 | n11460 ;
  assign n20231 = n12601 ^ n369 ^ 1'b0 ;
  assign n20232 = ~n9013 & n20231 ;
  assign n20233 = ~n1475 & n20232 ;
  assign n20234 = n2949 | n5618 ;
  assign n20235 = n20234 ^ n10885 ^ 1'b0 ;
  assign n20236 = n5539 ^ n2190 ^ 1'b0 ;
  assign n20237 = ( n3457 & ~n4710 ) | ( n3457 & n7629 ) | ( ~n4710 & n7629 ) ;
  assign n20238 = ~n1350 & n6010 ;
  assign n20239 = n2008 ^ x56 ^ 1'b0 ;
  assign n20240 = ~n359 & n6182 ;
  assign n20241 = n20239 & n20240 ;
  assign n20242 = ~n17976 & n20095 ;
  assign n20243 = ~n15900 & n20242 ;
  assign n20244 = n5339 & ~n16287 ;
  assign n20245 = ~n4406 & n20244 ;
  assign n20246 = n2214 & ~n3489 ;
  assign n20247 = n9413 & ~n20246 ;
  assign n20248 = n20247 ^ n5598 ^ 1'b0 ;
  assign n20249 = n4008 | n15247 ;
  assign n20250 = n1290 | n20249 ;
  assign n20251 = ~n148 & n12325 ;
  assign n20252 = n6400 ^ n2952 ^ 1'b0 ;
  assign n20253 = n20251 | n20252 ;
  assign n20254 = ( n2430 & n7245 ) | ( n2430 & ~n20253 ) | ( n7245 & ~n20253 ) ;
  assign n20255 = n4975 | n15426 ;
  assign n20256 = n2255 | n5491 ;
  assign n20257 = n20256 ^ n3668 ^ 1'b0 ;
  assign n20258 = n20257 ^ n7956 ^ 1'b0 ;
  assign n20260 = ~n1819 & n5335 ;
  assign n20259 = n1607 & ~n10815 ;
  assign n20261 = n20260 ^ n20259 ^ 1'b0 ;
  assign n20262 = n8216 ^ n2618 ^ 1'b0 ;
  assign n20263 = ~n1918 & n20262 ;
  assign n20264 = ~n607 & n2049 ;
  assign n20265 = ~n20263 & n20264 ;
  assign n20267 = n18517 ^ n5402 ^ 1'b0 ;
  assign n20266 = n15115 | n16100 ;
  assign n20268 = n20267 ^ n20266 ^ 1'b0 ;
  assign n20269 = n5747 & ~n16461 ;
  assign n20270 = n6371 & ~n20269 ;
  assign n20271 = ( n5896 & ~n12975 ) | ( n5896 & n14030 ) | ( ~n12975 & n14030 ) ;
  assign n20272 = n16176 ^ n6850 ^ 1'b0 ;
  assign n20273 = n3523 | n20272 ;
  assign n20274 = n9599 & n15515 ;
  assign n20275 = n20274 ^ n663 ^ 1'b0 ;
  assign n20276 = n8406 | n8692 ;
  assign n20277 = n7458 | n20276 ;
  assign n20278 = n892 & ~n7922 ;
  assign n20279 = ~n14438 & n20278 ;
  assign n20280 = n18351 & ~n20279 ;
  assign n20281 = n20280 ^ n8181 ^ 1'b0 ;
  assign n20282 = n6047 ^ n2364 ^ 1'b0 ;
  assign n20283 = ~n9159 & n20282 ;
  assign n20284 = ~n4303 & n20283 ;
  assign n20285 = n20284 ^ n6569 ^ 1'b0 ;
  assign n20286 = n20285 ^ n8476 ^ n3391 ;
  assign n20291 = ~n4062 & n10357 ;
  assign n20287 = ~n8068 & n8512 ;
  assign n20288 = ~n14212 & n20287 ;
  assign n20289 = n20288 ^ n1504 ^ 1'b0 ;
  assign n20290 = n9349 | n20289 ;
  assign n20292 = n20291 ^ n20290 ^ 1'b0 ;
  assign n20293 = n7054 ^ n3173 ^ 1'b0 ;
  assign n20294 = n6020 | n20293 ;
  assign n20295 = n5972 | n13955 ;
  assign n20296 = n1552 & ~n3519 ;
  assign n20297 = n2142 & n5185 ;
  assign n20298 = n20297 ^ n3468 ^ 1'b0 ;
  assign n20299 = ~n983 & n2268 ;
  assign n20300 = n20299 ^ n5602 ^ 1'b0 ;
  assign n20301 = ( n1998 & n12779 ) | ( n1998 & ~n20300 ) | ( n12779 & ~n20300 ) ;
  assign n20302 = ~n7190 & n20301 ;
  assign n20303 = n8552 ^ n4087 ^ 1'b0 ;
  assign n20304 = ~n6534 & n20303 ;
  assign n20305 = n20302 & n20304 ;
  assign n20306 = ~n840 & n5879 ;
  assign n20307 = n4714 & ~n20306 ;
  assign n20308 = n2532 | n11035 ;
  assign n20309 = n2478 & n12430 ;
  assign n20310 = n20309 ^ n15052 ^ 1'b0 ;
  assign n20311 = n17956 ^ n8581 ^ 1'b0 ;
  assign n20312 = n14902 & n20311 ;
  assign n20313 = n424 & n20312 ;
  assign n20314 = n19057 ^ n3766 ^ 1'b0 ;
  assign n20316 = n17370 ^ n12249 ^ 1'b0 ;
  assign n20317 = ~n2835 & n20316 ;
  assign n20315 = n14864 ^ n6566 ^ 1'b0 ;
  assign n20318 = n20317 ^ n20315 ^ 1'b0 ;
  assign n20319 = n6841 ^ n1109 ^ 1'b0 ;
  assign n20320 = n5664 & ~n20319 ;
  assign n20321 = ( ~n7914 & n12254 ) | ( ~n7914 & n20320 ) | ( n12254 & n20320 ) ;
  assign n20322 = n9001 ^ n6217 ^ 1'b0 ;
  assign n20323 = n15025 & ~n20322 ;
  assign n20324 = n4625 & n20323 ;
  assign n20325 = ~n454 & n20324 ;
  assign n20326 = n2897 ^ n1917 ^ 1'b0 ;
  assign n20327 = n1184 & n20326 ;
  assign n20328 = n20327 ^ n9971 ^ 1'b0 ;
  assign n20329 = n14178 ^ x106 ^ 1'b0 ;
  assign n20330 = ~n8458 & n9307 ;
  assign n20331 = n14149 & ~n19172 ;
  assign n20332 = ~n20330 & n20331 ;
  assign n20333 = n5188 | n13160 ;
  assign n20334 = n15241 & ~n20333 ;
  assign n20335 = n20334 ^ n20007 ^ n3900 ;
  assign n20336 = ( ~n2513 & n4155 ) | ( ~n2513 & n16931 ) | ( n4155 & n16931 ) ;
  assign n20337 = n6346 & n20336 ;
  assign n20338 = n8206 & n15125 ;
  assign n20339 = n20337 & n20338 ;
  assign n20340 = n6483 | n8914 ;
  assign n20341 = n20340 ^ n3724 ^ 1'b0 ;
  assign n20342 = n12084 ^ n8500 ^ 1'b0 ;
  assign n20343 = x3 & n20342 ;
  assign n20344 = n20343 ^ n10740 ^ 1'b0 ;
  assign n20345 = n20059 ^ n1592 ^ 1'b0 ;
  assign n20346 = n362 & n2055 ;
  assign n20347 = n20346 ^ n5464 ^ 1'b0 ;
  assign n20349 = n16372 ^ n8445 ^ n2214 ;
  assign n20350 = n2419 | n20349 ;
  assign n20351 = n6603 & ~n20350 ;
  assign n20348 = n6239 | n19325 ;
  assign n20352 = n20351 ^ n20348 ^ 1'b0 ;
  assign n20353 = n18210 ^ n4736 ^ 1'b0 ;
  assign n20354 = n4394 & ~n20353 ;
  assign n20355 = ( n2449 & n6514 ) | ( n2449 & ~n17649 ) | ( n6514 & ~n17649 ) ;
  assign n20356 = n5039 ^ n1371 ^ 1'b0 ;
  assign n20357 = n7888 ^ n6536 ^ 1'b0 ;
  assign n20358 = ~n9754 & n20357 ;
  assign n20359 = ( ~n5971 & n8727 ) | ( ~n5971 & n20358 ) | ( n8727 & n20358 ) ;
  assign n20360 = n7921 & n9657 ;
  assign n20361 = n20360 ^ n12591 ^ 1'b0 ;
  assign n20362 = ~n3376 & n17519 ;
  assign n20363 = n20362 ^ n3718 ^ 1'b0 ;
  assign n20364 = n3599 | n8481 ;
  assign n20365 = n5223 & n16063 ;
  assign n20366 = n16677 ^ n745 ^ 1'b0 ;
  assign n20367 = n16375 & ~n20366 ;
  assign n20368 = n3349 & n20367 ;
  assign n20369 = n19744 & n20368 ;
  assign n20370 = ~n1610 & n4115 ;
  assign n20371 = n20370 ^ n8900 ^ 1'b0 ;
  assign n20387 = n3587 & n10996 ;
  assign n20388 = n20387 ^ n17857 ^ 1'b0 ;
  assign n20385 = n14196 ^ n14115 ^ 1'b0 ;
  assign n20386 = n1046 & n20385 ;
  assign n20379 = ~n1597 & n9200 ;
  assign n20380 = n20379 ^ n7856 ^ 1'b0 ;
  assign n20381 = n2366 & n20380 ;
  assign n20382 = n20381 ^ n1690 ^ 1'b0 ;
  assign n20372 = n1401 | n9349 ;
  assign n20373 = n20372 ^ n11630 ^ 1'b0 ;
  assign n20374 = n12412 ^ n5995 ^ 1'b0 ;
  assign n20375 = n16124 ^ n13592 ^ 1'b0 ;
  assign n20376 = n5589 ^ n1277 ^ 1'b0 ;
  assign n20377 = ( n20374 & ~n20375 ) | ( n20374 & n20376 ) | ( ~n20375 & n20376 ) ;
  assign n20378 = n20373 & ~n20377 ;
  assign n20383 = n20382 ^ n20378 ^ 1'b0 ;
  assign n20384 = n20383 ^ n4447 ^ 1'b0 ;
  assign n20389 = n20388 ^ n20386 ^ n20384 ;
  assign n20390 = n19546 ^ n16135 ^ n3547 ;
  assign n20391 = ~n1457 & n11057 ;
  assign n20392 = ~n15760 & n20391 ;
  assign n20393 = n13930 | n20392 ;
  assign n20394 = n20393 ^ n2909 ^ 1'b0 ;
  assign n20395 = n4025 ^ n341 ^ 1'b0 ;
  assign n20396 = n7872 & n20395 ;
  assign n20397 = n20396 ^ n4455 ^ 1'b0 ;
  assign n20398 = n18073 ^ n2151 ^ n130 ;
  assign n20399 = n13828 ^ n650 ^ 1'b0 ;
  assign n20400 = n12304 ^ n3046 ^ 1'b0 ;
  assign n20401 = n1802 & n13749 ;
  assign n20402 = ~n3961 & n20401 ;
  assign n20403 = n2282 & n20402 ;
  assign n20404 = n564 & ~n1256 ;
  assign n20405 = n20404 ^ n4730 ^ 1'b0 ;
  assign n20406 = ~n4186 & n8552 ;
  assign n20407 = n20406 ^ n6241 ^ 1'b0 ;
  assign n20408 = n19169 ^ n11014 ^ 1'b0 ;
  assign n20409 = n20407 & ~n20408 ;
  assign n20410 = n20409 ^ n7816 ^ 1'b0 ;
  assign n20411 = n3861 ^ n2258 ^ 1'b0 ;
  assign n20412 = n18773 ^ n14848 ^ 1'b0 ;
  assign n20413 = n1057 & n20412 ;
  assign n20414 = n2897 & n20413 ;
  assign n20415 = n2118 | n17519 ;
  assign n20416 = n20415 ^ n14525 ^ 1'b0 ;
  assign n20417 = n20416 ^ n581 ^ 1'b0 ;
  assign n20418 = n17375 & n20417 ;
  assign n20419 = n14412 & n18099 ;
  assign n20420 = n333 & ~n6457 ;
  assign n20421 = ( ~n582 & n1348 ) | ( ~n582 & n5997 ) | ( n1348 & n5997 ) ;
  assign n20422 = n8279 & ~n20421 ;
  assign n20423 = ~n355 & n1017 ;
  assign n20424 = n20423 ^ n12858 ^ 1'b0 ;
  assign n20425 = ( n3617 & n20422 ) | ( n3617 & ~n20424 ) | ( n20422 & ~n20424 ) ;
  assign n20426 = n9388 & n9925 ;
  assign n20427 = n13901 ^ n4410 ^ 1'b0 ;
  assign n20428 = n15115 ^ x116 ^ 1'b0 ;
  assign n20429 = n3209 & ~n20428 ;
  assign n20430 = ~n20427 & n20429 ;
  assign n20433 = n3999 | n5490 ;
  assign n20432 = n1171 | n9481 ;
  assign n20431 = ( n6233 & ~n11481 ) | ( n6233 & n13948 ) | ( ~n11481 & n13948 ) ;
  assign n20434 = n20433 ^ n20432 ^ n20431 ;
  assign n20435 = n8733 & n20434 ;
  assign n20436 = n4820 ^ n2958 ^ 1'b0 ;
  assign n20438 = n276 & n1681 ;
  assign n20437 = n175 & n20380 ;
  assign n20439 = n20438 ^ n20437 ^ n17967 ;
  assign n20440 = n6773 & n8962 ;
  assign n20441 = n11476 | n20440 ;
  assign n20442 = n14926 ^ n1103 ^ 1'b0 ;
  assign n20443 = n17669 ^ n9209 ^ 1'b0 ;
  assign n20444 = n15263 ^ n5221 ^ 1'b0 ;
  assign n20445 = n20443 & n20444 ;
  assign n20446 = ~n3027 & n18746 ;
  assign n20447 = n7462 | n17242 ;
  assign n20448 = n20446 | n20447 ;
  assign n20449 = ( ~n3742 & n15815 ) | ( ~n3742 & n17763 ) | ( n15815 & n17763 ) ;
  assign n20450 = n4450 & n10680 ;
  assign n20451 = n4951 ^ n794 ^ n352 ;
  assign n20452 = n20451 ^ n6031 ^ n1459 ;
  assign n20453 = n20452 ^ n20074 ^ 1'b0 ;
  assign n20454 = n20450 & n20453 ;
  assign n20456 = ~x123 & n7118 ;
  assign n20455 = n6898 & n6996 ;
  assign n20457 = n20456 ^ n20455 ^ n7057 ;
  assign n20458 = n5528 & ~n11308 ;
  assign n20459 = ( n2182 & ~n7726 ) | ( n2182 & n15065 ) | ( ~n7726 & n15065 ) ;
  assign n20464 = n977 | n3978 ;
  assign n20465 = n20464 ^ n1222 ^ 1'b0 ;
  assign n20466 = n6786 & n20465 ;
  assign n20460 = n3021 | n6512 ;
  assign n20461 = n20460 ^ n3698 ^ 1'b0 ;
  assign n20462 = ( n1552 & ~n11055 ) | ( n1552 & n20461 ) | ( ~n11055 & n20461 ) ;
  assign n20463 = n20462 ^ n6266 ^ 1'b0 ;
  assign n20467 = n20466 ^ n20463 ^ 1'b0 ;
  assign n20468 = n10668 ^ n4827 ^ 1'b0 ;
  assign n20469 = n1231 & n8222 ;
  assign n20470 = n20469 ^ n11274 ^ 1'b0 ;
  assign n20473 = n4720 ^ n3605 ^ n3132 ;
  assign n20471 = n6097 | n6624 ;
  assign n20472 = n3767 | n20471 ;
  assign n20474 = n20473 ^ n20472 ^ 1'b0 ;
  assign n20475 = n10834 | n18480 ;
  assign n20476 = n20475 ^ n8505 ^ n2888 ;
  assign n20477 = n6288 ^ n1154 ^ 1'b0 ;
  assign n20478 = n19527 | n20477 ;
  assign n20479 = ( n3020 & n5108 ) | ( n3020 & n20478 ) | ( n5108 & n20478 ) ;
  assign n20480 = n4780 & n9050 ;
  assign n20481 = n20480 ^ x36 ^ 1'b0 ;
  assign n20492 = n2254 & ~n16755 ;
  assign n20491 = ~n563 & n1075 ;
  assign n20493 = n20492 ^ n20491 ^ 1'b0 ;
  assign n20482 = n14199 ^ n2926 ^ 1'b0 ;
  assign n20483 = ~n409 & n15900 ;
  assign n20484 = n20483 ^ n1650 ^ 1'b0 ;
  assign n20485 = ( ~n5039 & n20482 ) | ( ~n5039 & n20484 ) | ( n20482 & n20484 ) ;
  assign n20486 = n20485 ^ n11569 ^ 1'b0 ;
  assign n20487 = n18158 & ~n20486 ;
  assign n20488 = ~n4131 & n20487 ;
  assign n20489 = n20488 ^ n17383 ^ 1'b0 ;
  assign n20490 = ~n6498 & n20489 ;
  assign n20494 = n20493 ^ n20490 ^ 1'b0 ;
  assign n20495 = ( n8313 & n10513 ) | ( n8313 & ~n16509 ) | ( n10513 & ~n16509 ) ;
  assign n20496 = n20239 ^ n10456 ^ n2285 ;
  assign n20497 = n9856 & n20496 ;
  assign n20498 = n20497 ^ n1775 ^ 1'b0 ;
  assign n20499 = ( n14458 & n17996 ) | ( n14458 & ~n20498 ) | ( n17996 & ~n20498 ) ;
  assign n20500 = n10661 ^ n2522 ^ n1459 ;
  assign n20501 = n15312 & ~n20500 ;
  assign n20502 = n15751 ^ n6719 ^ 1'b0 ;
  assign n20503 = ~n14569 & n20502 ;
  assign n20504 = n20501 & n20503 ;
  assign n20505 = n11173 ^ n8894 ^ 1'b0 ;
  assign n20506 = ~n6633 & n20505 ;
  assign n20507 = n962 & n11277 ;
  assign n20508 = n20507 ^ n7367 ^ 1'b0 ;
  assign n20509 = ~n20506 & n20508 ;
  assign n20510 = n20509 ^ n15202 ^ n11592 ;
  assign n20511 = n11251 & ~n20510 ;
  assign n20512 = n18896 ^ n256 ^ 1'b0 ;
  assign n20513 = n1106 & n12091 ;
  assign n20514 = n5155 & n20513 ;
  assign n20515 = n20514 ^ n18289 ^ n17244 ;
  assign n20516 = n5119 & n6922 ;
  assign n20517 = n2289 & ~n8922 ;
  assign n20518 = n9765 & n12177 ;
  assign n20519 = n20518 ^ n19906 ^ 1'b0 ;
  assign n20520 = n15077 ^ n1985 ^ 1'b0 ;
  assign n20521 = n1968 ^ n202 ^ 1'b0 ;
  assign n20522 = n4291 ^ n984 ^ 1'b0 ;
  assign n20523 = n17058 ^ n13977 ^ n8146 ;
  assign n20524 = n17042 ^ n13200 ^ 1'b0 ;
  assign n20525 = n11865 ^ n7218 ^ 1'b0 ;
  assign n20526 = ~n1553 & n20525 ;
  assign n20527 = n7469 ^ n2089 ^ n1771 ;
  assign n20528 = n12816 ^ n3781 ^ 1'b0 ;
  assign n20529 = ~n20527 & n20528 ;
  assign n20530 = n20529 ^ n9390 ^ 1'b0 ;
  assign n20531 = ( ~n3087 & n3212 ) | ( ~n3087 & n6372 ) | ( n3212 & n6372 ) ;
  assign n20532 = n20531 ^ n7841 ^ 1'b0 ;
  assign n20533 = n1680 & n2638 ;
  assign n20534 = n20533 ^ n4655 ^ 1'b0 ;
  assign n20535 = n2190 | n11921 ;
  assign n20536 = n17565 ^ n13624 ^ 1'b0 ;
  assign n20537 = n10744 | n20536 ;
  assign n20538 = n14608 ^ n13633 ^ n4187 ;
  assign n20539 = n18973 ^ n1981 ^ 1'b0 ;
  assign n20540 = n20538 & ~n20539 ;
  assign n20541 = n8514 ^ n359 ^ 1'b0 ;
  assign n20542 = n8345 & ~n20541 ;
  assign n20543 = n3497 ^ n138 ^ 1'b0 ;
  assign n20544 = n502 & n20543 ;
  assign n20545 = n19749 ^ n14550 ^ n11592 ;
  assign n20546 = n20545 ^ n7759 ^ 1'b0 ;
  assign n20547 = ~n5554 & n14808 ;
  assign n20549 = ( n1195 & n9458 ) | ( n1195 & n10481 ) | ( n9458 & n10481 ) ;
  assign n20550 = n5398 ^ n2355 ^ 1'b0 ;
  assign n20551 = ~n20549 & n20550 ;
  assign n20548 = ~n1504 & n2331 ;
  assign n20552 = n20551 ^ n20548 ^ n9152 ;
  assign n20553 = n236 | n664 ;
  assign n20554 = n20553 ^ n261 ^ 1'b0 ;
  assign n20555 = ~n11025 & n20554 ;
  assign n20556 = n10768 & ~n20555 ;
  assign n20557 = ( n11085 & ~n11326 ) | ( n11085 & n20556 ) | ( ~n11326 & n20556 ) ;
  assign n20558 = n17383 ^ n11308 ^ 1'b0 ;
  assign n20559 = n2692 & n20558 ;
  assign n20560 = n3651 & n20559 ;
  assign n20561 = n20560 ^ n16422 ^ 1'b0 ;
  assign n20562 = n7969 & n11500 ;
  assign n20565 = ~n5677 & n6002 ;
  assign n20566 = n20565 ^ n436 ^ 1'b0 ;
  assign n20563 = n11553 & n15064 ;
  assign n20564 = n6314 | n20563 ;
  assign n20567 = n20566 ^ n20564 ^ 1'b0 ;
  assign n20568 = n20567 ^ n15385 ^ 1'b0 ;
  assign n20571 = ( n2569 & n7019 ) | ( n2569 & n13722 ) | ( n7019 & n13722 ) ;
  assign n20569 = n9156 & n16609 ;
  assign n20570 = n6099 & n20569 ;
  assign n20572 = n20571 ^ n20570 ^ n14554 ;
  assign n20573 = n3296 & ~n12765 ;
  assign n20574 = n8173 ^ n7453 ^ 1'b0 ;
  assign n20575 = n6410 ^ n5490 ^ 1'b0 ;
  assign n20576 = n5102 & ~n20575 ;
  assign n20577 = ~n5250 & n16718 ;
  assign n20578 = ( n2487 & n3886 ) | ( n2487 & ~n8104 ) | ( n3886 & ~n8104 ) ;
  assign n20579 = n20578 ^ n5066 ^ 1'b0 ;
  assign n20580 = n20577 & n20579 ;
  assign n20581 = ~n20576 & n20580 ;
  assign n20582 = n4749 & n5059 ;
  assign n20583 = ~n2020 & n8826 ;
  assign n20584 = n20582 & n20583 ;
  assign n20585 = n2408 & ~n2719 ;
  assign n20586 = n12895 & n20585 ;
  assign n20587 = ~n17681 & n20586 ;
  assign n20588 = n6839 & ~n11600 ;
  assign n20589 = n5980 ^ n3290 ^ n512 ;
  assign n20590 = ~n4987 & n7051 ;
  assign n20591 = ~n3037 & n14697 ;
  assign n20592 = n1994 & n20591 ;
  assign n20593 = n20592 ^ n4050 ^ 1'b0 ;
  assign n20594 = ~n20590 & n20593 ;
  assign n20595 = n7112 & ~n12767 ;
  assign n20596 = n20595 ^ n9081 ^ 1'b0 ;
  assign n20597 = n2596 | n20566 ;
  assign n20598 = n11542 ^ n9067 ^ n7808 ;
  assign n20602 = ~n4394 & n7999 ;
  assign n20599 = n12489 ^ n3538 ^ 1'b0 ;
  assign n20600 = ( ~n3576 & n9811 ) | ( ~n3576 & n20599 ) | ( n9811 & n20599 ) ;
  assign n20601 = n13346 | n20600 ;
  assign n20603 = n20602 ^ n20601 ^ n5981 ;
  assign n20604 = n505 & n10523 ;
  assign n20605 = n6359 & ~n18657 ;
  assign n20606 = n2064 & n20605 ;
  assign n20607 = n20606 ^ n18652 ^ 1'b0 ;
  assign n20608 = n20604 & ~n20607 ;
  assign n20609 = n612 & ~n9726 ;
  assign n20610 = n4552 & n20609 ;
  assign n20611 = n730 & ~n20610 ;
  assign n20612 = ~n1742 & n20611 ;
  assign n20613 = n8205 & n12964 ;
  assign n20614 = n250 & ~n2898 ;
  assign n20615 = ( n4529 & n4701 ) | ( n4529 & ~n20614 ) | ( n4701 & ~n20614 ) ;
  assign n20616 = n11995 | n20615 ;
  assign n20617 = n2299 | n4285 ;
  assign n20618 = n548 & ~n20617 ;
  assign n20619 = ~n6130 & n20618 ;
  assign n20620 = n1965 | n6547 ;
  assign n20621 = n20620 ^ n6332 ^ 1'b0 ;
  assign n20622 = n11050 | n20621 ;
  assign n20623 = n15612 ^ n12402 ^ 1'b0 ;
  assign n20624 = n20622 | n20623 ;
  assign n20625 = n18644 ^ n8713 ^ 1'b0 ;
  assign n20626 = n20624 | n20625 ;
  assign n20629 = n2747 | n17602 ;
  assign n20627 = n14879 ^ n4029 ^ 1'b0 ;
  assign n20628 = n20627 ^ n9887 ^ n438 ;
  assign n20630 = n20629 ^ n20628 ^ n18931 ;
  assign n20631 = n1266 & ~n15356 ;
  assign n20632 = n20631 ^ n2623 ^ 1'b0 ;
  assign n20633 = ~n17890 & n20632 ;
  assign n20634 = n11761 ^ n10253 ^ 1'b0 ;
  assign n20635 = ~n4929 & n16906 ;
  assign n20636 = n2353 & n14211 ;
  assign n20637 = n11476 ^ n1053 ^ 1'b0 ;
  assign n20638 = n16944 & ~n20637 ;
  assign n20639 = ~n3557 & n20638 ;
  assign n20640 = n18168 ^ n8750 ^ n5904 ;
  assign n20641 = ~n6430 & n20640 ;
  assign n20642 = n9971 & n14123 ;
  assign n20643 = n1610 & ~n3991 ;
  assign n20644 = ( ~n7328 & n13297 ) | ( ~n7328 & n20643 ) | ( n13297 & n20643 ) ;
  assign n20645 = n1416 & ~n6671 ;
  assign n20646 = ~n20644 & n20645 ;
  assign n20647 = ( x98 & ~n4782 ) | ( x98 & n16774 ) | ( ~n4782 & n16774 ) ;
  assign n20648 = n5652 & n20647 ;
  assign n20649 = ( n510 & n892 ) | ( n510 & n1700 ) | ( n892 & n1700 ) ;
  assign n20650 = n8252 & ~n16096 ;
  assign n20651 = n20650 ^ n2364 ^ 1'b0 ;
  assign n20652 = n20649 & n20651 ;
  assign n20653 = n6515 ^ n3264 ^ 1'b0 ;
  assign n20654 = n19144 ^ n11995 ^ n635 ;
  assign n20655 = ~n148 & n6286 ;
  assign n20656 = n20655 ^ n8914 ^ 1'b0 ;
  assign n20657 = ~n5926 & n17462 ;
  assign n20658 = n5527 & n20657 ;
  assign n20659 = ~n12121 & n20658 ;
  assign n20660 = n8481 ^ n7561 ^ 1'b0 ;
  assign n20661 = n12853 | n20660 ;
  assign n20662 = n5168 | n20661 ;
  assign n20663 = n6895 | n20662 ;
  assign n20664 = n13037 ^ n10626 ^ 1'b0 ;
  assign n20665 = n8617 & ~n20664 ;
  assign n20666 = n1520 ^ n1438 ^ 1'b0 ;
  assign n20667 = n17878 ^ n12369 ^ 1'b0 ;
  assign n20668 = n6141 | n20667 ;
  assign n20669 = n5185 & ~n20668 ;
  assign n20670 = n20666 & n20669 ;
  assign n20671 = n17761 ^ n14890 ^ 1'b0 ;
  assign n20672 = n13955 & ~n17892 ;
  assign n20673 = n11356 ^ n10448 ^ 1'b0 ;
  assign n20674 = n8845 | n20673 ;
  assign n20675 = ~n1179 & n16155 ;
  assign n20678 = ( n883 & ~n1950 ) | ( n883 & n3929 ) | ( ~n1950 & n3929 ) ;
  assign n20676 = ~n6665 & n16993 ;
  assign n20677 = ~n20554 & n20676 ;
  assign n20679 = n20678 ^ n20677 ^ n16693 ;
  assign n20680 = n13003 ^ n6758 ^ n3301 ;
  assign n20681 = ~n220 & n18275 ;
  assign n20682 = ~n1000 & n8466 ;
  assign n20683 = x83 & n20682 ;
  assign n20684 = ~n15964 & n20683 ;
  assign n20685 = n19488 ^ n6743 ^ n1452 ;
  assign n20686 = n13354 ^ n497 ^ 1'b0 ;
  assign n20687 = n20685 | n20686 ;
  assign n20688 = n10747 ^ n1025 ^ 1'b0 ;
  assign n20689 = n1762 & ~n20688 ;
  assign n20690 = n3363 | n13184 ;
  assign n20691 = n467 & n20690 ;
  assign n20692 = ~n20689 & n20691 ;
  assign n20693 = n3628 | n7462 ;
  assign n20694 = n14359 & ~n20693 ;
  assign n20695 = ~x71 & n4306 ;
  assign n20700 = n8966 | n17910 ;
  assign n20699 = n15633 ^ n4516 ^ 1'b0 ;
  assign n20697 = n4600 | n10769 ;
  assign n20696 = n997 & n11483 ;
  assign n20698 = n20697 ^ n20696 ^ 1'b0 ;
  assign n20701 = n20700 ^ n20699 ^ n20698 ;
  assign n20702 = n2833 ^ n1251 ^ 1'b0 ;
  assign n20703 = n17030 ^ n9017 ^ 1'b0 ;
  assign n20704 = n9649 ^ n1668 ^ 1'b0 ;
  assign n20705 = n922 & n6119 ;
  assign n20706 = n15201 ^ n14405 ^ n9198 ;
  assign n20707 = n12149 & ~n20706 ;
  assign n20708 = ~n10286 & n12149 ;
  assign n20709 = ( n2043 & n2146 ) | ( n2043 & ~n9068 ) | ( n2146 & ~n9068 ) ;
  assign n20710 = ( ~n6182 & n10426 ) | ( ~n6182 & n19842 ) | ( n10426 & n19842 ) ;
  assign n20713 = n20224 ^ n4247 ^ n3516 ;
  assign n20714 = ~n12893 & n20713 ;
  assign n20715 = n2428 & n20714 ;
  assign n20711 = n844 & n1827 ;
  assign n20712 = n442 & n20711 ;
  assign n20716 = n20715 ^ n20712 ^ 1'b0 ;
  assign n20717 = n4748 ^ n4626 ^ 1'b0 ;
  assign n20718 = n1185 | n19094 ;
  assign n20719 = n6763 & ~n18937 ;
  assign n20720 = n18112 ^ n3009 ^ 1'b0 ;
  assign n20721 = n14054 & n20720 ;
  assign n20722 = n13476 | n15633 ;
  assign n20723 = ~n1613 & n2457 ;
  assign n20724 = n5878 & n20723 ;
  assign n20725 = n6959 | n8886 ;
  assign n20726 = n20725 ^ x75 ^ 1'b0 ;
  assign n20727 = n3960 & ~n20726 ;
  assign n20729 = n10181 ^ n6201 ^ 1'b0 ;
  assign n20728 = n6983 & n10858 ;
  assign n20730 = n20729 ^ n20728 ^ 1'b0 ;
  assign n20731 = n8977 & ~n9832 ;
  assign n20732 = ~n11866 & n20731 ;
  assign n20733 = n1766 | n7031 ;
  assign n20734 = n12091 ^ n8603 ^ n6165 ;
  assign n20735 = n1183 & n20734 ;
  assign n20736 = n9031 & n20735 ;
  assign n20737 = n450 & n4085 ;
  assign n20738 = n19047 ^ n4151 ^ 1'b0 ;
  assign n20739 = ( n15880 & n18351 ) | ( n15880 & n20738 ) | ( n18351 & n20738 ) ;
  assign n20740 = n4771 ^ n4587 ^ n2169 ;
  assign n20741 = n20740 ^ n1040 ^ 1'b0 ;
  assign n20742 = n1418 & n5316 ;
  assign n20743 = n345 | n1041 ;
  assign n20744 = n9069 ^ n5888 ^ 1'b0 ;
  assign n20745 = n20743 & ~n20744 ;
  assign n20746 = ~n6117 & n14455 ;
  assign n20747 = n20746 ^ n7163 ^ 1'b0 ;
  assign n20748 = n3377 & ~n9327 ;
  assign n20749 = n20748 ^ n6940 ^ 1'b0 ;
  assign n20750 = n8678 & ~n20749 ;
  assign n20751 = ~n20747 & n20750 ;
  assign n20752 = n19888 ^ n8287 ^ 1'b0 ;
  assign n20753 = ~n14201 & n20752 ;
  assign n20754 = n20753 ^ n10395 ^ n1952 ;
  assign n20755 = n3580 & ~n3714 ;
  assign n20756 = n17733 & n20755 ;
  assign n20757 = n20756 ^ n7911 ^ n6407 ;
  assign n20758 = n3259 & n11328 ;
  assign n20759 = n6047 & n6526 ;
  assign n20760 = n15754 | n20759 ;
  assign n20761 = ~n7703 & n19652 ;
  assign n20762 = ~n19332 & n20761 ;
  assign n20763 = n2222 & n17487 ;
  assign n20764 = ( ~n13993 & n16289 ) | ( ~n13993 & n20763 ) | ( n16289 & n20763 ) ;
  assign n20765 = ~n6143 & n20764 ;
  assign n20766 = n15347 ^ n5061 ^ 1'b0 ;
  assign n20767 = n20765 & n20766 ;
  assign n20768 = n3006 & n12972 ;
  assign n20769 = ~n12536 & n20768 ;
  assign n20770 = n2487 & n3732 ;
  assign n20771 = ~n1758 & n20770 ;
  assign n20775 = n3714 & ~n5124 ;
  assign n20772 = n2112 ^ n1775 ^ 1'b0 ;
  assign n20773 = n13975 ^ n9020 ^ 1'b0 ;
  assign n20774 = ~n20772 & n20773 ;
  assign n20776 = n20775 ^ n20774 ^ n2605 ;
  assign n20777 = ( n2675 & ~n20771 ) | ( n2675 & n20776 ) | ( ~n20771 & n20776 ) ;
  assign n20778 = ( n5351 & ~n13733 ) | ( n5351 & n14738 ) | ( ~n13733 & n14738 ) ;
  assign n20779 = n1000 | n7622 ;
  assign n20780 = n3424 ^ n2581 ^ 1'b0 ;
  assign n20781 = n5448 & ~n20780 ;
  assign n20782 = n20781 ^ n10062 ^ 1'b0 ;
  assign n20783 = n1089 & n20782 ;
  assign n20784 = n13496 ^ n5909 ^ 1'b0 ;
  assign n20785 = ~n16645 & n20784 ;
  assign n20786 = ( ~n4097 & n14298 ) | ( ~n4097 & n16344 ) | ( n14298 & n16344 ) ;
  assign n20787 = n4779 & ~n9968 ;
  assign n20788 = n639 & n15951 ;
  assign n20789 = n9153 ^ n7022 ^ 1'b0 ;
  assign n20790 = n12932 ^ n12025 ^ 1'b0 ;
  assign n20791 = ~n20789 & n20790 ;
  assign n20792 = n8687 ^ n1360 ^ 1'b0 ;
  assign n20793 = n14308 ^ n13700 ^ n1059 ;
  assign n20794 = n20792 & n20793 ;
  assign n20795 = ~n13612 & n17044 ;
  assign n20796 = n15594 ^ n8471 ^ 1'b0 ;
  assign n20797 = n4827 & n13021 ;
  assign n20798 = n706 | n20797 ;
  assign n20799 = n10060 & ~n20798 ;
  assign n20800 = n20799 ^ n19614 ^ 1'b0 ;
  assign n20801 = n4611 & n20800 ;
  assign n20802 = ~n3374 & n20437 ;
  assign n20803 = n6223 & ~n12353 ;
  assign n20804 = n15946 ^ n5166 ^ 1'b0 ;
  assign n20805 = n562 | n20804 ;
  assign n20806 = n20805 ^ n3059 ^ 1'b0 ;
  assign n20807 = n11004 & ~n20806 ;
  assign n20808 = n13304 & n20807 ;
  assign n20809 = n20808 ^ n1407 ^ 1'b0 ;
  assign n20810 = n18690 ^ n4295 ^ 1'b0 ;
  assign n20811 = n8075 | n20810 ;
  assign n20812 = n2634 | n20811 ;
  assign n20813 = n14250 & ~n20812 ;
  assign n20814 = n306 & ~n5288 ;
  assign n20815 = n20814 ^ n13063 ^ 1'b0 ;
  assign n20816 = n13947 & ~n20815 ;
  assign n20817 = n497 & n16695 ;
  assign n20818 = ~n9555 & n20817 ;
  assign n20819 = ~n1683 & n20818 ;
  assign n20820 = ~n13361 & n17584 ;
  assign n20821 = n20820 ^ n18406 ^ 1'b0 ;
  assign n20822 = n12350 ^ n3529 ^ 1'b0 ;
  assign n20823 = n2197 ^ n1562 ^ 1'b0 ;
  assign n20824 = n20467 & n20823 ;
  assign n20825 = n20824 ^ n20689 ^ 1'b0 ;
  assign n20826 = n13510 & ~n16066 ;
  assign n20827 = n7936 & n20826 ;
  assign n20828 = n962 ^ n548 ^ x117 ;
  assign n20829 = n16120 & n16245 ;
  assign n20830 = ~n20828 & n20829 ;
  assign n20831 = n20830 ^ n2140 ^ 1'b0 ;
  assign n20832 = n809 | n1149 ;
  assign n20833 = n3931 | n20832 ;
  assign n20834 = n9464 ^ n8717 ^ 1'b0 ;
  assign n20835 = n20833 & n20834 ;
  assign n20836 = ( n4796 & n5552 ) | ( n4796 & ~n6867 ) | ( n5552 & ~n6867 ) ;
  assign n20837 = n3093 & n20836 ;
  assign n20838 = ~n3102 & n20837 ;
  assign n20839 = ~n2229 & n5963 ;
  assign n20841 = n7116 & n7358 ;
  assign n20842 = n20841 ^ n12772 ^ 1'b0 ;
  assign n20840 = n3935 | n7251 ;
  assign n20843 = n20842 ^ n20840 ^ 1'b0 ;
  assign n20844 = ~n159 & n691 ;
  assign n20845 = n3308 ^ n2011 ^ 1'b0 ;
  assign n20846 = n18947 ^ n7420 ^ 1'b0 ;
  assign n20847 = n2611 & n20846 ;
  assign n20850 = n746 & n16500 ;
  assign n20848 = n7260 & n9169 ;
  assign n20849 = ~n5453 & n20848 ;
  assign n20851 = n20850 ^ n20849 ^ 1'b0 ;
  assign n20852 = n8862 | n12066 ;
  assign n20853 = n20852 ^ n1123 ^ 1'b0 ;
  assign n20854 = ~n2925 & n7583 ;
  assign n20856 = ~n1039 & n13947 ;
  assign n20857 = n20856 ^ n8620 ^ 1'b0 ;
  assign n20855 = ~n3524 & n17315 ;
  assign n20858 = n20857 ^ n20855 ^ 1'b0 ;
  assign n20859 = ~n2527 & n6796 ;
  assign n20860 = ( ~n5538 & n5629 ) | ( ~n5538 & n20859 ) | ( n5629 & n20859 ) ;
  assign n20861 = n20428 ^ n17558 ^ n4204 ;
  assign n20862 = ~n5539 & n10153 ;
  assign n20863 = n11041 ^ n8500 ^ 1'b0 ;
  assign n20864 = ~n2958 & n20863 ;
  assign n20865 = n7566 & n20864 ;
  assign n20866 = n20865 ^ n13233 ^ 1'b0 ;
  assign n20867 = ~n2436 & n11925 ;
  assign n20868 = n11341 ^ n2667 ^ 1'b0 ;
  assign n20869 = n20867 & n20868 ;
  assign n20871 = n6998 & n12319 ;
  assign n20870 = n19804 ^ n8099 ^ 1'b0 ;
  assign n20872 = n20871 ^ n20870 ^ 1'b0 ;
  assign n20873 = n7653 ^ n3760 ^ 1'b0 ;
  assign n20874 = n13395 & ~n20873 ;
  assign n20875 = n20872 & n20874 ;
  assign n20876 = n7786 ^ n4745 ^ 1'b0 ;
  assign n20877 = ( ~n4999 & n5804 ) | ( ~n4999 & n15314 ) | ( n5804 & n15314 ) ;
  assign n20878 = n13158 ^ n5924 ^ 1'b0 ;
  assign n20879 = n3419 | n20878 ;
  assign n20880 = n16366 | n20879 ;
  assign n20881 = n3994 & ~n20880 ;
  assign n20882 = n7488 & ~n15641 ;
  assign n20883 = n16905 ^ n4449 ^ 1'b0 ;
  assign n20884 = n10296 & n20883 ;
  assign n20885 = n16005 & ~n20884 ;
  assign n20886 = n7573 & n20885 ;
  assign n20887 = n16267 & n20886 ;
  assign n20888 = n14662 ^ n8040 ^ 1'b0 ;
  assign n20889 = ~n2356 & n20888 ;
  assign n20893 = n4025 & ~n12771 ;
  assign n20890 = n5432 ^ n3347 ^ 1'b0 ;
  assign n20891 = n7453 & n20890 ;
  assign n20892 = ~n3175 & n20891 ;
  assign n20894 = n20893 ^ n20892 ^ 1'b0 ;
  assign n20895 = ~n12304 & n12544 ;
  assign n20896 = n20894 & n20895 ;
  assign n20897 = ~n4150 & n4665 ;
  assign n20898 = n20897 ^ n6612 ^ 1'b0 ;
  assign n20899 = n707 & ~n20898 ;
  assign n20900 = n10288 ^ n3306 ^ 1'b0 ;
  assign n20901 = n7413 & n14108 ;
  assign n20902 = n20901 ^ n15900 ^ 1'b0 ;
  assign n20903 = n20900 & n20902 ;
  assign n20904 = n13711 ^ n10125 ^ 1'b0 ;
  assign n20905 = n14920 ^ n7720 ^ 1'b0 ;
  assign n20906 = n20904 & ~n20905 ;
  assign n20909 = ~n2398 & n13084 ;
  assign n20910 = n4268 & ~n8154 ;
  assign n20911 = ~n20909 & n20910 ;
  assign n20907 = ~n6097 & n17686 ;
  assign n20908 = n3344 & n20907 ;
  assign n20912 = n20911 ^ n20908 ^ 1'b0 ;
  assign n20914 = n8994 & ~n20743 ;
  assign n20913 = n1906 & ~n2039 ;
  assign n20915 = n20914 ^ n20913 ^ 1'b0 ;
  assign n20916 = n3340 & n13575 ;
  assign n20917 = n20916 ^ n1385 ^ 1'b0 ;
  assign n20918 = n20917 ^ n6183 ^ 1'b0 ;
  assign n20919 = n6027 & ~n10533 ;
  assign n20920 = ( n3281 & n19995 ) | ( n3281 & ~n20919 ) | ( n19995 & ~n20919 ) ;
  assign n20921 = n7928 & ~n20337 ;
  assign n20922 = n13207 & ~n15612 ;
  assign n20923 = n20922 ^ n790 ^ 1'b0 ;
  assign n20924 = n6159 | n8288 ;
  assign n20925 = n20924 ^ n9945 ^ 1'b0 ;
  assign n20926 = n14308 ^ n2912 ^ 1'b0 ;
  assign n20927 = n16017 & ~n20926 ;
  assign n20928 = n7448 | n17838 ;
  assign n20929 = n10340 & ~n20928 ;
  assign n20931 = n12472 ^ n1169 ^ 1'b0 ;
  assign n20930 = x54 & n326 ;
  assign n20932 = n20931 ^ n20930 ^ n8977 ;
  assign n20933 = n17216 ^ n6075 ^ 1'b0 ;
  assign n20934 = ~n20932 & n20933 ;
  assign n20935 = n1929 & ~n12788 ;
  assign n20936 = ~n3518 & n13097 ;
  assign n20937 = n20936 ^ n7499 ^ 1'b0 ;
  assign n20938 = n20937 ^ n17266 ^ 1'b0 ;
  assign n20939 = ~n9498 & n10401 ;
  assign n20940 = n14340 & n20939 ;
  assign n20941 = n20940 ^ n5705 ^ 1'b0 ;
  assign n20942 = ~n3376 & n12522 ;
  assign n20943 = n9960 ^ n8599 ^ n5070 ;
  assign n20944 = ( n551 & ~n1654 ) | ( n551 & n20943 ) | ( ~n1654 & n20943 ) ;
  assign n20945 = ~n20330 & n20944 ;
  assign n20946 = n12019 & n20945 ;
  assign n20947 = n20946 ^ n1265 ^ 1'b0 ;
  assign n20948 = n2577 & n17788 ;
  assign n20949 = n8950 & n20948 ;
  assign n20950 = n20949 ^ n14235 ^ n4527 ;
  assign n20951 = n7971 ^ n932 ^ 1'b0 ;
  assign n20952 = n4779 & n20951 ;
  assign n20953 = ~n20951 & n20952 ;
  assign n20954 = x67 & ~n4270 ;
  assign n20955 = n8544 & n20954 ;
  assign n20956 = n15727 | n16207 ;
  assign n20957 = n16805 & ~n20956 ;
  assign n20958 = n8476 | n19359 ;
  assign n20959 = n577 & ~n2925 ;
  assign n20960 = ~n20644 & n20959 ;
  assign n20962 = n16290 ^ n6072 ^ 1'b0 ;
  assign n20961 = ( n4400 & n7358 ) | ( n4400 & n8657 ) | ( n7358 & n8657 ) ;
  assign n20963 = n20962 ^ n20961 ^ n5693 ;
  assign n20964 = n20963 ^ n16677 ^ n9321 ;
  assign n20965 = n8361 & ~n20218 ;
  assign n20966 = n2887 & n20965 ;
  assign n20967 = n20966 ^ n7717 ^ 1'b0 ;
  assign n20968 = n7425 ^ n6490 ^ n952 ;
  assign n20969 = ~n9012 & n11673 ;
  assign n20970 = n20969 ^ n2214 ^ 1'b0 ;
  assign n20971 = n3093 | n3550 ;
  assign n20974 = n1693 ^ x83 ^ 1'b0 ;
  assign n20972 = n6455 ^ n2803 ^ 1'b0 ;
  assign n20973 = n18846 & ~n20972 ;
  assign n20975 = n20974 ^ n20973 ^ 1'b0 ;
  assign n20976 = n2759 & ~n20975 ;
  assign n20977 = n20976 ^ n15316 ^ 1'b0 ;
  assign n20978 = n5263 & n20977 ;
  assign n20979 = n7234 ^ n4407 ^ n3538 ;
  assign n20980 = n20979 ^ n1168 ^ 1'b0 ;
  assign n20981 = n12560 & ~n20980 ;
  assign n20982 = n197 & n6921 ;
  assign n20983 = n20982 ^ n8169 ^ n7768 ;
  assign n20984 = n9562 ^ n1489 ^ 1'b0 ;
  assign n20985 = n11544 ^ n4610 ^ 1'b0 ;
  assign n20986 = ( n13060 & n20984 ) | ( n13060 & n20985 ) | ( n20984 & n20985 ) ;
  assign n20987 = ~n3896 & n11780 ;
  assign n20988 = n20987 ^ n13559 ^ 1'b0 ;
  assign n20989 = n20988 ^ n19062 ^ 1'b0 ;
  assign n20990 = n18373 ^ n11940 ^ 1'b0 ;
  assign n20991 = ( n8300 & ~n10835 ) | ( n8300 & n20990 ) | ( ~n10835 & n20990 ) ;
  assign n20992 = n8094 | n16443 ;
  assign n20993 = n12771 | n20992 ;
  assign n20994 = n4327 ^ n1686 ^ 1'b0 ;
  assign n20995 = n2243 & n20994 ;
  assign n20996 = n10888 & ~n20995 ;
  assign n20998 = ~n5291 & n7872 ;
  assign n20999 = n20998 ^ n3619 ^ 1'b0 ;
  assign n20997 = ( ~n9814 & n12150 ) | ( ~n9814 & n13186 ) | ( n12150 & n13186 ) ;
  assign n21000 = n20999 ^ n20997 ^ 1'b0 ;
  assign n21001 = n18871 | n21000 ;
  assign n21002 = n2059 & ~n8637 ;
  assign n21003 = n21002 ^ n1356 ^ 1'b0 ;
  assign n21006 = n4858 | n9717 ;
  assign n21005 = n6015 & n10449 ;
  assign n21007 = n21006 ^ n21005 ^ 1'b0 ;
  assign n21004 = n2831 | n14662 ;
  assign n21008 = n21007 ^ n21004 ^ 1'b0 ;
  assign n21009 = ~n1667 & n5736 ;
  assign n21010 = n21009 ^ n1511 ^ 1'b0 ;
  assign n21011 = n21010 ^ n7206 ^ 1'b0 ;
  assign n21012 = n1235 & ~n12274 ;
  assign n21013 = n7162 ^ n4879 ^ 1'b0 ;
  assign n21014 = ~n2334 & n5818 ;
  assign n21015 = n10241 ^ n8920 ^ n2770 ;
  assign n21016 = n8982 ^ n616 ^ 1'b0 ;
  assign n21017 = n6972 | n21016 ;
  assign n21018 = ( n7098 & ~n21015 ) | ( n7098 & n21017 ) | ( ~n21015 & n21017 ) ;
  assign n21019 = n4787 & ~n21018 ;
  assign n21020 = n20859 ^ n11870 ^ 1'b0 ;
  assign n21021 = n17514 & ~n21020 ;
  assign n21022 = ( n3005 & n4026 ) | ( n3005 & ~n5025 ) | ( n4026 & ~n5025 ) ;
  assign n21023 = n21022 ^ n11401 ^ 1'b0 ;
  assign n21024 = n8622 ^ n2613 ^ 1'b0 ;
  assign n21025 = n1217 & ~n21024 ;
  assign n21026 = ~n2417 & n21025 ;
  assign n21027 = n6694 ^ n6401 ^ 1'b0 ;
  assign n21028 = n21026 & ~n21027 ;
  assign n21029 = n6813 & n11787 ;
  assign n21030 = x110 & ~n20858 ;
  assign n21031 = n21029 & n21030 ;
  assign n21032 = n12921 ^ n7069 ^ n4174 ;
  assign n21033 = n21032 ^ n20066 ^ 1'b0 ;
  assign n21034 = ~n20288 & n21033 ;
  assign n21035 = n7761 | n21034 ;
  assign n21043 = ~n3025 & n7123 ;
  assign n21044 = n21043 ^ n11075 ^ 1'b0 ;
  assign n21042 = n510 & ~n1200 ;
  assign n21045 = n21044 ^ n21042 ^ 1'b0 ;
  assign n21037 = n8129 & n11929 ;
  assign n21038 = n21037 ^ n7448 ^ n5538 ;
  assign n21036 = ~n254 & n15000 ;
  assign n21039 = n21038 ^ n21036 ^ 1'b0 ;
  assign n21040 = n3793 ^ n1449 ^ 1'b0 ;
  assign n21041 = ~n21039 & n21040 ;
  assign n21046 = n21045 ^ n21041 ^ n16616 ;
  assign n21048 = n380 | n798 ;
  assign n21047 = n6802 | n20246 ;
  assign n21049 = n21048 ^ n21047 ^ 1'b0 ;
  assign n21050 = n21049 ^ n9731 ^ n827 ;
  assign n21051 = n3660 & n7754 ;
  assign n21052 = n15953 ^ n12619 ^ 1'b0 ;
  assign n21053 = n21051 | n21052 ;
  assign n21054 = n9327 | n11393 ;
  assign n21055 = ~n15831 & n18832 ;
  assign n21056 = ~n21054 & n21055 ;
  assign n21058 = n8582 ^ n7217 ^ 1'b0 ;
  assign n21059 = n1479 & ~n21058 ;
  assign n21057 = n13580 | n18788 ;
  assign n21060 = n21059 ^ n21057 ^ 1'b0 ;
  assign n21061 = n16185 ^ n271 ^ 1'b0 ;
  assign n21062 = n11265 & ~n21061 ;
  assign n21063 = n21062 ^ n17305 ^ n1451 ;
  assign n21064 = n5610 ^ n4211 ^ 1'b0 ;
  assign n21065 = ~x87 & n19431 ;
  assign n21066 = n2162 & n7107 ;
  assign n21067 = n21066 ^ n1762 ^ 1'b0 ;
  assign n21068 = n5485 ^ n2637 ^ n462 ;
  assign n21069 = n21068 ^ x10 ^ 1'b0 ;
  assign n21071 = n454 & ~n15668 ;
  assign n21072 = n21071 ^ n2204 ^ 1'b0 ;
  assign n21070 = x95 & ~n1621 ;
  assign n21073 = n21072 ^ n21070 ^ n9433 ;
  assign n21074 = ~n295 & n4277 ;
  assign n21075 = n21074 ^ n5900 ^ 1'b0 ;
  assign n21076 = n18502 | n21075 ;
  assign n21077 = n21076 ^ n11630 ^ 1'b0 ;
  assign n21078 = n7785 & n9950 ;
  assign n21079 = ~n7717 & n21078 ;
  assign n21080 = n615 | n1004 ;
  assign n21081 = n9270 | n21080 ;
  assign n21082 = n21081 ^ n2861 ^ 1'b0 ;
  assign n21083 = ( n2143 & n7561 ) | ( n2143 & ~n21082 ) | ( n7561 & ~n21082 ) ;
  assign n21084 = ( n908 & n1654 ) | ( n908 & ~n21083 ) | ( n1654 & ~n21083 ) ;
  assign n21085 = n10259 & ~n21084 ;
  assign n21086 = n21079 & n21085 ;
  assign n21087 = ( n527 & n19334 ) | ( n527 & ~n20961 ) | ( n19334 & ~n20961 ) ;
  assign n21088 = n9203 | n15438 ;
  assign n21089 = n403 | n10843 ;
  assign n21090 = n6792 | n9057 ;
  assign n21091 = ~n8912 & n17080 ;
  assign n21092 = n21091 ^ n20456 ^ 1'b0 ;
  assign n21093 = n16202 ^ n5765 ^ 1'b0 ;
  assign n21094 = n8994 & ~n21093 ;
  assign n21095 = ( n3865 & ~n10153 ) | ( n3865 & n21094 ) | ( ~n10153 & n21094 ) ;
  assign n21096 = n18209 ^ n16390 ^ 1'b0 ;
  assign n21097 = n7475 | n8598 ;
  assign n21098 = n12398 | n21097 ;
  assign n21099 = n6186 & n21098 ;
  assign n21100 = n1687 | n15167 ;
  assign n21101 = n19348 & ~n21100 ;
  assign n21102 = n19494 ^ n4552 ^ 1'b0 ;
  assign n21103 = ( ~n2997 & n17358 ) | ( ~n2997 & n21102 ) | ( n17358 & n21102 ) ;
  assign n21104 = n2719 | n20743 ;
  assign n21105 = n21104 ^ n13981 ^ n5452 ;
  assign n21106 = ( ~n3213 & n15787 ) | ( ~n3213 & n21105 ) | ( n15787 & n21105 ) ;
  assign n21107 = ~n4333 & n11569 ;
  assign n21108 = n21107 ^ n811 ^ 1'b0 ;
  assign n21109 = ~n8466 & n12274 ;
  assign n21110 = n3853 & n5837 ;
  assign n21111 = n21109 & n21110 ;
  assign n21112 = n18984 ^ n2431 ^ 1'b0 ;
  assign n21113 = n11449 | n14525 ;
  assign n21114 = n12317 ^ n7642 ^ 1'b0 ;
  assign n21115 = ~n14398 & n21114 ;
  assign n21116 = n18657 ^ n8148 ^ 1'b0 ;
  assign n21117 = ( ~n2431 & n13107 ) | ( ~n2431 & n21116 ) | ( n13107 & n21116 ) ;
  assign n21118 = n3904 ^ n146 ^ 1'b0 ;
  assign n21119 = ~n9009 & n21118 ;
  assign n21120 = n9278 ^ n8816 ^ 1'b0 ;
  assign n21121 = n10662 & ~n21120 ;
  assign n21122 = n650 | n5296 ;
  assign n21123 = n21121 | n21122 ;
  assign n21124 = n21123 ^ n3155 ^ 1'b0 ;
  assign n21125 = n13680 | n21124 ;
  assign n21126 = ( n630 & n4079 ) | ( n630 & n10526 ) | ( n4079 & n10526 ) ;
  assign n21127 = ( n1040 & n15226 ) | ( n1040 & n21126 ) | ( n15226 & n21126 ) ;
  assign n21128 = n12104 & n20128 ;
  assign n21129 = n12048 & n16421 ;
  assign n21130 = ( n2079 & ~n21128 ) | ( n2079 & n21129 ) | ( ~n21128 & n21129 ) ;
  assign n21131 = n14942 ^ n2035 ^ 1'b0 ;
  assign n21132 = n8974 & n21131 ;
  assign n21133 = n10649 & ~n18941 ;
  assign n21134 = ~n17614 & n17828 ;
  assign n21135 = n3439 | n9450 ;
  assign n21136 = n21135 ^ n696 ^ 1'b0 ;
  assign n21137 = n12535 & ~n21136 ;
  assign n21138 = n7908 & n21137 ;
  assign n21139 = n20224 ^ n6675 ^ 1'b0 ;
  assign n21140 = ( n2577 & n8886 ) | ( n2577 & ~n21139 ) | ( n8886 & ~n21139 ) ;
  assign n21141 = n5610 ^ n2223 ^ 1'b0 ;
  assign n21142 = n5277 & n21141 ;
  assign n21143 = ~n13496 & n21142 ;
  assign n21144 = n12571 ^ n8974 ^ n3347 ;
  assign n21145 = n21144 ^ n5217 ^ 1'b0 ;
  assign n21146 = n11019 | n21145 ;
  assign n21147 = n9768 & n17445 ;
  assign n21148 = ( n1559 & n2817 ) | ( n1559 & ~n21147 ) | ( n2817 & ~n21147 ) ;
  assign n21149 = n7978 & ~n9558 ;
  assign n21150 = n21149 ^ n2744 ^ 1'b0 ;
  assign n21151 = ( ~n5326 & n7104 ) | ( ~n5326 & n7559 ) | ( n7104 & n7559 ) ;
  assign n21152 = ( ~n10125 & n21150 ) | ( ~n10125 & n21151 ) | ( n21150 & n21151 ) ;
  assign n21153 = n2222 & n3979 ;
  assign n21154 = n21153 ^ n9735 ^ 1'b0 ;
  assign n21155 = n12487 & n21154 ;
  assign n21156 = ~n8931 & n21155 ;
  assign n21158 = n14184 ^ n9524 ^ 1'b0 ;
  assign n21159 = ~n13050 & n21158 ;
  assign n21157 = n14756 & ~n15223 ;
  assign n21160 = n21159 ^ n21157 ^ 1'b0 ;
  assign n21161 = ( n1681 & ~n11272 ) | ( n1681 & n18796 ) | ( ~n11272 & n18796 ) ;
  assign n21162 = ( x100 & ~n1305 ) | ( x100 & n3617 ) | ( ~n1305 & n3617 ) ;
  assign n21163 = n9518 | n11921 ;
  assign n21164 = n5217 | n21163 ;
  assign n21165 = ~n6607 & n10039 ;
  assign n21166 = n20562 ^ n4717 ^ 1'b0 ;
  assign n21167 = n5951 & ~n21166 ;
  assign n21168 = ~n4780 & n8232 ;
  assign n21169 = n21168 ^ n20312 ^ 1'b0 ;
  assign n21170 = ( n863 & n9737 ) | ( n863 & n14487 ) | ( n9737 & n14487 ) ;
  assign n21171 = n21170 ^ n10865 ^ 1'b0 ;
  assign n21172 = n803 & ~n21171 ;
  assign n21173 = n2333 | n8715 ;
  assign n21174 = n7924 & n21173 ;
  assign n21175 = n13012 & ~n15638 ;
  assign n21176 = ( ~n2173 & n4641 ) | ( ~n2173 & n11298 ) | ( n4641 & n11298 ) ;
  assign n21180 = n8163 | n10921 ;
  assign n21178 = n1305 | n14372 ;
  assign n21179 = ~n11696 & n21178 ;
  assign n21181 = n21180 ^ n21179 ^ 1'b0 ;
  assign n21177 = n844 & ~n4194 ;
  assign n21182 = n21181 ^ n21177 ^ 1'b0 ;
  assign n21183 = ~n4388 & n12621 ;
  assign n21184 = n7399 ^ n3404 ^ 1'b0 ;
  assign n21185 = n21183 & n21184 ;
  assign n21186 = n9385 & n17096 ;
  assign n21187 = n18672 ^ n1295 ^ 1'b0 ;
  assign n21188 = ~n8365 & n21187 ;
  assign n21189 = n20514 ^ n3158 ^ n584 ;
  assign n21190 = n1498 & n15157 ;
  assign n21191 = n21190 ^ n4648 ^ 1'b0 ;
  assign n21192 = ~n21189 & n21191 ;
  assign n21193 = n11568 ^ n3639 ^ 1'b0 ;
  assign n21194 = n5504 ^ n3255 ^ 1'b0 ;
  assign n21195 = n6274 & n21194 ;
  assign n21196 = ( n4420 & ~n11107 ) | ( n4420 & n12006 ) | ( ~n11107 & n12006 ) ;
  assign n21197 = n21196 ^ n12520 ^ 1'b0 ;
  assign n21198 = n18177 ^ n13471 ^ n7893 ;
  assign n21199 = n1414 & ~n4957 ;
  assign n21200 = ~n1414 & n21199 ;
  assign n21201 = n2113 | n19591 ;
  assign n21202 = n21201 ^ n10785 ^ 1'b0 ;
  assign n21203 = n21202 ^ n7223 ^ 1'b0 ;
  assign n21204 = n21203 ^ n19109 ^ 1'b0 ;
  assign n21205 = ~n21200 & n21204 ;
  assign n21206 = n11635 | n19053 ;
  assign n21207 = n14509 & ~n20797 ;
  assign n21208 = ~n11519 & n21207 ;
  assign n21209 = n6999 & ~n9210 ;
  assign n21210 = n21208 & n21209 ;
  assign n21211 = n8001 & n21210 ;
  assign n21213 = n9711 & ~n18801 ;
  assign n21214 = ~n16433 & n21213 ;
  assign n21212 = ~n2909 & n7620 ;
  assign n21215 = n21214 ^ n21212 ^ 1'b0 ;
  assign n21216 = n19325 | n19591 ;
  assign n21217 = n21216 ^ n13662 ^ 1'b0 ;
  assign n21218 = n9145 | n9263 ;
  assign n21219 = n21218 ^ n7796 ^ 1'b0 ;
  assign n21220 = n21219 ^ n5844 ^ 1'b0 ;
  assign n21221 = ~n12246 & n21220 ;
  assign n21222 = n7182 & n16662 ;
  assign n21223 = ( n7176 & n12166 ) | ( n7176 & n12728 ) | ( n12166 & n12728 ) ;
  assign n21224 = ~n2839 & n2980 ;
  assign n21225 = ~n2980 & n21224 ;
  assign n21226 = n3161 & n21225 ;
  assign n21227 = n21226 ^ n10499 ^ 1'b0 ;
  assign n21228 = n11184 & n21227 ;
  assign n21229 = ~n21227 & n21228 ;
  assign n21230 = n21229 ^ n13347 ^ n10729 ;
  assign n21231 = n1061 ^ n138 ^ 1'b0 ;
  assign n21232 = n21231 ^ n9008 ^ 1'b0 ;
  assign n21233 = n11475 & n21232 ;
  assign n21234 = n19270 & n21233 ;
  assign n21235 = n21234 ^ n13712 ^ 1'b0 ;
  assign n21236 = n9722 | n15346 ;
  assign n21237 = n21236 ^ n1785 ^ 1'b0 ;
  assign n21238 = n21237 ^ n7620 ^ 1'b0 ;
  assign n21239 = ~n4745 & n21238 ;
  assign n21240 = n21239 ^ n10549 ^ 1'b0 ;
  assign n21241 = n16320 ^ n9172 ^ 1'b0 ;
  assign n21242 = n18315 & n21241 ;
  assign n21243 = n21242 ^ n2112 ^ 1'b0 ;
  assign n21244 = n12695 | n21243 ;
  assign n21245 = n6515 & ~n21244 ;
  assign n21246 = n7172 ^ n309 ^ 1'b0 ;
  assign n21247 = n11524 & n16748 ;
  assign n21248 = ~n5400 & n21247 ;
  assign n21249 = n3308 & ~n21248 ;
  assign n21250 = n16542 ^ x60 ^ 1'b0 ;
  assign n21251 = n21249 | n21250 ;
  assign n21252 = n19031 & ~n21251 ;
  assign n21253 = n16505 ^ n3256 ^ n239 ;
  assign n21254 = n425 & ~n7698 ;
  assign n21255 = n1286 & n21254 ;
  assign n21257 = ~n6053 & n10840 ;
  assign n21256 = n701 & n6842 ;
  assign n21258 = n21257 ^ n21256 ^ 1'b0 ;
  assign n21259 = n21258 ^ n12025 ^ 1'b0 ;
  assign n21260 = n10619 & n10970 ;
  assign n21261 = n8122 & n21260 ;
  assign n21262 = n3538 & ~n9222 ;
  assign n21263 = n21261 & n21262 ;
  assign n21264 = n3957 ^ n398 ^ 1'b0 ;
  assign n21265 = n21263 | n21264 ;
  assign n21267 = n1123 & n19699 ;
  assign n21268 = n1135 & n21267 ;
  assign n21269 = x89 & n21268 ;
  assign n21266 = n10808 ^ n10623 ^ 1'b0 ;
  assign n21270 = n21269 ^ n21266 ^ n14198 ;
  assign n21271 = n7622 & n16191 ;
  assign n21272 = ( n6578 & ~n14718 ) | ( n6578 & n21271 ) | ( ~n14718 & n21271 ) ;
  assign n21273 = n19646 ^ n17478 ^ n13064 ;
  assign n21274 = n1721 | n9963 ;
  assign n21275 = n21274 ^ n5693 ^ 1'b0 ;
  assign n21276 = ~n20992 & n21275 ;
  assign n21277 = n21276 ^ n7899 ^ 1'b0 ;
  assign n21278 = ~n381 & n1765 ;
  assign n21279 = ~n9013 & n21278 ;
  assign n21280 = n10670 ^ n10279 ^ 1'b0 ;
  assign n21281 = n13304 & n21280 ;
  assign n21282 = ~n11998 & n21281 ;
  assign n21283 = ~n9670 & n21282 ;
  assign n21284 = n19097 ^ n398 ^ 1'b0 ;
  assign n21285 = ~n5610 & n21284 ;
  assign n21286 = n6251 ^ n1286 ^ n908 ;
  assign n21287 = n9672 ^ n505 ^ 1'b0 ;
  assign n21288 = n10651 ^ n3467 ^ 1'b0 ;
  assign n21289 = n4405 & n21288 ;
  assign n21290 = ~n9505 & n21289 ;
  assign n21297 = n3149 & ~n15742 ;
  assign n21298 = n454 & ~n21297 ;
  assign n21299 = n21298 ^ n7597 ^ 1'b0 ;
  assign n21300 = n11335 ^ n1115 ^ 1'b0 ;
  assign n21301 = n2282 & n21300 ;
  assign n21302 = ( n487 & ~n21299 ) | ( n487 & n21301 ) | ( ~n21299 & n21301 ) ;
  assign n21294 = n9289 ^ n2099 ^ 1'b0 ;
  assign n21295 = ~n9010 & n21294 ;
  assign n21296 = n12833 | n21295 ;
  assign n21303 = n21302 ^ n21296 ^ 1'b0 ;
  assign n21291 = n6211 & n16266 ;
  assign n21292 = n3777 ^ n3418 ^ 1'b0 ;
  assign n21293 = n21291 | n21292 ;
  assign n21304 = n21303 ^ n21293 ^ 1'b0 ;
  assign n21305 = n5841 & ~n10300 ;
  assign n21306 = n8779 & ~n21305 ;
  assign n21307 = n15332 ^ n2464 ^ 1'b0 ;
  assign n21308 = n11559 ^ n2643 ^ 1'b0 ;
  assign n21309 = n3281 & n21275 ;
  assign n21310 = n21309 ^ n7792 ^ 1'b0 ;
  assign n21311 = n7674 & ~n21310 ;
  assign n21316 = ~n1842 & n12443 ;
  assign n21317 = n21316 ^ n5519 ^ 1'b0 ;
  assign n21312 = n1550 ^ n1149 ^ n480 ;
  assign n21313 = n11280 | n13649 ;
  assign n21314 = n21313 ^ n883 ^ 1'b0 ;
  assign n21315 = ~n21312 & n21314 ;
  assign n21318 = n21317 ^ n21315 ^ 1'b0 ;
  assign n21319 = n21318 ^ n1683 ^ 1'b0 ;
  assign n21320 = ~n3887 & n21319 ;
  assign n21321 = n13943 ^ n9245 ^ 1'b0 ;
  assign n21322 = n1387 & ~n19451 ;
  assign n21323 = n6217 & n21322 ;
  assign n21324 = n7819 | n15954 ;
  assign n21325 = n21324 ^ n4893 ^ 1'b0 ;
  assign n21326 = n13577 ^ n8052 ^ 1'b0 ;
  assign n21327 = n4373 ^ n748 ^ n353 ;
  assign n21328 = n21327 ^ n16126 ^ 1'b0 ;
  assign n21329 = n18714 ^ n2841 ^ 1'b0 ;
  assign n21330 = n3658 & ~n21329 ;
  assign n21332 = n8606 & n15082 ;
  assign n21333 = n11070 & n21332 ;
  assign n21334 = ~n4025 & n21333 ;
  assign n21335 = n17179 & n21334 ;
  assign n21331 = n10326 & ~n12475 ;
  assign n21336 = n21335 ^ n21331 ^ 1'b0 ;
  assign n21337 = n6561 & ~n11961 ;
  assign n21338 = n13207 ^ n700 ^ 1'b0 ;
  assign n21339 = n1244 & ~n9489 ;
  assign n21348 = n5457 | n6867 ;
  assign n21349 = n1954 & ~n21348 ;
  assign n21344 = n7986 | n12440 ;
  assign n21345 = n7692 & ~n21344 ;
  assign n21341 = n5464 & n11872 ;
  assign n21342 = n11553 & n21341 ;
  assign n21340 = n3802 & n15985 ;
  assign n21343 = n21342 ^ n21340 ^ n7139 ;
  assign n21346 = n21345 ^ n21343 ^ n1832 ;
  assign n21347 = ~n10068 & n21346 ;
  assign n21350 = n21349 ^ n21347 ^ 1'b0 ;
  assign n21351 = n21350 ^ n17226 ^ n6765 ;
  assign n21352 = ~n6502 & n17344 ;
  assign n21353 = n21352 ^ n10134 ^ 1'b0 ;
  assign n21354 = n2905 | n15571 ;
  assign n21355 = n21354 ^ n2912 ^ 1'b0 ;
  assign n21356 = n1042 & ~n3429 ;
  assign n21357 = n306 & ~n21356 ;
  assign n21359 = ( n4518 & ~n7003 ) | ( n4518 & n10833 ) | ( ~n7003 & n10833 ) ;
  assign n21360 = ~n15488 & n21359 ;
  assign n21361 = n21360 ^ n8278 ^ 1'b0 ;
  assign n21358 = n653 & ~n17512 ;
  assign n21362 = n21361 ^ n21358 ^ 1'b0 ;
  assign n21363 = n5336 ^ n4108 ^ 1'b0 ;
  assign n21364 = n1549 & ~n3660 ;
  assign n21365 = n1236 & n21364 ;
  assign n21366 = ~n10484 & n21365 ;
  assign n21367 = n10393 | n16728 ;
  assign n21368 = n18617 ^ n12346 ^ 1'b0 ;
  assign n21369 = ( x108 & ~n3008 ) | ( x108 & n10307 ) | ( ~n3008 & n10307 ) ;
  assign n21370 = n21369 ^ n19174 ^ 1'b0 ;
  assign n21371 = n20997 ^ n16428 ^ n4497 ;
  assign n21372 = n9800 ^ n7439 ^ 1'b0 ;
  assign n21373 = n3725 & n21372 ;
  assign n21374 = n21373 ^ n8100 ^ n2535 ;
  assign n21375 = n21374 ^ n6555 ^ 1'b0 ;
  assign n21376 = ~n19033 & n20162 ;
  assign n21377 = n12707 ^ n1578 ^ 1'b0 ;
  assign n21378 = ~n21376 & n21377 ;
  assign n21379 = n5468 | n14205 ;
  assign n21380 = n21379 ^ n14182 ^ 1'b0 ;
  assign n21381 = n3853 & n10560 ;
  assign n21382 = ~n21380 & n21381 ;
  assign n21383 = n764 | n2965 ;
  assign n21384 = n13196 ^ n9564 ^ n1418 ;
  assign n21385 = ( n186 & n852 ) | ( n186 & n1231 ) | ( n852 & n1231 ) ;
  assign n21386 = n21385 ^ n14890 ^ 1'b0 ;
  assign n21387 = x104 & n6999 ;
  assign n21388 = n13992 & n21387 ;
  assign n21389 = n10786 ^ n9015 ^ 1'b0 ;
  assign n21390 = n2396 & n8753 ;
  assign n21391 = n21390 ^ n5971 ^ 1'b0 ;
  assign n21392 = n3319 | n17330 ;
  assign n21393 = n15227 | n21392 ;
  assign n21394 = n12185 ^ n8148 ^ n753 ;
  assign n21395 = n3751 ^ n2459 ^ 1'b0 ;
  assign n21396 = n2264 | n21395 ;
  assign n21397 = n252 & ~n3465 ;
  assign n21398 = n21396 & n21397 ;
  assign n21399 = ( n11265 & ~n21394 ) | ( n11265 & n21398 ) | ( ~n21394 & n21398 ) ;
  assign n21400 = n5356 ^ n2064 ^ 1'b0 ;
  assign n21401 = n1979 | n21400 ;
  assign n21402 = n4286 & ~n21401 ;
  assign n21403 = n21402 ^ n19599 ^ 1'b0 ;
  assign n21404 = ( n12872 & n21399 ) | ( n12872 & ~n21403 ) | ( n21399 & ~n21403 ) ;
  assign n21405 = n8279 ^ n1002 ^ 1'b0 ;
  assign n21407 = n16063 ^ n5030 ^ 1'b0 ;
  assign n21408 = ~n10721 & n21407 ;
  assign n21409 = n7358 & n21408 ;
  assign n21406 = ~n7885 & n8104 ;
  assign n21410 = n21409 ^ n21406 ^ 1'b0 ;
  assign n21411 = n4010 & n17871 ;
  assign n21412 = n1753 | n4932 ;
  assign n21413 = ~n6573 & n10550 ;
  assign n21414 = n11467 & n21413 ;
  assign n21415 = n16049 & n18829 ;
  assign n21416 = n21415 ^ n8336 ^ 1'b0 ;
  assign n21417 = n4497 & n4854 ;
  assign n21418 = n11031 ^ n2064 ^ 1'b0 ;
  assign n21419 = ~n9368 & n21418 ;
  assign n21420 = n21419 ^ n18935 ^ 1'b0 ;
  assign n21421 = n442 | n21173 ;
  assign n21422 = n4929 ^ n4625 ^ n4419 ;
  assign n21423 = n19328 ^ n12559 ^ n4884 ;
  assign n21424 = n21423 ^ n5107 ^ 1'b0 ;
  assign n21425 = n654 & n21424 ;
  assign n21426 = ( n8148 & ~n21422 ) | ( n8148 & n21425 ) | ( ~n21422 & n21425 ) ;
  assign n21427 = ( n9689 & n19031 ) | ( n9689 & ~n21426 ) | ( n19031 & ~n21426 ) ;
  assign n21428 = n2915 & n6557 ;
  assign n21429 = n21428 ^ n17737 ^ 1'b0 ;
  assign n21430 = n19387 & n21429 ;
  assign n21431 = n8317 & ~n16328 ;
  assign n21432 = n21431 ^ n2853 ^ 1'b0 ;
  assign n21433 = n4019 ^ n1455 ^ 1'b0 ;
  assign n21434 = ~n2255 & n14238 ;
  assign n21435 = ( n6174 & n17628 ) | ( n6174 & ~n20317 ) | ( n17628 & ~n20317 ) ;
  assign n21437 = n3499 & n4779 ;
  assign n21438 = n21437 ^ n4757 ^ 1'b0 ;
  assign n21436 = ( ~n9635 & n11025 ) | ( ~n9635 & n11718 ) | ( n11025 & n11718 ) ;
  assign n21439 = n21438 ^ n21436 ^ 1'b0 ;
  assign n21444 = n14504 ^ n10085 ^ 1'b0 ;
  assign n21440 = n1973 | n12307 ;
  assign n21441 = n17584 ^ n4933 ^ 1'b0 ;
  assign n21442 = n21441 ^ n20616 ^ 1'b0 ;
  assign n21443 = n21440 & n21442 ;
  assign n21445 = n21444 ^ n21443 ^ n5790 ;
  assign n21446 = n6937 ^ n3758 ^ 1'b0 ;
  assign n21447 = n2310 & ~n5205 ;
  assign n21448 = n1866 & n21447 ;
  assign n21449 = ~n8780 & n11768 ;
  assign n21450 = n21449 ^ n1692 ^ 1'b0 ;
  assign n21451 = ~n21448 & n21450 ;
  assign n21452 = n706 & n4470 ;
  assign n21453 = n21452 ^ n9982 ^ 1'b0 ;
  assign n21454 = ( ~n4199 & n12120 ) | ( ~n4199 & n21278 ) | ( n12120 & n21278 ) ;
  assign n21455 = n7341 ^ n1973 ^ 1'b0 ;
  assign n21456 = n8730 & ~n21455 ;
  assign n21457 = n21456 ^ n16634 ^ 1'b0 ;
  assign n21458 = n20914 ^ n12212 ^ 1'b0 ;
  assign n21459 = n7924 ^ n332 ^ 1'b0 ;
  assign n21460 = n2823 & ~n10538 ;
  assign n21461 = n3620 & n21460 ;
  assign n21462 = ~n793 & n2495 ;
  assign n21463 = n16274 & n21462 ;
  assign n21464 = n8457 ^ n2945 ^ 1'b0 ;
  assign n21465 = n21464 ^ n15937 ^ n7067 ;
  assign n21466 = n13158 & n21465 ;
  assign n21467 = n21466 ^ n8512 ^ n8392 ;
  assign n21468 = n908 & n5324 ;
  assign n21469 = n2622 ^ n273 ^ 1'b0 ;
  assign n21470 = ~n2750 & n21469 ;
  assign n21471 = ~n2692 & n21470 ;
  assign n21472 = n18769 ^ n15426 ^ 1'b0 ;
  assign n21473 = n10769 ^ n2647 ^ 1'b0 ;
  assign n21474 = ~n4456 & n21473 ;
  assign n21475 = ~n1617 & n21474 ;
  assign n21476 = n13310 & n21475 ;
  assign n21477 = n8079 & ~n18782 ;
  assign n21478 = n18782 & n21477 ;
  assign n21479 = n566 & ~n9773 ;
  assign n21480 = n21479 ^ n748 ^ 1'b0 ;
  assign n21481 = n1860 & ~n4008 ;
  assign n21482 = n21481 ^ n18910 ^ 1'b0 ;
  assign n21483 = ( n4660 & ~n11270 ) | ( n4660 & n14698 ) | ( ~n11270 & n14698 ) ;
  assign n21484 = n21483 ^ n10048 ^ n9543 ;
  assign n21485 = n19019 ^ x25 ^ 1'b0 ;
  assign n21486 = n16742 & n21485 ;
  assign n21487 = ~n17368 & n21486 ;
  assign n21488 = n8570 & ~n12651 ;
  assign n21489 = ~n9014 & n21488 ;
  assign n21491 = n16290 ^ n837 ^ 1'b0 ;
  assign n21490 = ~n8268 & n17893 ;
  assign n21492 = n21491 ^ n21490 ^ 1'b0 ;
  assign n21493 = n13626 ^ n9013 ^ 1'b0 ;
  assign n21494 = x58 & n21493 ;
  assign n21495 = n5002 & n9634 ;
  assign n21496 = n21495 ^ n1781 ^ 1'b0 ;
  assign n21497 = ( ~n2720 & n2774 ) | ( ~n2720 & n21496 ) | ( n2774 & n21496 ) ;
  assign n21500 = ~x21 & n950 ;
  assign n21498 = n6886 | n8768 ;
  assign n21499 = n21498 ^ n17818 ^ 1'b0 ;
  assign n21501 = n21500 ^ n21499 ^ n5432 ;
  assign n21502 = ( n5402 & n8403 ) | ( n5402 & n9953 ) | ( n8403 & n9953 ) ;
  assign n21503 = ~n4075 & n21502 ;
  assign n21504 = n9604 & ~n11914 ;
  assign n21505 = ( n681 & n9963 ) | ( n681 & n11745 ) | ( n9963 & n11745 ) ;
  assign n21506 = n6821 & n21505 ;
  assign n21507 = n21506 ^ n16005 ^ 1'b0 ;
  assign n21508 = n4144 & ~n14186 ;
  assign n21509 = n21508 ^ n5731 ^ 1'b0 ;
  assign n21510 = n21509 ^ n21017 ^ n5440 ;
  assign n21511 = n136 & ~n7882 ;
  assign n21512 = n8782 ^ n1264 ^ 1'b0 ;
  assign n21513 = x41 & ~n21512 ;
  assign n21514 = n1374 | n5613 ;
  assign n21515 = n21514 ^ n7262 ^ 1'b0 ;
  assign n21516 = n280 & ~n21515 ;
  assign n21517 = n21516 ^ n5375 ^ 1'b0 ;
  assign n21518 = n6073 & n17865 ;
  assign n21519 = n401 & n17686 ;
  assign n21520 = n21519 ^ x99 ^ 1'b0 ;
  assign n21521 = n6684 ^ n2692 ^ 1'b0 ;
  assign n21523 = ~n3299 & n7068 ;
  assign n21524 = n18109 & n21523 ;
  assign n21522 = n623 ^ x69 ^ 1'b0 ;
  assign n21525 = n21524 ^ n21522 ^ n10827 ;
  assign n21526 = n15247 ^ n7642 ^ 1'b0 ;
  assign n21527 = n11021 | n12693 ;
  assign n21528 = n5036 ^ n972 ^ 1'b0 ;
  assign n21529 = n15167 & ~n21528 ;
  assign n21530 = ( n567 & n12160 ) | ( n567 & n21529 ) | ( n12160 & n21529 ) ;
  assign n21531 = n21530 ^ n15460 ^ 1'b0 ;
  assign n21532 = ~n20260 & n21531 ;
  assign n21533 = n11255 | n17587 ;
  assign n21534 = n19703 | n21533 ;
  assign n21535 = n21275 ^ n18859 ^ n8775 ;
  assign n21536 = n13566 ^ n12147 ^ n5816 ;
  assign n21537 = n15987 & n21536 ;
  assign n21538 = n8877 ^ n547 ^ 1'b0 ;
  assign n21539 = n21538 ^ n14160 ^ n3297 ;
  assign n21540 = n14626 ^ n2083 ^ 1'b0 ;
  assign n21541 = n15340 ^ n218 ^ 1'b0 ;
  assign n21542 = n13063 & n21541 ;
  assign n21543 = n11881 & ~n15734 ;
  assign n21544 = ~n4351 & n16357 ;
  assign n21545 = n4467 ^ n986 ^ 1'b0 ;
  assign n21546 = ( n4998 & ~n10340 ) | ( n4998 & n21545 ) | ( ~n10340 & n21545 ) ;
  assign n21547 = n12521 ^ n227 ^ 1'b0 ;
  assign n21548 = n8042 | n21547 ;
  assign n21549 = ( n417 & n6765 ) | ( n417 & n8733 ) | ( n6765 & n8733 ) ;
  assign n21550 = n785 | n21168 ;
  assign n21551 = n21549 | n21550 ;
  assign n21552 = n8347 ^ n4272 ^ 1'b0 ;
  assign n21553 = n21552 ^ n20078 ^ 1'b0 ;
  assign n21554 = n4141 ^ n4082 ^ n576 ;
  assign n21555 = n21554 ^ n18898 ^ 1'b0 ;
  assign n21556 = ~n12104 & n13386 ;
  assign n21557 = n9963 ^ n3786 ^ 1'b0 ;
  assign n21558 = n1714 & n21557 ;
  assign n21559 = ~n10758 & n21558 ;
  assign n21560 = n3221 & ~n21559 ;
  assign n21561 = n21560 ^ n16609 ^ 1'b0 ;
  assign n21562 = n3956 & n15708 ;
  assign n21563 = ~n3705 & n8944 ;
  assign n21564 = n14375 & n16463 ;
  assign n21565 = ~n3113 & n20317 ;
  assign n21566 = n20926 ^ n6908 ^ 1'b0 ;
  assign n21567 = n3492 & ~n9827 ;
  assign n21568 = n12060 ^ n3276 ^ 1'b0 ;
  assign n21569 = ~n10704 & n21568 ;
  assign n21570 = ~n11942 & n19007 ;
  assign n21571 = ( n10551 & n14496 ) | ( n10551 & ~n21570 ) | ( n14496 & ~n21570 ) ;
  assign n21572 = n18337 ^ n6866 ^ 1'b0 ;
  assign n21573 = n21571 & n21572 ;
  assign n21574 = n5659 | n12437 ;
  assign n21575 = n19679 & n21574 ;
  assign n21576 = n7804 ^ n6026 ^ 1'b0 ;
  assign n21577 = n910 & n21576 ;
  assign n21578 = ( ~x19 & n4902 ) | ( ~x19 & n21577 ) | ( n4902 & n21577 ) ;
  assign n21579 = n2457 & n3139 ;
  assign n21580 = n3961 & n21579 ;
  assign n21581 = n21578 & n21580 ;
  assign n21582 = ( n3084 & n13826 ) | ( n3084 & n19860 ) | ( n13826 & n19860 ) ;
  assign n21583 = ~n4430 & n21582 ;
  assign n21584 = n20891 ^ n2861 ^ 1'b0 ;
  assign n21585 = n14933 ^ n10435 ^ n6145 ;
  assign n21586 = n21115 & ~n21585 ;
  assign n21587 = n7589 & n10738 ;
  assign n21588 = n21587 ^ n805 ^ 1'b0 ;
  assign n21589 = n2758 & n8497 ;
  assign n21590 = n14816 ^ n959 ^ 1'b0 ;
  assign n21591 = n13190 & n21590 ;
  assign n21592 = n2059 & n21591 ;
  assign n21602 = n5524 & n10935 ;
  assign n21597 = n7582 & n11903 ;
  assign n21598 = n2083 & n21597 ;
  assign n21595 = n6597 ^ n6430 ^ n671 ;
  assign n21593 = n9737 ^ n2721 ^ n1290 ;
  assign n21594 = n2981 & n21593 ;
  assign n21596 = n21595 ^ n21594 ^ 1'b0 ;
  assign n21599 = n21598 ^ n21596 ^ n644 ;
  assign n21600 = ~n10769 & n14639 ;
  assign n21601 = n21599 & n21600 ;
  assign n21603 = n21602 ^ n21601 ^ n3945 ;
  assign n21604 = n15299 | n17138 ;
  assign n21605 = n823 & ~n21604 ;
  assign n21606 = ( n6024 & ~n9183 ) | ( n6024 & n11714 ) | ( ~n9183 & n11714 ) ;
  assign n21607 = ~n7669 & n21606 ;
  assign n21608 = n8007 | n13031 ;
  assign n21609 = n21608 ^ n449 ^ 1'b0 ;
  assign n21610 = ~n6898 & n21609 ;
  assign n21611 = ~n4317 & n18245 ;
  assign n21612 = n14664 ^ n7772 ^ 1'b0 ;
  assign n21613 = n14138 ^ n9593 ^ 1'b0 ;
  assign n21614 = n17429 | n21613 ;
  assign n21615 = n21614 ^ n6530 ^ 1'b0 ;
  assign n21616 = n20624 | n21615 ;
  assign n21617 = n5933 ^ n5030 ^ 1'b0 ;
  assign n21618 = n12707 ^ n519 ^ 1'b0 ;
  assign n21619 = ~n2842 & n6362 ;
  assign n21620 = n21619 ^ n6802 ^ 1'b0 ;
  assign n21621 = ( n7385 & n14253 ) | ( n7385 & ~n21620 ) | ( n14253 & ~n21620 ) ;
  assign n21622 = n10658 ^ n4382 ^ 1'b0 ;
  assign n21623 = n4343 & ~n9900 ;
  assign n21624 = n3599 ^ n790 ^ 1'b0 ;
  assign n21625 = n886 & ~n21624 ;
  assign n21626 = ( n1082 & n9294 ) | ( n1082 & n16256 ) | ( n9294 & n16256 ) ;
  assign n21627 = n16848 ^ n8110 ^ n4655 ;
  assign n21628 = ( n9513 & n12205 ) | ( n9513 & ~n12207 ) | ( n12205 & ~n12207 ) ;
  assign n21629 = n12536 ^ n4171 ^ 1'b0 ;
  assign n21630 = n21628 & ~n21629 ;
  assign n21631 = n14193 ^ n166 ^ 1'b0 ;
  assign n21632 = n6916 & ~n21631 ;
  assign n21633 = x10 & ~n19254 ;
  assign n21634 = n15767 & n21633 ;
  assign n21635 = n11600 & ~n21634 ;
  assign n21636 = n20432 ^ n7865 ^ 1'b0 ;
  assign n21637 = n12964 | n21636 ;
  assign n21641 = ~n6114 & n13591 ;
  assign n21642 = n21641 ^ n865 ^ 1'b0 ;
  assign n21638 = n14156 ^ n11459 ^ 1'b0 ;
  assign n21639 = ~n12744 & n21638 ;
  assign n21640 = n21639 ^ n7883 ^ 1'b0 ;
  assign n21643 = n21642 ^ n21640 ^ n13899 ;
  assign n21644 = n21643 ^ n5925 ^ n1970 ;
  assign n21645 = n8143 & n19177 ;
  assign n21646 = ~n8143 & n21645 ;
  assign n21647 = ~n12015 & n13412 ;
  assign n21648 = n6346 ^ n5225 ^ 1'b0 ;
  assign n21649 = ~n14727 & n14970 ;
  assign n21650 = n10847 | n18127 ;
  assign n21651 = n21650 ^ n21588 ^ 1'b0 ;
  assign n21652 = ~n2304 & n21651 ;
  assign n21653 = n4632 | n7556 ;
  assign n21654 = n21653 ^ n17646 ^ 1'b0 ;
  assign n21655 = n13955 ^ n12171 ^ n8372 ;
  assign n21656 = n21655 ^ n3226 ^ 1'b0 ;
  assign n21657 = ~n20943 & n21656 ;
  assign n21658 = ~n3379 & n21657 ;
  assign n21659 = n15638 ^ n9977 ^ n6420 ;
  assign n21660 = n8152 & n21659 ;
  assign n21661 = n19850 ^ n15638 ^ 1'b0 ;
  assign n21662 = ( n4955 & n12847 ) | ( n4955 & n21661 ) | ( n12847 & n21661 ) ;
  assign n21663 = n21662 ^ n11505 ^ n664 ;
  assign n21664 = ~n3230 & n10858 ;
  assign n21665 = n18825 ^ n10647 ^ 1'b0 ;
  assign n21666 = n2558 & n5872 ;
  assign n21667 = n21665 & n21666 ;
  assign n21668 = ( n1034 & ~n9763 ) | ( n1034 & n21667 ) | ( ~n9763 & n21667 ) ;
  assign n21669 = n560 & ~n21668 ;
  assign n21670 = ~n1966 & n21669 ;
  assign n21671 = ( n3660 & n21664 ) | ( n3660 & ~n21670 ) | ( n21664 & ~n21670 ) ;
  assign n21672 = n10626 & n18124 ;
  assign n21673 = n14371 ^ n1560 ^ n879 ;
  assign n21674 = n21673 ^ n21275 ^ 1'b0 ;
  assign n21675 = n18898 & n21674 ;
  assign n21676 = ~n10199 & n21675 ;
  assign n21677 = n16721 ^ n7321 ^ 1'b0 ;
  assign n21678 = n20409 & ~n21677 ;
  assign n21679 = x35 | n16674 ;
  assign n21680 = n21679 ^ n1072 ^ 1'b0 ;
  assign n21681 = n5567 | n21680 ;
  assign n21682 = n21681 ^ n18046 ^ 1'b0 ;
  assign n21683 = n12207 ^ n463 ^ 1'b0 ;
  assign n21684 = n13926 & n21683 ;
  assign n21685 = ~n8317 & n16088 ;
  assign n21686 = ~n1652 & n18245 ;
  assign n21687 = ~n6387 & n17929 ;
  assign n21688 = ~n5901 & n7619 ;
  assign n21689 = n21688 ^ n14983 ^ 1'b0 ;
  assign n21690 = n2495 & n21689 ;
  assign n21692 = n10656 ^ n4342 ^ 1'b0 ;
  assign n21693 = n18628 | n21692 ;
  assign n21691 = n5606 & ~n21297 ;
  assign n21694 = n21693 ^ n21691 ^ 1'b0 ;
  assign n21695 = n21694 ^ n9514 ^ 1'b0 ;
  assign n21696 = n282 & ~n7949 ;
  assign n21697 = ~n19216 & n21696 ;
  assign n21698 = n21697 ^ n12192 ^ 1'b0 ;
  assign n21699 = n1724 | n21698 ;
  assign n21700 = n18269 ^ n8619 ^ n3349 ;
  assign n21701 = ~n1486 & n18339 ;
  assign n21702 = n21701 ^ n6512 ^ 1'b0 ;
  assign n21703 = n8608 | n12524 ;
  assign n21704 = n21702 | n21703 ;
  assign n21705 = ~n3882 & n21704 ;
  assign n21706 = ~n19419 & n21705 ;
  assign n21707 = n21706 ^ n9971 ^ 1'b0 ;
  assign n21708 = n15218 | n21707 ;
  assign n21709 = n13002 ^ n7340 ^ 1'b0 ;
  assign n21710 = n12261 | n21709 ;
  assign n21711 = n2026 & ~n5790 ;
  assign n21712 = n21711 ^ n250 ^ 1'b0 ;
  assign n21713 = n1501 & ~n1954 ;
  assign n21714 = n425 & n14412 ;
  assign n21715 = n21714 ^ n5901 ^ 1'b0 ;
  assign n21716 = n14889 | n17533 ;
  assign n21717 = n2487 ^ n875 ^ 1'b0 ;
  assign n21718 = n2829 | n21717 ;
  assign n21719 = n13602 ^ n2060 ^ 1'b0 ;
  assign n21720 = ( n5557 & n9935 ) | ( n5557 & ~n16329 ) | ( n9935 & ~n16329 ) ;
  assign n21721 = n12238 ^ n2926 ^ 1'b0 ;
  assign n21722 = n2489 & ~n16052 ;
  assign n21723 = ~n21721 & n21722 ;
  assign n21724 = n11809 & ~n21668 ;
  assign n21725 = n8776 | n8936 ;
  assign n21726 = n21725 ^ n7103 ^ 1'b0 ;
  assign n21727 = ~n700 & n18380 ;
  assign n21728 = n10186 & ~n21727 ;
  assign n21730 = n7162 & n10334 ;
  assign n21729 = n6430 | n16901 ;
  assign n21731 = n21730 ^ n21729 ^ 1'b0 ;
  assign n21732 = ( n9283 & n14375 ) | ( n9283 & n16170 ) | ( n14375 & n16170 ) ;
  assign n21734 = ~n5479 & n19208 ;
  assign n21735 = n21734 ^ n17612 ^ 1'b0 ;
  assign n21736 = n8432 & n21735 ;
  assign n21733 = n16362 & n20199 ;
  assign n21737 = n21736 ^ n21733 ^ n3918 ;
  assign n21738 = ~n10673 & n11813 ;
  assign n21739 = ~n3919 & n21738 ;
  assign n21740 = n5399 ^ n1172 ^ 1'b0 ;
  assign n21741 = ~n1692 & n21740 ;
  assign n21742 = n21741 ^ n3442 ^ 1'b0 ;
  assign n21743 = n21739 | n21742 ;
  assign n21744 = ( n13674 & n14040 ) | ( n13674 & ~n21743 ) | ( n14040 & ~n21743 ) ;
  assign n21749 = n2194 | n5695 ;
  assign n21745 = ~n3366 & n17365 ;
  assign n21746 = n4057 ^ n1892 ^ 1'b0 ;
  assign n21747 = ~n21745 & n21746 ;
  assign n21748 = ~n12309 & n21747 ;
  assign n21750 = n21749 ^ n21748 ^ 1'b0 ;
  assign n21751 = n8355 | n21750 ;
  assign n21752 = n4565 & n15687 ;
  assign n21753 = ~n4689 & n21752 ;
  assign n21754 = n11292 ^ n2007 ^ 1'b0 ;
  assign n21755 = n7575 | n21754 ;
  assign n21756 = n8090 | n21755 ;
  assign n21757 = n3881 & ~n4307 ;
  assign n21758 = n21756 & n21757 ;
  assign n21759 = n1226 | n10668 ;
  assign n21760 = n21759 ^ n5389 ^ 1'b0 ;
  assign n21761 = n12470 ^ n12061 ^ 1'b0 ;
  assign n21762 = x18 & ~n21761 ;
  assign n21763 = n1913 | n21762 ;
  assign n21764 = n946 & ~n10785 ;
  assign n21765 = n18648 & n21764 ;
  assign n21766 = n21765 ^ n8842 ^ 1'b0 ;
  assign n21767 = n7639 ^ n760 ^ 1'b0 ;
  assign n21768 = ~n12175 & n21767 ;
  assign n21769 = ~n9305 & n16514 ;
  assign n21770 = n20549 & n21769 ;
  assign n21771 = n14845 ^ n6303 ^ 1'b0 ;
  assign n21772 = ~n13465 & n17453 ;
  assign n21773 = n3627 ^ n1529 ^ 1'b0 ;
  assign n21774 = n176 & n21773 ;
  assign n21775 = x85 & ~n1072 ;
  assign n21776 = n21775 ^ n723 ^ 1'b0 ;
  assign n21777 = n6306 ^ n4157 ^ 1'b0 ;
  assign n21778 = ~n20982 & n21777 ;
  assign n21779 = n10809 & n21778 ;
  assign n21780 = n21779 ^ n7834 ^ 1'b0 ;
  assign n21781 = ~n21776 & n21780 ;
  assign n21782 = ( n2814 & n4723 ) | ( n2814 & ~n16265 ) | ( n4723 & ~n16265 ) ;
  assign n21783 = n1040 & n1981 ;
  assign n21784 = ~n3091 & n21783 ;
  assign n21785 = ( n4449 & n11003 ) | ( n4449 & n21784 ) | ( n11003 & n21784 ) ;
  assign n21786 = ~n5585 & n12218 ;
  assign n21788 = n2198 & ~n10905 ;
  assign n21787 = ~n1808 & n15408 ;
  assign n21789 = n21788 ^ n21787 ^ 1'b0 ;
  assign n21790 = n5499 ^ n3666 ^ 1'b0 ;
  assign n21791 = n21790 ^ n11676 ^ n10576 ;
  assign n21792 = n3147 ^ n1059 ^ 1'b0 ;
  assign n21793 = n314 & ~n15610 ;
  assign n21794 = ( n6569 & n7521 ) | ( n6569 & n16207 ) | ( n7521 & n16207 ) ;
  assign n21795 = n10046 | n21794 ;
  assign n21796 = n3765 & ~n21795 ;
  assign n21797 = n477 & n1302 ;
  assign n21798 = n21797 ^ n9698 ^ n7816 ;
  assign n21799 = n21798 ^ n16499 ^ n7484 ;
  assign n21800 = n21799 ^ n9682 ^ 1'b0 ;
  assign n21801 = n283 & n21800 ;
  assign n21802 = ~n6329 & n6979 ;
  assign n21803 = n18857 ^ n13928 ^ 1'b0 ;
  assign n21804 = n4038 & n21803 ;
  assign n21805 = n8610 ^ n303 ^ 1'b0 ;
  assign n21807 = n2964 | n5365 ;
  assign n21808 = n19463 | n21807 ;
  assign n21806 = n4442 ^ n3171 ^ n1730 ;
  assign n21809 = n21808 ^ n21806 ^ n18838 ;
  assign n21810 = n15298 ^ n14935 ^ 1'b0 ;
  assign n21811 = ~n2594 & n21810 ;
  assign n21812 = n19948 ^ n9710 ^ 1'b0 ;
  assign n21813 = ~n4757 & n21812 ;
  assign n21814 = n18802 & n21813 ;
  assign n21815 = n17607 ^ n4996 ^ 1'b0 ;
  assign n21824 = n4050 & ~n17868 ;
  assign n21816 = ( n623 & n1950 ) | ( n623 & ~n5189 ) | ( n1950 & ~n5189 ) ;
  assign n21817 = n7888 & ~n21816 ;
  assign n21818 = n21817 ^ n8984 ^ 1'b0 ;
  assign n21819 = n4082 & ~n18769 ;
  assign n21820 = n21819 ^ n4737 ^ 1'b0 ;
  assign n21821 = n21818 & n21820 ;
  assign n21822 = n21821 ^ n20954 ^ 1'b0 ;
  assign n21823 = n5598 & ~n21822 ;
  assign n21825 = n21824 ^ n21823 ^ 1'b0 ;
  assign n21826 = n14704 ^ n4178 ^ n2855 ;
  assign n21827 = n21826 ^ n1494 ^ 1'b0 ;
  assign n21828 = n21825 & n21827 ;
  assign n21829 = ( n13192 & n21815 ) | ( n13192 & ~n21828 ) | ( n21815 & ~n21828 ) ;
  assign n21831 = ~n1374 & n8889 ;
  assign n21832 = n371 | n21831 ;
  assign n21830 = n10394 ^ n1972 ^ 1'b0 ;
  assign n21833 = n21832 ^ n21830 ^ n7679 ;
  assign n21834 = n13531 ^ n10277 ^ 1'b0 ;
  assign n21835 = n4761 & ~n9781 ;
  assign n21836 = n21835 ^ n21249 ^ 1'b0 ;
  assign n21837 = n1215 | n15719 ;
  assign n21838 = n13815 & ~n21837 ;
  assign n21839 = n21838 ^ n5890 ^ 1'b0 ;
  assign n21840 = n18953 & n21839 ;
  assign n21842 = n1479 | n1987 ;
  assign n21843 = n21842 ^ n3875 ^ 1'b0 ;
  assign n21844 = ~n1874 & n21843 ;
  assign n21841 = ~n3820 & n5573 ;
  assign n21845 = n21844 ^ n21841 ^ 1'b0 ;
  assign n21846 = n21719 ^ n1268 ^ n665 ;
  assign n21847 = ~n338 & n8938 ;
  assign n21848 = n824 & ~n16693 ;
  assign n21849 = n14641 & ~n21848 ;
  assign n21851 = n12758 ^ n6438 ^ 1'b0 ;
  assign n21852 = n2108 & ~n21851 ;
  assign n21850 = ~n3740 & n10320 ;
  assign n21853 = n21852 ^ n21850 ^ n7491 ;
  assign n21854 = n21849 & ~n21853 ;
  assign n21855 = n2770 & n18980 ;
  assign n21856 = n6010 ^ n5947 ^ 1'b0 ;
  assign n21857 = n7287 | n21856 ;
  assign n21858 = n21857 ^ n12971 ^ n264 ;
  assign n21859 = n14793 ^ n10654 ^ 1'b0 ;
  assign n21860 = ( n11420 & n21661 ) | ( n11420 & n21859 ) | ( n21661 & n21859 ) ;
  assign n21861 = n422 & ~n4150 ;
  assign n21863 = n1682 & n6201 ;
  assign n21864 = n254 & n21863 ;
  assign n21862 = n134 & n1162 ;
  assign n21865 = n21864 ^ n21862 ^ 1'b0 ;
  assign n21866 = n490 & ~n3869 ;
  assign n21867 = ~n6149 & n21866 ;
  assign n21868 = n12291 & ~n21867 ;
  assign n21869 = n6102 ^ n530 ^ 1'b0 ;
  assign n21870 = n1099 | n21869 ;
  assign n21871 = ( ~n2275 & n16120 ) | ( ~n2275 & n21870 ) | ( n16120 & n21870 ) ;
  assign n21872 = n21871 ^ n20384 ^ 1'b0 ;
  assign n21873 = n13565 & ~n21872 ;
  assign n21874 = n2929 | n21873 ;
  assign n21876 = n4436 ^ n2790 ^ 1'b0 ;
  assign n21875 = ( n2343 & n2550 ) | ( n2343 & ~n6218 ) | ( n2550 & ~n6218 ) ;
  assign n21877 = n21876 ^ n21875 ^ n19751 ;
  assign n21878 = n651 & n6918 ;
  assign n21879 = n4948 & ~n10835 ;
  assign n21880 = n21878 & n21879 ;
  assign n21881 = n1154 ^ n297 ^ 1'b0 ;
  assign n21882 = n21375 ^ n14618 ^ 1'b0 ;
  assign n21883 = n8552 & n21882 ;
  assign n21885 = n13064 ^ n8086 ^ 1'b0 ;
  assign n21884 = n3725 | n6295 ;
  assign n21886 = n21885 ^ n21884 ^ n9771 ;
  assign n21887 = ~n6441 & n21886 ;
  assign n21888 = ~n13814 & n21887 ;
  assign n21889 = n12348 & ~n13457 ;
  assign n21890 = n8130 | n8914 ;
  assign n21891 = n21890 ^ n4174 ^ 1'b0 ;
  assign n21892 = n20450 & n21891 ;
  assign n21893 = n21892 ^ n7098 ^ n1487 ;
  assign n21894 = n12142 ^ n8515 ^ 1'b0 ;
  assign n21895 = n21314 ^ n10126 ^ 1'b0 ;
  assign n21896 = n14604 & n21895 ;
  assign n21897 = n21896 ^ n4369 ^ 1'b0 ;
  assign n21898 = n282 ^ x51 ^ 1'b0 ;
  assign n21899 = n12693 & ~n21898 ;
  assign n21900 = n21899 ^ n15654 ^ n8144 ;
  assign n21901 = n21900 ^ n21696 ^ n19877 ;
  assign n21902 = ( n11466 & ~n19649 ) | ( n11466 & n21901 ) | ( ~n19649 & n21901 ) ;
  assign n21903 = ~n4124 & n17079 ;
  assign n21904 = n21903 ^ n17640 ^ 1'b0 ;
  assign n21905 = n16515 & n21904 ;
  assign n21906 = n8353 & n21905 ;
  assign n21909 = n2668 & n3903 ;
  assign n21907 = n2167 | n14185 ;
  assign n21908 = n21907 ^ n2214 ^ 1'b0 ;
  assign n21910 = n21909 ^ n21908 ^ 1'b0 ;
  assign n21911 = n1095 & ~n11467 ;
  assign n21912 = ~n16329 & n21911 ;
  assign n21913 = n21910 & n21912 ;
  assign n21914 = n18894 & ~n21650 ;
  assign n21915 = n21914 ^ n10414 ^ 1'b0 ;
  assign n21916 = n3055 ^ n1837 ^ 1'b0 ;
  assign n21917 = n16650 ^ n9064 ^ 1'b0 ;
  assign n21918 = ~n21916 & n21917 ;
  assign n21919 = ( n499 & n5128 ) | ( n499 & ~n9635 ) | ( n5128 & ~n9635 ) ;
  assign n21920 = n9357 | n14900 ;
  assign n21921 = n9199 | n21920 ;
  assign n21922 = n21919 | n21921 ;
  assign n21923 = n16064 ^ n4261 ^ 1'b0 ;
  assign n21924 = n227 | n3067 ;
  assign n21925 = n227 & ~n21924 ;
  assign n21926 = n385 & n857 ;
  assign n21927 = n3470 & n21926 ;
  assign n21928 = ( n4605 & n21925 ) | ( n4605 & ~n21927 ) | ( n21925 & ~n21927 ) ;
  assign n21929 = n21928 ^ n14637 ^ n842 ;
  assign n21930 = n9830 & n17980 ;
  assign n21931 = n21930 ^ n21640 ^ 1'b0 ;
  assign n21932 = n5059 & ~n6609 ;
  assign n21933 = n3703 ^ n1117 ^ 1'b0 ;
  assign n21934 = n21932 | n21933 ;
  assign n21935 = n8345 & ~n21934 ;
  assign n21936 = n21935 ^ n4921 ^ 1'b0 ;
  assign n21937 = n19603 ^ n691 ^ 1'b0 ;
  assign n21938 = n4151 ^ n1627 ^ 1'b0 ;
  assign n21939 = n5285 & ~n21938 ;
  assign n21940 = n2214 & n21939 ;
  assign n21941 = n2429 & n3489 ;
  assign n21942 = n190 & n21941 ;
  assign n21943 = n770 & n3658 ;
  assign n21944 = n21943 ^ n1209 ^ 1'b0 ;
  assign n21945 = ~n21942 & n21944 ;
  assign n21946 = ( ~n5009 & n5885 ) | ( ~n5009 & n18142 ) | ( n5885 & n18142 ) ;
  assign n21947 = n510 & ~n4342 ;
  assign n21948 = n21946 & n21947 ;
  assign n21949 = ~n804 & n21948 ;
  assign n21950 = n1149 & n17768 ;
  assign n21951 = n9187 & ~n21950 ;
  assign n21952 = n21951 ^ n9366 ^ 1'b0 ;
  assign n21953 = n9424 & ~n11632 ;
  assign n21954 = n2441 & n18111 ;
  assign n21955 = n21954 ^ n15966 ^ 1'b0 ;
  assign n21956 = ~n16224 & n21955 ;
  assign n21957 = ~n5223 & n21956 ;
  assign n21958 = ~n1397 & n6815 ;
  assign n21959 = n6438 & ~n6461 ;
  assign n21960 = n21959 ^ n14542 ^ 1'b0 ;
  assign n21961 = ~n21958 & n21960 ;
  assign n21962 = n1955 | n5930 ;
  assign n21963 = n21962 ^ n7243 ^ 1'b0 ;
  assign n21964 = n12014 & ~n21963 ;
  assign n21965 = n21964 ^ n9870 ^ 1'b0 ;
  assign n21966 = n3301 ^ n1038 ^ 1'b0 ;
  assign n21967 = ~n8437 & n14908 ;
  assign n21968 = n1462 & n21967 ;
  assign n21969 = n21968 ^ n9567 ^ 1'b0 ;
  assign n21970 = n17789 & n21969 ;
  assign n21971 = n21970 ^ n16119 ^ 1'b0 ;
  assign n21972 = ( ~n1481 & n7033 ) | ( ~n1481 & n16063 ) | ( n7033 & n16063 ) ;
  assign n21973 = n9540 & n18254 ;
  assign n21974 = ~n4289 & n21973 ;
  assign n21975 = n3474 & n20040 ;
  assign n21976 = ~n3474 & n21975 ;
  assign n21977 = n320 | n21976 ;
  assign n21978 = n320 & ~n21977 ;
  assign n21979 = n21978 ^ n5551 ^ 1'b0 ;
  assign n21980 = n2431 & ~n21979 ;
  assign n21981 = n8641 & ~n21670 ;
  assign n21982 = n17686 ^ n3983 ^ 1'b0 ;
  assign n21983 = ~n12109 & n21982 ;
  assign n21984 = n11320 ^ n7639 ^ n6092 ;
  assign n21985 = n21984 ^ n15887 ^ 1'b0 ;
  assign n21986 = n21983 & n21985 ;
  assign n21987 = ~n10656 & n17975 ;
  assign n21988 = ( ~n1703 & n3396 ) | ( ~n1703 & n21987 ) | ( n3396 & n21987 ) ;
  assign n21989 = n18427 ^ n10649 ^ 1'b0 ;
  assign n21991 = n5063 ^ n2073 ^ 1'b0 ;
  assign n21992 = ~n10435 & n21991 ;
  assign n21993 = n21992 ^ n8768 ^ n5331 ;
  assign n21990 = n19571 ^ n2721 ^ 1'b0 ;
  assign n21994 = n21993 ^ n21990 ^ n11979 ;
  assign n21995 = n19169 | n21994 ;
  assign n21996 = n1948 & ~n13269 ;
  assign n21997 = n18353 ^ n14745 ^ n5942 ;
  assign n21998 = ( n1853 & n14181 ) | ( n1853 & ~n16185 ) | ( n14181 & ~n16185 ) ;
  assign n21999 = n13912 ^ n12520 ^ 1'b0 ;
  assign n22000 = x48 | n21999 ;
  assign n22001 = n8036 ^ n3380 ^ 1'b0 ;
  assign n22005 = n5289 ^ n3518 ^ n1067 ;
  assign n22006 = n4768 ^ n3562 ^ 1'b0 ;
  assign n22007 = ~n22005 & n22006 ;
  assign n22002 = ~n725 & n3349 ;
  assign n22003 = n9545 & n22002 ;
  assign n22004 = n15732 & ~n22003 ;
  assign n22008 = n22007 ^ n22004 ^ 1'b0 ;
  assign n22009 = n8437 ^ x78 ^ 1'b0 ;
  assign n22010 = n2119 & ~n16372 ;
  assign n22011 = n2355 ^ n908 ^ 1'b0 ;
  assign n22012 = ~n2285 & n22011 ;
  assign n22013 = n22012 ^ n4107 ^ 1'b0 ;
  assign n22014 = n2500 & ~n21007 ;
  assign n22015 = n4343 & n22014 ;
  assign n22016 = n819 ^ n510 ^ 1'b0 ;
  assign n22017 = n20168 & n22016 ;
  assign n22018 = n10348 & n21022 ;
  assign n22020 = ~n984 & n7609 ;
  assign n22021 = n22020 ^ n20224 ^ 1'b0 ;
  assign n22019 = n16063 ^ n8819 ^ n5785 ;
  assign n22022 = n22021 ^ n22019 ^ 1'b0 ;
  assign n22023 = n22018 & n22022 ;
  assign n22024 = ~n9884 & n20643 ;
  assign n22025 = ~n2642 & n9162 ;
  assign n22026 = n21679 & n22025 ;
  assign n22027 = n1915 & n9953 ;
  assign n22028 = n22027 ^ n4492 ^ n1196 ;
  assign n22029 = n6133 ^ n1281 ^ 1'b0 ;
  assign n22030 = ~n22028 & n22029 ;
  assign n22031 = n6867 & n14806 ;
  assign n22032 = n21449 ^ n3229 ^ 1'b0 ;
  assign n22033 = n1161 & n22032 ;
  assign n22034 = n16776 ^ n6523 ^ n2640 ;
  assign n22035 = ~n1777 & n4937 ;
  assign n22036 = n4534 ^ n2663 ^ n174 ;
  assign n22037 = n17454 & n22036 ;
  assign n22038 = n22037 ^ n16775 ^ 1'b0 ;
  assign n22039 = ~n22035 & n22038 ;
  assign n22040 = n5382 ^ n2550 ^ 1'b0 ;
  assign n22041 = n10353 | n22040 ;
  assign n22042 = n3980 | n4219 ;
  assign n22043 = n18858 | n22042 ;
  assign n22044 = n18858 ^ n14132 ^ 1'b0 ;
  assign n22045 = n22043 & ~n22044 ;
  assign n22046 = ~n6888 & n22045 ;
  assign n22047 = n3979 & ~n15042 ;
  assign n22048 = n13481 | n22047 ;
  assign n22049 = n14712 ^ x95 ^ 1'b0 ;
  assign n22050 = ~n2930 & n22049 ;
  assign n22051 = ( ~n4445 & n5046 ) | ( ~n4445 & n12660 ) | ( n5046 & n12660 ) ;
  assign n22052 = n22051 ^ n9982 ^ 1'b0 ;
  assign n22053 = ~n706 & n22052 ;
  assign n22054 = n1711 ^ n651 ^ 1'b0 ;
  assign n22055 = n17958 & ~n22054 ;
  assign n22056 = n22055 ^ n14975 ^ 1'b0 ;
  assign n22057 = n2861 & ~n4037 ;
  assign n22058 = n9939 & n22057 ;
  assign n22059 = n4034 & ~n16769 ;
  assign n22060 = n22059 ^ n9354 ^ 1'b0 ;
  assign n22061 = n10645 ^ n2085 ^ 1'b0 ;
  assign n22062 = ( n2583 & ~n21361 ) | ( n2583 & n22061 ) | ( ~n21361 & n22061 ) ;
  assign n22063 = n6482 ^ n4270 ^ 1'b0 ;
  assign n22064 = ( n13462 & n18719 ) | ( n13462 & ~n22063 ) | ( n18719 & ~n22063 ) ;
  assign n22065 = n9960 | n12943 ;
  assign n22066 = x104 & n2429 ;
  assign n22067 = n13527 ^ n1683 ^ 1'b0 ;
  assign n22068 = ~n19552 & n22067 ;
  assign n22069 = ~n22066 & n22068 ;
  assign n22070 = n8387 & n13200 ;
  assign n22071 = n22070 ^ n405 ^ 1'b0 ;
  assign n22072 = n2160 & ~n22071 ;
  assign n22073 = ~n4292 & n22072 ;
  assign n22074 = n4497 & ~n7594 ;
  assign n22075 = n22074 ^ n15622 ^ 1'b0 ;
  assign n22076 = n17413 ^ n9468 ^ 1'b0 ;
  assign n22077 = n13747 ^ n13133 ^ 1'b0 ;
  assign n22078 = n17446 ^ n7513 ^ n5137 ;
  assign n22079 = n14226 ^ n8860 ^ n4351 ;
  assign n22080 = ~n10686 & n15622 ;
  assign n22081 = n22079 | n22080 ;
  assign n22082 = n22081 ^ n18771 ^ 1'b0 ;
  assign n22083 = n7418 ^ n4095 ^ 1'b0 ;
  assign n22084 = n9273 & n22083 ;
  assign n22085 = ~n5235 & n22084 ;
  assign n22086 = n7383 & n14265 ;
  assign n22087 = ~n7023 & n22086 ;
  assign n22088 = n4739 | n22087 ;
  assign n22089 = n4916 & ~n22088 ;
  assign n22090 = ( n14042 & n17181 ) | ( n14042 & ~n21962 ) | ( n17181 & ~n21962 ) ;
  assign n22091 = n1319 ^ n612 ^ 1'b0 ;
  assign n22092 = n739 & ~n22091 ;
  assign n22093 = ( n16430 & n17570 ) | ( n16430 & ~n22092 ) | ( n17570 & ~n22092 ) ;
  assign n22094 = ( ~n11006 & n16734 ) | ( ~n11006 & n20466 ) | ( n16734 & n20466 ) ;
  assign n22095 = ~n10924 & n14194 ;
  assign n22096 = n22095 ^ n2369 ^ 1'b0 ;
  assign n22097 = n18549 & n22096 ;
  assign n22098 = n19264 & n22097 ;
  assign n22099 = n10081 ^ n9086 ^ 1'b0 ;
  assign n22100 = n16955 & ~n22099 ;
  assign n22101 = n19338 ^ n4522 ^ 1'b0 ;
  assign n22102 = n22100 | n22101 ;
  assign n22103 = n3781 ^ n642 ^ 1'b0 ;
  assign n22104 = n7578 & n22103 ;
  assign n22105 = n13504 ^ n2526 ^ 1'b0 ;
  assign n22106 = ( n3376 & ~n4610 ) | ( n3376 & n16185 ) | ( ~n4610 & n16185 ) ;
  assign n22107 = n12233 ^ n1481 ^ 1'b0 ;
  assign n22108 = n1175 & ~n17651 ;
  assign n22109 = n22108 ^ n19349 ^ 1'b0 ;
  assign n22110 = n9211 | n15588 ;
  assign n22111 = n1740 & n6916 ;
  assign n22112 = ~n16658 & n22111 ;
  assign n22113 = ( n8669 & n16420 ) | ( n8669 & n22112 ) | ( n16420 & n22112 ) ;
  assign n22114 = n19019 ^ n4320 ^ 1'b0 ;
  assign n22115 = ~n22113 & n22114 ;
  assign n22116 = n1713 | n3016 ;
  assign n22117 = n22116 ^ n2927 ^ 1'b0 ;
  assign n22118 = ( n17882 & n19271 ) | ( n17882 & n22117 ) | ( n19271 & n22117 ) ;
  assign n22119 = n13538 ^ n12823 ^ 1'b0 ;
  assign n22120 = ( n5585 & n6148 ) | ( n5585 & ~n7256 ) | ( n6148 & ~n7256 ) ;
  assign n22121 = ~n10426 & n13291 ;
  assign n22122 = n22121 ^ n2149 ^ 1'b0 ;
  assign n22123 = ~n13592 & n15900 ;
  assign n22124 = n15947 ^ n2929 ^ 1'b0 ;
  assign n22125 = n3585 ^ n1202 ^ 1'b0 ;
  assign n22126 = n22125 ^ n2623 ^ 1'b0 ;
  assign n22127 = n2091 & ~n3494 ;
  assign n22128 = n22127 ^ n9925 ^ n6530 ;
  assign n22129 = ~n2414 & n11364 ;
  assign n22130 = n22129 ^ n13111 ^ 1'b0 ;
  assign n22131 = n7931 ^ n5440 ^ 1'b0 ;
  assign n22132 = n1029 & n22131 ;
  assign n22133 = ~n7081 & n15843 ;
  assign n22134 = n22133 ^ n21984 ^ 1'b0 ;
  assign n22135 = ( n4984 & ~n22132 ) | ( n4984 & n22134 ) | ( ~n22132 & n22134 ) ;
  assign n22136 = ~n905 & n22135 ;
  assign n22137 = ~n1920 & n2632 ;
  assign n22138 = n22137 ^ n4749 ^ 1'b0 ;
  assign n22139 = n5282 & ~n20127 ;
  assign n22140 = ~n4565 & n22139 ;
  assign n22141 = n1319 & n22140 ;
  assign n22142 = ~n317 & n9796 ;
  assign n22143 = n22142 ^ n6164 ^ 1'b0 ;
  assign n22144 = n22143 ^ n10630 ^ 1'b0 ;
  assign n22145 = n20377 ^ n11601 ^ n6703 ;
  assign n22146 = ~n4594 & n7467 ;
  assign n22147 = n2014 & n22146 ;
  assign n22148 = n7416 & n22147 ;
  assign n22149 = n16909 & ~n17655 ;
  assign n22150 = n22149 ^ n14993 ^ 1'b0 ;
  assign n22151 = n3340 | n4883 ;
  assign n22152 = n17307 & ~n22151 ;
  assign n22153 = ~n193 & n7129 ;
  assign n22154 = n7227 & n21968 ;
  assign n22155 = ~n9138 & n22154 ;
  assign n22156 = n22155 ^ n10366 ^ 1'b0 ;
  assign n22157 = n22156 ^ n11883 ^ n6169 ;
  assign n22158 = n2151 & ~n18163 ;
  assign n22159 = n2997 | n4993 ;
  assign n22160 = n13749 | n22159 ;
  assign n22161 = ~n7792 & n17637 ;
  assign n22162 = n22161 ^ n7022 ^ 1'b0 ;
  assign n22163 = n22162 ^ n12399 ^ 1'b0 ;
  assign n22164 = n4085 ^ n2026 ^ 1'b0 ;
  assign n22165 = n12166 ^ n6002 ^ n5815 ;
  assign n22166 = n22164 | n22165 ;
  assign n22167 = n8865 ^ n6872 ^ n2292 ;
  assign n22168 = n5137 & ~n22167 ;
  assign n22169 = n22168 ^ n7744 ^ 1'b0 ;
  assign n22170 = n371 & n7491 ;
  assign n22171 = n19569 & n22170 ;
  assign n22172 = n22171 ^ n12906 ^ 1'b0 ;
  assign n22173 = n6539 ^ n2038 ^ 1'b0 ;
  assign n22174 = ( n348 & n4670 ) | ( n348 & ~n14415 ) | ( n4670 & ~n14415 ) ;
  assign n22175 = n1481 & ~n1829 ;
  assign n22176 = n18608 & n22175 ;
  assign n22177 = n9648 & ~n10977 ;
  assign n22178 = n20120 ^ n6691 ^ 1'b0 ;
  assign n22179 = ~n8170 & n22178 ;
  assign n22180 = n22179 ^ n19005 ^ 1'b0 ;
  assign n22181 = n22180 ^ n17123 ^ 1'b0 ;
  assign n22182 = n13682 ^ n3249 ^ 1'b0 ;
  assign n22183 = n6138 & ~n22182 ;
  assign n22184 = n15857 & n22183 ;
  assign n22185 = ( n1263 & n2053 ) | ( n1263 & n3332 ) | ( n2053 & n3332 ) ;
  assign n22186 = n7966 ^ n4858 ^ 1'b0 ;
  assign n22187 = ~n5257 & n22186 ;
  assign n22188 = n2908 & ~n22187 ;
  assign n22189 = n1928 | n4027 ;
  assign n22190 = n3254 & ~n22189 ;
  assign n22191 = n840 | n22190 ;
  assign n22192 = n282 | n11380 ;
  assign n22193 = n22192 ^ n11679 ^ 1'b0 ;
  assign n22194 = ~n377 & n6455 ;
  assign n22195 = n419 & n7872 ;
  assign n22196 = ~n3113 & n22195 ;
  assign n22197 = n10774 | n22196 ;
  assign n22198 = n22194 | n22197 ;
  assign n22199 = n21151 ^ n20202 ^ 1'b0 ;
  assign n22200 = ~n4700 & n22199 ;
  assign n22201 = ~n5852 & n6768 ;
  assign n22202 = ~n22200 & n22201 ;
  assign n22203 = n10504 & ~n11597 ;
  assign n22204 = n425 & ~n2169 ;
  assign n22205 = n22204 ^ n11898 ^ n1010 ;
  assign n22206 = n22205 ^ n21261 ^ 1'b0 ;
  assign n22207 = n15806 ^ n14151 ^ 1'b0 ;
  assign n22208 = ( n718 & ~n2060 ) | ( n718 & n19703 ) | ( ~n2060 & n19703 ) ;
  assign n22209 = n22208 ^ n15536 ^ 1'b0 ;
  assign n22210 = ~n7367 & n8931 ;
  assign n22211 = n22210 ^ n1966 ^ 1'b0 ;
  assign n22212 = n22211 ^ n16222 ^ 1'b0 ;
  assign n22213 = n6114 & ~n19816 ;
  assign n22214 = ~n7325 & n18782 ;
  assign n22215 = n1108 | n15863 ;
  assign n22216 = n22215 ^ n5563 ^ 1'b0 ;
  assign n22217 = n2574 | n4475 ;
  assign n22218 = n22217 ^ n4354 ^ 1'b0 ;
  assign n22219 = n9198 & n22218 ;
  assign n22220 = n6687 & n18545 ;
  assign n22221 = ( ~n20128 & n22219 ) | ( ~n20128 & n22220 ) | ( n22219 & n22220 ) ;
  assign n22222 = n22216 & ~n22221 ;
  assign n22223 = n3022 & n5696 ;
  assign n22224 = n22223 ^ n17390 ^ 1'b0 ;
  assign n22228 = n5641 | n9724 ;
  assign n22225 = ~n1511 & n3676 ;
  assign n22226 = n15810 ^ n740 ^ 1'b0 ;
  assign n22227 = n22225 & n22226 ;
  assign n22229 = n22228 ^ n22227 ^ n1521 ;
  assign n22230 = ( n7723 & n11530 ) | ( n7723 & n17069 ) | ( n11530 & n17069 ) ;
  assign n22231 = n15847 ^ n8716 ^ 1'b0 ;
  assign n22232 = n3615 & n22231 ;
  assign n22233 = n22232 ^ n6563 ^ 1'b0 ;
  assign n22234 = n22233 ^ n8929 ^ 1'b0 ;
  assign n22235 = n22234 ^ n2840 ^ n2422 ;
  assign n22236 = n18201 ^ n8089 ^ 1'b0 ;
  assign n22237 = n10101 ^ n1133 ^ 1'b0 ;
  assign n22238 = n12207 & n22237 ;
  assign n22239 = n18251 ^ n10658 ^ 1'b0 ;
  assign n22240 = n21040 | n22239 ;
  assign n22241 = n4131 ^ n1675 ^ 1'b0 ;
  assign n22242 = n3702 ^ n3301 ^ 1'b0 ;
  assign n22243 = ~n22241 & n22242 ;
  assign n22244 = n3653 ^ n3647 ^ 1'b0 ;
  assign n22245 = n1853 & n4955 ;
  assign n22246 = n16894 & n22245 ;
  assign n22247 = ( ~n716 & n3214 ) | ( ~n716 & n19376 ) | ( n3214 & n19376 ) ;
  assign n22248 = n15337 ^ n10179 ^ 1'b0 ;
  assign n22249 = n20228 | n22248 ;
  assign n22250 = n4382 & n10670 ;
  assign n22251 = n8680 ^ n7795 ^ n2505 ;
  assign n22252 = n8476 | n22251 ;
  assign n22253 = n22252 ^ n12413 ^ 1'b0 ;
  assign n22254 = n3424 & ~n17694 ;
  assign n22255 = n7642 & n8856 ;
  assign n22256 = n4699 ^ n1815 ^ 1'b0 ;
  assign n22257 = n7022 ^ n4652 ^ 1'b0 ;
  assign n22262 = n2870 & ~n4589 ;
  assign n22263 = n4589 & n22262 ;
  assign n22261 = n3590 | n9412 ;
  assign n22264 = n22263 ^ n22261 ^ 1'b0 ;
  assign n22258 = x106 & ~n3036 ;
  assign n22259 = ~x106 & n22258 ;
  assign n22260 = n10747 & ~n22259 ;
  assign n22265 = n22264 ^ n22260 ^ 1'b0 ;
  assign n22266 = n619 & n1583 ;
  assign n22267 = n22266 ^ n11120 ^ 1'b0 ;
  assign n22268 = n8994 ^ n6859 ^ 1'b0 ;
  assign n22269 = ~n19680 & n22268 ;
  assign n22272 = ~n1044 & n13864 ;
  assign n22273 = n3563 & n22272 ;
  assign n22270 = n3853 & ~n4407 ;
  assign n22271 = n22270 ^ n10721 ^ n7804 ;
  assign n22274 = n22273 ^ n22271 ^ n17441 ;
  assign n22275 = n13668 | n22274 ;
  assign n22276 = n14735 ^ n5743 ^ 1'b0 ;
  assign n22277 = n6095 | n18648 ;
  assign n22278 = n3604 & ~n22277 ;
  assign n22279 = n1276 & n16402 ;
  assign n22280 = n22279 ^ n12265 ^ 1'b0 ;
  assign n22281 = n4420 & ~n16860 ;
  assign n22282 = n9583 ^ n8862 ^ 1'b0 ;
  assign n22283 = n7647 | n22282 ;
  assign n22284 = n886 & ~n11955 ;
  assign n22285 = n22283 & n22284 ;
  assign n22286 = ( ~n5509 & n13720 ) | ( ~n5509 & n22285 ) | ( n13720 & n22285 ) ;
  assign n22289 = n6319 & n7490 ;
  assign n22287 = n12407 ^ n11810 ^ 1'b0 ;
  assign n22288 = n14141 | n22287 ;
  assign n22290 = n22289 ^ n22288 ^ 1'b0 ;
  assign n22291 = n4857 | n15877 ;
  assign n22292 = n3528 & ~n22291 ;
  assign n22293 = ~n2248 & n14510 ;
  assign n22294 = n22293 ^ n801 ^ 1'b0 ;
  assign n22295 = n2304 & ~n22294 ;
  assign n22296 = n16831 & n22295 ;
  assign n22297 = n11101 & n20359 ;
  assign n22298 = ~n1680 & n19544 ;
  assign n22299 = ( n1860 & n5008 ) | ( n1860 & n6048 ) | ( n5008 & n6048 ) ;
  assign n22300 = n1283 & n3752 ;
  assign n22301 = n22300 ^ n4263 ^ 1'b0 ;
  assign n22302 = n5861 | n22301 ;
  assign n22303 = n22299 | n22302 ;
  assign n22305 = n15826 ^ n1081 ^ 1'b0 ;
  assign n22304 = n2313 & ~n17490 ;
  assign n22306 = n22305 ^ n22304 ^ 1'b0 ;
  assign n22307 = n2537 & ~n13802 ;
  assign n22308 = n22307 ^ n4028 ^ 1'b0 ;
  assign n22309 = n14678 ^ n10095 ^ 1'b0 ;
  assign n22310 = n8832 ^ n4808 ^ 1'b0 ;
  assign n22311 = ~n8185 & n22310 ;
  assign n22312 = n19243 | n21923 ;
  assign n22313 = n14229 | n22312 ;
  assign n22314 = ~n3950 & n7955 ;
  assign n22315 = n22314 ^ n8425 ^ 1'b0 ;
  assign n22316 = n22315 ^ n19297 ^ 1'b0 ;
  assign n22317 = n17517 | n22316 ;
  assign n22318 = n14163 ^ n9919 ^ 1'b0 ;
  assign n22319 = n20871 & n22318 ;
  assign n22320 = n22319 ^ n8011 ^ n3757 ;
  assign n22321 = n19546 ^ n6041 ^ 1'b0 ;
  assign n22322 = n3948 & n14015 ;
  assign n22323 = n22322 ^ n21177 ^ 1'b0 ;
  assign n22324 = x96 | n15753 ;
  assign n22325 = n15617 ^ n610 ^ 1'b0 ;
  assign n22326 = n22324 | n22325 ;
  assign n22327 = n1150 | n22326 ;
  assign n22328 = n10709 | n19179 ;
  assign n22329 = n3767 & n11611 ;
  assign n22330 = ( n6651 & ~n15634 ) | ( n6651 & n22329 ) | ( ~n15634 & n22329 ) ;
  assign n22331 = ( ~n13633 & n19818 ) | ( ~n13633 & n22330 ) | ( n19818 & n22330 ) ;
  assign n22332 = ( ~n3560 & n8786 ) | ( ~n3560 & n12987 ) | ( n8786 & n12987 ) ;
  assign n22333 = ~n884 & n1494 ;
  assign n22334 = n22333 ^ n17602 ^ 1'b0 ;
  assign n22335 = ( n6063 & n9167 ) | ( n6063 & n22334 ) | ( n9167 & n22334 ) ;
  assign n22336 = n22335 ^ n5356 ^ 1'b0 ;
  assign n22337 = n1089 & n22336 ;
  assign n22338 = n18771 ^ n1181 ^ 1'b0 ;
  assign n22339 = n1581 | n22338 ;
  assign n22340 = n5788 & ~n13232 ;
  assign n22341 = ~n18022 & n21429 ;
  assign n22342 = n5896 | n7693 ;
  assign n22343 = n22341 & ~n22342 ;
  assign n22344 = n5092 | n7429 ;
  assign n22345 = n346 & ~n22344 ;
  assign n22346 = n10472 & ~n12258 ;
  assign n22347 = ~n11686 & n22346 ;
  assign n22348 = n10436 & n16082 ;
  assign n22349 = ( n3067 & ~n22347 ) | ( n3067 & n22348 ) | ( ~n22347 & n22348 ) ;
  assign n22350 = n4285 & n15271 ;
  assign n22351 = n22350 ^ n21655 ^ 1'b0 ;
  assign n22352 = ~x70 & n11490 ;
  assign n22353 = n22352 ^ n2790 ^ 1'b0 ;
  assign n22354 = ~n20251 & n22353 ;
  assign n22355 = n14744 & n22354 ;
  assign n22356 = n22351 | n22355 ;
  assign n22357 = n19405 ^ n6751 ^ 1'b0 ;
  assign n22360 = n7899 ^ n2705 ^ 1'b0 ;
  assign n22359 = ~n1256 & n6164 ;
  assign n22358 = n17611 ^ x63 ^ x26 ;
  assign n22361 = n22360 ^ n22359 ^ n22358 ;
  assign n22362 = n2483 ^ n1154 ^ 1'b0 ;
  assign n22363 = n22362 ^ n6164 ^ 1'b0 ;
  assign n22364 = n15668 ^ n7379 ^ n7016 ;
  assign n22365 = ( n4456 & ~n8249 ) | ( n4456 & n22364 ) | ( ~n8249 & n22364 ) ;
  assign n22366 = ( n8895 & ~n22363 ) | ( n8895 & n22365 ) | ( ~n22363 & n22365 ) ;
  assign n22367 = n15401 ^ n7288 ^ 1'b0 ;
  assign n22368 = ~n4279 & n22367 ;
  assign n22369 = n22368 ^ n18726 ^ 1'b0 ;
  assign n22370 = n4946 ^ n1313 ^ 1'b0 ;
  assign n22371 = n14398 | n22370 ;
  assign n22372 = n3999 & ~n5829 ;
  assign n22373 = n22372 ^ n5018 ^ 1'b0 ;
  assign n22374 = n9331 ^ n8621 ^ 1'b0 ;
  assign n22375 = n6517 ^ n1753 ^ n322 ;
  assign n22376 = n8574 & n22375 ;
  assign n22377 = n22374 & n22376 ;
  assign n22378 = n8259 & ~n17190 ;
  assign n22379 = n22378 ^ n12592 ^ 1'b0 ;
  assign n22380 = n4180 & ~n12132 ;
  assign n22381 = ~n10951 & n22380 ;
  assign n22382 = n11419 & ~n18938 ;
  assign n22383 = n8738 & n22382 ;
  assign n22384 = n16186 ^ n13724 ^ 1'b0 ;
  assign n22385 = n9090 ^ n9045 ^ 1'b0 ;
  assign n22386 = n3395 | n5025 ;
  assign n22387 = n22386 ^ n5633 ^ n2742 ;
  assign n22388 = n6768 & n18126 ;
  assign n22389 = ~n11524 & n22388 ;
  assign n22390 = n10448 | n22389 ;
  assign n22391 = ~n488 & n13449 ;
  assign n22392 = n13052 ^ n9356 ^ 1'b0 ;
  assign n22393 = ( x33 & n235 ) | ( x33 & n571 ) | ( n235 & n571 ) ;
  assign n22394 = n22393 ^ n1856 ^ x87 ;
  assign n22395 = n6448 | n22394 ;
  assign n22396 = n14815 ^ n8075 ^ 1'b0 ;
  assign n22397 = n16977 ^ n8438 ^ n500 ;
  assign n22398 = ~n4113 & n5941 ;
  assign n22399 = n22398 ^ n19118 ^ 1'b0 ;
  assign n22401 = n6919 & n22196 ;
  assign n22400 = n4227 & n5868 ;
  assign n22402 = n22401 ^ n22400 ^ 1'b0 ;
  assign n22403 = n18625 ^ n925 ^ 1'b0 ;
  assign n22404 = ( x111 & n4358 ) | ( x111 & n22403 ) | ( n4358 & n22403 ) ;
  assign n22405 = n14946 & ~n22404 ;
  assign n22406 = ~n5330 & n7796 ;
  assign n22407 = n3599 & ~n22406 ;
  assign n22408 = ~n2435 & n3172 ;
  assign n22409 = n22408 ^ n6701 ^ 1'b0 ;
  assign n22410 = n571 | n3352 ;
  assign n22411 = n22410 ^ n1293 ^ 1'b0 ;
  assign n22412 = ~n2847 & n22411 ;
  assign n22413 = n22412 ^ n1721 ^ 1'b0 ;
  assign n22414 = n22409 | n22413 ;
  assign n22415 = n12463 ^ n12023 ^ 1'b0 ;
  assign n22416 = n9366 | n22415 ;
  assign n22417 = n15699 | n22416 ;
  assign n22418 = n16512 ^ n14105 ^ n3653 ;
  assign n22419 = n3985 ^ n3128 ^ 1'b0 ;
  assign n22420 = n22418 & ~n22419 ;
  assign n22421 = n22420 ^ n18150 ^ n13553 ;
  assign n22423 = n3969 & n15229 ;
  assign n22422 = n6631 & n10327 ;
  assign n22424 = n22423 ^ n22422 ^ 1'b0 ;
  assign n22425 = n1680 | n14920 ;
  assign n22426 = n9720 & n22425 ;
  assign n22427 = n11584 & n19603 ;
  assign n22428 = n2304 ^ n1578 ^ n1036 ;
  assign n22429 = n19015 ^ n9229 ^ 1'b0 ;
  assign n22430 = x19 & ~n22429 ;
  assign n22431 = n22430 ^ n533 ^ 1'b0 ;
  assign n22432 = n19485 | n22431 ;
  assign n22433 = n15062 | n22432 ;
  assign n22434 = n4981 & ~n22433 ;
  assign n22435 = n1256 ^ n435 ^ 1'b0 ;
  assign n22436 = n12786 & n22435 ;
  assign n22437 = n20032 ^ n14354 ^ n2024 ;
  assign n22438 = ~n3939 & n22437 ;
  assign n22439 = n20984 ^ n17099 ^ 1'b0 ;
  assign n22440 = n22439 ^ n10459 ^ 1'b0 ;
  assign n22441 = n4597 & n22440 ;
  assign n22442 = n22441 ^ n702 ^ 1'b0 ;
  assign n22443 = n6451 ^ n5723 ^ n3658 ;
  assign n22444 = n9979 & ~n15820 ;
  assign n22445 = n1097 & ~n22444 ;
  assign n22446 = n22445 ^ n7594 ^ 1'b0 ;
  assign n22447 = n22446 ^ n5407 ^ 1'b0 ;
  assign n22448 = n10212 ^ n3920 ^ 1'b0 ;
  assign n22449 = ~n15149 & n20232 ;
  assign n22450 = ~n22448 & n22449 ;
  assign n22451 = n15199 ^ n6539 ^ n210 ;
  assign n22452 = ( n1627 & n3066 ) | ( n1627 & ~n21025 ) | ( n3066 & ~n21025 ) ;
  assign n22453 = n22452 ^ n9542 ^ 1'b0 ;
  assign n22454 = n9426 | n22453 ;
  assign n22455 = ( x37 & ~n14511 ) | ( x37 & n15824 ) | ( ~n14511 & n15824 ) ;
  assign n22456 = n20932 ^ n14265 ^ n1922 ;
  assign n22457 = ~n668 & n11284 ;
  assign n22459 = n373 | n9927 ;
  assign n22458 = n4534 | n9304 ;
  assign n22460 = n22459 ^ n22458 ^ 1'b0 ;
  assign n22461 = ( n1198 & n3290 ) | ( n1198 & n16530 ) | ( n3290 & n16530 ) ;
  assign n22462 = n5425 & n22461 ;
  assign n22463 = n5339 | n9935 ;
  assign n22464 = ~n4528 & n12351 ;
  assign n22465 = n22464 ^ n12647 ^ 1'b0 ;
  assign n22466 = n9037 & ~n22465 ;
  assign n22467 = ~n22463 & n22466 ;
  assign n22468 = ~n10631 & n19707 ;
  assign n22469 = n865 | n4497 ;
  assign n22470 = n15190 ^ n7804 ^ 1'b0 ;
  assign n22471 = n20734 ^ n14958 ^ n5027 ;
  assign n22472 = n16083 ^ n14421 ^ 1'b0 ;
  assign n22473 = n1555 | n8230 ;
  assign n22474 = n22473 ^ n2002 ^ 1'b0 ;
  assign n22475 = n22474 ^ n9144 ^ n7547 ;
  assign n22476 = n22475 ^ n18719 ^ 1'b0 ;
  assign n22477 = n19351 | n22476 ;
  assign n22478 = n16517 ^ n14828 ^ 1'b0 ;
  assign n22479 = n11212 ^ n10113 ^ x101 ;
  assign n22480 = ~n14667 & n22479 ;
  assign n22481 = ~n22478 & n22480 ;
  assign n22482 = n4144 & n11190 ;
  assign n22483 = n19819 & n22482 ;
  assign n22484 = n8148 & ~n22483 ;
  assign n22485 = n22484 ^ n18820 ^ n6672 ;
  assign n22486 = n2325 & n21579 ;
  assign n22487 = n22486 ^ n5648 ^ 1'b0 ;
  assign n22488 = n13970 & n22487 ;
  assign n22489 = n22488 ^ n5922 ^ 1'b0 ;
  assign n22490 = n5900 & ~n22489 ;
  assign n22491 = n5218 ^ n619 ^ 1'b0 ;
  assign n22492 = n19031 | n22491 ;
  assign n22493 = n5183 & n8495 ;
  assign n22494 = n1205 & n22493 ;
  assign n22495 = n22494 ^ n6830 ^ 1'b0 ;
  assign n22496 = n2882 | n3030 ;
  assign n22497 = n22495 | n22496 ;
  assign n22498 = n3457 & n7641 ;
  assign n22499 = ~n5139 & n22498 ;
  assign n22500 = n17404 ^ n12673 ^ 1'b0 ;
  assign n22501 = ~n13593 & n22500 ;
  assign n22502 = n14655 & ~n20022 ;
  assign n22503 = n6959 & n22502 ;
  assign n22504 = ~n3340 & n6970 ;
  assign n22505 = n4456 | n22504 ;
  assign n22506 = ~n2800 & n10572 ;
  assign n22507 = ~n2868 & n5818 ;
  assign n22508 = n4382 & ~n22507 ;
  assign n22509 = n13119 ^ n12872 ^ n12224 ;
  assign n22510 = n15201 ^ n8144 ^ 1'b0 ;
  assign n22511 = ~n22509 & n22510 ;
  assign n22512 = n22508 | n22511 ;
  assign n22513 = n6558 ^ n729 ^ 1'b0 ;
  assign n22514 = n8942 | n22513 ;
  assign n22516 = ~n8877 & n12333 ;
  assign n22517 = n12132 & n22516 ;
  assign n22515 = ~x3 & n9862 ;
  assign n22518 = n22517 ^ n22515 ^ 1'b0 ;
  assign n22519 = n9874 | n11594 ;
  assign n22520 = n12683 & ~n22519 ;
  assign n22521 = n8469 | n22520 ;
  assign n22522 = n16558 | n22521 ;
  assign n22523 = n8170 ^ n2007 ^ 1'b0 ;
  assign n22524 = n5425 ^ n969 ^ 1'b0 ;
  assign n22525 = n5420 & ~n22524 ;
  assign n22526 = n22525 ^ n17211 ^ 1'b0 ;
  assign n22527 = ~n22523 & n22526 ;
  assign n22528 = n20283 ^ n7240 ^ 1'b0 ;
  assign n22529 = n2292 | n22528 ;
  assign n22530 = n22529 ^ n12652 ^ 1'b0 ;
  assign n22531 = n4564 & ~n22530 ;
  assign n22532 = n22527 & n22531 ;
  assign n22533 = n5805 | n10334 ;
  assign n22534 = n22533 ^ n1487 ^ 1'b0 ;
  assign n22535 = n10254 & n22534 ;
  assign n22536 = n8606 ^ n7240 ^ 1'b0 ;
  assign n22537 = ~n20606 & n22536 ;
  assign n22538 = ~n736 & n5693 ;
  assign n22539 = n4987 & n22538 ;
  assign n22540 = n9745 & ~n22539 ;
  assign n22541 = n1762 & ~n7900 ;
  assign n22542 = n22540 & n22541 ;
  assign n22543 = n20772 | n22542 ;
  assign n22544 = n18518 | n22543 ;
  assign n22545 = n10250 | n12469 ;
  assign n22546 = n11380 & n22545 ;
  assign n22547 = n9636 & n9735 ;
  assign n22548 = ~n21010 & n22547 ;
  assign n22549 = n21462 ^ n7934 ^ n6810 ;
  assign n22550 = ~n346 & n12018 ;
  assign n22551 = ( n3128 & n6829 ) | ( n3128 & ~n22550 ) | ( n6829 & ~n22550 ) ;
  assign n22552 = x24 & n3135 ;
  assign n22553 = ~n22551 & n22552 ;
  assign n22554 = ~n1484 & n3482 ;
  assign n22555 = ~n4751 & n22554 ;
  assign n22556 = x34 & n16961 ;
  assign n22557 = n7139 ^ n2850 ^ 1'b0 ;
  assign n22558 = n8198 & ~n22557 ;
  assign n22559 = ~n4907 & n22558 ;
  assign n22560 = n11419 ^ n2229 ^ 1'b0 ;
  assign n22561 = n7458 ^ n4213 ^ 1'b0 ;
  assign n22562 = ( n6984 & n18926 ) | ( n6984 & n22561 ) | ( n18926 & n22561 ) ;
  assign n22563 = x41 | n3012 ;
  assign n22564 = n19362 & ~n22563 ;
  assign n22565 = n22564 ^ n3864 ^ 1'b0 ;
  assign n22566 = x13 & n12812 ;
  assign n22567 = n22566 ^ n8872 ^ 1'b0 ;
  assign n22568 = n19051 ^ n8349 ^ 1'b0 ;
  assign n22569 = n22567 | n22568 ;
  assign n22570 = n8044 & n16191 ;
  assign n22571 = n4307 & n22570 ;
  assign n22572 = n10436 & ~n10701 ;
  assign n22573 = ~n6245 & n22572 ;
  assign n22583 = n3098 ^ n2785 ^ 1'b0 ;
  assign n22584 = n8495 & n22583 ;
  assign n22578 = ~n569 & n3103 ;
  assign n22579 = n22578 ^ n6442 ^ 1'b0 ;
  assign n22580 = n5681 & n22579 ;
  assign n22581 = ~x38 & n22580 ;
  assign n22574 = n4073 | n5041 ;
  assign n22575 = x33 & n4946 ;
  assign n22576 = n22575 ^ n7391 ^ 1'b0 ;
  assign n22577 = ( ~n712 & n22574 ) | ( ~n712 & n22576 ) | ( n22574 & n22576 ) ;
  assign n22582 = n22581 ^ n22577 ^ n21305 ;
  assign n22585 = n22584 ^ n22582 ^ 1'b0 ;
  assign n22586 = ~n13720 & n22585 ;
  assign n22587 = n1321 | n22003 ;
  assign n22588 = n15713 & ~n22587 ;
  assign n22589 = n8574 & ~n14371 ;
  assign n22590 = n11899 | n22589 ;
  assign n22591 = n1860 | n3340 ;
  assign n22592 = ( ~n1953 & n19769 ) | ( ~n1953 & n22591 ) | ( n19769 & n22591 ) ;
  assign n22593 = n22592 ^ n7756 ^ 1'b0 ;
  assign n22594 = n1168 | n4614 ;
  assign n22595 = n5548 | n22594 ;
  assign n22596 = n5064 & ~n22595 ;
  assign n22597 = n22596 ^ n12589 ^ 1'b0 ;
  assign n22598 = n15956 & ~n22597 ;
  assign n22599 = n19975 ^ n5946 ^ 1'b0 ;
  assign n22600 = ~n14412 & n22599 ;
  assign n22601 = x104 & ~n910 ;
  assign n22602 = n6436 & ~n11444 ;
  assign n22603 = n22602 ^ n3915 ^ 1'b0 ;
  assign n22604 = n8185 | n22603 ;
  assign n22605 = n15216 & ~n22604 ;
  assign n22606 = n2572 | n18811 ;
  assign n22607 = n22606 ^ n11696 ^ 1'b0 ;
  assign n22608 = n13733 ^ n8900 ^ n2487 ;
  assign n22609 = ~n8231 & n12562 ;
  assign n22610 = ( n7320 & ~n8622 ) | ( n7320 & n22609 ) | ( ~n8622 & n22609 ) ;
  assign n22611 = n1810 ^ n1711 ^ 1'b0 ;
  assign n22612 = n6217 | n22611 ;
  assign n22613 = n8779 ^ n2966 ^ 1'b0 ;
  assign n22614 = ~n22612 & n22613 ;
  assign n22615 = n597 & n3753 ;
  assign n22616 = n22615 ^ n3740 ^ 1'b0 ;
  assign n22617 = n22616 ^ n8040 ^ 1'b0 ;
  assign n22618 = n361 | n22617 ;
  assign n22619 = n9371 ^ n3591 ^ 1'b0 ;
  assign n22620 = ~n22618 & n22619 ;
  assign n22621 = ( n2369 & ~n11389 ) | ( n2369 & n11482 ) | ( ~n11389 & n11482 ) ;
  assign n22622 = n9655 | n10460 ;
  assign n22623 = n22622 ^ n3019 ^ 1'b0 ;
  assign n22624 = n15219 ^ n1481 ^ 1'b0 ;
  assign n22625 = ( n2074 & n22623 ) | ( n2074 & ~n22624 ) | ( n22623 & ~n22624 ) ;
  assign n22629 = n6005 ^ n1086 ^ 1'b0 ;
  assign n22630 = n22194 & n22629 ;
  assign n22626 = n6012 & ~n8128 ;
  assign n22627 = n22626 ^ n2157 ^ 1'b0 ;
  assign n22628 = ~n16501 & n22627 ;
  assign n22631 = n22630 ^ n22628 ^ n5657 ;
  assign n22632 = ~n5561 & n6063 ;
  assign n22633 = n16775 ^ n9535 ^ 1'b0 ;
  assign n22634 = n10250 & ~n22633 ;
  assign n22635 = n21385 ^ n7639 ^ 1'b0 ;
  assign n22636 = n22635 ^ n9210 ^ 1'b0 ;
  assign n22637 = n7524 | n9379 ;
  assign n22638 = n22637 ^ n18563 ^ 1'b0 ;
  assign n22639 = ~n3617 & n3849 ;
  assign n22640 = ~n1019 & n22639 ;
  assign n22641 = n2073 | n22640 ;
  assign n22642 = n1000 | n12209 ;
  assign n22643 = n22641 | n22642 ;
  assign n22644 = ( n148 & n405 ) | ( n148 & n655 ) | ( n405 & n655 ) ;
  assign n22645 = n22644 ^ n6864 ^ n5400 ;
  assign n22646 = ( n1542 & ~n3728 ) | ( n1542 & n17725 ) | ( ~n3728 & n17725 ) ;
  assign n22647 = n4844 & ~n10416 ;
  assign n22648 = ~n5581 & n22647 ;
  assign n22649 = n13749 ^ n8320 ^ n3900 ;
  assign n22650 = n22649 ^ n2312 ^ 1'b0 ;
  assign n22651 = n7833 | n22650 ;
  assign n22652 = ~n20809 & n22651 ;
  assign n22653 = n764 & ~n5355 ;
  assign n22654 = ~n20508 & n22653 ;
  assign n22655 = n1088 & n2444 ;
  assign n22656 = n196 & n22655 ;
  assign n22657 = ~n6941 & n22656 ;
  assign n22658 = n22657 ^ n8755 ^ n1378 ;
  assign n22659 = n1097 & n19037 ;
  assign n22660 = n22659 ^ n4308 ^ 1'b0 ;
  assign n22661 = n11024 & ~n19804 ;
  assign n22662 = n2102 & n22661 ;
  assign n22663 = ( ~n5155 & n22660 ) | ( ~n5155 & n22662 ) | ( n22660 & n22662 ) ;
  assign n22664 = n1835 & n10241 ;
  assign n22665 = ( n2929 & n17782 ) | ( n2929 & ~n18105 ) | ( n17782 & ~n18105 ) ;
  assign n22666 = n13692 & ~n22665 ;
  assign n22667 = n17458 ^ n1030 ^ 1'b0 ;
  assign n22672 = n16845 ^ n553 ^ 1'b0 ;
  assign n22668 = n9203 ^ n8849 ^ 1'b0 ;
  assign n22669 = ~n14186 & n22668 ;
  assign n22670 = n9567 & n22669 ;
  assign n22671 = n16299 & n22670 ;
  assign n22673 = n22672 ^ n22671 ^ 1'b0 ;
  assign n22674 = ( n588 & n21984 ) | ( n588 & n22228 ) | ( n21984 & n22228 ) ;
  assign n22675 = n18824 ^ n1722 ^ 1'b0 ;
  assign n22676 = n5747 ^ n4122 ^ 1'b0 ;
  assign n22677 = ~n2802 & n22676 ;
  assign n22678 = n6576 ^ n6569 ^ n5829 ;
  assign n22679 = n7296 & n22678 ;
  assign n22680 = n1106 | n6211 ;
  assign n22681 = n478 & n5923 ;
  assign n22682 = ~n306 & n22681 ;
  assign n22683 = n22680 | n22682 ;
  assign n22684 = n14202 ^ n1886 ^ 1'b0 ;
  assign n22685 = n11474 | n22684 ;
  assign n22686 = n2297 ^ n190 ^ 1'b0 ;
  assign n22687 = n17898 ^ n2640 ^ 1'b0 ;
  assign n22688 = ~n22686 & n22687 ;
  assign n22689 = n22688 ^ n1371 ^ 1'b0 ;
  assign n22690 = n19944 ^ n10542 ^ 1'b0 ;
  assign n22691 = n22507 ^ n22409 ^ n15843 ;
  assign n22693 = n11419 & ~n22673 ;
  assign n22692 = n4662 ^ n1805 ^ n868 ;
  assign n22694 = n22693 ^ n22692 ^ 1'b0 ;
  assign n22695 = n2079 & ~n19839 ;
  assign n22696 = n22695 ^ n14794 ^ 1'b0 ;
  assign n22697 = n1771 & n3156 ;
  assign n22698 = ~n2981 & n22697 ;
  assign n22699 = n7780 | n22698 ;
  assign n22700 = n22699 ^ n9093 ^ 1'b0 ;
  assign n22701 = n22700 ^ n22420 ^ 1'b0 ;
  assign n22702 = n8165 | n22701 ;
  assign n22703 = n22702 ^ n11389 ^ 1'b0 ;
  assign n22704 = n2866 & ~n3754 ;
  assign n22705 = n802 & ~n22704 ;
  assign n22706 = ~n14289 & n22705 ;
  assign n22707 = n13791 ^ n12900 ^ n2751 ;
  assign n22708 = n15190 ^ n1236 ^ 1'b0 ;
  assign n22709 = n312 | n10744 ;
  assign n22710 = n4650 ^ n3576 ^ 1'b0 ;
  assign n22711 = n12877 | n22710 ;
  assign n22712 = n6004 | n22711 ;
  assign n22713 = n15139 & n22712 ;
  assign n22714 = n15664 & n19861 ;
  assign n22715 = n7797 & n22714 ;
  assign n22716 = n14574 & ~n22715 ;
  assign n22717 = n22716 ^ n8541 ^ 1'b0 ;
  assign n22718 = ( n615 & n21802 ) | ( n615 & ~n22717 ) | ( n21802 & ~n22717 ) ;
  assign n22719 = n9634 & n21219 ;
  assign n22720 = n22719 ^ n4603 ^ 1'b0 ;
  assign n22721 = n3107 | n7674 ;
  assign n22722 = ~n4281 & n22721 ;
  assign n22723 = n22722 ^ n3304 ^ 1'b0 ;
  assign n22724 = n22723 ^ n5090 ^ 1'b0 ;
  assign n22725 = n13816 & ~n22724 ;
  assign n22726 = n2958 & n7442 ;
  assign n22727 = ~x37 & n22726 ;
  assign n22728 = n6819 & n22727 ;
  assign n22729 = ~n4570 & n15034 ;
  assign n22730 = n9020 & n22729 ;
  assign n22731 = n22730 ^ n7161 ^ n4197 ;
  assign n22732 = n1791 & n2526 ;
  assign n22733 = n22732 ^ n17329 ^ n4039 ;
  assign n22734 = n2875 & ~n16328 ;
  assign n22735 = n3109 | n3617 ;
  assign n22736 = n22735 ^ n1143 ^ 1'b0 ;
  assign n22737 = n17828 ^ n17255 ^ 1'b0 ;
  assign n22738 = n18844 & n22737 ;
  assign n22739 = n22738 ^ n20062 ^ 1'b0 ;
  assign n22740 = n5774 | n9142 ;
  assign n22741 = n7484 & ~n19757 ;
  assign n22742 = ~n3977 & n6304 ;
  assign n22743 = n3415 & n22742 ;
  assign n22744 = n22743 ^ n4452 ^ 1'b0 ;
  assign n22745 = ~n7555 & n16164 ;
  assign n22746 = ~n21091 & n22745 ;
  assign n22747 = n22744 | n22746 ;
  assign n22748 = n9974 & n16803 ;
  assign n22749 = ( n805 & ~n9594 ) | ( n805 & n16627 ) | ( ~n9594 & n16627 ) ;
  assign n22750 = n21526 & ~n22749 ;
  assign n22751 = n22750 ^ n1888 ^ 1'b0 ;
  assign n22754 = n5240 | n7225 ;
  assign n22755 = n2980 | n22754 ;
  assign n22752 = ( n4044 & n10982 ) | ( n4044 & ~n15029 ) | ( n10982 & ~n15029 ) ;
  assign n22753 = n22618 | n22752 ;
  assign n22756 = n22755 ^ n22753 ^ 1'b0 ;
  assign n22757 = n2189 | n4599 ;
  assign n22758 = n12779 & ~n22757 ;
  assign n22759 = n322 & n22758 ;
  assign n22760 = ~n6647 & n10499 ;
  assign n22761 = n7434 & n22760 ;
  assign n22762 = n19909 ^ n17697 ^ 1'b0 ;
  assign n22763 = ( ~n12893 & n13048 ) | ( ~n12893 & n15461 ) | ( n13048 & n15461 ) ;
  assign n22764 = ~n6776 & n7905 ;
  assign n22765 = n13335 & n22764 ;
  assign n22766 = n22765 ^ n22612 ^ 1'b0 ;
  assign n22767 = n6322 & n22766 ;
  assign n22768 = n5169 ^ n3250 ^ 1'b0 ;
  assign n22769 = n22767 & n22768 ;
  assign n22770 = n697 | n6860 ;
  assign n22771 = ~n22181 & n22770 ;
  assign n22773 = n3686 ^ n3374 ^ 1'b0 ;
  assign n22772 = n10686 & ~n14944 ;
  assign n22774 = n22773 ^ n22772 ^ 1'b0 ;
  assign n22775 = ( n3199 & ~n4923 ) | ( n3199 & n7680 ) | ( ~n4923 & n7680 ) ;
  assign n22776 = n22775 ^ n11982 ^ 1'b0 ;
  assign n22777 = n12592 & ~n22776 ;
  assign n22778 = n22777 ^ n2007 ^ 1'b0 ;
  assign n22779 = n22778 ^ n8146 ^ 1'b0 ;
  assign n22780 = n764 & n15144 ;
  assign n22782 = n6903 ^ n6411 ^ n2331 ;
  assign n22781 = n7222 & n15931 ;
  assign n22783 = n22782 ^ n22781 ^ 1'b0 ;
  assign n22784 = n16558 ^ n10216 ^ n165 ;
  assign n22785 = ( n3126 & n7781 ) | ( n3126 & n22784 ) | ( n7781 & n22784 ) ;
  assign n22786 = n1017 & ~n7575 ;
  assign n22787 = n22786 ^ n1173 ^ 1'b0 ;
  assign n22788 = n1064 ^ x91 ^ 1'b0 ;
  assign n22789 = n22787 | n22788 ;
  assign n22790 = ~n1966 & n15042 ;
  assign n22791 = n8841 ^ n3424 ^ 1'b0 ;
  assign n22792 = n15837 | n22791 ;
  assign n22793 = n22792 ^ n13504 ^ n567 ;
  assign n22794 = n3679 & ~n22793 ;
  assign n22795 = n22794 ^ n19873 ^ 1'b0 ;
  assign n22796 = n3773 & n9340 ;
  assign n22797 = n22796 ^ n16295 ^ 1'b0 ;
  assign n22800 = n10562 ^ n9691 ^ 1'b0 ;
  assign n22801 = ~n14716 & n22800 ;
  assign n22798 = n5862 & n16288 ;
  assign n22799 = n11835 & ~n22798 ;
  assign n22802 = n22801 ^ n22799 ^ n4789 ;
  assign n22803 = ( n452 & n4061 ) | ( n452 & ~n21736 ) | ( n4061 & ~n21736 ) ;
  assign n22804 = n2523 & n19414 ;
  assign n22805 = n1522 ^ n515 ^ 1'b0 ;
  assign n22806 = n16099 | n22805 ;
  assign n22807 = n22806 ^ n14331 ^ 1'b0 ;
  assign n22808 = n10863 | n22807 ;
  assign n22809 = n8740 & ~n12999 ;
  assign n22810 = n14064 ^ n215 ^ 1'b0 ;
  assign n22811 = ~n324 & n22810 ;
  assign n22812 = n2462 & ~n2801 ;
  assign n22813 = n19819 | n22812 ;
  assign n22814 = n4858 | n8331 ;
  assign n22815 = n22814 ^ n8956 ^ n2992 ;
  assign n22817 = n14354 ^ n9684 ^ n4325 ;
  assign n22816 = n2811 ^ x110 ^ 1'b0 ;
  assign n22818 = n22817 ^ n22816 ^ 1'b0 ;
  assign n22819 = ~n9289 & n18110 ;
  assign n22820 = n22819 ^ n3565 ^ 1'b0 ;
  assign n22821 = ( n3983 & n9162 ) | ( n3983 & n22037 ) | ( n9162 & n22037 ) ;
  assign n22822 = ~n1461 & n14236 ;
  assign n22823 = n3633 & n6136 ;
  assign n22824 = ~n17453 & n22823 ;
  assign n22825 = n22824 ^ n15969 ^ n14103 ;
  assign n22826 = ~n5517 & n22825 ;
  assign n22827 = n11731 ^ n5103 ^ 1'b0 ;
  assign n22828 = n8834 & ~n22827 ;
  assign n22829 = n2593 & ~n5359 ;
  assign n22830 = n22829 ^ n11753 ^ 1'b0 ;
  assign n22831 = n21458 & n22830 ;
  assign n22832 = n17341 ^ n12875 ^ 1'b0 ;
  assign n22833 = ~n9388 & n22832 ;
  assign n22834 = n22833 ^ n7240 ^ 1'b0 ;
  assign n22835 = n19325 | n22834 ;
  assign n22836 = n765 & ~n2755 ;
  assign n22837 = n3983 & n22836 ;
  assign n22838 = n7551 & n22837 ;
  assign n22839 = n1601 & n22838 ;
  assign n22840 = n22839 ^ n11597 ^ 1'b0 ;
  assign n22841 = n22840 ^ n12090 ^ 1'b0 ;
  assign n22842 = n1010 & n4071 ;
  assign n22843 = n2285 & n22842 ;
  assign n22844 = ( ~n3509 & n18477 ) | ( ~n3509 & n22843 ) | ( n18477 & n22843 ) ;
  assign n22845 = n11819 ^ n1335 ^ 1'b0 ;
  assign n22846 = ~n13692 & n22845 ;
  assign n22847 = n11053 ^ n805 ^ 1'b0 ;
  assign n22848 = n10668 & ~n22847 ;
  assign n22849 = ~n13393 & n22848 ;
  assign n22850 = n19666 | n22618 ;
  assign n22851 = n22850 ^ n16964 ^ 1'b0 ;
  assign n22852 = n15728 ^ n2648 ^ 1'b0 ;
  assign n22853 = n22852 ^ n10977 ^ 1'b0 ;
  assign n22854 = n6694 | n22853 ;
  assign n22855 = n12021 & ~n22854 ;
  assign n22856 = n11378 | n19153 ;
  assign n22857 = ~n2749 & n6520 ;
  assign n22859 = n8044 & n14440 ;
  assign n22858 = n2944 | n9349 ;
  assign n22860 = n22859 ^ n22858 ^ 1'b0 ;
  assign n22861 = n8349 ^ n7181 ^ 1'b0 ;
  assign n22862 = n4667 & n8616 ;
  assign n22863 = ( n19209 & n22861 ) | ( n19209 & n22862 ) | ( n22861 & n22862 ) ;
  assign n22864 = n9898 ^ n6566 ^ 1'b0 ;
  assign n22865 = n22864 ^ n4122 ^ 1'b0 ;
  assign n22866 = ( n5347 & n11149 ) | ( n5347 & n22865 ) | ( n11149 & n22865 ) ;
  assign n22867 = n4639 ^ n4547 ^ 1'b0 ;
  assign n22868 = n4460 & ~n6636 ;
  assign n22869 = ~n4460 & n22868 ;
  assign n22870 = ( n7894 & n8887 ) | ( n7894 & n22869 ) | ( n8887 & n22869 ) ;
  assign n22871 = n1972 & n2331 ;
  assign n22872 = n22871 ^ n939 ^ 1'b0 ;
  assign n22873 = ~n22870 & n22872 ;
  assign n22874 = n20531 ^ n6634 ^ 1'b0 ;
  assign n22875 = n13918 & n22874 ;
  assign n22876 = n22875 ^ n20885 ^ 1'b0 ;
  assign n22877 = n3269 & n20930 ;
  assign n22878 = n11351 & n22877 ;
  assign n22879 = n3624 & n12136 ;
  assign n22880 = n22879 ^ n7780 ^ 1'b0 ;
  assign n22881 = n7982 & ~n22880 ;
  assign n22882 = n12227 ^ n3439 ^ 1'b0 ;
  assign n22883 = n11509 & ~n22882 ;
  assign n22884 = n22883 ^ n12721 ^ n9933 ;
  assign n22885 = ~n3991 & n11483 ;
  assign n22886 = n22885 ^ n10121 ^ 1'b0 ;
  assign n22887 = n12515 & n16063 ;
  assign n22888 = ( n3919 & n11662 ) | ( n3919 & ~n22887 ) | ( n11662 & ~n22887 ) ;
  assign n22889 = ( n17259 & n22886 ) | ( n17259 & n22888 ) | ( n22886 & n22888 ) ;
  assign n22890 = ( ~n3919 & n11736 ) | ( ~n3919 & n16425 ) | ( n11736 & n16425 ) ;
  assign n22891 = n9229 & n10874 ;
  assign n22892 = n22891 ^ n6599 ^ 1'b0 ;
  assign n22893 = n5154 ^ n1248 ^ 1'b0 ;
  assign n22894 = n6045 & ~n8967 ;
  assign n22895 = ~n22893 & n22894 ;
  assign n22897 = n1639 | n6908 ;
  assign n22896 = n13735 | n15864 ;
  assign n22898 = n22897 ^ n22896 ^ 1'b0 ;
  assign n22899 = n22895 & n22898 ;
  assign n22900 = n17707 ^ n16533 ^ n15882 ;
  assign n22901 = n673 | n9866 ;
  assign n22902 = n3157 | n22901 ;
  assign n22903 = n1578 | n22902 ;
  assign n22904 = n22903 ^ n16137 ^ 1'b0 ;
  assign n22905 = n22900 & ~n22904 ;
  assign n22906 = x111 & n8850 ;
  assign n22907 = ~n2354 & n22906 ;
  assign n22908 = n1592 | n2401 ;
  assign n22909 = n5093 ^ n1452 ^ 1'b0 ;
  assign n22910 = ~n4462 & n22909 ;
  assign n22911 = n8114 & n22910 ;
  assign n22912 = ~n22908 & n22911 ;
  assign n22913 = n22912 ^ n15580 ^ n2178 ;
  assign n22914 = ~n4361 & n11921 ;
  assign n22915 = n1467 & n12587 ;
  assign n22916 = n22915 ^ n543 ^ 1'b0 ;
  assign n22917 = n9413 & ~n19607 ;
  assign n22918 = n827 | n14727 ;
  assign n22919 = n3012 & ~n22918 ;
  assign n22920 = n22919 ^ x23 ^ 1'b0 ;
  assign n22921 = n2719 | n10040 ;
  assign n22922 = n22921 ^ n13117 ^ n5863 ;
  assign n22923 = x47 & ~n16753 ;
  assign n22924 = n9257 & ~n18033 ;
  assign n22925 = n14979 & n22924 ;
  assign n22926 = n1265 & n1318 ;
  assign n22927 = n6546 & n22926 ;
  assign n22928 = n22927 ^ n6933 ^ 1'b0 ;
  assign n22929 = n22928 ^ n9720 ^ 1'b0 ;
  assign n22930 = n8212 | n22929 ;
  assign n22931 = n4785 & ~n13947 ;
  assign n22932 = n6271 & ~n22931 ;
  assign n22933 = n21045 ^ n5647 ^ 1'b0 ;
  assign n22934 = ~n22932 & n22933 ;
  assign n22935 = ~n3213 & n4285 ;
  assign n22936 = n5439 | n18009 ;
  assign n22937 = n5241 & ~n22936 ;
  assign n22938 = n11860 ^ n2218 ^ 1'b0 ;
  assign n22939 = ~n17791 & n22938 ;
  assign n22940 = ( ~x21 & n3087 ) | ( ~x21 & n22939 ) | ( n3087 & n22939 ) ;
  assign n22941 = ( n7471 & ~n18589 ) | ( n7471 & n20153 ) | ( ~n18589 & n20153 ) ;
  assign n22942 = n7915 ^ n2645 ^ 1'b0 ;
  assign n22943 = n6240 & ~n22942 ;
  assign n22944 = n11749 | n16486 ;
  assign n22945 = n10158 | n13467 ;
  assign n22946 = n9986 ^ n9455 ^ 1'b0 ;
  assign n22947 = n5363 & ~n22946 ;
  assign n22948 = n16655 ^ n3883 ^ 1'b0 ;
  assign n22949 = n22947 & n22948 ;
  assign n22950 = n1397 ^ n1203 ^ 1'b0 ;
  assign n22951 = n22950 ^ n14835 ^ 1'b0 ;
  assign n22952 = n20698 ^ n6140 ^ 1'b0 ;
  assign n22953 = n22033 & ~n22952 ;
  assign n22954 = n16435 ^ n7577 ^ 1'b0 ;
  assign n22955 = n14641 & n22954 ;
  assign n22956 = n3475 & ~n14793 ;
  assign n22957 = ~n18650 & n22956 ;
  assign n22958 = n22957 ^ n15843 ^ 1'b0 ;
  assign n22959 = n15822 ^ n12374 ^ 1'b0 ;
  assign n22960 = n2419 & ~n14708 ;
  assign n22961 = n7359 | n10467 ;
  assign n22962 = n22961 ^ n4075 ^ 1'b0 ;
  assign n22963 = ~n5457 & n12989 ;
  assign n22964 = n22963 ^ n13003 ^ 1'b0 ;
  assign n22965 = n11790 | n22964 ;
  assign n22966 = n18741 ^ n3528 ^ 1'b0 ;
  assign n22967 = n22787 | n22966 ;
  assign n22970 = n10627 & n18228 ;
  assign n22968 = n10030 ^ n6936 ^ 1'b0 ;
  assign n22969 = n13346 | n22968 ;
  assign n22971 = n22970 ^ n22969 ^ 1'b0 ;
  assign n22972 = n22971 ^ n10981 ^ n7496 ;
  assign n22973 = n10547 | n22972 ;
  assign n22974 = n828 & n18651 ;
  assign n22975 = n17519 ^ n5340 ^ n3023 ;
  assign n22976 = n12018 | n16689 ;
  assign n22977 = n487 & ~n10279 ;
  assign n22978 = n22977 ^ n2958 ^ 1'b0 ;
  assign n22979 = ~n8967 & n22978 ;
  assign n22980 = n22976 & n22979 ;
  assign n22981 = n5142 | n18440 ;
  assign n22982 = n5474 ^ n570 ^ 1'b0 ;
  assign n22983 = ~n22981 & n22982 ;
  assign n22984 = ~n4070 & n19566 ;
  assign n22985 = n6215 & n8861 ;
  assign n22986 = n2417 | n18736 ;
  assign n22987 = n15610 & ~n22986 ;
  assign n22988 = n2421 & n10551 ;
  assign n22989 = ~n4419 & n22988 ;
  assign n22990 = n5383 & ~n22989 ;
  assign n22992 = n1343 & n2192 ;
  assign n22991 = ~n859 & n1967 ;
  assign n22993 = n22992 ^ n22991 ^ 1'b0 ;
  assign n22994 = n22993 ^ n6498 ^ n6280 ;
  assign n22995 = n4138 ^ n2907 ^ 1'b0 ;
  assign n22996 = n3017 & ~n22995 ;
  assign n22997 = n22996 ^ n10594 ^ 1'b0 ;
  assign n22998 = n14810 ^ n8515 ^ 1'b0 ;
  assign n22999 = n11177 & ~n22998 ;
  assign n23000 = n1791 & ~n15918 ;
  assign n23001 = ~n7035 & n23000 ;
  assign n23002 = n11066 ^ n2411 ^ n1080 ;
  assign n23003 = n6918 | n23002 ;
  assign n23006 = ( n2070 & n15007 ) | ( n2070 & ~n18079 ) | ( n15007 & ~n18079 ) ;
  assign n23004 = n1088 & ~n2863 ;
  assign n23005 = n23004 ^ n4942 ^ 1'b0 ;
  assign n23007 = n23006 ^ n23005 ^ 1'b0 ;
  assign n23008 = ( n4942 & n10649 ) | ( n4942 & ~n17088 ) | ( n10649 & ~n17088 ) ;
  assign n23009 = n2461 & ~n5145 ;
  assign n23010 = ( n1151 & ~n17424 ) | ( n1151 & n23009 ) | ( ~n17424 & n23009 ) ;
  assign n23011 = n23008 & n23010 ;
  assign n23012 = n3978 ^ n2471 ^ 1'b0 ;
  assign n23013 = ~n3465 & n4667 ;
  assign n23014 = n23012 & ~n23013 ;
  assign n23015 = n6439 ^ n6264 ^ n3149 ;
  assign n23016 = n18954 ^ n1150 ^ 1'b0 ;
  assign n23017 = n4727 & n7368 ;
  assign n23018 = n23017 ^ n5783 ^ 1'b0 ;
  assign n23019 = n7567 & ~n8328 ;
  assign n23020 = n23018 & n23019 ;
  assign n23021 = n13896 & n15126 ;
  assign n23022 = n3328 | n4868 ;
  assign n23023 = n2742 | n23022 ;
  assign n23024 = n20474 ^ n3440 ^ 1'b0 ;
  assign n23025 = n23023 & ~n23024 ;
  assign n23026 = n175 & n8966 ;
  assign n23027 = ( ~n2090 & n15512 ) | ( ~n2090 & n21798 ) | ( n15512 & n21798 ) ;
  assign n23028 = n1713 | n8573 ;
  assign n23029 = n23028 ^ n22970 ^ 1'b0 ;
  assign n23030 = n19527 ^ n8415 ^ 1'b0 ;
  assign n23031 = n16805 & n23030 ;
  assign n23032 = ( ~n18698 & n23029 ) | ( ~n18698 & n23031 ) | ( n23029 & n23031 ) ;
  assign n23033 = n9271 | n20400 ;
  assign n23034 = n6696 & ~n16144 ;
  assign n23035 = n15584 & n23034 ;
  assign n23036 = n988 & n2079 ;
  assign n23037 = ~n3562 & n12772 ;
  assign n23038 = n23037 ^ n830 ^ 1'b0 ;
  assign n23039 = n4714 & ~n7197 ;
  assign n23040 = n23039 ^ n4686 ^ 1'b0 ;
  assign n23041 = n23040 ^ n12121 ^ 1'b0 ;
  assign n23042 = n22623 ^ n15583 ^ n3834 ;
  assign n23043 = n2690 & ~n10609 ;
  assign n23044 = n11760 | n15911 ;
  assign n23045 = n23044 ^ n607 ^ 1'b0 ;
  assign n23046 = n8432 & n8809 ;
  assign n23047 = n23046 ^ n10448 ^ 1'b0 ;
  assign n23048 = n22110 ^ n16587 ^ 1'b0 ;
  assign n23051 = n2243 & ~n6804 ;
  assign n23052 = n3352 & n23051 ;
  assign n23049 = n8142 & n13803 ;
  assign n23050 = n21246 & n23049 ;
  assign n23053 = n23052 ^ n23050 ^ 1'b0 ;
  assign n23054 = n19957 ^ n9455 ^ 1'b0 ;
  assign n23055 = ~n12779 & n23054 ;
  assign n23056 = ( n12907 & n12916 ) | ( n12907 & ~n23055 ) | ( n12916 & ~n23055 ) ;
  assign n23057 = n3181 & n12479 ;
  assign n23058 = n23057 ^ n20791 ^ 1'b0 ;
  assign n23059 = n6257 & ~n16648 ;
  assign n23060 = n6998 & n11579 ;
  assign n23061 = ~n3277 & n23060 ;
  assign n23062 = ~n12573 & n17191 ;
  assign n23063 = n23062 ^ n6728 ^ 1'b0 ;
  assign n23064 = n9409 & n17162 ;
  assign n23065 = ~n10218 & n23064 ;
  assign n23066 = n11926 & n20358 ;
  assign n23067 = ~n23065 & n23066 ;
  assign n23068 = n1982 | n6358 ;
  assign n23069 = n23068 ^ n7275 ^ 1'b0 ;
  assign n23070 = n3838 | n23069 ;
  assign n23071 = n14289 ^ n7090 ^ 1'b0 ;
  assign n23072 = n20251 ^ n8096 ^ 1'b0 ;
  assign n23073 = n14908 ^ n7117 ^ 1'b0 ;
  assign n23074 = ~n20658 & n23073 ;
  assign n23075 = n14837 ^ n933 ^ n725 ;
  assign n23076 = n5980 | n23075 ;
  assign n23077 = ~n8484 & n11536 ;
  assign n23078 = ~n11471 & n23077 ;
  assign n23079 = n1970 | n8331 ;
  assign n23081 = n990 | n1632 ;
  assign n23082 = n23081 ^ n11130 ^ n6610 ;
  assign n23080 = n7359 ^ n7135 ^ 1'b0 ;
  assign n23083 = n23082 ^ n23080 ^ n18911 ;
  assign n23084 = n23083 ^ n8355 ^ 1'b0 ;
  assign n23085 = n17866 ^ n11542 ^ 1'b0 ;
  assign n23086 = ~n15174 & n23085 ;
  assign n23087 = n4277 & ~n6539 ;
  assign n23088 = n10412 & n21102 ;
  assign n23089 = n3404 | n23088 ;
  assign n23090 = n23087 | n23089 ;
  assign n23091 = n7920 ^ n5324 ^ 1'b0 ;
  assign n23092 = n19145 ^ n16499 ^ 1'b0 ;
  assign n23096 = ( n1318 & n1432 ) | ( n1318 & n3085 ) | ( n1432 & n3085 ) ;
  assign n23093 = n1630 | n14674 ;
  assign n23094 = n23093 ^ n20867 ^ 1'b0 ;
  assign n23095 = n10502 & n23094 ;
  assign n23097 = n23096 ^ n23095 ^ 1'b0 ;
  assign n23098 = n12493 ^ n10772 ^ 1'b0 ;
  assign n23099 = n5443 | n23098 ;
  assign n23100 = ( n11984 & ~n20382 ) | ( n11984 & n20690 ) | ( ~n20382 & n20690 ) ;
  assign n23101 = n4961 & n19193 ;
  assign n23102 = n7973 & ~n19426 ;
  assign n23103 = ~n7251 & n19604 ;
  assign n23104 = ~n19975 & n23103 ;
  assign n23105 = ~n1795 & n19806 ;
  assign n23106 = n5413 & n12252 ;
  assign n23107 = n5796 & ~n23106 ;
  assign n23108 = n22682 & n23107 ;
  assign n23109 = ( ~n1358 & n9498 ) | ( ~n1358 & n22180 ) | ( n9498 & n22180 ) ;
  assign n23110 = n4272 ^ n406 ^ 1'b0 ;
  assign n23111 = n18298 & n23110 ;
  assign n23112 = n8676 & n23111 ;
  assign n23115 = n11780 ^ n1100 ^ 1'b0 ;
  assign n23113 = n1643 & ~n4678 ;
  assign n23114 = n8732 & n23113 ;
  assign n23116 = n23115 ^ n23114 ^ n7654 ;
  assign n23117 = x46 & ~n10631 ;
  assign n23118 = n23117 ^ n10395 ^ 1'b0 ;
  assign n23119 = n14888 ^ n3325 ^ 1'b0 ;
  assign n23120 = n14784 | n23119 ;
  assign n23121 = n14338 ^ n11320 ^ 1'b0 ;
  assign n23122 = n23121 ^ n5371 ^ 1'b0 ;
  assign n23123 = n7879 ^ n1788 ^ 1'b0 ;
  assign n23124 = n4090 & ~n23123 ;
  assign n23125 = n5156 & n16087 ;
  assign n23126 = ~n23124 & n23125 ;
  assign n23127 = n17821 ^ n5752 ^ 1'b0 ;
  assign n23128 = n9477 | n23127 ;
  assign n23129 = n2189 & n23128 ;
  assign n23130 = ( n7836 & ~n14810 ) | ( n7836 & n18083 ) | ( ~n14810 & n18083 ) ;
  assign n23131 = n11014 ^ n4502 ^ 1'b0 ;
  assign n23132 = n20435 & ~n23131 ;
  assign n23133 = n9222 & n23132 ;
  assign n23134 = n2478 & n14791 ;
  assign n23135 = n1436 & n2819 ;
  assign n23136 = ~n9297 & n10941 ;
  assign n23137 = n12631 & ~n23136 ;
  assign n23138 = n9026 ^ n1074 ^ 1'b0 ;
  assign n23139 = ~n3297 & n23138 ;
  assign n23140 = n2892 ^ n1929 ^ 1'b0 ;
  assign n23141 = n345 & ~n23140 ;
  assign n23142 = ~n19094 & n23141 ;
  assign n23143 = n20465 ^ n9832 ^ n6923 ;
  assign n23144 = n2622 & n3908 ;
  assign n23145 = ~n4459 & n9610 ;
  assign n23146 = ( n20099 & ~n23144 ) | ( n20099 & n23145 ) | ( ~n23144 & n23145 ) ;
  assign n23147 = n13723 ^ n11530 ^ 1'b0 ;
  assign n23148 = n22033 & ~n23147 ;
  assign n23149 = n5620 & n16534 ;
  assign n23150 = ~n352 & n23149 ;
  assign n23151 = n20579 ^ n14056 ^ 1'b0 ;
  assign n23152 = ~n23150 & n23151 ;
  assign n23153 = n7681 | n20283 ;
  assign n23154 = n22205 ^ n6743 ^ 1'b0 ;
  assign n23155 = n7529 | n23154 ;
  assign n23156 = n23155 ^ n22812 ^ 1'b0 ;
  assign n23157 = n22793 | n23156 ;
  assign n23158 = n22167 ^ n5217 ^ 1'b0 ;
  assign n23159 = n5990 ^ n433 ^ 1'b0 ;
  assign n23160 = n6631 & n23159 ;
  assign n23161 = n14060 ^ n135 ^ 1'b0 ;
  assign n23162 = n10624 ^ n3547 ^ 1'b0 ;
  assign n23163 = n23162 ^ n9917 ^ n1766 ;
  assign n23164 = n9039 ^ n3591 ^ 1'b0 ;
  assign n23165 = n18752 ^ n791 ^ 1'b0 ;
  assign n23166 = n7797 | n18296 ;
  assign n23167 = n5845 | n23166 ;
  assign n23168 = ~n18217 & n23167 ;
  assign n23169 = ~n3282 & n23168 ;
  assign n23170 = x121 & n14442 ;
  assign n23171 = n23170 ^ n18702 ^ 1'b0 ;
  assign n23172 = n3617 ^ n1599 ^ 1'b0 ;
  assign n23173 = n2940 & ~n23172 ;
  assign n23174 = ~n20685 & n23173 ;
  assign n23175 = n23174 ^ n337 ^ 1'b0 ;
  assign n23176 = n7623 | n23175 ;
  assign n23177 = n23176 ^ n9989 ^ 1'b0 ;
  assign n23178 = n13862 ^ n6747 ^ 1'b0 ;
  assign n23179 = n7172 | n23178 ;
  assign n23180 = n4449 & n4693 ;
  assign n23181 = ~n19189 & n23180 ;
  assign n23182 = ~n16482 & n20312 ;
  assign n23183 = n23181 & n23182 ;
  assign n23185 = n10707 ^ n3916 ^ 1'b0 ;
  assign n23186 = n8730 & n23185 ;
  assign n23184 = n6553 & ~n7836 ;
  assign n23187 = n23186 ^ n23184 ^ 1'b0 ;
  assign n23188 = n5519 ^ n3538 ^ 1'b0 ;
  assign n23189 = n20262 ^ n519 ^ 1'b0 ;
  assign n23190 = n6220 | n23189 ;
  assign n23191 = n20285 ^ n1033 ^ 1'b0 ;
  assign n23192 = x3 & ~n23191 ;
  assign n23193 = ~n16003 & n23192 ;
  assign n23194 = n19395 ^ n5277 ^ 1'b0 ;
  assign n23195 = ~n6428 & n23194 ;
  assign n23196 = n4273 & n23118 ;
  assign n23197 = n646 & n17234 ;
  assign n23198 = n23197 ^ n2802 ^ 1'b0 ;
  assign n23203 = ~n1309 & n4044 ;
  assign n23201 = n20805 ^ n12205 ^ 1'b0 ;
  assign n23202 = n733 | n23201 ;
  assign n23199 = ( n3640 & ~n4564 ) | ( n3640 & n9178 ) | ( ~n4564 & n9178 ) ;
  assign n23200 = n6114 & n23199 ;
  assign n23204 = n23203 ^ n23202 ^ n23200 ;
  assign n23205 = n22154 ^ n12287 ^ n7881 ;
  assign n23206 = n15337 ^ n2926 ^ 1'b0 ;
  assign n23207 = ~n310 & n1205 ;
  assign n23208 = n23207 ^ n3547 ^ 1'b0 ;
  assign n23209 = ~n4456 & n8500 ;
  assign n23210 = ~n23208 & n23209 ;
  assign n23211 = ( n6148 & n14152 ) | ( n6148 & ~n23210 ) | ( n14152 & ~n23210 ) ;
  assign n23212 = n9341 | n16953 ;
  assign n23213 = n23211 & ~n23212 ;
  assign n23214 = n11713 | n21461 ;
  assign n23215 = n23214 ^ n19197 ^ 1'b0 ;
  assign n23216 = n11542 | n20765 ;
  assign n23217 = n19308 & ~n23216 ;
  assign n23218 = n5654 & ~n7646 ;
  assign n23219 = n13912 & n23218 ;
  assign n23220 = n1145 | n4532 ;
  assign n23223 = n484 & n2570 ;
  assign n23224 = n23223 ^ n19035 ^ 1'b0 ;
  assign n23221 = n12015 | n16179 ;
  assign n23222 = n8028 & ~n23221 ;
  assign n23225 = n23224 ^ n23222 ^ n14647 ;
  assign n23226 = n22208 ^ n8341 ^ 1'b0 ;
  assign n23227 = n1680 | n16436 ;
  assign n23228 = n10749 | n23227 ;
  assign n23229 = n16083 ^ n13604 ^ 1'b0 ;
  assign n23230 = n19865 ^ n8417 ^ 1'b0 ;
  assign n23231 = n4097 & ~n23230 ;
  assign n23232 = n18909 ^ n4528 ^ 1'b0 ;
  assign n23233 = n22796 ^ n3447 ^ 1'b0 ;
  assign n23234 = n12438 ^ n2649 ^ 1'b0 ;
  assign n23235 = ~n3409 & n23234 ;
  assign n23236 = n9413 & n23235 ;
  assign n23237 = ~n1290 & n23236 ;
  assign n23238 = ( n2194 & n9007 ) | ( n2194 & ~n22928 ) | ( n9007 & ~n22928 ) ;
  assign n23239 = n15804 ^ n8537 ^ 1'b0 ;
  assign n23240 = ~n7031 & n13549 ;
  assign n23241 = n5223 & n23240 ;
  assign n23242 = n15253 & n23241 ;
  assign n23243 = n6937 & ~n10134 ;
  assign n23244 = n4452 & ~n22425 ;
  assign n23245 = n4858 ^ n1475 ^ 1'b0 ;
  assign n23246 = n19819 ^ n14173 ^ 1'b0 ;
  assign n23247 = n23245 & n23246 ;
  assign n23248 = ~n3159 & n6359 ;
  assign n23249 = n23248 ^ n975 ^ 1'b0 ;
  assign n23250 = n7048 & n23249 ;
  assign n23251 = ( n1615 & n4946 ) | ( n1615 & ~n23250 ) | ( n4946 & ~n23250 ) ;
  assign n23252 = ~n9164 & n10540 ;
  assign n23253 = n19778 ^ n6841 ^ 1'b0 ;
  assign n23254 = n9582 ^ n2399 ^ 1'b0 ;
  assign n23255 = ~n8190 & n23254 ;
  assign n23256 = n20030 ^ n4131 ^ 1'b0 ;
  assign n23257 = ~n23255 & n23256 ;
  assign n23258 = n15569 | n23257 ;
  assign n23259 = n18710 ^ n10223 ^ 1'b0 ;
  assign n23260 = n17478 | n23259 ;
  assign n23261 = n6170 ^ n6156 ^ n4439 ;
  assign n23262 = n23261 ^ n9572 ^ 1'b0 ;
  assign n23263 = n17987 | n23262 ;
  assign n23264 = n11987 & n16119 ;
  assign n23265 = n23264 ^ n9237 ^ 1'b0 ;
  assign n23266 = n23265 ^ n19335 ^ n17555 ;
  assign n23267 = ( n9048 & ~n10478 ) | ( n9048 & n14673 ) | ( ~n10478 & n14673 ) ;
  assign n23268 = n4308 | n23267 ;
  assign n23269 = n2243 | n23268 ;
  assign n23270 = ( n3156 & ~n7872 ) | ( n3156 & n8207 ) | ( ~n7872 & n8207 ) ;
  assign n23271 = n23270 ^ n14084 ^ n7594 ;
  assign n23272 = n12109 & n23271 ;
  assign n23273 = n14810 ^ n6799 ^ x116 ;
  assign n23274 = ( n7626 & ~n22019 ) | ( n7626 & n23273 ) | ( ~n22019 & n23273 ) ;
  assign n23275 = n23274 ^ n18558 ^ 1'b0 ;
  assign n23276 = n18325 & ~n23275 ;
  assign n23277 = n2706 & n10341 ;
  assign n23278 = n5485 & ~n12522 ;
  assign n23279 = ( n13316 & n16911 ) | ( n13316 & ~n21040 ) | ( n16911 & ~n21040 ) ;
  assign n23280 = ~n2167 & n14512 ;
  assign n23281 = n23280 ^ n7490 ^ 1'b0 ;
  assign n23282 = n1970 & ~n23281 ;
  assign n23283 = n654 ^ x51 ^ 1'b0 ;
  assign n23284 = n493 & n23283 ;
  assign n23285 = n23284 ^ n20258 ^ 1'b0 ;
  assign n23286 = n23285 ^ n18871 ^ n8187 ;
  assign n23287 = n13920 ^ n6199 ^ n5147 ;
  assign n23288 = n14306 ^ n13367 ^ 1'b0 ;
  assign n23289 = ~n8487 & n23288 ;
  assign n23290 = n23289 ^ n19809 ^ 1'b0 ;
  assign n23291 = ~n23287 & n23290 ;
  assign n23292 = n2184 & ~n13987 ;
  assign n23293 = n764 | n6247 ;
  assign n23294 = n23292 & ~n23293 ;
  assign n23297 = n10339 & ~n17429 ;
  assign n23298 = ~n11002 & n23297 ;
  assign n23295 = n18698 ^ n1615 ^ 1'b0 ;
  assign n23296 = ~n18820 & n23295 ;
  assign n23299 = n23298 ^ n23296 ^ 1'b0 ;
  assign n23300 = ~n6432 & n11683 ;
  assign n23301 = n23300 ^ n7462 ^ 1'b0 ;
  assign n23305 = n7550 & ~n14267 ;
  assign n23302 = n15620 ^ n3044 ^ 1'b0 ;
  assign n23303 = ~n4951 & n23302 ;
  assign n23304 = ~n16688 & n23303 ;
  assign n23306 = n23305 ^ n23304 ^ 1'b0 ;
  assign n23307 = n23306 ^ n22912 ^ n6717 ;
  assign n23308 = n10862 ^ n9900 ^ n7727 ;
  assign n23309 = n13341 ^ n6384 ^ 1'b0 ;
  assign n23310 = n16636 ^ n4075 ^ 1'b0 ;
  assign n23311 = n19839 ^ n12224 ^ 1'b0 ;
  assign n23312 = n23310 & ~n23311 ;
  assign n23313 = ~n6335 & n11070 ;
  assign n23314 = ~n12132 & n16216 ;
  assign n23315 = ~n23313 & n23314 ;
  assign n23316 = n6745 & n20030 ;
  assign n23317 = n575 & ~n2026 ;
  assign n23318 = n23317 ^ n10999 ^ 1'b0 ;
  assign n23319 = n20917 ^ n6828 ^ 1'b0 ;
  assign n23320 = ~n21755 & n23319 ;
  assign n23321 = n22603 ^ n1424 ^ 1'b0 ;
  assign n23322 = n5575 & ~n14718 ;
  assign n23323 = n3204 | n23322 ;
  assign n23324 = n23323 ^ n7705 ^ 1'b0 ;
  assign n23330 = ~n6457 & n12880 ;
  assign n23331 = n23330 ^ n8181 ^ 1'b0 ;
  assign n23326 = n5419 ^ n163 ^ 1'b0 ;
  assign n23325 = n7156 | n19649 ;
  assign n23327 = n23326 ^ n23325 ^ 1'b0 ;
  assign n23328 = n23327 ^ n2706 ^ 1'b0 ;
  assign n23329 = n23036 & n23328 ;
  assign n23332 = n23331 ^ n23329 ^ 1'b0 ;
  assign n23333 = n19591 ^ n12665 ^ 1'b0 ;
  assign n23334 = ~n9534 & n23333 ;
  assign n23335 = n20860 & n23334 ;
  assign n23336 = n20230 & n23335 ;
  assign n23337 = n619 & ~n6036 ;
  assign n23338 = n9515 & n23337 ;
  assign n23339 = n13186 | n23338 ;
  assign n23340 = n9149 ^ n4348 ^ 1'b0 ;
  assign n23341 = n12969 | n23340 ;
  assign n23353 = ( n182 & ~n2329 ) | ( n182 & n4041 ) | ( ~n2329 & n4041 ) ;
  assign n23345 = n691 & n1206 ;
  assign n23346 = ~n1206 & n23345 ;
  assign n23347 = ~n480 & n23346 ;
  assign n23348 = n2825 | n23347 ;
  assign n23349 = n23347 & ~n23348 ;
  assign n23350 = n10609 ^ n4819 ^ 1'b0 ;
  assign n23351 = ~n23349 & n23350 ;
  assign n23342 = n5326 & n9346 ;
  assign n23343 = n23342 ^ n10783 ^ 1'b0 ;
  assign n23344 = ~n2225 & n23343 ;
  assign n23352 = n23351 ^ n23344 ^ 1'b0 ;
  assign n23354 = n23353 ^ n23352 ^ 1'b0 ;
  assign n23355 = n11957 | n22529 ;
  assign n23356 = n23355 ^ n9381 ^ 1'b0 ;
  assign n23357 = ~n7410 & n23356 ;
  assign n23358 = n11686 & n14859 ;
  assign n23359 = n23358 ^ n6701 ^ 1'b0 ;
  assign n23360 = n21153 ^ n14119 ^ n2656 ;
  assign n23361 = ( n5680 & ~n10770 ) | ( n5680 & n17010 ) | ( ~n10770 & n17010 ) ;
  assign n23362 = n1500 | n3626 ;
  assign n23363 = n23362 ^ n3109 ^ 1'b0 ;
  assign n23364 = n2065 & n15863 ;
  assign n23365 = n18580 ^ n7142 ^ 1'b0 ;
  assign n23366 = n3738 & ~n9379 ;
  assign n23367 = ~n18057 & n23366 ;
  assign n23368 = n23326 ^ n1730 ^ 1'b0 ;
  assign n23369 = ( ~n2696 & n6963 ) | ( ~n2696 & n12238 ) | ( n6963 & n12238 ) ;
  assign n23370 = n2326 & n3662 ;
  assign n23371 = ~n23369 & n23370 ;
  assign n23372 = ~n7181 & n11579 ;
  assign n23373 = ( n805 & ~n3016 ) | ( n805 & n3617 ) | ( ~n3016 & n3617 ) ;
  assign n23374 = n14621 ^ n11382 ^ 1'b0 ;
  assign n23375 = ~n8427 & n23374 ;
  assign n23376 = n11525 | n20521 ;
  assign n23377 = n18226 | n23376 ;
  assign n23378 = n19354 ^ n14391 ^ 1'b0 ;
  assign n23379 = n23377 & n23378 ;
  assign n23380 = n1175 & n6223 ;
  assign n23381 = ~n19057 & n23380 ;
  assign n23382 = n12871 | n21086 ;
  assign n23383 = n23382 ^ n13307 ^ 1'b0 ;
  assign n23384 = n23383 ^ n16613 ^ n5955 ;
  assign n23385 = n4071 & ~n5014 ;
  assign n23386 = n23385 ^ n1412 ^ 1'b0 ;
  assign n23387 = n23386 ^ n5882 ^ 1'b0 ;
  assign n23388 = n5236 ^ n3930 ^ 1'b0 ;
  assign n23389 = n23387 & ~n23388 ;
  assign n23390 = n7560 & ~n13869 ;
  assign n23391 = n11391 ^ n2914 ^ 1'b0 ;
  assign n23392 = ~n17002 & n23391 ;
  assign n23393 = ( n7021 & n11736 ) | ( n7021 & n13199 ) | ( n11736 & n13199 ) ;
  assign n23394 = n23393 ^ n4727 ^ 1'b0 ;
  assign n23395 = x80 & n6349 ;
  assign n23396 = n5805 & n23395 ;
  assign n23397 = ( n7567 & n8865 ) | ( n7567 & n23396 ) | ( n8865 & n23396 ) ;
  assign n23398 = n22618 ^ n7597 ^ 1'b0 ;
  assign n23399 = n636 & ~n1610 ;
  assign n23400 = n23399 ^ n13548 ^ 1'b0 ;
  assign n23401 = n12685 & n21423 ;
  assign n23402 = n7469 | n23401 ;
  assign n23403 = n7172 & ~n23402 ;
  assign n23404 = n8338 | n12536 ;
  assign n23405 = n4395 | n14219 ;
  assign n23406 = n23404 | n23405 ;
  assign n23407 = n2451 & n7480 ;
  assign n23408 = ~n4614 & n5629 ;
  assign n23409 = ~n3649 & n23408 ;
  assign n23410 = n20947 & ~n23409 ;
  assign n23411 = ( n20133 & n23407 ) | ( n20133 & n23410 ) | ( n23407 & n23410 ) ;
  assign n23412 = n225 | n6724 ;
  assign n23413 = n23412 ^ n11894 ^ 1'b0 ;
  assign n23414 = ~n986 & n23413 ;
  assign n23415 = ( n730 & n1286 ) | ( n730 & ~n23414 ) | ( n1286 & ~n23414 ) ;
  assign n23416 = ( n3181 & n6586 ) | ( n3181 & ~n11780 ) | ( n6586 & ~n11780 ) ;
  assign n23420 = n10050 ^ n3706 ^ 1'b0 ;
  assign n23421 = x110 & ~n23420 ;
  assign n23417 = ~n5817 & n8116 ;
  assign n23418 = n23417 ^ n5517 ^ 1'b0 ;
  assign n23419 = n15263 | n23418 ;
  assign n23422 = n23421 ^ n23419 ^ 1'b0 ;
  assign n23423 = n8845 & ~n15540 ;
  assign n23424 = n3564 & ~n6073 ;
  assign n23425 = ~n14462 & n23424 ;
  assign n23426 = n12083 | n21864 ;
  assign n23427 = n20396 ^ n17077 ^ 1'b0 ;
  assign n23428 = n2365 | n23427 ;
  assign n23429 = ( ~n5852 & n6996 ) | ( ~n5852 & n23428 ) | ( n6996 & n23428 ) ;
  assign n23434 = ( ~n2654 & n4757 ) | ( ~n2654 & n17490 ) | ( n4757 & n17490 ) ;
  assign n23430 = n4683 & ~n5507 ;
  assign n23431 = ~n6212 & n23430 ;
  assign n23432 = n7692 | n23431 ;
  assign n23433 = n23432 ^ n20279 ^ 1'b0 ;
  assign n23435 = n23434 ^ n23433 ^ n8049 ;
  assign n23436 = ~n8310 & n16313 ;
  assign n23437 = ~n2851 & n23436 ;
  assign n23438 = ~n4186 & n4637 ;
  assign n23439 = n4059 ^ n2453 ^ 1'b0 ;
  assign n23440 = n2089 | n23439 ;
  assign n23441 = n21068 ^ n5546 ^ 1'b0 ;
  assign n23442 = ~n23440 & n23441 ;
  assign n23443 = n6473 & n19629 ;
  assign n23444 = n13827 & n23443 ;
  assign n23445 = n18774 ^ n13260 ^ n1272 ;
  assign n23446 = n23445 ^ n411 ^ 1'b0 ;
  assign n23449 = n2508 ^ n612 ^ 1'b0 ;
  assign n23450 = n17935 & ~n23449 ;
  assign n23448 = n14412 ^ n3563 ^ 1'b0 ;
  assign n23447 = n12338 ^ n12116 ^ n5010 ;
  assign n23451 = n23450 ^ n23448 ^ n23447 ;
  assign n23452 = n6148 | n8743 ;
  assign n23453 = n17138 & ~n23452 ;
  assign n23454 = n11168 | n14018 ;
  assign n23455 = ( n8654 & n23453 ) | ( n8654 & n23454 ) | ( n23453 & n23454 ) ;
  assign n23456 = n12308 & ~n21667 ;
  assign n23457 = n23456 ^ n6581 ^ 1'b0 ;
  assign n23458 = n12374 & n23457 ;
  assign n23459 = n1046 & n2278 ;
  assign n23460 = ~n3515 & n14105 ;
  assign n23461 = n23459 & n23460 ;
  assign n23462 = n15503 ^ n3674 ^ n557 ;
  assign n23463 = n4097 & n7798 ;
  assign n23464 = ~n9898 & n23463 ;
  assign n23465 = n23464 ^ n13001 ^ 1'b0 ;
  assign n23466 = n23450 ^ n11549 ^ n1528 ;
  assign n23467 = ~n23465 & n23466 ;
  assign n23468 = n1088 & n3480 ;
  assign n23469 = n13873 & n23468 ;
  assign n23470 = n6564 & ~n23469 ;
  assign n23471 = n6365 & n23470 ;
  assign n23472 = n13014 | n23471 ;
  assign n23473 = n23472 ^ n12379 ^ 1'b0 ;
  assign n23474 = ( n7814 & n8673 ) | ( n7814 & ~n17972 ) | ( n8673 & ~n17972 ) ;
  assign n23475 = n23474 ^ n20482 ^ n7253 ;
  assign n23476 = n1031 & ~n7143 ;
  assign n23477 = n22688 ^ n8775 ^ 1'b0 ;
  assign n23478 = n9294 ^ n5149 ^ 1'b0 ;
  assign n23479 = n10384 & ~n23478 ;
  assign n23480 = n13021 | n23479 ;
  assign n23481 = ( ~n5874 & n14053 ) | ( ~n5874 & n21219 ) | ( n14053 & n21219 ) ;
  assign n23482 = n12193 ^ n10609 ^ n1965 ;
  assign n23483 = n2197 & n2713 ;
  assign n23484 = ~x112 & n23483 ;
  assign n23485 = ( n3281 & n7391 ) | ( n3281 & n23484 ) | ( n7391 & n23484 ) ;
  assign n23486 = n4378 & n11225 ;
  assign n23487 = n9149 | n11370 ;
  assign n23488 = n15285 ^ n7816 ^ 1'b0 ;
  assign n23489 = ~n23487 & n23488 ;
  assign n23490 = n7845 & ~n7986 ;
  assign n23491 = n2858 & ~n23490 ;
  assign n23492 = ~n13747 & n23491 ;
  assign n23493 = n6228 & ~n14343 ;
  assign n23494 = n1897 & ~n4602 ;
  assign n23495 = n11379 & n23494 ;
  assign n23497 = n2419 & n11600 ;
  assign n23496 = n4564 | n22864 ;
  assign n23498 = n23497 ^ n23496 ^ 1'b0 ;
  assign n23499 = ~n6529 & n7130 ;
  assign n23500 = n23499 ^ n1314 ^ 1'b0 ;
  assign n23501 = ~n5077 & n17161 ;
  assign n23503 = n8206 | n20805 ;
  assign n23504 = n23503 ^ n3816 ^ n330 ;
  assign n23502 = n424 & n17826 ;
  assign n23505 = n23504 ^ n23502 ^ 1'b0 ;
  assign n23506 = ~n3924 & n23505 ;
  assign n23507 = ( n7865 & ~n8144 ) | ( n7865 & n17242 ) | ( ~n8144 & n17242 ) ;
  assign n23508 = n3658 ^ n683 ^ 1'b0 ;
  assign n23509 = n12591 | n16231 ;
  assign n23510 = n23508 | n23509 ;
  assign n23511 = n615 | n23510 ;
  assign n23512 = n5689 & n22294 ;
  assign n23513 = n23512 ^ n2935 ^ 1'b0 ;
  assign n23514 = n8006 & n23513 ;
  assign n23515 = ~n2712 & n22553 ;
  assign n23516 = n252 & ~n4817 ;
  assign n23517 = n23516 ^ n1974 ^ 1'b0 ;
  assign n23518 = n8277 ^ n5567 ^ 1'b0 ;
  assign n23519 = n20792 & ~n23518 ;
  assign n23520 = n23118 & ~n23519 ;
  assign n23521 = n23517 & n23520 ;
  assign n23522 = n6174 ^ n4178 ^ 1'b0 ;
  assign n23523 = n13723 & ~n23522 ;
  assign n23524 = n23523 ^ n22482 ^ 1'b0 ;
  assign n23525 = n6798 & ~n7637 ;
  assign n23526 = n12558 ^ n1999 ^ 1'b0 ;
  assign n23527 = n9339 & n23526 ;
  assign n23528 = n909 | n18431 ;
  assign n23529 = n13235 & ~n23528 ;
  assign n23530 = n10263 ^ n5393 ^ 1'b0 ;
  assign n23531 = n2589 & ~n23530 ;
  assign n23534 = ~n7099 & n8863 ;
  assign n23535 = n23534 ^ n5962 ^ 1'b0 ;
  assign n23533 = n14315 | n20566 ;
  assign n23536 = n23535 ^ n23533 ^ 1'b0 ;
  assign n23532 = n18635 & n20702 ;
  assign n23537 = n23536 ^ n23532 ^ 1'b0 ;
  assign n23538 = x122 | n4161 ;
  assign n23539 = n23538 ^ n6046 ^ 1'b0 ;
  assign n23540 = n9516 | n17390 ;
  assign n23541 = n23540 ^ n17967 ^ 1'b0 ;
  assign n23542 = ~n630 & n5077 ;
  assign n23543 = ~n2697 & n23542 ;
  assign n23544 = n20715 | n23543 ;
  assign n23545 = n3856 & ~n23544 ;
  assign n23546 = ( n2236 & ~n11074 ) | ( n2236 & n12691 ) | ( ~n11074 & n12691 ) ;
  assign n23547 = n23546 ^ n4450 ^ 1'b0 ;
  assign n23548 = n6387 | n20171 ;
  assign n23549 = n16665 ^ n642 ^ 1'b0 ;
  assign n23550 = ~n12767 & n13052 ;
  assign n23551 = n4698 & n23550 ;
  assign n23552 = n3562 & n23551 ;
  assign n23553 = ~n8738 & n10986 ;
  assign n23554 = n1061 & ~n23553 ;
  assign n23555 = n23554 ^ n4521 ^ 1'b0 ;
  assign n23556 = n17774 ^ n308 ^ 1'b0 ;
  assign n23557 = n17549 ^ n9461 ^ 1'b0 ;
  assign n23558 = n2958 & n23557 ;
  assign n23559 = ~n12734 & n23558 ;
  assign n23560 = n23559 ^ n11444 ^ 1'b0 ;
  assign n23561 = n23560 ^ n14363 ^ n6824 ;
  assign n23562 = n6075 & ~n17080 ;
  assign n23563 = n23562 ^ n4020 ^ 1'b0 ;
  assign n23564 = n22391 ^ n5145 ^ 1'b0 ;
  assign n23565 = ( n1492 & ~n14619 ) | ( n1492 & n21444 ) | ( ~n14619 & n21444 ) ;
  assign n23566 = n15601 ^ n7386 ^ 1'b0 ;
  assign n23567 = n485 | n23566 ;
  assign n23568 = n23567 ^ n14740 ^ 1'b0 ;
  assign n23569 = n5433 & n12281 ;
  assign n23570 = ~n2671 & n7701 ;
  assign n23571 = n23570 ^ n5039 ^ 1'b0 ;
  assign n23572 = n2135 | n23005 ;
  assign n23573 = n3195 & ~n11485 ;
  assign n23574 = n23573 ^ n16979 ^ 1'b0 ;
  assign n23575 = n12754 & ~n23574 ;
  assign n23576 = n5453 ^ n3453 ^ 1'b0 ;
  assign n23577 = n1568 & ~n23576 ;
  assign n23578 = n23577 ^ n9759 ^ 1'b0 ;
  assign n23579 = ~n15239 & n23578 ;
  assign n23580 = n6308 | n21601 ;
  assign n23581 = n10062 & n18469 ;
  assign n23582 = n2805 | n7847 ;
  assign n23583 = n23582 ^ n4768 ^ 1'b0 ;
  assign n23584 = n23583 ^ n13853 ^ 1'b0 ;
  assign n23585 = n15325 ^ n12082 ^ 1'b0 ;
  assign n23586 = ( ~n1086 & n20199 ) | ( ~n1086 & n22430 ) | ( n20199 & n22430 ) ;
  assign n23587 = n22187 ^ n1821 ^ 1'b0 ;
  assign n23588 = n19264 | n23587 ;
  assign n23589 = n13758 ^ n2159 ^ 1'b0 ;
  assign n23590 = ~n18415 & n21458 ;
  assign n23591 = n23590 ^ n21559 ^ 1'b0 ;
  assign n23592 = n11684 ^ n8138 ^ 1'b0 ;
  assign n23593 = x22 & ~n6867 ;
  assign n23594 = n6867 & n23593 ;
  assign n23595 = n16304 | n20759 ;
  assign n23596 = n23594 & ~n23595 ;
  assign n23597 = n16686 ^ n5589 ^ n4121 ;
  assign n23598 = ~n19813 & n23597 ;
  assign n23599 = n23596 | n23598 ;
  assign n23600 = n23599 ^ n13795 ^ 1'b0 ;
  assign n23601 = n6346 | n10179 ;
  assign n23602 = n904 | n23601 ;
  assign n23603 = n12497 & ~n21189 ;
  assign n23604 = n5651 & n23603 ;
  assign n23605 = n23604 ^ n11857 ^ 1'b0 ;
  assign n23606 = n13112 | n20504 ;
  assign n23607 = n7177 | n23606 ;
  assign n23608 = n15634 ^ n4259 ^ 1'b0 ;
  assign n23609 = ~n1414 & n8917 ;
  assign n23611 = ( ~n1034 & n13765 ) | ( ~n1034 & n17219 ) | ( n13765 & n17219 ) ;
  assign n23610 = n9375 & n15900 ;
  assign n23612 = n23611 ^ n23610 ^ 1'b0 ;
  assign n23613 = n5312 & n23612 ;
  assign n23614 = n23613 ^ n10175 ^ 1'b0 ;
  assign n23615 = n14928 | n17374 ;
  assign n23616 = n23615 ^ n9017 ^ 1'b0 ;
  assign n23617 = n19020 ^ n18503 ^ 1'b0 ;
  assign n23618 = n23617 ^ n18922 ^ n6159 ;
  assign n23619 = n9825 & ~n16122 ;
  assign n23620 = n7908 ^ n7348 ^ 1'b0 ;
  assign n23621 = ~n3191 & n16425 ;
  assign n23622 = n23620 & n23621 ;
  assign n23623 = n1394 | n23622 ;
  assign n23624 = n12929 ^ n5855 ^ 1'b0 ;
  assign n23625 = n6240 | n6581 ;
  assign n23626 = n23625 ^ n12386 ^ 1'b0 ;
  assign n23627 = n9684 & ~n23626 ;
  assign n23628 = n7802 & n13894 ;
  assign n23629 = n6164 & ~n15470 ;
  assign n23630 = n6435 | n13711 ;
  assign n23631 = n23630 ^ n15530 ^ 1'b0 ;
  assign n23632 = n9486 ^ n7286 ^ 1'b0 ;
  assign n23633 = x6 & n23632 ;
  assign n23634 = ( n935 & ~n2464 ) | ( n935 & n3135 ) | ( ~n2464 & n3135 ) ;
  assign n23635 = n23634 ^ n12858 ^ 1'b0 ;
  assign n23636 = ( n2353 & n14900 ) | ( n2353 & ~n23635 ) | ( n14900 & ~n23635 ) ;
  assign n23637 = ~n5475 & n18518 ;
  assign n23638 = n23637 ^ n872 ^ 1'b0 ;
  assign n23639 = n1560 & ~n23638 ;
  assign n23640 = n23639 ^ n2341 ^ 1'b0 ;
  assign n23641 = n1671 & n23640 ;
  assign n23642 = n23584 ^ n6522 ^ 1'b0 ;
  assign n23643 = n21920 | n23642 ;
  assign n23644 = n193 | n21984 ;
  assign n23645 = n1422 | n23644 ;
  assign n23646 = n23645 ^ n890 ^ 1'b0 ;
  assign n23647 = n10799 ^ n8645 ^ n967 ;
  assign n23648 = n10419 & ~n23647 ;
  assign n23649 = n5950 ^ n4596 ^ 1'b0 ;
  assign n23650 = ~n186 & n23649 ;
  assign n23651 = ~n23649 & n23650 ;
  assign n23652 = n4578 & ~n14412 ;
  assign n23653 = n18539 ^ n6722 ^ n750 ;
  assign n23654 = ~n10164 & n14698 ;
  assign n23655 = n23654 ^ n17744 ^ 1'b0 ;
  assign n23656 = n23655 ^ n10580 ^ 1'b0 ;
  assign n23658 = n802 ^ n701 ^ 1'b0 ;
  assign n23657 = ~n6020 & n20057 ;
  assign n23659 = n23658 ^ n23657 ^ 1'b0 ;
  assign n23660 = n16017 ^ n15242 ^ 1'b0 ;
  assign n23661 = n2041 | n6833 ;
  assign n23662 = ( n218 & n15234 ) | ( n218 & ~n23661 ) | ( n15234 & ~n23661 ) ;
  assign n23663 = n13658 ^ n235 ^ 1'b0 ;
  assign n23664 = n13231 & n23663 ;
  assign n23665 = n2353 & n12761 ;
  assign n23666 = n14552 ^ n10126 ^ 1'b0 ;
  assign n23667 = n9677 | n15966 ;
  assign n23668 = n1324 | n23667 ;
  assign n23669 = n2417 | n15410 ;
  assign n23670 = n8328 | n23669 ;
  assign n23671 = n23670 ^ n7103 ^ 1'b0 ;
  assign n23672 = n23671 ^ n11306 ^ 1'b0 ;
  assign n23673 = n1182 | n23672 ;
  assign n23674 = n23673 ^ n1080 ^ 1'b0 ;
  assign n23675 = n3468 ^ n1463 ^ 1'b0 ;
  assign n23676 = n2223 & n23675 ;
  assign n23677 = n18565 ^ n8733 ^ n769 ;
  assign n23678 = ( n1374 & ~n4214 ) | ( n1374 & n11836 ) | ( ~n4214 & n11836 ) ;
  assign n23679 = n13651 ^ n1364 ^ 1'b0 ;
  assign n23680 = n13880 & ~n23679 ;
  assign n23681 = x86 & n23680 ;
  assign n23682 = n3102 | n8308 ;
  assign n23683 = n13605 ^ n3537 ^ 1'b0 ;
  assign n23684 = n23682 | n23683 ;
  assign n23685 = n5937 & n14576 ;
  assign n23686 = x41 & n5626 ;
  assign n23687 = n4785 ^ n4764 ^ 1'b0 ;
  assign n23688 = n4778 & ~n17697 ;
  assign n23689 = n23688 ^ n17759 ^ 1'b0 ;
  assign n23690 = ~n7824 & n16641 ;
  assign n23691 = n4975 & n23690 ;
  assign n23692 = ( ~n2146 & n11435 ) | ( ~n2146 & n18463 ) | ( n11435 & n18463 ) ;
  assign n23693 = n7391 & ~n8464 ;
  assign n23694 = ~n12979 & n23693 ;
  assign n23695 = n1116 & ~n9048 ;
  assign n23696 = n10835 & n23695 ;
  assign n23698 = ( n1656 & n1869 ) | ( n1656 & ~n15610 ) | ( n1869 & ~n15610 ) ;
  assign n23697 = ~n9090 & n11177 ;
  assign n23699 = n23698 ^ n23697 ^ 1'b0 ;
  assign n23700 = ( n13320 & ~n19310 ) | ( n13320 & n23002 ) | ( ~n19310 & n23002 ) ;
  assign n23701 = n22220 & ~n23257 ;
  assign n23702 = ~n1888 & n3103 ;
  assign n23703 = ~n16164 & n23702 ;
  assign n23704 = n19491 ^ n2212 ^ n231 ;
  assign n23705 = ( n3413 & n23703 ) | ( n3413 & n23704 ) | ( n23703 & n23704 ) ;
  assign n23706 = n9870 | n16114 ;
  assign n23707 = n835 | n23706 ;
  assign n23708 = n10454 & ~n17463 ;
  assign n23709 = ~n4812 & n23708 ;
  assign n23714 = n10260 | n19568 ;
  assign n23710 = ~n4367 & n9323 ;
  assign n23711 = n23710 ^ n5298 ^ 1'b0 ;
  assign n23712 = n1627 & n23711 ;
  assign n23713 = n12540 & n23712 ;
  assign n23715 = n23714 ^ n23713 ^ 1'b0 ;
  assign n23716 = n20608 ^ n20373 ^ 1'b0 ;
  assign n23717 = ~n3979 & n23716 ;
  assign n23718 = n4354 & ~n6916 ;
  assign n23719 = n8347 & n23010 ;
  assign n23720 = n4116 | n4616 ;
  assign n23721 = n14021 ^ n6195 ^ 1'b0 ;
  assign n23722 = n7139 & ~n23721 ;
  assign n23723 = ( n20649 & ~n23720 ) | ( n20649 & n23722 ) | ( ~n23720 & n23722 ) ;
  assign n23725 = n5283 ^ n836 ^ 1'b0 ;
  assign n23724 = n7254 | n12902 ;
  assign n23726 = n23725 ^ n23724 ^ 1'b0 ;
  assign n23727 = ( n1374 & n7305 ) | ( n1374 & n23726 ) | ( n7305 & n23726 ) ;
  assign n23728 = n23727 ^ n8271 ^ n867 ;
  assign n23729 = n23447 ^ n10625 ^ 1'b0 ;
  assign n23730 = n6043 | n20960 ;
  assign n23731 = n23730 ^ n9171 ^ 1'b0 ;
  assign n23732 = n757 & n1718 ;
  assign n23733 = n1570 & ~n1855 ;
  assign n23734 = n23732 & n23733 ;
  assign n23735 = n3634 & ~n10424 ;
  assign n23736 = n10424 & n23735 ;
  assign n23737 = n5702 & n6051 ;
  assign n23738 = n23736 & n23737 ;
  assign n23739 = n4803 & ~n15133 ;
  assign n23740 = n10306 & n23739 ;
  assign n23741 = n5958 ^ n5179 ^ n977 ;
  assign n23742 = n12921 & n16588 ;
  assign n23743 = n23742 ^ n22021 ^ 1'b0 ;
  assign n23744 = ( n14071 & n23741 ) | ( n14071 & ~n23743 ) | ( n23741 & ~n23743 ) ;
  assign n23745 = n13907 ^ n9376 ^ 1'b0 ;
  assign n23746 = n11622 | n23745 ;
  assign n23747 = n4478 | n10111 ;
  assign n23748 = n11115 & n23747 ;
  assign n23749 = n4099 & n22584 ;
  assign n23750 = n23749 ^ n16178 ^ 1'b0 ;
  assign n23751 = ~n837 & n14773 ;
  assign n23752 = n2868 & n23751 ;
  assign n23753 = n3684 & ~n16238 ;
  assign n23754 = ( n664 & n6349 ) | ( n664 & n13264 ) | ( n6349 & n13264 ) ;
  assign n23755 = n17943 ^ n9571 ^ n6079 ;
  assign n23756 = n7705 & n13900 ;
  assign n23757 = n23756 ^ n5144 ^ 1'b0 ;
  assign n23758 = n2800 ^ n2341 ^ 1'b0 ;
  assign n23759 = n16370 & n23758 ;
  assign n23760 = n2307 | n3232 ;
  assign n23761 = n4225 | n23760 ;
  assign n23762 = n3281 & ~n5628 ;
  assign n23763 = n6676 & n11447 ;
  assign n23764 = n20713 & n23763 ;
  assign n23771 = n1069 | n15277 ;
  assign n23765 = ~n3155 & n5517 ;
  assign n23766 = n23765 ^ n3148 ^ 1'b0 ;
  assign n23767 = n23766 ^ n14533 ^ n6753 ;
  assign n23768 = n1135 | n9069 ;
  assign n23769 = n23767 | n23768 ;
  assign n23770 = ~n5243 & n23769 ;
  assign n23772 = n23771 ^ n23770 ^ 1'b0 ;
  assign n23773 = n8437 ^ n4991 ^ 1'b0 ;
  assign n23774 = ~n15970 & n17281 ;
  assign n23775 = n13184 ^ n11286 ^ n288 ;
  assign n23776 = ~n6665 & n10627 ;
  assign n23777 = ~n23775 & n23776 ;
  assign n23778 = n5780 | n15853 ;
  assign n23779 = n5304 | n11721 ;
  assign n23780 = n23779 ^ n22461 ^ 1'b0 ;
  assign n23781 = n13856 ^ n10811 ^ n8287 ;
  assign n23782 = ( ~n6784 & n7328 ) | ( ~n6784 & n11419 ) | ( n7328 & n11419 ) ;
  assign n23783 = n3245 & n8582 ;
  assign n23784 = ~n9059 & n23783 ;
  assign n23785 = n2021 | n23784 ;
  assign n23786 = n23785 ^ n8185 ^ 1'b0 ;
  assign n23787 = n11530 ^ n8667 ^ 1'b0 ;
  assign n23788 = x89 & ~n23787 ;
  assign n23789 = n1734 & n23788 ;
  assign n23790 = n23789 ^ n5594 ^ 1'b0 ;
  assign n23791 = ~n4476 & n23401 ;
  assign n23792 = n619 & ~n5712 ;
  assign n23793 = n23792 ^ n6837 ^ 1'b0 ;
  assign n23794 = n10978 ^ n7759 ^ 1'b0 ;
  assign n23795 = ~n14685 & n23794 ;
  assign n23798 = n19682 ^ n14350 ^ 1'b0 ;
  assign n23799 = n16141 | n23798 ;
  assign n23797 = n4880 | n8478 ;
  assign n23796 = ~n12531 & n13084 ;
  assign n23800 = n23799 ^ n23797 ^ n23796 ;
  assign n23801 = ~n1354 & n6543 ;
  assign n23802 = n4025 & ~n12509 ;
  assign n23803 = n23802 ^ n2564 ^ 1'b0 ;
  assign n23804 = n12814 & n23803 ;
  assign n23805 = n9182 ^ n2634 ^ 1'b0 ;
  assign n23806 = ~n8256 & n23805 ;
  assign n23807 = ~n10438 & n23806 ;
  assign n23808 = n5499 | n8991 ;
  assign n23809 = n12728 ^ n3664 ^ 1'b0 ;
  assign n23810 = n6124 & n23809 ;
  assign n23811 = n6346 | n17625 ;
  assign n23812 = n17972 ^ n17239 ^ 1'b0 ;
  assign n23813 = n15704 ^ n10668 ^ 1'b0 ;
  assign n23814 = n23812 & n23813 ;
  assign n23815 = n11452 ^ n490 ^ 1'b0 ;
  assign n23816 = ~n19749 & n23815 ;
  assign n23817 = n10195 ^ n10168 ^ 1'b0 ;
  assign n23818 = n20235 & ~n23817 ;
  assign n23819 = n5063 & n23818 ;
  assign n23820 = n23139 ^ n4757 ^ 1'b0 ;
  assign n23822 = n3216 & n12744 ;
  assign n23821 = x58 & n341 ;
  assign n23823 = n23822 ^ n23821 ^ 1'b0 ;
  assign n23824 = ( n9331 & ~n12374 ) | ( n9331 & n22656 ) | ( ~n12374 & n22656 ) ;
  assign n23825 = n20870 ^ n20230 ^ 1'b0 ;
  assign n23826 = n1200 | n23825 ;
  assign n23827 = n21253 ^ n10662 ^ 1'b0 ;
  assign n23828 = n7619 & ~n22205 ;
  assign n23829 = n23828 ^ n7810 ^ n6000 ;
  assign n23830 = n23465 ^ n5212 ^ 1'b0 ;
  assign n23831 = n5295 ^ n3666 ^ 1'b0 ;
  assign n23832 = n5715 & n12309 ;
  assign n23833 = ( n3972 & ~n18121 ) | ( n3972 & n23832 ) | ( ~n18121 & n23832 ) ;
  assign n23834 = n23831 | n23833 ;
  assign n23835 = n6362 ^ n4502 ^ 1'b0 ;
  assign n23836 = n6760 | n23835 ;
  assign n23837 = ( n8833 & ~n9366 ) | ( n8833 & n23836 ) | ( ~n9366 & n23836 ) ;
  assign n23838 = n14030 & n23837 ;
  assign n23839 = n19933 & n23838 ;
  assign n23840 = ~n22542 & n23839 ;
  assign n23841 = n2577 & ~n11553 ;
  assign n23842 = ~n7697 & n23841 ;
  assign n23843 = ( n607 & n7219 ) | ( n607 & n14972 ) | ( n7219 & n14972 ) ;
  assign n23844 = x108 & ~n7497 ;
  assign n23845 = ( n3640 & n6771 ) | ( n3640 & ~n23844 ) | ( n6771 & ~n23844 ) ;
  assign n23846 = n14817 & ~n22651 ;
  assign n23847 = n23846 ^ n9971 ^ 1'b0 ;
  assign n23848 = x16 & n1499 ;
  assign n23849 = n23848 ^ n23612 ^ 1'b0 ;
  assign n23850 = n17896 ^ n801 ^ 1'b0 ;
  assign n23851 = n6689 | n23850 ;
  assign n23852 = n15555 & ~n21521 ;
  assign n23853 = n17230 ^ n6090 ^ 1'b0 ;
  assign n23854 = n651 | n23853 ;
  assign n23855 = n23854 ^ n14107 ^ n12927 ;
  assign n23856 = n18228 | n20508 ;
  assign n23857 = n23856 ^ n8667 ^ n7234 ;
  assign n23858 = n8652 ^ n471 ^ 1'b0 ;
  assign n23859 = n23858 ^ n7516 ^ 1'b0 ;
  assign n23860 = n5475 ^ n3304 ^ n2972 ;
  assign n23861 = n23860 ^ n5952 ^ 1'b0 ;
  assign n23862 = n20327 ^ n4663 ^ n4520 ;
  assign n23863 = n23862 ^ n16235 ^ n13374 ;
  assign n23873 = n1387 & ~n1421 ;
  assign n23870 = n718 | n2607 ;
  assign n23871 = n10308 | n23870 ;
  assign n23872 = ( n10761 & ~n23645 ) | ( n10761 & n23871 ) | ( ~n23645 & n23871 ) ;
  assign n23874 = n23873 ^ n23872 ^ n2779 ;
  assign n23875 = ( n299 & ~n8830 ) | ( n299 & n23874 ) | ( ~n8830 & n23874 ) ;
  assign n23868 = n9450 ^ n3014 ^ 1'b0 ;
  assign n23869 = n23868 ^ n10873 ^ n2825 ;
  assign n23864 = n5006 & ~n8835 ;
  assign n23865 = n4239 & ~n8730 ;
  assign n23866 = n22335 & n23865 ;
  assign n23867 = n23864 & n23866 ;
  assign n23876 = n23875 ^ n23869 ^ n23867 ;
  assign n23887 = n1244 & n1669 ;
  assign n23888 = ~n1244 & n23887 ;
  assign n23889 = ~x110 & n23888 ;
  assign n23877 = ~n2417 & n12360 ;
  assign n23878 = n2417 & n23877 ;
  assign n23879 = n11298 & ~n23878 ;
  assign n23880 = n23878 & n23879 ;
  assign n23881 = n3012 | n4650 ;
  assign n23882 = n23881 ^ n12482 ^ 1'b0 ;
  assign n23883 = n23880 & n23882 ;
  assign n23884 = n7582 ^ n7031 ^ 1'b0 ;
  assign n23885 = n674 & ~n23884 ;
  assign n23886 = ~n23883 & n23885 ;
  assign n23890 = n23889 ^ n23886 ^ 1'b0 ;
  assign n23891 = x20 | n23890 ;
  assign n23892 = n2429 & ~n23891 ;
  assign n23893 = n13215 & n23892 ;
  assign n23894 = n10634 | n15752 ;
  assign n23895 = n23894 ^ n4291 ^ 1'b0 ;
  assign n23896 = n15328 & ~n15347 ;
  assign n23897 = ~n10906 & n23896 ;
  assign n23899 = n4610 & ~n9096 ;
  assign n23900 = n9403 & n23899 ;
  assign n23901 = ~n467 & n13903 ;
  assign n23902 = ~n23900 & n23901 ;
  assign n23898 = n858 & n1034 ;
  assign n23903 = n23902 ^ n23898 ^ n1140 ;
  assign n23904 = ( n11631 & ~n13012 ) | ( n11631 & n18773 ) | ( ~n13012 & n18773 ) ;
  assign n23905 = n18095 & n22837 ;
  assign n23906 = n15306 ^ n909 ^ 1'b0 ;
  assign n23907 = ~n13128 & n23906 ;
  assign n23908 = n4289 & ~n10922 ;
  assign n23909 = ~n23907 & n23908 ;
  assign n23910 = n21599 ^ n5673 ^ 1'b0 ;
  assign n23911 = ~n5077 & n9008 ;
  assign n23912 = n23911 ^ n17020 ^ 1'b0 ;
  assign n23913 = n5012 & n23912 ;
  assign n23914 = ~n7255 & n8222 ;
  assign n23915 = n23914 ^ n2634 ^ 1'b0 ;
  assign n23916 = n12559 ^ n5412 ^ 1'b0 ;
  assign n23917 = n9910 & ~n23916 ;
  assign n23918 = n23917 ^ n14550 ^ 1'b0 ;
  assign n23919 = n273 ^ x84 ^ 1'b0 ;
  assign n23920 = n23919 ^ n15034 ^ 1'b0 ;
  assign n23921 = n1053 & n14374 ;
  assign n23922 = ~n23920 & n23921 ;
  assign n23923 = n16141 ^ n2935 ^ 1'b0 ;
  assign n23924 = ~n10379 & n23923 ;
  assign n23925 = n23924 ^ n11196 ^ 1'b0 ;
  assign n23926 = ( n5681 & n23922 ) | ( n5681 & ~n23925 ) | ( n23922 & ~n23925 ) ;
  assign n23927 = n3268 | n9758 ;
  assign n23928 = n23927 ^ n10396 ^ 1'b0 ;
  assign n23929 = n1300 | n13567 ;
  assign n23930 = n720 & n3701 ;
  assign n23931 = n21287 | n23930 ;
  assign n23933 = n11768 ^ n8492 ^ n7323 ;
  assign n23934 = n13240 & n23933 ;
  assign n23932 = ~n16354 & n20841 ;
  assign n23935 = n23934 ^ n23932 ^ 1'b0 ;
  assign n23936 = n5883 ^ n5760 ^ 1'b0 ;
  assign n23937 = n3354 & ~n23936 ;
  assign n23938 = n23937 ^ n17167 ^ 1'b0 ;
  assign n23939 = n8499 ^ n1430 ^ 1'b0 ;
  assign n23940 = n16052 | n23939 ;
  assign n23941 = ~n6691 & n23940 ;
  assign n23942 = n2970 & n23941 ;
  assign n23943 = n1040 & n9981 ;
  assign n23944 = n6600 ^ n3525 ^ 1'b0 ;
  assign n23945 = n20741 ^ n9243 ^ 1'b0 ;
  assign n23946 = n20592 ^ n3552 ^ 1'b0 ;
  assign n23947 = n21373 & ~n23946 ;
  assign n23948 = n12180 ^ n6385 ^ 1'b0 ;
  assign n23949 = ~n14719 & n23948 ;
  assign n23951 = n1670 & n1861 ;
  assign n23950 = ( n8933 & n13706 ) | ( n8933 & n16818 ) | ( n13706 & n16818 ) ;
  assign n23952 = n23951 ^ n23950 ^ 1'b0 ;
  assign n23953 = n23952 ^ n1819 ^ 1'b0 ;
  assign n23954 = n23355 ^ n3903 ^ 1'b0 ;
  assign n23956 = ( n6966 & n15783 ) | ( n6966 & n17543 ) | ( n15783 & n17543 ) ;
  assign n23955 = x51 | n21066 ;
  assign n23957 = n23956 ^ n23955 ^ n6198 ;
  assign n23958 = n3386 ^ n2339 ^ 1'b0 ;
  assign n23959 = n23958 ^ n12079 ^ 1'b0 ;
  assign n23960 = n7075 | n23959 ;
  assign n23961 = n8979 & n23960 ;
  assign n23962 = ~n9811 & n20704 ;
  assign n23963 = n23962 ^ n15116 ^ 1'b0 ;
  assign n23964 = ( n469 & n933 ) | ( n469 & n15498 ) | ( n933 & n15498 ) ;
  assign n23965 = n23964 ^ n19078 ^ 1'b0 ;
  assign n23966 = ~n6644 & n23965 ;
  assign n23968 = ~n10460 & n19328 ;
  assign n23969 = n10610 & n23968 ;
  assign n23967 = n4317 | n22514 ;
  assign n23970 = n23969 ^ n23967 ^ 1'b0 ;
  assign n23971 = n779 & n3265 ;
  assign n23972 = ~n10234 & n23971 ;
  assign n23973 = n15058 | n19918 ;
  assign n23974 = n23972 & ~n23973 ;
  assign n23975 = n17010 ^ n4664 ^ 1'b0 ;
  assign n23976 = n2103 & ~n23975 ;
  assign n23977 = n23976 ^ n17374 ^ n7604 ;
  assign n23978 = ~n11114 & n14098 ;
  assign n23980 = n17699 ^ n9333 ^ 1'b0 ;
  assign n23979 = n3834 & n4253 ;
  assign n23981 = n23980 ^ n23979 ^ x92 ;
  assign n23982 = ~n12734 & n20283 ;
  assign n23983 = n23982 ^ n16407 ^ 1'b0 ;
  assign n23984 = n508 | n1171 ;
  assign n23985 = n22901 & ~n23984 ;
  assign n23986 = n4966 & ~n14458 ;
  assign n23987 = n938 & n23986 ;
  assign n23988 = ~x114 & n16088 ;
  assign n23989 = n6171 & n23988 ;
  assign n23990 = n13095 ^ n6876 ^ 1'b0 ;
  assign n23991 = n7042 ^ n1027 ^ 1'b0 ;
  assign n23992 = ~n6431 & n23991 ;
  assign n23993 = ( n7691 & ~n9206 ) | ( n7691 & n23992 ) | ( ~n9206 & n23992 ) ;
  assign n23994 = n9037 ^ n4859 ^ 1'b0 ;
  assign n23995 = n23994 ^ n3546 ^ 1'b0 ;
  assign n23996 = n3158 | n18186 ;
  assign n23997 = n6431 & n12437 ;
  assign n23998 = n23997 ^ n4474 ^ 1'b0 ;
  assign n23999 = n19993 | n23998 ;
  assign n24000 = n9271 | n14690 ;
  assign n24001 = n5326 | n24000 ;
  assign n24002 = n1462 & ~n6707 ;
  assign n24003 = n24002 ^ n19614 ^ 1'b0 ;
  assign n24004 = n3254 ^ x91 ^ 1'b0 ;
  assign n24005 = n5981 & n7167 ;
  assign n24006 = n24005 ^ n867 ^ 1'b0 ;
  assign n24007 = n8313 & n24006 ;
  assign n24008 = n17888 ^ n11309 ^ n2355 ;
  assign n24009 = n24008 ^ n18736 ^ n13576 ;
  assign n24010 = ~n6295 & n9985 ;
  assign n24015 = n4601 | n20700 ;
  assign n24011 = ~n5096 & n11159 ;
  assign n24012 = n24011 ^ n6399 ^ 1'b0 ;
  assign n24013 = n4018 & ~n24012 ;
  assign n24014 = n4214 & n24013 ;
  assign n24016 = n24015 ^ n24014 ^ 1'b0 ;
  assign n24017 = n3057 | n7845 ;
  assign n24018 = n12011 ^ n8819 ^ 1'b0 ;
  assign n24019 = n24017 | n24018 ;
  assign n24020 = n13816 ^ n11552 ^ n4787 ;
  assign n24021 = n19744 & n24020 ;
  assign n24022 = n4470 | n8769 ;
  assign n24023 = n17543 ^ n8931 ^ 1'b0 ;
  assign n24024 = ~n14928 & n24023 ;
  assign n24025 = ( n2677 & n4757 ) | ( n2677 & ~n9941 ) | ( n4757 & ~n9941 ) ;
  assign n24026 = n2322 ^ n2219 ^ 1'b0 ;
  assign n24027 = ( ~n16083 & n19771 ) | ( ~n16083 & n24026 ) | ( n19771 & n24026 ) ;
  assign n24029 = n22368 ^ n12512 ^ 1'b0 ;
  assign n24028 = n16025 ^ n3554 ^ 1'b0 ;
  assign n24030 = n24029 ^ n24028 ^ n8164 ;
  assign n24031 = n18121 | n19591 ;
  assign n24032 = n24031 ^ n8120 ^ 1'b0 ;
  assign n24033 = n21099 ^ n17791 ^ 1'b0 ;
  assign n24034 = n7799 ^ n2102 ^ n1649 ;
  assign n24035 = n4223 ^ n1950 ^ 1'b0 ;
  assign n24036 = n24035 ^ n9917 ^ n1033 ;
  assign n24037 = ~n1165 & n24036 ;
  assign n24038 = n5722 ^ n5638 ^ n1266 ;
  assign n24039 = ~n12205 & n23837 ;
  assign n24040 = n5695 & n24039 ;
  assign n24041 = n3856 | n16329 ;
  assign n24042 = n381 & n15622 ;
  assign n24043 = n425 & n9969 ;
  assign n24044 = n12397 ^ n10941 ^ 1'b0 ;
  assign n24045 = n21688 ^ n2554 ^ 1'b0 ;
  assign n24046 = n18269 & n24045 ;
  assign n24047 = n7473 ^ n4832 ^ 1'b0 ;
  assign n24048 = n15581 ^ n4576 ^ 1'b0 ;
  assign n24049 = ( n12197 & n24047 ) | ( n12197 & n24048 ) | ( n24047 & n24048 ) ;
  assign n24050 = n15432 ^ n4714 ^ 1'b0 ;
  assign n24051 = n10251 & ~n24050 ;
  assign n24052 = ~n10184 & n24051 ;
  assign n24053 = n24052 ^ n12588 ^ 1'b0 ;
  assign n24054 = ~n2272 & n24053 ;
  assign n24055 = n8965 & n24054 ;
  assign n24056 = n14598 ^ n1195 ^ 1'b0 ;
  assign n24057 = n14567 ^ n5739 ^ 1'b0 ;
  assign n24058 = ~n21743 & n24057 ;
  assign n24059 = ~n628 & n8162 ;
  assign n24060 = n24059 ^ n1462 ^ 1'b0 ;
  assign n24061 = n20949 ^ n11274 ^ n7069 ;
  assign n24062 = n6363 ^ n5531 ^ 1'b0 ;
  assign n24063 = n12968 | n14879 ;
  assign n24064 = ~n13829 & n13910 ;
  assign n24065 = n24064 ^ n16817 ^ 1'b0 ;
  assign n24066 = ~n5991 & n13630 ;
  assign n24067 = n18226 & n24066 ;
  assign n24068 = n177 | n13711 ;
  assign n24069 = n24068 ^ n11096 ^ 1'b0 ;
  assign n24070 = ~n293 & n2800 ;
  assign n24071 = n8080 | n8536 ;
  assign n24072 = n24071 ^ n22640 ^ n2035 ;
  assign n24073 = n18498 | n24072 ;
  assign n24074 = n7442 | n24073 ;
  assign n24075 = n5263 & ~n24074 ;
  assign n24076 = n11017 ^ n4564 ^ n661 ;
  assign n24077 = ( n8478 & n15803 ) | ( n8478 & n24076 ) | ( n15803 & n24076 ) ;
  assign n24078 = ( x16 & ~n2436 ) | ( x16 & n14813 ) | ( ~n2436 & n14813 ) ;
  assign n24079 = n301 | n10259 ;
  assign n24080 = ~n2509 & n7999 ;
  assign n24081 = n24080 ^ n4650 ^ 1'b0 ;
  assign n24082 = n1042 ^ x57 ^ 1'b0 ;
  assign n24083 = n24048 ^ n22574 ^ 1'b0 ;
  assign n24084 = n11647 & n24083 ;
  assign n24085 = ~n2825 & n24084 ;
  assign n24086 = n24085 ^ n5463 ^ 1'b0 ;
  assign n24087 = n7093 | n24086 ;
  assign n24088 = n24082 & ~n24087 ;
  assign n24089 = n1040 & n7891 ;
  assign n24090 = n24089 ^ n20288 ^ n4683 ;
  assign n24091 = n9263 & n24090 ;
  assign n24092 = ~n4662 & n10138 ;
  assign n24093 = n1321 & ~n20501 ;
  assign n24094 = n1514 & n24093 ;
  assign n24095 = n1565 & n9440 ;
  assign n24096 = n24095 ^ n3528 ^ 1'b0 ;
  assign n24097 = ( n256 & n3494 ) | ( n256 & ~n3994 ) | ( n3494 & ~n3994 ) ;
  assign n24098 = n5293 | n24097 ;
  assign n24099 = n24098 ^ n9709 ^ 1'b0 ;
  assign n24100 = n6908 & ~n9107 ;
  assign n24101 = n9107 & n24100 ;
  assign n24102 = n8422 | n24101 ;
  assign n24103 = n8422 & ~n24102 ;
  assign n24104 = n6435 ^ n640 ^ 1'b0 ;
  assign n24105 = ( n14439 & n24103 ) | ( n14439 & ~n24104 ) | ( n24103 & ~n24104 ) ;
  assign n24106 = n14978 & ~n21349 ;
  assign n24107 = n20482 ^ n15351 ^ 1'b0 ;
  assign n24109 = n14618 ^ n1092 ^ 1'b0 ;
  assign n24110 = n3269 & ~n24109 ;
  assign n24108 = n9364 & n16961 ;
  assign n24111 = n24110 ^ n24108 ^ 1'b0 ;
  assign n24112 = n830 | n5492 ;
  assign n24113 = n12445 & ~n24112 ;
  assign n24114 = n4904 & n8390 ;
  assign n24115 = n24114 ^ n6678 ^ 1'b0 ;
  assign n24116 = n12592 ^ n6815 ^ 1'b0 ;
  assign n24117 = n24115 & n24116 ;
  assign n24118 = n7092 | n7347 ;
  assign n24119 = n2112 | n20811 ;
  assign n24120 = n5096 & ~n24119 ;
  assign n24121 = n24120 ^ n15865 ^ 1'b0 ;
  assign n24122 = ( ~n13578 & n24118 ) | ( ~n13578 & n24121 ) | ( n24118 & n24121 ) ;
  assign n24123 = n23295 ^ n17303 ^ n8158 ;
  assign n24125 = n1033 | n18351 ;
  assign n24126 = n12858 ^ n9964 ^ 1'b0 ;
  assign n24127 = n24125 & ~n24126 ;
  assign n24124 = ~n8682 & n21145 ;
  assign n24128 = n24127 ^ n24124 ^ 1'b0 ;
  assign n24129 = n865 | n3113 ;
  assign n24130 = n13439 ^ n10515 ^ 1'b0 ;
  assign n24131 = n24130 ^ n20165 ^ 1'b0 ;
  assign n24132 = ~n24129 & n24131 ;
  assign n24133 = n14129 & n24132 ;
  assign n24134 = n7845 & n14105 ;
  assign n24135 = n11085 | n13414 ;
  assign n24136 = n24135 ^ n22770 ^ n13467 ;
  assign n24138 = n9979 ^ n3195 ^ 1'b0 ;
  assign n24137 = n13891 ^ n2166 ^ x6 ;
  assign n24139 = n24138 ^ n24137 ^ n21822 ;
  assign n24141 = n12983 ^ n9830 ^ 1'b0 ;
  assign n24142 = n6982 & ~n24141 ;
  assign n24140 = n7161 | n9635 ;
  assign n24143 = n24142 ^ n24140 ^ 1'b0 ;
  assign n24144 = n3135 & n19615 ;
  assign n24145 = n24144 ^ n19161 ^ 1'b0 ;
  assign n24146 = n671 & ~n8198 ;
  assign n24147 = ~n9761 & n24146 ;
  assign n24148 = n10519 ^ n9282 ^ 1'b0 ;
  assign n24150 = ( ~n819 & n6581 ) | ( ~n819 & n10927 ) | ( n6581 & n10927 ) ;
  assign n24149 = ~n8887 & n9540 ;
  assign n24151 = n24150 ^ n24149 ^ 1'b0 ;
  assign n24152 = n8776 ^ n6885 ^ 1'b0 ;
  assign n24153 = n4019 & n24152 ;
  assign n24154 = n3791 & n13208 ;
  assign n24155 = n7953 & ~n24154 ;
  assign n24156 = n24155 ^ x13 ^ 1'b0 ;
  assign n24157 = n6992 ^ n1295 ^ 1'b0 ;
  assign n24158 = n19777 ^ n16400 ^ 1'b0 ;
  assign n24159 = ~n4664 & n17774 ;
  assign n24160 = n5797 ^ n4435 ^ 1'b0 ;
  assign n24161 = n19280 & ~n24160 ;
  assign n24162 = n12661 ^ n8823 ^ 1'b0 ;
  assign n24163 = n24162 ^ n15126 ^ 1'b0 ;
  assign n24164 = n8836 | n24163 ;
  assign n24165 = n7187 | n9516 ;
  assign n24166 = n12987 | n24165 ;
  assign n24167 = n22721 ^ n11630 ^ 1'b0 ;
  assign n24168 = n3853 & n9843 ;
  assign n24169 = ~x110 & n24168 ;
  assign n24170 = n24169 ^ n5231 ^ 1'b0 ;
  assign n24171 = n13615 & ~n24170 ;
  assign n24172 = ( n1730 & n4351 ) | ( n1730 & ~n10623 ) | ( n4351 & ~n10623 ) ;
  assign n24173 = n12043 ^ n361 ^ 1'b0 ;
  assign n24174 = n24172 | n24173 ;
  assign n24175 = ( n17084 & ~n24171 ) | ( n17084 & n24174 ) | ( ~n24171 & n24174 ) ;
  assign n24176 = n9062 & n16472 ;
  assign n24177 = ~n2702 & n22992 ;
  assign n24178 = ( ~n4589 & n7969 ) | ( ~n4589 & n24177 ) | ( n7969 & n24177 ) ;
  assign n24179 = n13943 ^ n11708 ^ n707 ;
  assign n24180 = ~n381 & n4184 ;
  assign n24181 = n24180 ^ n12660 ^ 1'b0 ;
  assign n24182 = n24181 ^ n4419 ^ 1'b0 ;
  assign n24183 = ~n1594 & n24182 ;
  assign n24184 = n12120 | n24183 ;
  assign n24185 = n24184 ^ n245 ^ 1'b0 ;
  assign n24186 = n929 & n15848 ;
  assign n24187 = n24186 ^ n6759 ^ 1'b0 ;
  assign n24188 = n12464 | n24187 ;
  assign n24189 = n19683 ^ n16901 ^ 1'b0 ;
  assign n24190 = n24188 | n24189 ;
  assign n24191 = n4903 & ~n10860 ;
  assign n24192 = n10500 & ~n12916 ;
  assign n24193 = n8139 ^ n305 ^ 1'b0 ;
  assign n24194 = n24192 & n24193 ;
  assign n24195 = n24191 & n24194 ;
  assign n24196 = n6977 | n19898 ;
  assign n24197 = ( ~n8733 & n15983 ) | ( ~n8733 & n24196 ) | ( n15983 & n24196 ) ;
  assign n24198 = ~n2751 & n15714 ;
  assign n24199 = ~n19538 & n24198 ;
  assign n24200 = n20689 | n24199 ;
  assign n24201 = n7083 & ~n15048 ;
  assign n24202 = n24201 ^ n16422 ^ 1'b0 ;
  assign n24203 = n24202 ^ n15112 ^ n3792 ;
  assign n24204 = n17805 ^ n8504 ^ 1'b0 ;
  assign n24205 = ~n5093 & n17701 ;
  assign n24206 = ~n2317 & n24205 ;
  assign n24207 = n24206 ^ n5661 ^ 1'b0 ;
  assign n24208 = n9209 ^ n2390 ^ n1016 ;
  assign n24209 = n21305 & n24208 ;
  assign n24211 = ~n11748 & n17977 ;
  assign n24212 = n24211 ^ n19400 ^ 1'b0 ;
  assign n24210 = ~n12239 & n23508 ;
  assign n24213 = n24212 ^ n24210 ^ 1'b0 ;
  assign n24214 = ( n8204 & ~n24209 ) | ( n8204 & n24213 ) | ( ~n24209 & n24213 ) ;
  assign n24215 = n13550 | n18650 ;
  assign n24216 = n4246 ^ n3243 ^ 1'b0 ;
  assign n24217 = n1849 ^ n1040 ^ n603 ;
  assign n24218 = n10704 ^ n7245 ^ 1'b0 ;
  assign n24219 = n8530 ^ n5968 ^ n1520 ;
  assign n24220 = n6759 ^ n2225 ^ 1'b0 ;
  assign n24221 = ~n8767 & n24220 ;
  assign n24222 = n7189 & ~n24221 ;
  assign n24223 = n24222 ^ n8730 ^ 1'b0 ;
  assign n24224 = n24219 & n24223 ;
  assign n24225 = ( ~n2510 & n4770 ) | ( ~n2510 & n8230 ) | ( n4770 & n8230 ) ;
  assign n24226 = n5369 | n24225 ;
  assign n24227 = n893 & n23153 ;
  assign n24228 = n3959 & n18338 ;
  assign n24229 = n7328 & ~n9464 ;
  assign n24230 = n1438 | n13047 ;
  assign n24231 = n24229 | n24230 ;
  assign n24232 = ~n16994 & n24231 ;
  assign n24233 = n4044 | n15806 ;
  assign n24234 = n6845 & ~n21756 ;
  assign n24235 = n24234 ^ n11669 ^ 1'b0 ;
  assign n24236 = n17409 & n24235 ;
  assign n24237 = ~n24233 & n24236 ;
  assign n24238 = n19599 ^ n7251 ^ n817 ;
  assign n24239 = n18879 ^ n14285 ^ 1'b0 ;
  assign n24240 = ~n24238 & n24239 ;
  assign n24241 = n19590 ^ n14197 ^ 1'b0 ;
  assign n24242 = ~n18394 & n24241 ;
  assign n24243 = ~n4306 & n24242 ;
  assign n24244 = n2061 | n11028 ;
  assign n24245 = n24244 ^ n13703 ^ 1'b0 ;
  assign n24246 = n24245 ^ n2464 ^ 1'b0 ;
  assign n24247 = ( ~n3831 & n3958 ) | ( ~n3831 & n4469 ) | ( n3958 & n4469 ) ;
  assign n24248 = ~n702 & n9062 ;
  assign n24249 = n1440 & n24248 ;
  assign n24250 = n21949 | n24249 ;
  assign n24251 = n24247 & ~n24250 ;
  assign n24252 = n1021 & n5938 ;
  assign n24253 = n24252 ^ n145 ^ 1'b0 ;
  assign n24254 = n15913 & n24253 ;
  assign n24255 = n13604 ^ n7606 ^ 1'b0 ;
  assign n24256 = n7189 | n24255 ;
  assign n24257 = n24256 ^ n23442 ^ 1'b0 ;
  assign n24258 = n4029 & n24257 ;
  assign n24259 = n24258 ^ n17519 ^ 1'b0 ;
  assign n24260 = ~n2868 & n5730 ;
  assign n24261 = n8567 & n24260 ;
  assign n24262 = n7258 | n20396 ;
  assign n24263 = n285 & n20066 ;
  assign n24264 = n24262 & n24263 ;
  assign n24265 = n10761 ^ n2090 ^ 1'b0 ;
  assign n24266 = n1036 & n24265 ;
  assign n24267 = n19557 | n24266 ;
  assign n24268 = n11187 & ~n13076 ;
  assign n24269 = n17356 & n24268 ;
  assign n24270 = n4233 | n5613 ;
  assign n24271 = n24270 ^ n20811 ^ 1'b0 ;
  assign n24272 = n14210 ^ n551 ^ 1'b0 ;
  assign n24273 = n7439 ^ n3538 ^ 1'b0 ;
  assign n24274 = ~n17399 & n21846 ;
  assign n24275 = n24273 & n24274 ;
  assign n24276 = ~n18920 & n20710 ;
  assign n24277 = n24276 ^ n9203 ^ 1'b0 ;
  assign n24278 = n16548 ^ n6497 ^ n3939 ;
  assign n24279 = ( n6709 & ~n12205 ) | ( n6709 & n19693 ) | ( ~n12205 & n19693 ) ;
  assign n24280 = n8038 & n22721 ;
  assign n24281 = n24280 ^ n2032 ^ 1'b0 ;
  assign n24282 = n4042 ^ n815 ^ 1'b0 ;
  assign n24283 = n20966 ^ n997 ^ 1'b0 ;
  assign n24285 = n5257 & n16548 ;
  assign n24284 = n15607 & n16374 ;
  assign n24286 = n24285 ^ n24284 ^ 1'b0 ;
  assign n24287 = n16894 ^ n9094 ^ 1'b0 ;
  assign n24288 = n11628 & n24287 ;
  assign n24289 = n7425 & ~n8158 ;
  assign n24290 = n5862 | n17597 ;
  assign n24291 = ( n791 & n4618 ) | ( n791 & n24290 ) | ( n4618 & n24290 ) ;
  assign n24292 = n4222 & n8480 ;
  assign n24293 = n6474 ^ n5400 ^ 1'b0 ;
  assign n24294 = ~n2011 & n24293 ;
  assign n24295 = ~n20724 & n24294 ;
  assign n24296 = n24295 ^ n9182 ^ 1'b0 ;
  assign n24297 = n4108 | n15458 ;
  assign n24298 = n3391 & n5544 ;
  assign n24299 = n21808 ^ n2591 ^ 1'b0 ;
  assign n24300 = n3000 | n24299 ;
  assign n24301 = n24298 & ~n24300 ;
  assign n24302 = n6239 & ~n8900 ;
  assign n24303 = n24302 ^ n6563 ^ n1109 ;
  assign n24304 = n19491 ^ n5357 ^ 1'b0 ;
  assign n24305 = n1860 & ~n19148 ;
  assign n24306 = n24305 ^ n19336 ^ 1'b0 ;
  assign n24307 = n7488 ^ n3235 ^ 1'b0 ;
  assign n24308 = n13969 & ~n24307 ;
  assign n24309 = n11751 & n24308 ;
  assign n24310 = n24309 ^ n502 ^ 1'b0 ;
  assign n24311 = ~n16982 & n20427 ;
  assign n24312 = n24311 ^ n21094 ^ 1'b0 ;
  assign n24313 = n20775 ^ n12830 ^ 1'b0 ;
  assign n24314 = n5271 | n24313 ;
  assign n24315 = n4490 & ~n24314 ;
  assign n24316 = n14054 ^ n312 ^ 1'b0 ;
  assign n24317 = x93 & ~n290 ;
  assign n24318 = n24317 ^ n4420 ^ 1'b0 ;
  assign n24319 = ~n206 & n1643 ;
  assign n24320 = n13671 ^ n4860 ^ n2104 ;
  assign n24321 = n24320 ^ n17579 ^ n13732 ;
  assign n24322 = ( n801 & n6526 ) | ( n801 & n12588 ) | ( n6526 & n12588 ) ;
  assign n24323 = ~n8055 & n24322 ;
  assign n24324 = n24323 ^ n23080 ^ 1'b0 ;
  assign n24325 = n14552 ^ n10617 ^ 1'b0 ;
  assign n24326 = n23543 ^ n12940 ^ 1'b0 ;
  assign n24327 = n24325 | n24326 ;
  assign n24328 = n7057 | n24327 ;
  assign n24329 = n12695 ^ n2077 ^ 1'b0 ;
  assign n24330 = ~n20629 & n24329 ;
  assign n24331 = n9612 | n21599 ;
  assign n24332 = n6184 | n24331 ;
  assign n24333 = n2355 & n9450 ;
  assign n24334 = n20128 | n24333 ;
  assign n24335 = n17044 & ~n21168 ;
  assign n24336 = n24335 ^ n7999 ^ 1'b0 ;
  assign n24337 = n24336 ^ n16984 ^ n555 ;
  assign n24338 = n24337 ^ n23111 ^ 1'b0 ;
  assign n24339 = n22079 ^ n1476 ^ 1'b0 ;
  assign n24340 = n3456 | n24339 ;
  assign n24341 = n5790 & ~n23564 ;
  assign n24342 = n3741 & n24341 ;
  assign n24343 = ~n8519 & n13512 ;
  assign n24344 = n20682 ^ n8030 ^ 1'b0 ;
  assign n24345 = n623 | n24344 ;
  assign n24346 = n7723 & n24345 ;
  assign n24347 = ~n11567 & n17055 ;
  assign n24348 = n24347 ^ n15568 ^ 1'b0 ;
  assign n24349 = x31 & n7142 ;
  assign n24350 = n15879 & n24349 ;
  assign n24351 = n21981 ^ n14274 ^ 1'b0 ;
  assign n24352 = ~n24350 & n24351 ;
  assign n24353 = n1507 & n6359 ;
  assign n24354 = n4632 | n22710 ;
  assign n24355 = n24354 ^ n5719 ^ 1'b0 ;
  assign n24356 = ( n18645 & ~n19748 ) | ( n18645 & n24355 ) | ( ~n19748 & n24355 ) ;
  assign n24357 = n19317 ^ n2595 ^ 1'b0 ;
  assign n24358 = ~n5662 & n24357 ;
  assign n24359 = n1086 & n24358 ;
  assign n24361 = n2208 ^ n1407 ^ 1'b0 ;
  assign n24362 = n24361 ^ n1248 ^ 1'b0 ;
  assign n24363 = ~n1399 & n24362 ;
  assign n24364 = n24363 ^ n9662 ^ 1'b0 ;
  assign n24360 = n319 | n9463 ;
  assign n24365 = n24364 ^ n24360 ^ 1'b0 ;
  assign n24366 = ~n10658 & n17528 ;
  assign n24367 = n15440 ^ n667 ^ 1'b0 ;
  assign n24368 = n6034 | n24367 ;
  assign n24369 = n24368 ^ n1307 ^ 1'b0 ;
  assign n24370 = n24369 ^ n20120 ^ 1'b0 ;
  assign n24371 = n6518 & n11796 ;
  assign n24372 = n19033 ^ n1323 ^ 1'b0 ;
  assign n24373 = n17775 | n24372 ;
  assign n24374 = n16256 ^ n2829 ^ 1'b0 ;
  assign n24375 = n24373 & ~n24374 ;
  assign n24376 = ~n2996 & n16041 ;
  assign n24377 = ~n21639 & n24376 ;
  assign n24378 = n24377 ^ n4727 ^ 1'b0 ;
  assign n24379 = n6570 | n15332 ;
  assign n24380 = n23946 ^ n2921 ^ 1'b0 ;
  assign n24381 = ( n8185 & n24379 ) | ( n8185 & n24380 ) | ( n24379 & n24380 ) ;
  assign n24382 = n5722 ^ n5476 ^ 1'b0 ;
  assign n24383 = n13448 & ~n24382 ;
  assign n24384 = n8220 & ~n11575 ;
  assign n24385 = n3684 & n8499 ;
  assign n24386 = n24384 & n24385 ;
  assign n24387 = n7032 | n18101 ;
  assign n24388 = ( n3997 & n8748 ) | ( n3997 & ~n11088 ) | ( n8748 & ~n11088 ) ;
  assign n24392 = n150 & n151 ;
  assign n24389 = ( n4560 & ~n12877 ) | ( n4560 & n15711 ) | ( ~n12877 & n15711 ) ;
  assign n24390 = n24389 ^ n8999 ^ 1'b0 ;
  assign n24391 = n12328 & ~n24390 ;
  assign n24393 = n24392 ^ n24391 ^ n6657 ;
  assign n24394 = ~n4900 & n14058 ;
  assign n24395 = n22774 ^ n21915 ^ n2192 ;
  assign n24396 = n3955 & ~n24395 ;
  assign n24397 = n467 & n14470 ;
  assign n24398 = n24397 ^ n9090 ^ 1'b0 ;
  assign n24399 = n16984 ^ n2146 ^ 1'b0 ;
  assign n24400 = n24399 ^ n13803 ^ n2472 ;
  assign n24401 = n9400 & ~n10317 ;
  assign n24402 = n9326 ^ n5544 ^ 1'b0 ;
  assign n24403 = n9307 & n24402 ;
  assign n24404 = n19370 ^ n13504 ^ 1'b0 ;
  assign n24405 = n24403 & ~n24404 ;
  assign n24406 = n7217 & ~n11945 ;
  assign n24407 = ~n9896 & n15177 ;
  assign n24408 = n24407 ^ n967 ^ 1'b0 ;
  assign n24409 = n5244 & n15269 ;
  assign n24410 = ~n24408 & n24409 ;
  assign n24411 = n5567 | n10618 ;
  assign n24412 = n16830 ^ n13993 ^ 1'b0 ;
  assign n24413 = n4059 & n24412 ;
  assign n24414 = n20833 ^ n4167 ^ 1'b0 ;
  assign n24415 = n24414 ^ n6933 ^ n1364 ;
  assign n24416 = n9065 ^ n7458 ^ 1'b0 ;
  assign n24417 = n8298 & n24416 ;
  assign n24418 = n1613 | n24417 ;
  assign n24419 = n10277 & ~n11389 ;
  assign n24420 = n24419 ^ n21838 ^ 1'b0 ;
  assign n24421 = ( n1985 & ~n24418 ) | ( n1985 & n24420 ) | ( ~n24418 & n24420 ) ;
  assign n24422 = n17626 ^ n8733 ^ 1'b0 ;
  assign n24423 = n10563 & ~n24422 ;
  assign n24424 = ~n16318 & n20833 ;
  assign n24425 = n2194 | n9528 ;
  assign n24426 = n24425 ^ n20615 ^ 1'b0 ;
  assign n24427 = n17314 ^ n2811 ^ 1'b0 ;
  assign n24428 = n5511 | n20578 ;
  assign n24429 = ( ~n6211 & n7854 ) | ( ~n6211 & n21797 ) | ( n7854 & n21797 ) ;
  assign n24431 = n17462 ^ n6148 ^ n503 ;
  assign n24430 = ~n3709 & n4285 ;
  assign n24432 = n24431 ^ n24430 ^ n15025 ;
  assign n24433 = n1824 | n21020 ;
  assign n24434 = n18247 & n18938 ;
  assign n24435 = ( n21908 & n24433 ) | ( n21908 & n24434 ) | ( n24433 & n24434 ) ;
  assign n24436 = ( ~n3034 & n5854 ) | ( ~n3034 & n18658 ) | ( n5854 & n18658 ) ;
  assign n24437 = ~n2414 & n2666 ;
  assign n24438 = n21848 & n24437 ;
  assign n24439 = n6784 | n13649 ;
  assign n24440 = n13649 & ~n24439 ;
  assign n24441 = n10234 ^ n1485 ^ 1'b0 ;
  assign n24442 = ~n306 & n17611 ;
  assign n24443 = n19743 ^ n4895 ^ 1'b0 ;
  assign n24444 = n2214 & ~n24443 ;
  assign n24445 = x46 & n7983 ;
  assign n24446 = n24445 ^ n19030 ^ 1'b0 ;
  assign n24447 = ~n1135 & n24446 ;
  assign n24448 = n24444 & n24447 ;
  assign n24449 = n1358 & ~n21978 ;
  assign n24450 = n21978 & n24449 ;
  assign n24451 = n12474 ^ n4467 ^ 1'b0 ;
  assign n24452 = n24450 | n24451 ;
  assign n24453 = n1860 & n3038 ;
  assign n24454 = ~n3398 & n24453 ;
  assign n24455 = n24454 ^ n8089 ^ 1'b0 ;
  assign n24456 = ( n14160 & n24452 ) | ( n14160 & n24455 ) | ( n24452 & n24455 ) ;
  assign n24457 = ( n2715 & n4578 ) | ( n2715 & ~n18896 ) | ( n4578 & ~n18896 ) ;
  assign n24458 = n24457 ^ n9233 ^ n5603 ;
  assign n24459 = ( ~n1001 & n11184 ) | ( ~n1001 & n22942 ) | ( n11184 & n22942 ) ;
  assign n24460 = n13101 ^ n13066 ^ 1'b0 ;
  assign n24461 = n24459 & n24460 ;
  assign n24462 = n6716 ^ n2105 ^ 1'b0 ;
  assign n24463 = n373 & ~n24462 ;
  assign n24464 = n24463 ^ n19450 ^ 1'b0 ;
  assign n24465 = n3031 ^ n987 ^ 1'b0 ;
  assign n24466 = ~n1842 & n9681 ;
  assign n24467 = n24466 ^ n11745 ^ 1'b0 ;
  assign n24468 = n24467 ^ n17196 ^ 1'b0 ;
  assign n24469 = n7401 & n10703 ;
  assign n24470 = n24469 ^ n12120 ^ n2875 ;
  assign n24471 = n22943 ^ n9591 ^ n9587 ;
  assign n24472 = n311 ^ x3 ^ 1'b0 ;
  assign n24475 = n15971 ^ n1476 ^ 1'b0 ;
  assign n24476 = n3172 & n24475 ;
  assign n24473 = n15616 ^ n4581 ^ 1'b0 ;
  assign n24474 = n15957 | n24473 ;
  assign n24477 = n24476 ^ n24474 ^ 1'b0 ;
  assign n24478 = n20872 ^ n6097 ^ 1'b0 ;
  assign n24479 = n18509 & n24478 ;
  assign n24480 = n7762 ^ n4634 ^ 1'b0 ;
  assign n24481 = n7967 & ~n24480 ;
  assign n24482 = n4942 & n24481 ;
  assign n24483 = n24482 ^ n10099 ^ 1'b0 ;
  assign n24484 = n415 & n11292 ;
  assign n24485 = n24484 ^ n2920 ^ 1'b0 ;
  assign n24486 = ~n14320 & n24485 ;
  assign n24487 = n24486 ^ n9382 ^ 1'b0 ;
  assign n24488 = n4477 & n9184 ;
  assign n24489 = n16643 & ~n20992 ;
  assign n24492 = n8834 | n11376 ;
  assign n24491 = n1212 & n10491 ;
  assign n24493 = n24492 ^ n24491 ^ 1'b0 ;
  assign n24490 = n9142 & ~n13815 ;
  assign n24494 = n24493 ^ n24490 ^ n18226 ;
  assign n24495 = n23124 & ~n24160 ;
  assign n24496 = ( n16658 & ~n24369 ) | ( n16658 & n24495 ) | ( ~n24369 & n24495 ) ;
  assign n24497 = n3749 ^ n3235 ^ 1'b0 ;
  assign n24498 = ~n1318 & n24497 ;
  assign n24499 = n7231 | n14435 ;
  assign n24500 = n7795 & ~n13685 ;
  assign n24501 = n1046 | n5965 ;
  assign n24502 = n24501 ^ n13216 ^ 1'b0 ;
  assign n24503 = n18496 ^ n15722 ^ n9221 ;
  assign n24504 = n603 & ~n14603 ;
  assign n24505 = ~n3770 & n24504 ;
  assign n24506 = ~n2243 & n24505 ;
  assign n24507 = ( ~n11085 & n22947 ) | ( ~n11085 & n24506 ) | ( n22947 & n24506 ) ;
  assign n24508 = n21026 ^ n612 ^ 1'b0 ;
  assign n24509 = n6548 & n24508 ;
  assign n24510 = n10594 & n24509 ;
  assign n24511 = n2379 ^ n873 ^ 1'b0 ;
  assign n24512 = n3634 & n24511 ;
  assign n24513 = n5277 & n24512 ;
  assign n24514 = n24513 ^ n14342 ^ 1'b0 ;
  assign n24517 = n12169 ^ n425 ^ 1'b0 ;
  assign n24515 = ~n891 & n24454 ;
  assign n24516 = ~n18342 & n24515 ;
  assign n24518 = n24517 ^ n24516 ^ 1'b0 ;
  assign n24519 = ~n547 & n2543 ;
  assign n24520 = ~n3230 & n24519 ;
  assign n24521 = n24520 ^ n10616 ^ n3297 ;
  assign n24522 = n3152 | n24521 ;
  assign n24523 = n15284 | n24522 ;
  assign n24524 = n20019 ^ n11079 ^ 1'b0 ;
  assign n24525 = n1675 & n24524 ;
  assign n24526 = n10581 ^ n1387 ^ 1'b0 ;
  assign n24527 = ~n2463 & n24526 ;
  assign n24528 = n8664 & ~n12747 ;
  assign n24529 = n24528 ^ n2337 ^ 1'b0 ;
  assign n24530 = n20067 ^ n8919 ^ n6348 ;
  assign n24531 = n7185 & n24530 ;
  assign n24532 = n15150 ^ n8022 ^ 1'b0 ;
  assign n24533 = n7558 & n22815 ;
  assign n24534 = ~n24532 & n24533 ;
  assign n24536 = n12785 ^ n9010 ^ 1'b0 ;
  assign n24537 = ~n18168 & n24536 ;
  assign n24538 = n24537 ^ n1260 ^ 1'b0 ;
  assign n24535 = n1637 ^ n1081 ^ 1'b0 ;
  assign n24539 = n24538 ^ n24535 ^ n10935 ;
  assign n24540 = n24539 ^ n2654 ^ 1'b0 ;
  assign n24541 = n2355 & n24540 ;
  assign n24542 = n13842 ^ n1886 ^ 1'b0 ;
  assign n24543 = n24541 & ~n24542 ;
  assign n24544 = n16643 ^ n5355 ^ 1'b0 ;
  assign n24545 = n18858 & n24544 ;
  assign n24546 = ( n10047 & n20137 ) | ( n10047 & n20246 ) | ( n20137 & n20246 ) ;
  assign n24547 = ~n11419 & n19881 ;
  assign n24548 = ( n3886 & n13144 ) | ( n3886 & ~n24547 ) | ( n13144 & ~n24547 ) ;
  assign n24549 = ~n7689 & n8287 ;
  assign n24550 = n11203 ^ n6016 ^ 1'b0 ;
  assign n24551 = ~n24549 & n24550 ;
  assign n24552 = ~n13777 & n14580 ;
  assign n24553 = n24552 ^ n10948 ^ 1'b0 ;
  assign n24554 = n2219 & n18417 ;
  assign n24555 = n13085 & ~n24554 ;
  assign n24556 = n24553 & n24555 ;
  assign n24558 = n3770 ^ n1480 ^ 1'b0 ;
  assign n24559 = ~n1747 & n24558 ;
  assign n24557 = n8974 & ~n16708 ;
  assign n24560 = n24559 ^ n24557 ^ 1'b0 ;
  assign n24561 = n2717 & ~n10048 ;
  assign n24562 = n9428 | n21601 ;
  assign n24563 = n24562 ^ n10473 ^ 1'b0 ;
  assign n24565 = n12942 ^ n11298 ^ n536 ;
  assign n24564 = n9865 & n11792 ;
  assign n24566 = n24565 ^ n24564 ^ n9923 ;
  assign n24567 = n18164 & n24566 ;
  assign n24568 = n7814 ^ n3585 ^ 1'b0 ;
  assign n24569 = n8329 & n8330 ;
  assign n24570 = n21906 ^ n2107 ^ 1'b0 ;
  assign n24571 = n5836 & ~n24570 ;
  assign n24572 = n3269 & ~n8063 ;
  assign n24573 = ~n1603 & n8437 ;
  assign n24574 = n24573 ^ n388 ^ 1'b0 ;
  assign n24575 = n6407 | n17143 ;
  assign n24576 = n24574 & ~n24575 ;
  assign n24577 = n8377 ^ n5662 ^ 1'b0 ;
  assign n24578 = n14437 ^ n12728 ^ n5645 ;
  assign n24579 = n22384 | n24578 ;
  assign n24580 = n24579 ^ n21242 ^ 1'b0 ;
  assign n24581 = ( ~n757 & n4747 ) | ( ~n757 & n5340 ) | ( n4747 & n5340 ) ;
  assign n24582 = n11058 ^ n6789 ^ 1'b0 ;
  assign n24583 = n24581 & ~n24582 ;
  assign n24584 = ~n515 & n17549 ;
  assign n24585 = n18585 & n24584 ;
  assign n24586 = ( n3582 & n12412 ) | ( n3582 & n19998 ) | ( n12412 & n19998 ) ;
  assign n24587 = ( n5201 & n9457 ) | ( n5201 & ~n13022 ) | ( n9457 & ~n13022 ) ;
  assign n24588 = n14856 & ~n18442 ;
  assign n24589 = n1853 & n16641 ;
  assign n24590 = n24589 ^ n14750 ^ 1'b0 ;
  assign n24592 = n11420 ^ n2264 ^ 1'b0 ;
  assign n24591 = n1370 | n12034 ;
  assign n24593 = n24592 ^ n24591 ^ 1'b0 ;
  assign n24594 = n2621 & n16844 ;
  assign n24595 = ~n8776 & n24594 ;
  assign n24596 = n24595 ^ n23514 ^ 1'b0 ;
  assign n24597 = n11420 & n24596 ;
  assign n24598 = ~n7549 & n7691 ;
  assign n24599 = n12897 ^ n11519 ^ n11518 ;
  assign n24600 = ~n1592 & n5554 ;
  assign n24601 = ~n5554 & n24600 ;
  assign n24602 = n24601 ^ n2236 ^ 1'b0 ;
  assign n24603 = ( n11463 & n21082 ) | ( n11463 & ~n24602 ) | ( n21082 & ~n24602 ) ;
  assign n24604 = n10150 & ~n23442 ;
  assign n24605 = n3571 & n7994 ;
  assign n24606 = n15704 ^ n11428 ^ 1'b0 ;
  assign n24607 = n24605 | n24606 ;
  assign n24608 = ~n1979 & n9339 ;
  assign n24609 = n24607 & n24608 ;
  assign n24610 = ( ~n24603 & n24604 ) | ( ~n24603 & n24609 ) | ( n24604 & n24609 ) ;
  assign n24611 = n10045 ^ n1382 ^ 1'b0 ;
  assign n24612 = ~n7938 & n24611 ;
  assign n24613 = n11343 ^ n10428 ^ 1'b0 ;
  assign n24614 = ~n6241 & n8962 ;
  assign n24615 = n24614 ^ n1844 ^ 1'b0 ;
  assign n24616 = n15229 & n16275 ;
  assign n24617 = n24616 ^ n21317 ^ 1'b0 ;
  assign n24618 = n5135 ^ n3308 ^ 1'b0 ;
  assign n24619 = n1237 & ~n24618 ;
  assign n24620 = n24619 ^ n9438 ^ 1'b0 ;
  assign n24621 = ( n6353 & n10229 ) | ( n6353 & ~n12546 ) | ( n10229 & ~n12546 ) ;
  assign n24622 = n4689 | n11762 ;
  assign n24623 = n753 | n24622 ;
  assign n24624 = n9910 | n24623 ;
  assign n24625 = n13940 ^ n12273 ^ 1'b0 ;
  assign n24626 = ~n15327 & n24625 ;
  assign n24627 = n14306 ^ n7748 ^ 1'b0 ;
  assign n24628 = n8187 | n24627 ;
  assign n24632 = n20465 ^ n15879 ^ 1'b0 ;
  assign n24633 = n3783 & n24632 ;
  assign n24629 = ~n10060 & n19723 ;
  assign n24630 = n24629 ^ n7083 ^ 1'b0 ;
  assign n24631 = n21961 & ~n24630 ;
  assign n24634 = n24633 ^ n24631 ^ 1'b0 ;
  assign n24635 = n24430 ^ n11230 ^ n5947 ;
  assign n24636 = n24635 ^ n12812 ^ 1'b0 ;
  assign n24637 = n3391 ^ n3040 ^ 1'b0 ;
  assign n24638 = n24637 ^ n5945 ^ n2279 ;
  assign n24639 = n3760 & ~n9145 ;
  assign n24640 = n24639 ^ n17052 ^ 1'b0 ;
  assign n24641 = ~n3117 & n6998 ;
  assign n24642 = n24641 ^ n8788 ^ 1'b0 ;
  assign n24643 = n24642 ^ n381 ^ 1'b0 ;
  assign n24644 = ~n3979 & n20024 ;
  assign n24645 = n24644 ^ n12121 ^ 1'b0 ;
  assign n24646 = n24645 ^ n5924 ^ 1'b0 ;
  assign n24647 = n14422 & ~n24646 ;
  assign n24648 = n18432 ^ n16178 ^ 1'b0 ;
  assign n24649 = n24648 ^ n3275 ^ 1'b0 ;
  assign n24650 = n2844 | n11882 ;
  assign n24651 = n24650 ^ n3624 ^ n2376 ;
  assign n24652 = ~n9169 & n11611 ;
  assign n24653 = n19820 ^ n13550 ^ n12037 ;
  assign n24654 = n1191 | n5754 ;
  assign n24655 = ( n2014 & ~n19652 ) | ( n2014 & n24654 ) | ( ~n19652 & n24654 ) ;
  assign n24656 = n24655 ^ n12518 ^ n8528 ;
  assign n24657 = ( ~n3576 & n7908 ) | ( ~n3576 & n13713 ) | ( n7908 & n13713 ) ;
  assign n24658 = ~n2317 & n8505 ;
  assign n24659 = n24658 ^ n188 ^ 1'b0 ;
  assign n24660 = ~n1467 & n13052 ;
  assign n24661 = n1083 & ~n24660 ;
  assign n24662 = n4281 ^ n1229 ^ 1'b0 ;
  assign n24663 = n9043 & n24662 ;
  assign n24664 = ~n5741 & n10729 ;
  assign n24665 = n24664 ^ n21639 ^ 1'b0 ;
  assign n24666 = n4993 | n24665 ;
  assign n24667 = n1683 & ~n24666 ;
  assign n24668 = n3111 ^ x111 ^ 1'b0 ;
  assign n24669 = n24668 ^ n21524 ^ 1'b0 ;
  assign n24670 = n14054 & n15713 ;
  assign n24671 = ~n12171 & n24670 ;
  assign n24672 = n19975 ^ n11684 ^ 1'b0 ;
  assign n24673 = n14073 & ~n20823 ;
  assign n24674 = n15290 ^ n9957 ^ 1'b0 ;
  assign n24675 = n134 & n8106 ;
  assign n24676 = n24675 ^ n19678 ^ 1'b0 ;
  assign n24677 = n7703 | n24676 ;
  assign n24678 = n24677 ^ n4644 ^ 1'b0 ;
  assign n24679 = ~n7496 & n16517 ;
  assign n24680 = ~n13527 & n24679 ;
  assign n24681 = n8273 ^ n1046 ^ 1'b0 ;
  assign n24682 = n8198 ^ n7379 ^ n2861 ;
  assign n24683 = n6964 & n8202 ;
  assign n24684 = n5826 & n24683 ;
  assign n24685 = n24684 ^ n7368 ^ 1'b0 ;
  assign n24686 = n10863 | n24685 ;
  assign n24687 = ~n8090 & n11651 ;
  assign n24688 = n5225 ^ n717 ^ 1'b0 ;
  assign n24689 = ~n5673 & n19340 ;
  assign n24690 = n24183 ^ n4025 ^ 1'b0 ;
  assign n24691 = n6265 & n15303 ;
  assign n24692 = n3372 & ~n11212 ;
  assign n24693 = ~n4757 & n24692 ;
  assign n24694 = n24693 ^ n10530 ^ 1'b0 ;
  assign n24695 = ~n2812 & n24694 ;
  assign n24696 = ~n6428 & n24695 ;
  assign n24697 = n12226 & n18706 ;
  assign n24698 = n24697 ^ n16057 ^ 1'b0 ;
  assign n24699 = x12 & n2505 ;
  assign n24700 = n24698 & n24699 ;
  assign n24701 = ( n7566 & n13021 ) | ( n7566 & ~n24700 ) | ( n13021 & ~n24700 ) ;
  assign n24702 = n10971 ^ n956 ^ 1'b0 ;
  assign n24703 = n24701 & ~n24702 ;
  assign n24704 = n6087 ^ n4429 ^ 1'b0 ;
  assign n24705 = n9417 & n24704 ;
  assign n24706 = ~n23225 & n24705 ;
  assign n24707 = n5338 & n24706 ;
  assign n24708 = n10188 & n23285 ;
  assign n24709 = n9558 ^ n5447 ^ n5340 ;
  assign n24710 = n15336 & ~n24709 ;
  assign n24711 = n4223 & ~n6202 ;
  assign n24712 = n3845 & n24711 ;
  assign n24713 = n6494 | n17913 ;
  assign n24714 = n20221 & n24713 ;
  assign n24715 = n24714 ^ n8845 ^ 1'b0 ;
  assign n24717 = n1169 & ~n5973 ;
  assign n24718 = n24717 ^ n2315 ^ 1'b0 ;
  assign n24716 = n5730 & ~n10517 ;
  assign n24719 = n24718 ^ n24716 ^ n18373 ;
  assign n24720 = n6134 & ~n24719 ;
  assign n24723 = n5486 ^ n1041 ^ n129 ;
  assign n24724 = n5185 & n24723 ;
  assign n24725 = n3656 | n24724 ;
  assign n24721 = n10325 & n16677 ;
  assign n24722 = n12230 | n24721 ;
  assign n24726 = n24725 ^ n24722 ^ n1738 ;
  assign n24727 = n14766 ^ n4268 ^ n2863 ;
  assign n24728 = n235 & n22744 ;
  assign n24729 = n2969 | n15194 ;
  assign n24730 = n398 & ~n21385 ;
  assign n24731 = ~n13997 & n24730 ;
  assign n24732 = n4685 & n20446 ;
  assign n24733 = n24732 ^ n237 ^ 1'b0 ;
  assign n24734 = n14748 | n16971 ;
  assign n24735 = n14267 & ~n24734 ;
  assign n24736 = n6931 & ~n24735 ;
  assign n24737 = n19954 ^ n14056 ^ n3567 ;
  assign n24738 = n9800 ^ n9605 ^ 1'b0 ;
  assign n24739 = n7416 | n24738 ;
  assign n24740 = n24739 ^ n24252 ^ n16330 ;
  assign n24741 = n16328 | n22326 ;
  assign n24742 = n11193 | n24741 ;
  assign n24743 = ~n19627 & n24742 ;
  assign n24744 = ~n8382 & n24743 ;
  assign n24745 = n8845 | n20421 ;
  assign n24746 = n4246 | n24745 ;
  assign n24749 = ~n4907 & n9322 ;
  assign n24750 = ~n8231 & n24749 ;
  assign n24747 = n7562 ^ n5711 ^ 1'b0 ;
  assign n24748 = n1504 & n24747 ;
  assign n24751 = n24750 ^ n24748 ^ 1'b0 ;
  assign n24752 = n24751 ^ n17799 ^ 1'b0 ;
  assign n24753 = n4410 & n20579 ;
  assign n24754 = ~n17673 & n24753 ;
  assign n24755 = n1423 & n7238 ;
  assign n24756 = n4532 ^ n2850 ^ 1'b0 ;
  assign n24757 = n14749 | n24756 ;
  assign n24758 = n24757 ^ n6363 ^ n5081 ;
  assign n24759 = n23497 ^ n8102 ^ n2951 ;
  assign n24760 = n153 & n691 ;
  assign n24761 = n13758 & n24760 ;
  assign n24762 = ( n6448 & ~n13966 ) | ( n6448 & n24761 ) | ( ~n13966 & n24761 ) ;
  assign n24763 = n4801 ^ x63 ^ 1'b0 ;
  assign n24764 = n2485 & n24763 ;
  assign n24765 = n9657 | n13022 ;
  assign n24766 = n24764 & n24765 ;
  assign n24767 = ~n5970 & n11767 ;
  assign n24768 = n24767 ^ n3259 ^ 1'b0 ;
  assign n24769 = n15800 & n16150 ;
  assign n24770 = n7558 & n15734 ;
  assign n24771 = n24770 ^ n4006 ^ 1'b0 ;
  assign n24772 = n6845 & ~n24771 ;
  assign n24773 = ~n13212 & n24772 ;
  assign n24774 = n20317 ^ n4693 ^ 1'b0 ;
  assign n24775 = n24773 | n24774 ;
  assign n24776 = n7731 | n16662 ;
  assign n24777 = n19252 & ~n20815 ;
  assign n24778 = n1109 | n2835 ;
  assign n24779 = n24778 ^ n5585 ^ 1'b0 ;
  assign n24780 = n7865 & ~n24779 ;
  assign n24781 = n24780 ^ n9950 ^ 1'b0 ;
  assign n24785 = n10482 ^ n9068 ^ n3866 ;
  assign n24782 = n18331 ^ n10801 ^ 1'b0 ;
  assign n24783 = n7920 & n24782 ;
  assign n24784 = n4055 | n24783 ;
  assign n24786 = n24785 ^ n24784 ^ 1'b0 ;
  assign n24787 = n24774 ^ n7796 ^ 1'b0 ;
  assign n24788 = ( ~n3281 & n12772 ) | ( ~n3281 & n14829 ) | ( n12772 & n14829 ) ;
  assign n24789 = n12588 ^ n10580 ^ 1'b0 ;
  assign n24790 = n7781 & n24789 ;
  assign n24791 = n20232 ^ n523 ^ 1'b0 ;
  assign n24792 = n2519 & n9787 ;
  assign n24793 = n24792 ^ n20690 ^ 1'b0 ;
  assign n24794 = ~n3681 & n6265 ;
  assign n24795 = n24794 ^ n4316 ^ 1'b0 ;
  assign n24796 = n24795 ^ n950 ^ 1'b0 ;
  assign n24797 = ~n13685 & n24796 ;
  assign n24798 = ( ~n2253 & n4428 ) | ( ~n2253 & n7716 ) | ( n4428 & n7716 ) ;
  assign n24799 = n24798 ^ n3900 ^ n2640 ;
  assign n24800 = n24799 ^ n19691 ^ 1'b0 ;
  assign n24801 = n22700 ^ n7787 ^ 1'b0 ;
  assign n24802 = n24801 ^ n2291 ^ n2216 ;
  assign n24803 = ( ~n299 & n3594 ) | ( ~n299 & n18440 ) | ( n3594 & n18440 ) ;
  assign n24804 = n24803 ^ n18846 ^ n4285 ;
  assign n24805 = n3741 | n7444 ;
  assign n24806 = n24805 ^ n4297 ^ 1'b0 ;
  assign n24807 = ~n700 & n24806 ;
  assign n24808 = ~n267 & n892 ;
  assign n24809 = n267 & n24808 ;
  assign n24810 = n1364 & ~n24809 ;
  assign n24811 = ~n1364 & n24810 ;
  assign n24812 = n2603 & ~n2897 ;
  assign n24813 = n24811 & n24812 ;
  assign n24814 = n521 & n4689 ;
  assign n24815 = ~n4689 & n24814 ;
  assign n24816 = n24813 | n24815 ;
  assign n24817 = n24813 & ~n24816 ;
  assign n24818 = n2333 | n4720 ;
  assign n24819 = n24817 & ~n24818 ;
  assign n24820 = n4691 & ~n24819 ;
  assign n24821 = n24819 & n24820 ;
  assign n24822 = n4937 | n24821 ;
  assign n24823 = n24822 ^ n14032 ^ 1'b0 ;
  assign n24824 = ~n3999 & n24823 ;
  assign n24825 = n24824 ^ n2801 ^ 1'b0 ;
  assign n24826 = n23635 & n24825 ;
  assign n24827 = n16537 ^ n9096 ^ 1'b0 ;
  assign n24828 = n16025 & ~n24827 ;
  assign n24829 = n6015 ^ n1909 ^ 1'b0 ;
  assign n24830 = n24828 & n24829 ;
  assign n24831 = n17978 ^ n7604 ^ 1'b0 ;
  assign n24832 = ~n23327 & n24831 ;
  assign n24833 = ~n1163 & n22173 ;
  assign n24834 = ~n24832 & n24833 ;
  assign n24835 = n6916 & ~n9228 ;
  assign n24836 = n24835 ^ n1276 ^ 1'b0 ;
  assign n24837 = ~n1104 & n7639 ;
  assign n24838 = n632 | n923 ;
  assign n24839 = n11729 | n24838 ;
  assign n24840 = n18078 & ~n21595 ;
  assign n24841 = ~n258 & n21346 ;
  assign n24842 = ( n6187 & ~n8697 ) | ( n6187 & n24841 ) | ( ~n8697 & n24841 ) ;
  assign n24843 = ( n3758 & ~n5771 ) | ( n3758 & n24536 ) | ( ~n5771 & n24536 ) ;
  assign n24844 = n5189 ^ n4778 ^ 1'b0 ;
  assign n24845 = ( ~n8848 & n24843 ) | ( ~n8848 & n24844 ) | ( n24843 & n24844 ) ;
  assign n24846 = n7111 & ~n12516 ;
  assign n24847 = ~n10419 & n24846 ;
  assign n24848 = n24847 ^ n6195 ^ 1'b0 ;
  assign n24849 = n23690 ^ n18164 ^ 1'b0 ;
  assign n24850 = ~n8805 & n20961 ;
  assign n24851 = n1977 ^ x39 ^ 1'b0 ;
  assign n24852 = n901 & n24851 ;
  assign n24853 = n24852 ^ n12386 ^ 1'b0 ;
  assign n24854 = n9284 ^ n8050 ^ 1'b0 ;
  assign n24855 = n6765 | n24854 ;
  assign n24856 = n24855 ^ n10888 ^ 1'b0 ;
  assign n24857 = n21020 ^ n10040 ^ n3947 ;
  assign n24858 = n24857 ^ n21210 ^ n4014 ;
  assign n24859 = n2912 ^ n2128 ^ 1'b0 ;
  assign n24860 = n11001 ^ n2861 ^ 1'b0 ;
  assign n24861 = n895 & ~n24860 ;
  assign n24862 = n10640 ^ n4143 ^ 1'b0 ;
  assign n24863 = n581 & n2528 ;
  assign n24864 = n6517 & ~n24863 ;
  assign n24865 = ~n6488 & n24864 ;
  assign n24866 = n11230 | n18465 ;
  assign n24871 = ~n6046 & n16628 ;
  assign n24872 = n24871 ^ n18219 ^ 1'b0 ;
  assign n24867 = ~n4819 & n12487 ;
  assign n24868 = ~n3899 & n24867 ;
  assign n24869 = n7666 & n24868 ;
  assign n24870 = n24869 ^ n6632 ^ 1'b0 ;
  assign n24873 = n24872 ^ n24870 ^ n8026 ;
  assign n24874 = ~n928 & n11474 ;
  assign n24875 = n7396 ^ n3342 ^ 1'b0 ;
  assign n24876 = n1633 & n24875 ;
  assign n24877 = n24874 & n24876 ;
  assign n24878 = n9908 ^ n840 ^ 1'b0 ;
  assign n24879 = n24877 | n24878 ;
  assign n24880 = n7883 & n12305 ;
  assign n24881 = ~n24879 & n24880 ;
  assign n24883 = n15997 ^ n10266 ^ n928 ;
  assign n24884 = n3561 & ~n24883 ;
  assign n24882 = ~n1866 & n12210 ;
  assign n24885 = n24884 ^ n24882 ^ 1'b0 ;
  assign n24886 = ~n6899 & n7562 ;
  assign n24887 = n24886 ^ n7463 ^ 1'b0 ;
  assign n24888 = n5156 & ~n24887 ;
  assign n24889 = ~n13970 & n24888 ;
  assign n24890 = n1360 ^ n698 ^ 1'b0 ;
  assign n24891 = n19769 ^ n10740 ^ 1'b0 ;
  assign n24892 = ~n1200 & n15367 ;
  assign n24893 = ~n2672 & n24892 ;
  assign n24894 = n24893 ^ n16685 ^ 1'b0 ;
  assign n24895 = n21465 ^ n12660 ^ n10673 ;
  assign n24896 = n24895 ^ n23283 ^ 1'b0 ;
  assign n24897 = n24129 ^ n16534 ^ n11954 ;
  assign n24898 = n1559 & ~n6231 ;
  assign n24899 = n2276 & n24898 ;
  assign n24900 = n8097 & ~n22096 ;
  assign n24901 = n4011 & ~n24900 ;
  assign n24902 = ~n1776 & n24901 ;
  assign n24903 = ( n5383 & ~n6781 ) | ( n5383 & n7124 ) | ( ~n6781 & n7124 ) ;
  assign n24904 = n9485 & ~n24903 ;
  assign n24905 = n13977 ^ n9425 ^ n1261 ;
  assign n24906 = n3947 | n24905 ;
  assign n24907 = ~n6907 & n13433 ;
  assign n24908 = ( ~n7587 & n13548 ) | ( ~n7587 & n23189 ) | ( n13548 & n23189 ) ;
  assign n24909 = n8130 & n24908 ;
  assign n24910 = n24909 ^ n22700 ^ n296 ;
  assign n24911 = n18535 ^ n6826 ^ 1'b0 ;
  assign n24912 = n24911 ^ n19703 ^ n3732 ;
  assign n24913 = n4946 & ~n9184 ;
  assign n24914 = n3537 & ~n17764 ;
  assign n24915 = n24914 ^ n10181 ^ 1'b0 ;
  assign n24916 = ~n6400 & n13685 ;
  assign n24917 = n13113 | n18592 ;
  assign n24918 = n24916 | n24917 ;
  assign n24919 = n614 & n803 ;
  assign n24920 = ~n1436 & n24919 ;
  assign n24921 = n24920 ^ n13624 ^ 1'b0 ;
  assign n24922 = n17969 ^ n1590 ^ 1'b0 ;
  assign n24925 = n7197 & ~n8052 ;
  assign n24923 = n7877 & n19199 ;
  assign n24924 = n24923 ^ x3 ^ 1'b0 ;
  assign n24926 = n24925 ^ n24924 ^ n1589 ;
  assign n24927 = ~n11344 & n16185 ;
  assign n24928 = n24927 ^ n683 ^ 1'b0 ;
  assign n24929 = n19306 & n21332 ;
  assign n24930 = ( ~n5259 & n24928 ) | ( ~n5259 & n24929 ) | ( n24928 & n24929 ) ;
  assign n24931 = n4806 | n14585 ;
  assign n24932 = n10436 | n24931 ;
  assign n24933 = n20402 | n24932 ;
  assign n24934 = n18024 ^ x83 ^ 1'b0 ;
  assign n24935 = n16044 | n24934 ;
  assign n24936 = n19174 | n24935 ;
  assign n24937 = n19097 ^ n12293 ^ 1'b0 ;
  assign n24938 = ~n4443 & n24937 ;
  assign n24939 = n13733 & ~n24938 ;
  assign n24940 = ~n5826 & n19773 ;
  assign n24941 = ~n4528 & n24940 ;
  assign n24942 = n1203 | n4361 ;
  assign n24943 = n24942 ^ n9027 ^ 1'b0 ;
  assign n24944 = n16326 & ~n24943 ;
  assign n24945 = n838 & n24944 ;
  assign n24946 = n8231 ^ n3350 ^ 1'b0 ;
  assign n24947 = n1846 & n24946 ;
  assign n24948 = n14882 ^ n6153 ^ 1'b0 ;
  assign n24949 = n14274 & n24948 ;
  assign n24950 = ( x49 & ~n24947 ) | ( x49 & n24949 ) | ( ~n24947 & n24949 ) ;
  assign n24955 = ~n846 & n22099 ;
  assign n24951 = n7894 ^ n352 ^ 1'b0 ;
  assign n24952 = n23018 ^ n4092 ^ 1'b0 ;
  assign n24953 = n13424 | n24952 ;
  assign n24954 = ( n20450 & n24951 ) | ( n20450 & n24953 ) | ( n24951 & n24953 ) ;
  assign n24956 = n24955 ^ n24954 ^ 1'b0 ;
  assign n24957 = n18778 & ~n21388 ;
  assign n24958 = ( n6907 & ~n8261 ) | ( n6907 & n24957 ) | ( ~n8261 & n24957 ) ;
  assign n24959 = ( n2789 & ~n18127 ) | ( n2789 & n24958 ) | ( ~n18127 & n24958 ) ;
  assign n24960 = n18658 ^ n10888 ^ 1'b0 ;
  assign n24961 = ~n254 & n12177 ;
  assign n24962 = ~n11173 & n24961 ;
  assign n24963 = n919 & ~n3800 ;
  assign n24964 = ~n15312 & n24963 ;
  assign n24965 = ( ~n4721 & n7607 ) | ( ~n4721 & n16263 ) | ( n7607 & n16263 ) ;
  assign n24966 = n7976 & ~n8120 ;
  assign n24967 = n24966 ^ n10306 ^ 1'b0 ;
  assign n24968 = ~n229 & n24967 ;
  assign n24969 = n24965 & n24968 ;
  assign n24970 = n12812 & n13818 ;
  assign n24971 = n6703 ^ n3976 ^ 1'b0 ;
  assign n24972 = ( n4283 & ~n21144 ) | ( n4283 & n24718 ) | ( ~n21144 & n24718 ) ;
  assign n24973 = n24972 ^ n13965 ^ 1'b0 ;
  assign n24974 = n13566 | n24973 ;
  assign n24975 = ~n1461 & n9857 ;
  assign n24976 = n24975 ^ n23469 ^ 1'b0 ;
  assign n24977 = ( n24971 & n24974 ) | ( n24971 & n24976 ) | ( n24974 & n24976 ) ;
  assign n24978 = n11176 ^ n9602 ^ n9141 ;
  assign n24980 = ~n1309 & n12687 ;
  assign n24981 = ~x49 & n24980 ;
  assign n24979 = n21844 ^ n13551 ^ n7866 ;
  assign n24982 = n24981 ^ n24979 ^ n9988 ;
  assign n24983 = n9663 ^ n1157 ^ 1'b0 ;
  assign n24984 = n1147 & ~n24983 ;
  assign n24985 = n24984 ^ n16986 ^ 1'b0 ;
  assign n24986 = n4511 | n24985 ;
  assign n24987 = n3503 | n3996 ;
  assign n24988 = n9085 & ~n10445 ;
  assign n24989 = n13870 ^ n7764 ^ n6126 ;
  assign n24990 = ( n3176 & n4951 ) | ( n3176 & ~n24989 ) | ( n4951 & ~n24989 ) ;
  assign n24991 = n5920 ^ n1815 ^ 1'b0 ;
  assign n24992 = ( n3315 & n3411 ) | ( n3315 & n13786 ) | ( n3411 & n13786 ) ;
  assign n24993 = n10214 | n24992 ;
  assign n24994 = n13034 | n24993 ;
  assign n24995 = ~n155 & n24994 ;
  assign n24996 = n24995 ^ n11230 ^ 1'b0 ;
  assign n24997 = n10922 | n24996 ;
  assign n24998 = n11557 ^ n1994 ^ 1'b0 ;
  assign n24999 = n24998 ^ n12731 ^ 1'b0 ;
  assign n25000 = n1244 & ~n3217 ;
  assign n25001 = n24999 & n25000 ;
  assign n25002 = n17623 ^ n4082 ^ 1'b0 ;
  assign n25003 = n6464 ^ n3484 ^ 1'b0 ;
  assign n25004 = ~n25002 & n25003 ;
  assign n25005 = n1692 & ~n2306 ;
  assign n25006 = ( n1261 & n17115 ) | ( n1261 & ~n20168 ) | ( n17115 & ~n20168 ) ;
  assign n25007 = n1728 & ~n4667 ;
  assign n25008 = ( n9999 & n16433 ) | ( n9999 & n25007 ) | ( n16433 & n25007 ) ;
  assign n25009 = n20330 ^ n17898 ^ 1'b0 ;
  assign n25010 = ( n4219 & n4307 ) | ( n4219 & n11191 ) | ( n4307 & n11191 ) ;
  assign n25011 = n2663 & ~n25010 ;
  assign n25012 = ~n4371 & n15711 ;
  assign n25013 = ~n15554 & n25012 ;
  assign n25014 = n5265 & ~n25013 ;
  assign n25015 = n25014 ^ n21441 ^ 1'b0 ;
  assign n25016 = n3691 & ~n5236 ;
  assign n25017 = n9909 & n25016 ;
  assign n25018 = n1133 | n7463 ;
  assign n25019 = ~n12374 & n14950 ;
  assign n25020 = n25019 ^ n12880 ^ 1'b0 ;
  assign n25021 = ( n6451 & n18491 ) | ( n6451 & ~n23381 ) | ( n18491 & ~n23381 ) ;
  assign n25022 = ~n16294 & n19719 ;
  assign n25023 = n25022 ^ n19571 ^ n6023 ;
  assign n25024 = n13940 ^ n6384 ^ n731 ;
  assign n25025 = n8118 ^ n6891 ^ 1'b0 ;
  assign n25026 = n2523 & ~n25025 ;
  assign n25028 = n676 & n6133 ;
  assign n25029 = n25028 ^ n4717 ^ 1'b0 ;
  assign n25027 = n1675 & ~n9268 ;
  assign n25030 = n25029 ^ n25027 ^ 1'b0 ;
  assign n25031 = n8795 & n25030 ;
  assign n25032 = n4454 & ~n21409 ;
  assign n25033 = n22589 ^ n12318 ^ 1'b0 ;
  assign n25034 = n22691 ^ n9152 ^ 1'b0 ;
  assign n25035 = ~n1169 & n25034 ;
  assign n25036 = n22341 ^ n18380 ^ n3935 ;
  assign n25037 = n19388 ^ n14531 ^ 1'b0 ;
  assign n25038 = ( n2581 & n4076 ) | ( n2581 & ~n25037 ) | ( n4076 & ~n25037 ) ;
  assign n25039 = n899 & ~n7071 ;
  assign n25040 = n9088 ^ n6371 ^ 1'b0 ;
  assign n25041 = ~n15057 & n25040 ;
  assign n25042 = n25041 ^ n12817 ^ 1'b0 ;
  assign n25043 = n3800 ^ n3652 ^ n1307 ;
  assign n25044 = n2081 | n25043 ;
  assign n25045 = n18940 | n21466 ;
  assign n25046 = n1476 & ~n1927 ;
  assign n25047 = n18065 | n25046 ;
  assign n25048 = n19574 ^ n18939 ^ n9285 ;
  assign n25049 = n8137 ^ n949 ^ 1'b0 ;
  assign n25050 = n6214 & n25049 ;
  assign n25051 = ~n25048 & n25050 ;
  assign n25053 = n9863 ^ n2510 ^ x16 ;
  assign n25054 = n11010 & ~n25053 ;
  assign n25052 = n865 & ~n3540 ;
  assign n25055 = n25054 ^ n25052 ^ 1'b0 ;
  assign n25056 = n6145 ^ n1025 ^ 1'b0 ;
  assign n25057 = n24181 ^ n3694 ^ 1'b0 ;
  assign n25058 = n2417 ^ n1542 ^ 1'b0 ;
  assign n25059 = n25058 ^ n17763 ^ n6955 ;
  assign n25060 = ~n7772 & n19526 ;
  assign n25061 = n6439 ^ n4456 ^ 1'b0 ;
  assign n25062 = n25060 | n25061 ;
  assign n25066 = n9052 | n9634 ;
  assign n25063 = n10763 ^ n7850 ^ 1'b0 ;
  assign n25064 = n15800 & n25063 ;
  assign n25065 = ~n7365 & n25064 ;
  assign n25067 = n25066 ^ n25065 ^ 1'b0 ;
  assign n25068 = n9176 ^ n1839 ^ 1'b0 ;
  assign n25069 = n6569 ^ n3350 ^ 1'b0 ;
  assign n25070 = n21082 | n25069 ;
  assign n25071 = n25070 ^ n9679 ^ 1'b0 ;
  assign n25072 = n1230 | n25071 ;
  assign n25073 = n11163 ^ n2173 ^ 1'b0 ;
  assign n25074 = n4039 & ~n25073 ;
  assign n25075 = ( n652 & ~n12434 ) | ( n652 & n25074 ) | ( ~n12434 & n25074 ) ;
  assign n25076 = n25075 ^ n13602 ^ 1'b0 ;
  assign n25077 = n16442 ^ n10497 ^ 1'b0 ;
  assign n25078 = n7004 & ~n25077 ;
  assign n25079 = ( n3065 & ~n17087 ) | ( n3065 & n25078 ) | ( ~n17087 & n25078 ) ;
  assign n25080 = n6943 ^ n1307 ^ 1'b0 ;
  assign n25081 = n15906 & ~n25080 ;
  assign n25082 = ~n25010 & n25081 ;
  assign n25083 = ( n681 & n1008 ) | ( n681 & ~n1181 ) | ( n1008 & ~n1181 ) ;
  assign n25084 = n5786 ^ n4966 ^ 1'b0 ;
  assign n25085 = n25083 & ~n25084 ;
  assign n25086 = ~n7695 & n25085 ;
  assign n25087 = n13142 & n25086 ;
  assign n25088 = n7778 | n15804 ;
  assign n25089 = n8191 & ~n25088 ;
  assign n25090 = n10084 & n19928 ;
  assign n25091 = n25090 ^ n12653 ^ 1'b0 ;
  assign n25101 = n4181 | n7311 ;
  assign n25097 = n3680 ^ n2807 ^ 1'b0 ;
  assign n25098 = n5573 & ~n25097 ;
  assign n25099 = n1887 & n25098 ;
  assign n25100 = n5685 & ~n25099 ;
  assign n25092 = n350 & ~n1841 ;
  assign n25093 = n25092 ^ n16810 ^ 1'b0 ;
  assign n25094 = n20128 & ~n23265 ;
  assign n25095 = n25093 & n25094 ;
  assign n25096 = n25095 ^ n10990 ^ n4375 ;
  assign n25102 = n25101 ^ n25100 ^ n25096 ;
  assign n25103 = n3212 ^ n2608 ^ n2500 ;
  assign n25104 = n25103 ^ n6320 ^ 1'b0 ;
  assign n25105 = ( n7480 & n22805 ) | ( n7480 & ~n25104 ) | ( n22805 & ~n25104 ) ;
  assign n25110 = ( ~n1265 & n14588 ) | ( ~n1265 & n24362 ) | ( n14588 & n24362 ) ;
  assign n25111 = n25110 ^ n23960 ^ 1'b0 ;
  assign n25112 = ~n22981 & n25111 ;
  assign n25106 = n597 & ~n12464 ;
  assign n25107 = n25106 ^ n436 ^ 1'b0 ;
  assign n25108 = n25107 ^ n19646 ^ n14308 ;
  assign n25109 = n25108 ^ n14119 ^ 1'b0 ;
  assign n25113 = n25112 ^ n25109 ^ n23167 ;
  assign n25114 = ~x51 & n7990 ;
  assign n25115 = ~n1550 & n25114 ;
  assign n25116 = n1354 | n6557 ;
  assign n25117 = ~n9060 & n13540 ;
  assign n25118 = ~n14683 & n25117 ;
  assign n25119 = n6931 & n8376 ;
  assign n25120 = n25119 ^ n7808 ^ 1'b0 ;
  assign n25121 = ~n817 & n2700 ;
  assign n25122 = n25121 ^ n9409 ^ 1'b0 ;
  assign n25123 = n8711 | n25122 ;
  assign n25124 = n9881 & ~n14933 ;
  assign n25125 = ~n24032 & n25124 ;
  assign n25126 = n16664 ^ n6070 ^ 1'b0 ;
  assign n25127 = n23698 ^ n8353 ^ n1677 ;
  assign n25128 = n758 & ~n3036 ;
  assign n25129 = ~n778 & n25128 ;
  assign n25130 = n15255 & ~n25129 ;
  assign n25131 = n25130 ^ n11931 ^ 1'b0 ;
  assign n25133 = ( ~n379 & n6571 ) | ( ~n379 & n17171 ) | ( n6571 & n17171 ) ;
  assign n25132 = n5845 & n23577 ;
  assign n25134 = n25133 ^ n25132 ^ 1'b0 ;
  assign n25135 = n3962 & ~n14734 ;
  assign n25136 = n15388 & n24002 ;
  assign n25137 = n25136 ^ n7939 ^ 1'b0 ;
  assign n25138 = n10619 ^ n2623 ^ 1'b0 ;
  assign n25139 = n17411 & n25138 ;
  assign n25140 = n3240 ^ n254 ^ 1'b0 ;
  assign n25141 = n25139 & n25140 ;
  assign n25143 = n20629 ^ n14957 ^ 1'b0 ;
  assign n25142 = n12281 ^ n8983 ^ n4714 ;
  assign n25144 = n25143 ^ n25142 ^ 1'b0 ;
  assign n25145 = ~n640 & n23343 ;
  assign n25146 = ( ~n6192 & n19668 ) | ( ~n6192 & n23508 ) | ( n19668 & n23508 ) ;
  assign n25147 = n21116 & n25146 ;
  assign n25148 = ~n7900 & n18156 ;
  assign n25149 = n25148 ^ n4959 ^ 1'b0 ;
  assign n25150 = n14959 & ~n20763 ;
  assign n25151 = ~n24857 & n25150 ;
  assign n25153 = ( n1734 & ~n3684 ) | ( n1734 & n4497 ) | ( ~n3684 & n4497 ) ;
  assign n25152 = n2098 & n9077 ;
  assign n25154 = n25153 ^ n25152 ^ 1'b0 ;
  assign n25155 = n5389 & ~n16294 ;
  assign n25156 = n25155 ^ n20263 ^ 1'b0 ;
  assign n25157 = n24905 ^ n5233 ^ 1'b0 ;
  assign n25158 = n24512 ^ n14835 ^ n4721 ;
  assign n25159 = n3228 ^ n974 ^ 1'b0 ;
  assign n25160 = ~n6687 & n25159 ;
  assign n25161 = n4362 ^ n873 ^ 1'b0 ;
  assign n25162 = ~n7196 & n8482 ;
  assign n25163 = n25162 ^ n4575 ^ 1'b0 ;
  assign n25164 = n25163 ^ n7491 ^ 1'b0 ;
  assign n25165 = n5910 | n20655 ;
  assign n25166 = n12217 & n25165 ;
  assign n25167 = n19037 & ~n19419 ;
  assign n25168 = ( n16938 & n22665 ) | ( n16938 & n22898 ) | ( n22665 & n22898 ) ;
  assign n25169 = n5381 & ~n25168 ;
  assign n25170 = n11559 ^ n1309 ^ 1'b0 ;
  assign n25171 = n1281 & n14359 ;
  assign n25175 = ~n4543 & n14836 ;
  assign n25176 = n25175 ^ n2553 ^ 1'b0 ;
  assign n25173 = ~n1260 & n5990 ;
  assign n25174 = n20643 & n25173 ;
  assign n25172 = ~n673 & n1674 ;
  assign n25177 = n25176 ^ n25174 ^ n25172 ;
  assign n25178 = n2951 & n25177 ;
  assign n25179 = n25178 ^ n14911 ^ 1'b0 ;
  assign n25180 = n19203 | n19878 ;
  assign n25181 = n12765 | n25180 ;
  assign n25182 = n25066 ^ n12451 ^ 1'b0 ;
  assign n25183 = n12025 & ~n14697 ;
  assign n25184 = ~n3637 & n22021 ;
  assign n25185 = n9026 & n14729 ;
  assign n25186 = ( n19351 & n19861 ) | ( n19351 & n24538 ) | ( n19861 & n24538 ) ;
  assign n25187 = ~n5246 & n16063 ;
  assign n25188 = n2442 & n25187 ;
  assign n25189 = n11003 | n25188 ;
  assign n25190 = ~n833 & n22658 ;
  assign n25191 = n8541 & n25190 ;
  assign n25192 = n14231 | n16041 ;
  assign n25193 = n22370 ^ n442 ^ 1'b0 ;
  assign n25194 = n2007 | n25193 ;
  assign n25195 = n12050 & ~n25194 ;
  assign n25196 = n8818 & ~n15216 ;
  assign n25197 = n25196 ^ n15399 ^ 1'b0 ;
  assign n25198 = n25195 & ~n25197 ;
  assign n25199 = n25198 ^ n14819 ^ x121 ;
  assign n25200 = n5950 & ~n9211 ;
  assign n25201 = n2005 & ~n25200 ;
  assign n25202 = n25201 ^ n19724 ^ n18804 ;
  assign n25203 = n14748 ^ n13561 ^ 1'b0 ;
  assign n25204 = n15911 | n25203 ;
  assign n25205 = n25204 ^ n13744 ^ n4466 ;
  assign n25206 = n2809 & ~n11460 ;
  assign n25207 = n25206 ^ n10675 ^ 1'b0 ;
  assign n25208 = ~n1040 & n12275 ;
  assign n25209 = ~n555 & n21123 ;
  assign n25210 = x38 & n19576 ;
  assign n25211 = n25210 ^ n7094 ^ 1'b0 ;
  assign n25212 = ( x3 & ~n436 ) | ( x3 & n12536 ) | ( ~n436 & n12536 ) ;
  assign n25213 = n11114 ^ n8344 ^ 1'b0 ;
  assign n25214 = n25212 | n25213 ;
  assign n25215 = ~n11235 & n25214 ;
  assign n25216 = n3070 & n14322 ;
  assign n25217 = n5997 ^ n3438 ^ 1'b0 ;
  assign n25218 = n25217 ^ n13731 ^ 1'b0 ;
  assign n25219 = n15816 ^ n12696 ^ n8152 ;
  assign n25220 = n14997 & ~n21670 ;
  assign n25221 = ( ~n17135 & n17672 ) | ( ~n17135 & n25220 ) | ( n17672 & n25220 ) ;
  assign n25222 = n16690 ^ n9564 ^ 1'b0 ;
  assign n25223 = n16136 ^ n791 ^ 1'b0 ;
  assign n25224 = n14699 | n25223 ;
  assign n25225 = n25224 ^ n1989 ^ 1'b0 ;
  assign n25226 = ~n9653 & n25225 ;
  assign n25227 = n5872 & n10436 ;
  assign n25228 = ~n5723 & n25227 ;
  assign n25229 = n3979 ^ n3249 ^ 1'b0 ;
  assign n25230 = n8344 & ~n25229 ;
  assign n25231 = n10487 & n25230 ;
  assign n25232 = n9525 & n25231 ;
  assign n25233 = n4915 ^ n1669 ^ 1'b0 ;
  assign n25234 = n20600 ^ n11042 ^ n6176 ;
  assign n25235 = n3985 ^ n764 ^ 1'b0 ;
  assign n25236 = n10691 ^ n9746 ^ n6131 ;
  assign n25237 = n25236 ^ n19852 ^ 1'b0 ;
  assign n25238 = n2958 & ~n10188 ;
  assign n25239 = n21485 ^ n21269 ^ n8408 ;
  assign n25240 = ~n1051 & n25239 ;
  assign n25241 = ~n19177 & n25240 ;
  assign n25242 = n314 & ~n17648 ;
  assign n25243 = n25242 ^ n9222 ^ 1'b0 ;
  assign n25244 = n25243 ^ n7109 ^ x2 ;
  assign n25245 = n25244 ^ n16623 ^ 1'b0 ;
  assign n25246 = n10054 ^ n1621 ^ 1'b0 ;
  assign n25247 = n9754 | n25246 ;
  assign n25248 = ~n5449 & n13097 ;
  assign n25249 = n25248 ^ n17593 ^ n3593 ;
  assign n25250 = ( n3612 & n11485 ) | ( n3612 & n21301 ) | ( n11485 & n21301 ) ;
  assign n25251 = n22125 | n25250 ;
  assign n25252 = n8900 ^ n7328 ^ 1'b0 ;
  assign n25253 = n3567 | n25252 ;
  assign n25254 = n708 & ~n18210 ;
  assign n25255 = n25253 & n25254 ;
  assign n25256 = n3270 & n24648 ;
  assign n25257 = n25256 ^ n12314 ^ 1'b0 ;
  assign n25258 = n480 ^ n220 ^ 1'b0 ;
  assign n25259 = n25258 ^ n12121 ^ 1'b0 ;
  assign n25260 = n9152 & ~n17138 ;
  assign n25261 = n25260 ^ n24389 ^ 1'b0 ;
  assign n25262 = n5025 & ~n10229 ;
  assign n25263 = n15769 ^ n3546 ^ 1'b0 ;
  assign n25264 = n5773 | n20303 ;
  assign n25265 = n2972 & ~n25264 ;
  assign n25266 = n912 & n15906 ;
  assign n25267 = n25266 ^ n2101 ^ 1'b0 ;
  assign n25268 = n18728 & ~n25267 ;
  assign n25269 = n14582 | n22027 ;
  assign n25270 = n20545 ^ n18376 ^ 1'b0 ;
  assign n25271 = ~n7353 & n25270 ;
  assign n25272 = n25269 | n25271 ;
  assign n25273 = ~n8269 & n15739 ;
  assign n25274 = n11468 ^ n8487 ^ 1'b0 ;
  assign n25275 = n22206 & ~n25274 ;
  assign n25276 = ~n6227 & n22446 ;
  assign n25277 = ~n24463 & n25276 ;
  assign n25278 = n24755 ^ n10481 ^ 1'b0 ;
  assign n25279 = n18289 & n25278 ;
  assign n25280 = n16309 ^ n3037 ^ 1'b0 ;
  assign n25281 = n4252 & ~n25280 ;
  assign n25282 = n5258 & n5383 ;
  assign n25283 = ~n11061 & n25282 ;
  assign n25284 = n840 | n25283 ;
  assign n25285 = n21248 ^ n3105 ^ 1'b0 ;
  assign n25286 = ~n25284 & n25285 ;
  assign n25287 = n2386 & n7558 ;
  assign n25288 = n20768 ^ n2190 ^ n599 ;
  assign n25289 = ( n4755 & ~n25287 ) | ( n4755 & n25288 ) | ( ~n25287 & n25288 ) ;
  assign n25290 = n10971 ^ n5373 ^ n1373 ;
  assign n25291 = n1240 & n8134 ;
  assign n25292 = n967 | n25100 ;
  assign n25293 = n1062 | n25292 ;
  assign n25294 = ( n10273 & ~n25291 ) | ( n10273 & n25293 ) | ( ~n25291 & n25293 ) ;
  assign n25295 = n25290 | n25294 ;
  assign n25296 = n2710 & ~n20107 ;
  assign n25297 = ~n2886 & n25296 ;
  assign n25298 = n25297 ^ n5243 ^ 1'b0 ;
  assign n25299 = ( n10210 & ~n13142 ) | ( n10210 & n25298 ) | ( ~n13142 & n25298 ) ;
  assign n25300 = x51 & ~n5089 ;
  assign n25301 = n8534 | n25300 ;
  assign n25302 = n3491 | n25301 ;
  assign n25303 = n25302 ^ n9960 ^ 1'b0 ;
  assign n25304 = n14306 | n15263 ;
  assign n25305 = n25304 ^ n12443 ^ 1'b0 ;
  assign n25306 = n9778 ^ x44 ^ 1'b0 ;
  assign n25307 = ~n25305 & n25306 ;
  assign n25308 = n2243 & n19269 ;
  assign n25309 = n25308 ^ n1009 ^ 1'b0 ;
  assign n25310 = ( n5293 & ~n11190 ) | ( n5293 & n12032 ) | ( ~n11190 & n12032 ) ;
  assign n25311 = n25310 ^ n16559 ^ 1'b0 ;
  assign n25312 = ~n25309 & n25311 ;
  assign n25318 = ~n6255 & n6497 ;
  assign n25313 = n2608 ^ n1615 ^ 1'b0 ;
  assign n25314 = n280 & ~n25313 ;
  assign n25315 = ~n11420 & n25314 ;
  assign n25316 = n6283 ^ x46 ^ 1'b0 ;
  assign n25317 = n25315 | n25316 ;
  assign n25319 = n25318 ^ n25317 ^ n17623 ;
  assign n25320 = n10577 & n19226 ;
  assign n25321 = n25320 ^ n10668 ^ 1'b0 ;
  assign n25322 = n13215 ^ n12084 ^ 1'b0 ;
  assign n25323 = n24496 ^ n1333 ^ 1'b0 ;
  assign n25324 = n3048 & n15192 ;
  assign n25325 = n9790 & n25324 ;
  assign n25326 = n8382 & ~n25325 ;
  assign n25327 = n11441 & n25326 ;
  assign n25328 = n8727 ^ n1693 ^ 1'b0 ;
  assign n25329 = n11556 & ~n15937 ;
  assign n25330 = n25329 ^ n4770 ^ 1'b0 ;
  assign n25331 = n21822 ^ n20791 ^ 1'b0 ;
  assign n25332 = n25330 | n25331 ;
  assign n25333 = n17074 & ~n22640 ;
  assign n25334 = n10939 ^ x105 ^ 1'b0 ;
  assign n25335 = n21466 ^ n6478 ^ 1'b0 ;
  assign n25336 = n3291 | n14540 ;
  assign n25337 = n1169 | n8780 ;
  assign n25338 = n25337 ^ n4847 ^ 1'b0 ;
  assign n25339 = n7444 | n25338 ;
  assign n25340 = n2761 & ~n25339 ;
  assign n25341 = n2647 & n25340 ;
  assign n25342 = n2649 ^ n1473 ^ 1'b0 ;
  assign n25343 = n4490 & ~n25342 ;
  assign n25344 = n1722 | n19849 ;
  assign n25345 = n25343 & n25344 ;
  assign n25346 = n8608 & ~n25345 ;
  assign n25347 = n25346 ^ n6906 ^ 1'b0 ;
  assign n25348 = n4472 | n23769 ;
  assign n25349 = ~n10946 & n25348 ;
  assign n25350 = n5247 ^ n929 ^ 1'b0 ;
  assign n25351 = n8640 | n25350 ;
  assign n25352 = n6813 ^ n5274 ^ 1'b0 ;
  assign n25353 = ( n5082 & n8565 ) | ( n5082 & ~n19574 ) | ( n8565 & ~n19574 ) ;
  assign n25354 = ( n22439 & ~n25352 ) | ( n22439 & n25353 ) | ( ~n25352 & n25353 ) ;
  assign n25355 = n3475 & ~n17954 ;
  assign n25356 = n8358 | n25355 ;
  assign n25359 = x85 & ~n2923 ;
  assign n25360 = n25359 ^ n1185 ^ 1'b0 ;
  assign n25357 = n8195 ^ n8120 ^ 1'b0 ;
  assign n25358 = n7182 & n25357 ;
  assign n25361 = n25360 ^ n25358 ^ n4443 ;
  assign n25362 = n1966 & n5598 ;
  assign n25363 = ~n25361 & n25362 ;
  assign n25364 = n14675 & ~n15296 ;
  assign n25365 = n6295 | n7558 ;
  assign n25366 = n4085 | n13701 ;
  assign n25367 = n10504 ^ n8269 ^ 1'b0 ;
  assign n25368 = ~n8249 & n25367 ;
  assign n25369 = ( ~n265 & n2612 ) | ( ~n265 & n20147 ) | ( n2612 & n20147 ) ;
  assign n25370 = n21038 & ~n25369 ;
  assign n25371 = n22738 ^ n17346 ^ n4087 ;
  assign n25372 = ( n427 & n3995 ) | ( n427 & ~n18388 ) | ( n3995 & ~n18388 ) ;
  assign n25373 = n7454 & ~n25372 ;
  assign n25374 = n21029 & n25373 ;
  assign n25375 = n13598 ^ n7698 ^ 1'b0 ;
  assign n25376 = n9667 | n25375 ;
  assign n25377 = n10622 & n13212 ;
  assign n25378 = ~n4085 & n15267 ;
  assign n25379 = n17043 & n25378 ;
  assign n25380 = n25379 ^ n9209 ^ 1'b0 ;
  assign n25381 = n14725 ^ n3208 ^ 1'b0 ;
  assign n25383 = n2199 & ~n3376 ;
  assign n25382 = n20682 ^ n18123 ^ 1'b0 ;
  assign n25384 = n25383 ^ n25382 ^ n5705 ;
  assign n25385 = ( n1459 & n17729 ) | ( n1459 & ~n19488 ) | ( n17729 & ~n19488 ) ;
  assign n25386 = n4884 | n25385 ;
  assign n25387 = n17771 ^ n2049 ^ 1'b0 ;
  assign n25388 = n11300 ^ n4264 ^ 1'b0 ;
  assign n25389 = n19404 & ~n25388 ;
  assign n25390 = ~n3998 & n25389 ;
  assign n25391 = n6182 & n25390 ;
  assign n25392 = n25391 ^ n10185 ^ n8122 ;
  assign n25393 = n1800 & n4927 ;
  assign n25394 = n25393 ^ n1432 ^ 1'b0 ;
  assign n25395 = n18547 | n20156 ;
  assign n25396 = ( n11520 & ~n25394 ) | ( n11520 & n25395 ) | ( ~n25394 & n25395 ) ;
  assign n25397 = ~n5790 & n24131 ;
  assign n25398 = n23203 ^ n6431 ^ 1'b0 ;
  assign n25399 = ~n18338 & n23082 ;
  assign n25400 = ~n25398 & n25399 ;
  assign n25401 = n9376 & ~n25400 ;
  assign n25402 = ~n4812 & n8523 ;
  assign n25403 = n25402 ^ n17757 ^ 1'b0 ;
  assign n25404 = ~n11320 & n25403 ;
  assign n25405 = n3497 & ~n10916 ;
  assign n25406 = n25405 ^ n13282 ^ 1'b0 ;
  assign n25407 = n141 ^ x86 ^ 1'b0 ;
  assign n25408 = n8838 | n17587 ;
  assign n25410 = ~n4047 & n21469 ;
  assign n25409 = n12752 & ~n19450 ;
  assign n25411 = n25410 ^ n25409 ^ 1'b0 ;
  assign n25413 = n8390 | n10312 ;
  assign n25414 = n25413 ^ n17999 ^ 1'b0 ;
  assign n25415 = ~n22817 & n25414 ;
  assign n25412 = n6344 | n10324 ;
  assign n25416 = n25415 ^ n25412 ^ 1'b0 ;
  assign n25417 = n10430 ^ n2262 ^ 1'b0 ;
  assign n25418 = n3061 & ~n25417 ;
  assign n25419 = n25418 ^ n13532 ^ 1'b0 ;
  assign n25420 = ( n14526 & n16426 ) | ( n14526 & n25419 ) | ( n16426 & n25419 ) ;
  assign n25421 = n7169 | n25420 ;
  assign n25422 = n6617 & ~n23831 ;
  assign n25423 = ( ~n5885 & n16427 ) | ( ~n5885 & n25422 ) | ( n16427 & n25422 ) ;
  assign n25424 = n18109 ^ n3618 ^ 1'b0 ;
  assign n25425 = n25424 ^ n11790 ^ n3189 ;
  assign n25426 = n25425 ^ n14735 ^ 1'b0 ;
  assign n25427 = n4029 & ~n25426 ;
  assign n25428 = ( ~n730 & n21505 ) | ( ~n730 & n25427 ) | ( n21505 & n25427 ) ;
  assign n25429 = ( n1669 & ~n3028 ) | ( n1669 & n3124 ) | ( ~n3028 & n3124 ) ;
  assign n25430 = n14114 & ~n25429 ;
  assign n25431 = n2299 & n25430 ;
  assign n25432 = n4951 | n15438 ;
  assign n25433 = n25432 ^ n19763 ^ n9239 ;
  assign n25434 = x96 & n9981 ;
  assign n25435 = ~x122 & n25434 ;
  assign n25436 = n1970 | n4940 ;
  assign n25437 = n13869 & ~n25436 ;
  assign n25438 = n2489 & n3240 ;
  assign n25439 = n25438 ^ n6015 ^ 1'b0 ;
  assign n25440 = n2450 & ~n6756 ;
  assign n25441 = n15902 | n25440 ;
  assign n25442 = n13787 & ~n25441 ;
  assign n25443 = n24868 ^ n11165 ^ 1'b0 ;
  assign n25444 = n25443 ^ n1006 ^ n513 ;
  assign n25445 = n1971 | n6866 ;
  assign n25446 = n25195 | n25445 ;
  assign n25447 = n25446 ^ n9823 ^ 1'b0 ;
  assign n25448 = ~n442 & n25447 ;
  assign n25449 = ( n411 & n17463 ) | ( n411 & n25448 ) | ( n17463 & n25448 ) ;
  assign n25450 = n20407 ^ n7069 ^ 1'b0 ;
  assign n25451 = n3609 & n18537 ;
  assign n25452 = ~n4667 & n6579 ;
  assign n25453 = n25452 ^ n19177 ^ 1'b0 ;
  assign n25454 = n14745 ^ n11446 ^ 1'b0 ;
  assign n25455 = ~n3738 & n5655 ;
  assign n25456 = ~n11363 & n25455 ;
  assign n25457 = ~n25454 & n25456 ;
  assign n25458 = n6522 & ~n10662 ;
  assign n25459 = n2285 ^ n2011 ^ n2005 ;
  assign n25460 = n25459 ^ n5324 ^ 1'b0 ;
  assign n25461 = n25460 ^ n7778 ^ 1'b0 ;
  assign n25462 = n19443 ^ n9518 ^ 1'b0 ;
  assign n25463 = ~n5881 & n25462 ;
  assign n25464 = ( n2256 & n12571 ) | ( n2256 & n23181 ) | ( n12571 & n23181 ) ;
  assign n25465 = n7853 ^ n5848 ^ 1'b0 ;
  assign n25466 = ~n25464 & n25465 ;
  assign n25468 = ~n5032 & n6849 ;
  assign n25467 = ~n4506 & n12136 ;
  assign n25469 = n25468 ^ n25467 ^ 1'b0 ;
  assign n25470 = ~x3 & n9857 ;
  assign n25471 = ~n2122 & n25470 ;
  assign n25472 = ( n1652 & n11760 ) | ( n1652 & n25471 ) | ( n11760 & n25471 ) ;
  assign n25473 = n25472 ^ n9144 ^ n4880 ;
  assign n25474 = ( n1680 & ~n3626 ) | ( n1680 & n25473 ) | ( ~n3626 & n25473 ) ;
  assign n25475 = n17686 ^ n10522 ^ n6933 ;
  assign n25476 = n21336 & n24463 ;
  assign n25477 = n6899 & n25476 ;
  assign n25478 = n218 & ~n20228 ;
  assign n25479 = n25478 ^ n22581 ^ 1'b0 ;
  assign n25480 = n23664 ^ n13666 ^ 1'b0 ;
  assign n25481 = ( ~n2371 & n2965 ) | ( ~n2371 & n8257 ) | ( n2965 & n8257 ) ;
  assign n25484 = n8217 ^ n3214 ^ 1'b0 ;
  assign n25485 = n2574 | n25484 ;
  assign n25482 = ~n202 & n13481 ;
  assign n25483 = n25482 ^ n8719 ^ 1'b0 ;
  assign n25486 = n25485 ^ n25483 ^ n24086 ;
  assign n25487 = n7941 & ~n17635 ;
  assign n25488 = n25487 ^ n17869 ^ 1'b0 ;
  assign n25489 = ( ~n977 & n4008 ) | ( ~n977 & n25488 ) | ( n4008 & n25488 ) ;
  assign n25490 = n14373 ^ n240 ^ 1'b0 ;
  assign n25491 = n15580 | n25490 ;
  assign n25492 = ~n10533 & n21006 ;
  assign n25493 = n25492 ^ n10060 ^ 1'b0 ;
  assign n25495 = n14275 & n18887 ;
  assign n25494 = n16814 & ~n17264 ;
  assign n25496 = n25495 ^ n25494 ^ 1'b0 ;
  assign n25497 = n20995 ^ n6291 ^ 1'b0 ;
  assign n25498 = n25497 ^ n15706 ^ 1'b0 ;
  assign n25499 = n22784 ^ n19707 ^ n5067 ;
  assign n25500 = n22483 ^ n13214 ^ n7067 ;
  assign n25501 = n18168 & n25500 ;
  assign n25502 = ~n2133 & n19761 ;
  assign n25503 = n25502 ^ n15211 ^ 1'b0 ;
  assign n25504 = n10461 ^ n665 ^ 1'b0 ;
  assign n25505 = n3040 & n9840 ;
  assign n25506 = n17732 | n25505 ;
  assign n25507 = n25506 ^ n21602 ^ n8181 ;
  assign n25508 = n24273 ^ n10753 ^ n2637 ;
  assign n25509 = ( ~n17860 & n20867 ) | ( ~n17860 & n20909 ) | ( n20867 & n20909 ) ;
  assign n25510 = ~n10741 & n25509 ;
  assign n25511 = n9647 ^ n7955 ^ 1'b0 ;
  assign n25512 = ~n21097 & n25511 ;
  assign n25513 = n25512 ^ n22033 ^ 1'b0 ;
  assign n25514 = n25510 & ~n25513 ;
  assign n25515 = n18773 ^ n1806 ^ 1'b0 ;
  assign n25516 = n22881 ^ n17860 ^ 1'b0 ;
  assign n25517 = ~n25515 & n25516 ;
  assign n25518 = ~n3024 & n5307 ;
  assign n25519 = ~n380 & n2414 ;
  assign n25520 = n9287 & ~n25519 ;
  assign n25521 = n25518 & n25520 ;
  assign n25522 = n25521 ^ n1870 ^ 1'b0 ;
  assign n25523 = n1131 | n25522 ;
  assign n25524 = n7251 & n9540 ;
  assign n25525 = ( ~n9971 & n17609 ) | ( ~n9971 & n17799 ) | ( n17609 & n17799 ) ;
  assign n25526 = ( n601 & n1343 ) | ( n601 & n3503 ) | ( n1343 & n3503 ) ;
  assign n25527 = n25526 ^ n4035 ^ n2920 ;
  assign n25528 = ~n3166 & n25527 ;
  assign n25529 = ~n612 & n11677 ;
  assign n25530 = n25529 ^ n17744 ^ 1'b0 ;
  assign n25531 = n5662 & n25121 ;
  assign n25532 = n8438 | n8653 ;
  assign n25533 = n25532 ^ n6991 ^ n1410 ;
  assign n25534 = ~n4419 & n5968 ;
  assign n25535 = n18615 ^ n9216 ^ 1'b0 ;
  assign n25536 = n17270 | n25535 ;
  assign n25537 = n8401 | n16931 ;
  assign n25538 = n5542 & ~n25537 ;
  assign n25539 = n25538 ^ n23772 ^ 1'b0 ;
  assign n25540 = n24744 ^ n17712 ^ 1'b0 ;
  assign n25541 = ~n7381 & n8004 ;
  assign n25542 = n7263 | n25541 ;
  assign n25543 = n19795 & ~n25542 ;
  assign n25544 = n1424 & n6018 ;
  assign n25545 = n25358 ^ n5409 ^ 1'b0 ;
  assign n25546 = n25230 & n25545 ;
  assign n25547 = n19105 ^ n3765 ^ n3307 ;
  assign n25548 = n13808 | n23922 ;
  assign n25549 = n3950 & ~n25548 ;
  assign n25550 = n25549 ^ n24953 ^ n6518 ;
  assign n25551 = n2844 | n14967 ;
  assign n25552 = n12092 ^ n4311 ^ 1'b0 ;
  assign n25553 = n22520 | n25552 ;
  assign n25554 = n7084 ^ n6002 ^ 1'b0 ;
  assign n25555 = n9756 | n25554 ;
  assign n25556 = n3528 ^ n422 ^ 1'b0 ;
  assign n25557 = n8401 | n25556 ;
  assign n25558 = n25557 ^ n3940 ^ 1'b0 ;
  assign n25560 = n182 | n22698 ;
  assign n25561 = n10229 & ~n25560 ;
  assign n25559 = ~n7309 & n25098 ;
  assign n25562 = n25561 ^ n25559 ^ 1'b0 ;
  assign n25563 = ~n6633 & n13207 ;
  assign n25564 = n6011 & n25563 ;
  assign n25565 = n25564 ^ x23 ^ 1'b0 ;
  assign n25566 = ~n11128 & n15349 ;
  assign n25568 = n18953 & n22680 ;
  assign n25569 = n640 & n25568 ;
  assign n25567 = ~n5285 & n10723 ;
  assign n25570 = n25569 ^ n25567 ^ 1'b0 ;
  assign n25571 = n1819 & ~n22494 ;
  assign n25572 = n25571 ^ n11731 ^ 1'b0 ;
  assign n25573 = n25572 ^ n3794 ^ 1'b0 ;
  assign n25574 = n12835 & n15664 ;
  assign n25575 = ( ~n7265 & n11003 ) | ( ~n7265 & n25574 ) | ( n11003 & n25574 ) ;
  assign n25576 = n7154 & ~n10204 ;
  assign n25577 = n6555 & n25576 ;
  assign n25578 = n5201 & n11704 ;
  assign n25579 = n6705 & n25578 ;
  assign n25580 = n2146 | n5078 ;
  assign n25581 = n20698 | n25580 ;
  assign n25582 = n18167 ^ n10438 ^ 1'b0 ;
  assign n25583 = n23920 & ~n25582 ;
  assign n25584 = n1079 & n25583 ;
  assign n25585 = n18625 & n25584 ;
  assign n25586 = n1492 | n13153 ;
  assign n25587 = n370 & ~n1278 ;
  assign n25588 = n25587 ^ n1677 ^ 1'b0 ;
  assign n25589 = ( n18309 & n22287 ) | ( n18309 & ~n25588 ) | ( n22287 & ~n25588 ) ;
  assign n25590 = n10547 ^ n3997 ^ 1'b0 ;
  assign n25591 = n20127 | n25590 ;
  assign n25592 = n4489 | n14149 ;
  assign n25593 = n350 | n15525 ;
  assign n25594 = n25593 ^ n1713 ^ 1'b0 ;
  assign n25595 = n7326 | n10581 ;
  assign n25596 = n25594 & ~n25595 ;
  assign n25597 = n13538 ^ n1530 ^ 1'b0 ;
  assign n25599 = n4001 & ~n15576 ;
  assign n25600 = n25599 ^ n23832 ^ 1'b0 ;
  assign n25598 = n4582 & ~n7935 ;
  assign n25601 = n25600 ^ n25598 ^ 1'b0 ;
  assign n25602 = n6482 | n25601 ;
  assign n25603 = n3073 | n8795 ;
  assign n25604 = ~n9350 & n25603 ;
  assign n25605 = n697 & ~n23391 ;
  assign n25606 = n6367 | n13043 ;
  assign n25607 = n25606 ^ n14565 ^ 1'b0 ;
  assign n25612 = n5316 & n14697 ;
  assign n25609 = ~n8911 & n13135 ;
  assign n25610 = n25609 ^ n6040 ^ 1'b0 ;
  assign n25611 = ( ~n7258 & n15655 ) | ( ~n7258 & n25610 ) | ( n15655 & n25610 ) ;
  assign n25613 = n25612 ^ n25611 ^ n9137 ;
  assign n25608 = n210 & n8231 ;
  assign n25614 = n25613 ^ n25608 ^ 1'b0 ;
  assign n25615 = ~n7451 & n10781 ;
  assign n25616 = n8878 | n25615 ;
  assign n25617 = n20719 ^ n4029 ^ 1'b0 ;
  assign n25618 = ( n10800 & n17088 ) | ( n10800 & ~n20638 ) | ( n17088 & ~n20638 ) ;
  assign n25621 = n9803 & ~n12968 ;
  assign n25619 = n8532 ^ n7018 ^ 1'b0 ;
  assign n25620 = n25619 ^ n24665 ^ 1'b0 ;
  assign n25622 = n25621 ^ n25620 ^ n1099 ;
  assign n25623 = n10805 ^ n1521 ^ 1'b0 ;
  assign n25624 = n1338 & ~n21251 ;
  assign n25625 = ~n25623 & n25624 ;
  assign n25626 = n3953 & n9805 ;
  assign n25627 = n24876 ^ n828 ^ 1'b0 ;
  assign n25628 = n2611 & ~n25627 ;
  assign n25629 = n8818 & ~n15896 ;
  assign n25630 = n5333 & ~n12078 ;
  assign n25631 = n5267 & ~n13930 ;
  assign n25632 = n17331 & n25631 ;
  assign n25633 = ( n6685 & n16433 ) | ( n6685 & n25632 ) | ( n16433 & n25632 ) ;
  assign n25634 = n13503 ^ n12539 ^ n12379 ;
  assign n25635 = ~n5614 & n21526 ;
  assign n25636 = n25635 ^ n6189 ^ 1'b0 ;
  assign n25637 = n3823 ^ n407 ^ 1'b0 ;
  assign n25638 = n25637 ^ n12571 ^ 1'b0 ;
  assign n25639 = ~n5335 & n9713 ;
  assign n25640 = ( n235 & n4028 ) | ( n235 & n25639 ) | ( n4028 & n25639 ) ;
  assign n25641 = n25638 & n25640 ;
  assign n25642 = n6769 ^ n3212 ^ 1'b0 ;
  assign n25643 = ~n9074 & n16427 ;
  assign n25644 = n25643 ^ n6075 ^ 1'b0 ;
  assign n25645 = n25644 ^ n11380 ^ 1'b0 ;
  assign n25646 = n7328 & ~n25645 ;
  assign n25647 = n21015 ^ n6072 ^ 1'b0 ;
  assign n25648 = n21401 ^ n7172 ^ 1'b0 ;
  assign n25649 = n3859 & ~n25648 ;
  assign n25650 = n6878 ^ n6644 ^ 1'b0 ;
  assign n25651 = n899 | n22642 ;
  assign n25652 = n18309 & n19508 ;
  assign n25653 = n6245 & n10312 ;
  assign n25654 = n770 | n25653 ;
  assign n25655 = n25652 & ~n25654 ;
  assign n25656 = n22727 ^ n2853 ^ 1'b0 ;
  assign n25657 = ~n1808 & n25656 ;
  assign n25658 = n6858 ^ n763 ^ 1'b0 ;
  assign n25659 = n25657 & n25658 ;
  assign n25660 = n10368 ^ n130 ^ 1'b0 ;
  assign n25661 = n2507 | n25660 ;
  assign n25662 = n1914 & ~n10366 ;
  assign n25663 = n6217 | n10018 ;
  assign n25664 = n25663 ^ n7384 ^ 1'b0 ;
  assign n25665 = n3576 & n23767 ;
  assign n25666 = n9068 ^ n1408 ^ n285 ;
  assign n25667 = n8738 ^ n2647 ^ 1'b0 ;
  assign n25668 = n5217 & ~n25667 ;
  assign n25669 = n8471 & n25668 ;
  assign n25670 = n25666 & n25669 ;
  assign n25671 = n12227 & ~n14186 ;
  assign n25672 = ( n25665 & ~n25670 ) | ( n25665 & n25671 ) | ( ~n25670 & n25671 ) ;
  assign n25673 = n2333 & n18909 ;
  assign n25674 = n25673 ^ n23640 ^ 1'b0 ;
  assign n25675 = n23065 ^ n15135 ^ n3488 ;
  assign n25676 = n18118 ^ n6558 ^ 1'b0 ;
  assign n25677 = ~n171 & n5096 ;
  assign n25678 = n9088 & n12308 ;
  assign n25679 = n3910 | n24300 ;
  assign n25680 = n4044 | n11832 ;
  assign n25681 = n25680 ^ n17927 ^ n6139 ;
  assign n25682 = n2065 & n15861 ;
  assign n25683 = n2940 & ~n5066 ;
  assign n25684 = n24763 ^ n9702 ^ 1'b0 ;
  assign n25685 = n250 & ~n25684 ;
  assign n25686 = ( n2682 & n7028 ) | ( n2682 & n25685 ) | ( n7028 & n25685 ) ;
  assign n25687 = n25642 ^ n10183 ^ 1'b0 ;
  assign n25688 = n11225 ^ n6804 ^ 1'b0 ;
  assign n25689 = ~n3656 & n25688 ;
  assign n25690 = n19823 ^ n4337 ^ 1'b0 ;
  assign n25691 = n18591 & n25690 ;
  assign n25692 = n13612 & n23289 ;
  assign n25693 = ~n11236 & n12417 ;
  assign n25694 = ~n14412 & n25693 ;
  assign n25695 = ~n7778 & n25694 ;
  assign n25696 = n17584 ^ n7072 ^ 1'b0 ;
  assign n25697 = n17961 ^ n1843 ^ n190 ;
  assign n25699 = n2693 ^ n2216 ^ 1'b0 ;
  assign n25700 = n6325 | n25699 ;
  assign n25698 = n1813 | n5633 ;
  assign n25701 = n25700 ^ n25698 ^ 1'b0 ;
  assign n25702 = n18228 & ~n18863 ;
  assign n25703 = n2364 | n11101 ;
  assign n25704 = n25703 ^ n11524 ^ 1'b0 ;
  assign n25705 = ~n13681 & n20698 ;
  assign n25706 = ~n25704 & n25705 ;
  assign n25707 = ~n1082 & n3426 ;
  assign n25708 = ~n8622 & n17242 ;
  assign n25709 = n10440 & n10626 ;
  assign n25710 = n25709 ^ n13520 ^ 1'b0 ;
  assign n25711 = n3687 ^ n2073 ^ 1'b0 ;
  assign n25712 = n25710 & ~n25711 ;
  assign n25713 = n3389 & n3395 ;
  assign n25714 = ( ~n3870 & n11958 ) | ( ~n3870 & n25713 ) | ( n11958 & n25713 ) ;
  assign n25715 = n20012 ^ n239 ^ 1'b0 ;
  assign n25716 = n7794 ^ n4298 ^ 1'b0 ;
  assign n25717 = n8587 | n25716 ;
  assign n25718 = x25 & n2668 ;
  assign n25719 = ~n5548 & n25718 ;
  assign n25720 = n13419 & n25719 ;
  assign n25722 = n4358 | n13815 ;
  assign n25721 = n6394 & n12776 ;
  assign n25723 = n25722 ^ n25721 ^ 1'b0 ;
  assign n25724 = n9031 | n13243 ;
  assign n25725 = n25724 ^ n20666 ^ 1'b0 ;
  assign n25726 = n25725 ^ n13640 ^ 1'b0 ;
  assign n25727 = n8491 ^ n5003 ^ 1'b0 ;
  assign n25728 = ~n8288 & n25727 ;
  assign n25729 = ~n13070 & n19856 ;
  assign n25730 = ( n19902 & n25728 ) | ( n19902 & n25729 ) | ( n25728 & n25729 ) ;
  assign n25731 = n13093 ^ n11673 ^ n11046 ;
  assign n25732 = ( n12872 & n13814 ) | ( n12872 & ~n25731 ) | ( n13814 & ~n25731 ) ;
  assign n25733 = n6381 | n24733 ;
  assign n25734 = n12008 ^ n9370 ^ 1'b0 ;
  assign n25735 = n2969 | n25734 ;
  assign n25736 = ~n11111 & n25735 ;
  assign n25737 = n16078 ^ n7842 ^ 1'b0 ;
  assign n25738 = ~n21749 & n25737 ;
  assign n25739 = n21044 ^ n4938 ^ 1'b0 ;
  assign n25740 = n24204 | n25739 ;
  assign n25741 = n5074 ^ n1240 ^ 1'b0 ;
  assign n25742 = n4750 & ~n25741 ;
  assign n25743 = n17547 ^ n11746 ^ n6768 ;
  assign n25744 = n25742 & n25743 ;
  assign n25745 = n25744 ^ n4805 ^ 1'b0 ;
  assign n25746 = n9821 | n25745 ;
  assign n25747 = n24541 ^ n18844 ^ 1'b0 ;
  assign n25748 = n4376 & ~n25121 ;
  assign n25749 = ~n8204 & n11736 ;
  assign n25750 = n2840 | n13153 ;
  assign n25751 = n25749 & ~n25750 ;
  assign n25752 = n4294 ^ n2262 ^ n1935 ;
  assign n25753 = n4693 & ~n25752 ;
  assign n25754 = n25753 ^ n11399 ^ 1'b0 ;
  assign n25755 = n10199 & n10547 ;
  assign n25756 = ~n13085 & n25755 ;
  assign n25757 = n5944 ^ n3055 ^ 1'b0 ;
  assign n25758 = n12802 ^ n6927 ^ 1'b0 ;
  assign n25761 = n4260 ^ n2151 ^ 1'b0 ;
  assign n25759 = n3265 & n3434 ;
  assign n25760 = n25759 ^ n15433 ^ 1'b0 ;
  assign n25762 = n25761 ^ n25760 ^ n5718 ;
  assign n25763 = n9210 & n25762 ;
  assign n25765 = n2455 & ~n7400 ;
  assign n25766 = ( n5191 & ~n5530 ) | ( n5191 & n25765 ) | ( ~n5530 & n25765 ) ;
  assign n25764 = ~n7791 & n22225 ;
  assign n25767 = n25766 ^ n25764 ^ 1'b0 ;
  assign n25768 = n24182 ^ n6668 ^ 1'b0 ;
  assign n25769 = n159 | n13180 ;
  assign n25770 = ~n8552 & n22457 ;
  assign n25771 = n4655 | n6223 ;
  assign n25772 = n15489 & ~n25771 ;
  assign n25773 = n6052 | n9814 ;
  assign n25774 = n10789 & ~n25773 ;
  assign n25775 = ~n14957 & n25774 ;
  assign n25776 = ~n4993 & n14930 ;
  assign n25777 = n25776 ^ n6927 ^ 1'b0 ;
  assign n25778 = n1239 & n2313 ;
  assign n25779 = n1542 & n25778 ;
  assign n25780 = n25779 ^ n16714 ^ n5346 ;
  assign n25781 = ~n1139 & n24305 ;
  assign n25782 = n8530 & n25781 ;
  assign n25783 = n18243 ^ n2656 ^ 1'b0 ;
  assign n25784 = ~n4387 & n25783 ;
  assign n25785 = n510 | n5166 ;
  assign n25786 = n9822 & n14207 ;
  assign n25787 = n25786 ^ n1876 ^ 1'b0 ;
  assign n25788 = n8091 & ~n25787 ;
  assign n25789 = ~n2005 & n25788 ;
  assign n25790 = n24433 ^ n23112 ^ 1'b0 ;
  assign n25791 = n25789 & ~n25790 ;
  assign n25792 = x9 & ~n16805 ;
  assign n25794 = n17104 ^ n3374 ^ 1'b0 ;
  assign n25793 = x3 & ~n12493 ;
  assign n25795 = n25794 ^ n25793 ^ 1'b0 ;
  assign n25796 = n6176 | n25795 ;
  assign n25799 = ( n895 & n1239 ) | ( n895 & n3374 ) | ( n1239 & n3374 ) ;
  assign n25797 = n497 & n22903 ;
  assign n25798 = n25797 ^ n11854 ^ 1'b0 ;
  assign n25800 = n25799 ^ n25798 ^ n16745 ;
  assign n25801 = n6770 | n8899 ;
  assign n25802 = n25801 ^ n5656 ^ 1'b0 ;
  assign n25803 = ( n9482 & n23295 ) | ( n9482 & ~n25802 ) | ( n23295 & ~n25802 ) ;
  assign n25804 = n17888 ^ n13311 ^ n13307 ;
  assign n25805 = n7484 & n21039 ;
  assign n25806 = n11116 | n13327 ;
  assign n25807 = n9045 | n25806 ;
  assign n25808 = n15241 ^ n11265 ^ 1'b0 ;
  assign n25809 = ~n21706 & n23556 ;
  assign n25810 = ~n881 & n17382 ;
  assign n25811 = n1654 | n18961 ;
  assign n25812 = n25811 ^ n12588 ^ 1'b0 ;
  assign n25813 = n1645 ^ n1231 ^ 1'b0 ;
  assign n25814 = ~n1667 & n6392 ;
  assign n25815 = n25814 ^ n2081 ^ 1'b0 ;
  assign n25816 = n7258 ^ n3948 ^ n512 ;
  assign n25817 = n25815 & n25816 ;
  assign n25818 = n821 | n2596 ;
  assign n25819 = n25817 | n25818 ;
  assign n25820 = n12848 ^ n167 ^ x110 ;
  assign n25821 = n4448 & n25820 ;
  assign n25822 = n25821 ^ n19019 ^ 1'b0 ;
  assign n25823 = ~n2292 & n4429 ;
  assign n25824 = ~n345 & n25823 ;
  assign n25825 = n11187 ^ n5474 ^ 1'b0 ;
  assign n25826 = ( n383 & n21546 ) | ( n383 & n25825 ) | ( n21546 & n25825 ) ;
  assign n25827 = n25826 ^ n11526 ^ 1'b0 ;
  assign n25828 = n1134 & ~n5569 ;
  assign n25829 = n9615 | n25828 ;
  assign n25831 = n4700 | n7374 ;
  assign n25830 = n24177 ^ n15512 ^ n2892 ;
  assign n25832 = n25831 ^ n25830 ^ n10480 ;
  assign n25833 = n7919 ^ n6283 ^ n5295 ;
  assign n25834 = n4151 | n10188 ;
  assign n25835 = n25834 ^ n350 ^ 1'b0 ;
  assign n25836 = n25835 ^ n5831 ^ 1'b0 ;
  assign n25837 = n962 & n25836 ;
  assign n25838 = ~n3565 & n4526 ;
  assign n25839 = n25838 ^ n13659 ^ 1'b0 ;
  assign n25840 = ~n4916 & n15227 ;
  assign n25841 = n25840 ^ n8594 ^ 1'b0 ;
  assign n25842 = x63 & n1029 ;
  assign n25843 = n25841 & n25842 ;
  assign n25844 = n25843 ^ n7044 ^ 1'b0 ;
  assign n25845 = n22036 & n25844 ;
  assign n25846 = n6790 & n21177 ;
  assign n25847 = n25846 ^ n22125 ^ 1'b0 ;
  assign n25848 = n10878 & n25847 ;
  assign n25849 = n1761 | n14669 ;
  assign n25850 = n25849 ^ n10771 ^ 1'b0 ;
  assign n25853 = n5052 & ~n6028 ;
  assign n25854 = ~n9503 & n25853 ;
  assign n25851 = n9162 ^ n9002 ^ n8919 ;
  assign n25852 = n25851 ^ n8794 ^ 1'b0 ;
  assign n25855 = n25854 ^ n25852 ^ 1'b0 ;
  assign n25858 = ~n4282 & n15984 ;
  assign n25856 = n399 & n20650 ;
  assign n25857 = n6197 & n25856 ;
  assign n25859 = n25858 ^ n25857 ^ 1'b0 ;
  assign n25860 = n10355 | n25859 ;
  assign n25861 = n1085 & n23412 ;
  assign n25862 = n3387 & n20226 ;
  assign n25863 = n10660 ^ n950 ^ 1'b0 ;
  assign n25864 = n9239 ^ n1970 ^ 1'b0 ;
  assign n25865 = n5719 | n25864 ;
  assign n25866 = ( n6974 & n14806 ) | ( n6974 & ~n25865 ) | ( n14806 & ~n25865 ) ;
  assign n25867 = n908 & ~n4793 ;
  assign n25868 = ~n18388 & n25867 ;
  assign n25869 = ~n2262 & n4610 ;
  assign n25870 = n25869 ^ n8900 ^ 1'b0 ;
  assign n25871 = n1654 & n19560 ;
  assign n25872 = n8641 ^ n7099 ^ 1'b0 ;
  assign n25873 = n22420 & n25872 ;
  assign n25874 = n25873 ^ n2008 ^ 1'b0 ;
  assign n25875 = n1130 & n25874 ;
  assign n25876 = n22018 ^ n1481 ^ 1'b0 ;
  assign n25877 = n631 & n25876 ;
  assign n25878 = n6765 ^ n2836 ^ 1'b0 ;
  assign n25879 = n1706 | n18431 ;
  assign n25880 = n25879 ^ n17917 ^ n159 ;
  assign n25881 = ( n12776 & n21401 ) | ( n12776 & n25880 ) | ( n21401 & n25880 ) ;
  assign n25882 = n2222 & ~n6748 ;
  assign n25883 = n25882 ^ n4337 ^ 1'b0 ;
  assign n25884 = ~n9164 & n25883 ;
  assign n25885 = n25884 ^ n21003 ^ 1'b0 ;
  assign n25886 = ~n3361 & n25885 ;
  assign n25887 = n8261 & ~n11666 ;
  assign n25888 = n19423 & n25887 ;
  assign n25889 = n1867 | n15267 ;
  assign n25890 = ~n6617 & n17397 ;
  assign n25891 = ~n25889 & n25890 ;
  assign n25892 = n10668 ^ n1780 ^ 1'b0 ;
  assign n25893 = n7451 | n25892 ;
  assign n25894 = n25893 ^ n15580 ^ n5336 ;
  assign n25895 = n25894 ^ n5039 ^ n892 ;
  assign n25898 = n11406 | n21528 ;
  assign n25896 = n18029 ^ n1124 ^ 1'b0 ;
  assign n25897 = n3509 & ~n25896 ;
  assign n25899 = n25898 ^ n25897 ^ n1172 ;
  assign n25900 = n13946 ^ n6557 ^ 1'b0 ;
  assign n25901 = n13691 ^ n12149 ^ 1'b0 ;
  assign n25902 = n5562 | n25901 ;
  assign n25903 = n19262 ^ n336 ^ 1'b0 ;
  assign n25904 = n25902 | n25903 ;
  assign n25905 = n9176 ^ n2840 ^ n2422 ;
  assign n25906 = n8680 ^ n1613 ^ 1'b0 ;
  assign n25907 = n25905 & ~n25906 ;
  assign n25908 = n4314 | n24155 ;
  assign n25909 = n25642 | n25908 ;
  assign n25912 = ( n9977 & n13527 ) | ( n9977 & ~n18189 ) | ( n13527 & ~n18189 ) ;
  assign n25910 = n6162 ^ n4241 ^ 1'b0 ;
  assign n25911 = n8652 | n25910 ;
  assign n25913 = n25912 ^ n25911 ^ 1'b0 ;
  assign n25915 = n12659 ^ x3 ^ 1'b0 ;
  assign n25914 = ~n891 & n3245 ;
  assign n25916 = n25915 ^ n25914 ^ 1'b0 ;
  assign n25917 = n4202 & n21045 ;
  assign n25918 = n3556 ^ n1055 ^ 1'b0 ;
  assign n25919 = n6488 & ~n25918 ;
  assign n25920 = ~n5904 & n17908 ;
  assign n25921 = ( ~n3734 & n25919 ) | ( ~n3734 & n25920 ) | ( n25919 & n25920 ) ;
  assign n25922 = n4167 & n6030 ;
  assign n25923 = n3935 & n25922 ;
  assign n25924 = n6392 & ~n19903 ;
  assign n25925 = ( n3371 & ~n25923 ) | ( n3371 & n25924 ) | ( ~n25923 & n25924 ) ;
  assign n25926 = n6390 & ~n25621 ;
  assign n25927 = n25926 ^ n2790 ^ 1'b0 ;
  assign n25928 = n25927 ^ n17609 ^ n5281 ;
  assign n25930 = n12582 | n20179 ;
  assign n25931 = n21916 & ~n25930 ;
  assign n25929 = n1869 | n12475 ;
  assign n25932 = n25931 ^ n25929 ^ 1'b0 ;
  assign n25933 = n4674 & n14658 ;
  assign n25934 = n24665 & n25933 ;
  assign n25935 = n8917 ^ n980 ^ 1'b0 ;
  assign n25936 = ~n8187 & n25935 ;
  assign n25937 = n12469 | n17285 ;
  assign n25938 = ( ~n8899 & n9877 ) | ( ~n8899 & n25937 ) | ( n9877 & n25937 ) ;
  assign n25939 = n7733 & ~n25938 ;
  assign n25940 = n7439 & ~n20235 ;
  assign n25941 = n17587 ^ n13827 ^ 1'b0 ;
  assign n25942 = n16044 | n25941 ;
  assign n25943 = n25940 | n25942 ;
  assign n25944 = ~n2888 & n9933 ;
  assign n25945 = n11028 | n18648 ;
  assign n25946 = n25945 ^ n15754 ^ 1'b0 ;
  assign n25947 = n25946 ^ n9724 ^ n8885 ;
  assign n25948 = ( n1036 & n3626 ) | ( n1036 & n16805 ) | ( n3626 & n16805 ) ;
  assign n25949 = ~n6087 & n18556 ;
  assign n25950 = n13279 ^ n7902 ^ 1'b0 ;
  assign n25951 = n9085 & n25950 ;
  assign n25952 = n14793 ^ n9060 ^ n8786 ;
  assign n25953 = n25951 & n25952 ;
  assign n25954 = n3024 & n25953 ;
  assign n25955 = ~n3110 & n25954 ;
  assign n25956 = n1230 & n19318 ;
  assign n25957 = n12616 & ~n25956 ;
  assign n25958 = n11435 & n13525 ;
  assign n25959 = ~n842 & n25958 ;
  assign n25960 = n3315 & ~n7833 ;
  assign n25961 = n25960 ^ n8422 ^ 1'b0 ;
  assign n25962 = n25961 ^ n10946 ^ 1'b0 ;
  assign n25963 = n25959 | n25962 ;
  assign n25964 = n13252 ^ n1800 ^ n1791 ;
  assign n25965 = n2443 & ~n6700 ;
  assign n25966 = n25965 ^ n5955 ^ 1'b0 ;
  assign n25967 = n3499 & ~n25966 ;
  assign n25968 = n10108 & n25967 ;
  assign n25969 = ~n3006 & n25968 ;
  assign n25970 = n9573 & ~n25969 ;
  assign n25971 = n25964 & n25970 ;
  assign n25972 = n1451 | n25971 ;
  assign n25973 = ( n18057 & n23131 ) | ( n18057 & n25972 ) | ( n23131 & n25972 ) ;
  assign n25974 = n23181 ^ n8654 ^ 1'b0 ;
  assign n25975 = n5545 ^ n4736 ^ 1'b0 ;
  assign n25976 = n11269 | n25975 ;
  assign n25977 = n3292 & ~n25976 ;
  assign n25978 = n6874 ^ n707 ^ 1'b0 ;
  assign n25979 = n11080 | n21136 ;
  assign n25980 = n750 & n9971 ;
  assign n25981 = ( n6052 & ~n12074 ) | ( n6052 & n25980 ) | ( ~n12074 & n25980 ) ;
  assign n25982 = n1815 & n3172 ;
  assign n25983 = n5633 & n25982 ;
  assign n25984 = n13105 | n25983 ;
  assign n25985 = n6668 & ~n25984 ;
  assign n25986 = n3668 ^ n3076 ^ 1'b0 ;
  assign n25987 = n20127 | n25986 ;
  assign n25988 = n17032 ^ n8081 ^ 1'b0 ;
  assign n25989 = n5705 | n25988 ;
  assign n25990 = n12326 ^ n11020 ^ 1'b0 ;
  assign n25991 = n15306 & n25990 ;
  assign n25992 = n24174 ^ n14309 ^ n5925 ;
  assign n25993 = ~n3814 & n21499 ;
  assign n25994 = n3080 | n8185 ;
  assign n25995 = n25994 ^ n130 ^ 1'b0 ;
  assign n25996 = n8616 & ~n11263 ;
  assign n25997 = n10867 | n25996 ;
  assign n25998 = n25997 ^ n4902 ^ 1'b0 ;
  assign n25999 = n4450 & n7894 ;
  assign n26000 = n15773 ^ n15597 ^ 1'b0 ;
  assign n26001 = n1954 & ~n26000 ;
  assign n26002 = n9857 ^ n7385 ^ 1'b0 ;
  assign n26003 = n4736 | n9832 ;
  assign n26004 = ( n2553 & ~n4442 ) | ( n2553 & n12347 ) | ( ~n4442 & n12347 ) ;
  assign n26005 = ( n12296 & ~n22758 ) | ( n12296 & n26004 ) | ( ~n22758 & n26004 ) ;
  assign n26006 = ~n24123 & n26005 ;
  assign n26007 = ~n11057 & n26006 ;
  assign n26008 = n2254 | n6178 ;
  assign n26009 = n18091 | n26008 ;
  assign n26010 = x2 & n1439 ;
  assign n26011 = n7986 | n24614 ;
  assign n26012 = n11941 & n13856 ;
  assign n26013 = ~n26011 & n26012 ;
  assign n26014 = n1779 ^ x62 ^ 1'b0 ;
  assign n26015 = ~n1023 & n26014 ;
  assign n26016 = n26015 ^ n10881 ^ n7022 ;
  assign n26017 = n15591 ^ n8861 ^ 1'b0 ;
  assign n26018 = n18947 ^ n17735 ^ 1'b0 ;
  assign n26019 = n26018 ^ n17722 ^ n1680 ;
  assign n26020 = n1433 & n5647 ;
  assign n26021 = n6680 ^ n794 ^ 1'b0 ;
  assign n26022 = n16400 ^ n681 ^ 1'b0 ;
  assign n26023 = n243 | n11691 ;
  assign n26024 = n26023 ^ n15568 ^ 1'b0 ;
  assign n26025 = n2498 ^ n703 ^ n271 ;
  assign n26026 = ~n2419 & n15580 ;
  assign n26027 = n26026 ^ n19885 ^ 1'b0 ;
  assign n26028 = n1151 | n26027 ;
  assign n26029 = n17099 ^ n1743 ^ 1'b0 ;
  assign n26030 = ~n7352 & n15704 ;
  assign n26031 = n15887 & n26030 ;
  assign n26032 = ( n1833 & n2348 ) | ( n1833 & n17548 ) | ( n2348 & n17548 ) ;
  assign n26033 = n26032 ^ n907 ^ 1'b0 ;
  assign n26034 = n978 & n20710 ;
  assign n26035 = n4799 & ~n15222 ;
  assign n26036 = n4911 ^ n4094 ^ n2328 ;
  assign n26037 = n1033 & ~n26036 ;
  assign n26038 = n26037 ^ n323 ^ 1'b0 ;
  assign n26039 = n13545 ^ n8818 ^ 1'b0 ;
  assign n26040 = n26039 ^ n23418 ^ 1'b0 ;
  assign n26041 = n18459 ^ n8804 ^ 1'b0 ;
  assign n26042 = ~n4207 & n26041 ;
  assign n26043 = n4824 & ~n13553 ;
  assign n26044 = ~n26042 & n26043 ;
  assign n26045 = n7460 & ~n9630 ;
  assign n26046 = n750 | n13221 ;
  assign n26047 = n26046 ^ n24377 ^ 1'b0 ;
  assign n26048 = n191 & n26047 ;
  assign n26049 = n26045 & ~n26048 ;
  assign n26050 = n12869 & ~n15511 ;
  assign n26051 = ~n13025 & n26050 ;
  assign n26052 = n15477 ^ n1909 ^ 1'b0 ;
  assign n26053 = n1382 & ~n6156 ;
  assign n26054 = n10436 & ~n26053 ;
  assign n26055 = n26052 & n26054 ;
  assign n26056 = ( n4506 & n7295 ) | ( n4506 & ~n21388 ) | ( n7295 & ~n21388 ) ;
  assign n26057 = ( ~n11020 & n24149 ) | ( ~n11020 & n26056 ) | ( n24149 & n26056 ) ;
  assign n26058 = n17234 ^ n3559 ^ 1'b0 ;
  assign n26059 = n6135 | n26058 ;
  assign n26060 = n2021 & ~n4495 ;
  assign n26061 = n26060 ^ n8440 ^ 1'b0 ;
  assign n26062 = n4783 & n6789 ;
  assign n26063 = n26062 ^ n1974 ^ 1'b0 ;
  assign n26064 = ~n2157 & n26063 ;
  assign n26065 = n26064 ^ n479 ^ 1'b0 ;
  assign n26066 = n1188 | n17292 ;
  assign n26067 = n26065 | n26066 ;
  assign n26068 = n7969 & n21509 ;
  assign n26069 = n26068 ^ n2562 ^ 1'b0 ;
  assign n26070 = n19855 & n24174 ;
  assign n26071 = n22391 ^ n717 ^ 1'b0 ;
  assign n26072 = n6068 & ~n10198 ;
  assign n26073 = n8303 | n22273 ;
  assign n26074 = n26073 ^ n4373 ^ 1'b0 ;
  assign n26075 = n424 & ~n26074 ;
  assign n26076 = n10178 ^ n2236 ^ 1'b0 ;
  assign n26077 = n26075 & n26076 ;
  assign n26078 = n7047 | n26077 ;
  assign n26079 = ( ~n5470 & n5848 ) | ( ~n5470 & n12682 ) | ( n5848 & n12682 ) ;
  assign n26080 = ( ~n10147 & n22261 ) | ( ~n10147 & n26079 ) | ( n22261 & n26079 ) ;
  assign n26081 = ~n7547 & n15734 ;
  assign n26082 = ~n387 & n26081 ;
  assign n26083 = n7018 & ~n26082 ;
  assign n26085 = ~n11658 & n19199 ;
  assign n26086 = n26085 ^ n23274 ^ 1'b0 ;
  assign n26084 = n14179 | n14851 ;
  assign n26087 = n26086 ^ n26084 ^ 1'b0 ;
  assign n26088 = n5544 ^ n3192 ^ 1'b0 ;
  assign n26089 = n9703 & ~n26088 ;
  assign n26090 = n18115 ^ n2441 ^ 1'b0 ;
  assign n26091 = n16549 & ~n26090 ;
  assign n26092 = ~n26089 & n26091 ;
  assign n26093 = n9182 & n15512 ;
  assign n26094 = ~n3881 & n5832 ;
  assign n26095 = n10139 & ~n26094 ;
  assign n26096 = n26095 ^ n6566 ^ 1'b0 ;
  assign n26101 = n24928 ^ n10339 ^ 1'b0 ;
  assign n26097 = n510 | n3515 ;
  assign n26098 = n26097 ^ n2762 ^ 1'b0 ;
  assign n26099 = n26098 ^ n21066 ^ n11281 ;
  assign n26100 = n2063 & n26099 ;
  assign n26102 = n26101 ^ n26100 ^ 1'b0 ;
  assign n26103 = x9 & ~n5924 ;
  assign n26104 = n6360 & n26103 ;
  assign n26105 = ~n1578 & n10201 ;
  assign n26106 = ( n14069 & n23980 ) | ( n14069 & n26105 ) | ( n23980 & n26105 ) ;
  assign n26107 = n14432 ^ n5541 ^ 1'b0 ;
  assign n26108 = n8807 | n23487 ;
  assign n26109 = n26108 ^ n24463 ^ n9356 ;
  assign n26110 = n5051 & n11755 ;
  assign n26111 = n13760 ^ n4222 ^ 1'b0 ;
  assign n26112 = ~n21890 & n26111 ;
  assign n26114 = ( x80 & n8165 ) | ( x80 & ~n9596 ) | ( n8165 & ~n9596 ) ;
  assign n26113 = n8134 & ~n13733 ;
  assign n26115 = n26114 ^ n26113 ^ 1'b0 ;
  assign n26116 = ( n15172 & n18968 ) | ( n15172 & n26115 ) | ( n18968 & n26115 ) ;
  assign n26117 = n26116 ^ n14554 ^ 1'b0 ;
  assign n26118 = n23083 & n26117 ;
  assign n26119 = n8875 | n10774 ;
  assign n26120 = n4939 | n25440 ;
  assign n26121 = n26120 ^ n18530 ^ 1'b0 ;
  assign n26122 = n16081 & ~n26121 ;
  assign n26123 = ~n5874 & n10571 ;
  assign n26124 = n21688 ^ n1479 ^ 1'b0 ;
  assign n26125 = n14178 & ~n26124 ;
  assign n26126 = n14631 ^ n9513 ^ 1'b0 ;
  assign n26127 = n1264 ^ n725 ^ 1'b0 ;
  assign n26128 = n26126 & ~n26127 ;
  assign n26129 = n1283 & ~n16329 ;
  assign n26130 = n26129 ^ x119 ^ 1'b0 ;
  assign n26131 = n15530 ^ n9593 ^ 1'b0 ;
  assign n26132 = ( ~n1671 & n3315 ) | ( ~n1671 & n6190 ) | ( n3315 & n6190 ) ;
  assign n26133 = n12404 ^ n945 ^ 1'b0 ;
  assign n26134 = n8924 & ~n26133 ;
  assign n26135 = n5940 & ~n13819 ;
  assign n26136 = ~n13429 & n26135 ;
  assign n26137 = n26136 ^ n12109 ^ 1'b0 ;
  assign n26138 = n10377 ^ n8175 ^ 1'b0 ;
  assign n26139 = ~n8621 & n26138 ;
  assign n26140 = n20807 & n26139 ;
  assign n26141 = n7362 ^ n1585 ^ 1'b0 ;
  assign n26142 = ~n1877 & n26141 ;
  assign n26143 = n26142 ^ n411 ^ 1'b0 ;
  assign n26144 = n11493 | n26143 ;
  assign n26145 = n25378 ^ n9754 ^ 1'b0 ;
  assign n26146 = n17399 ^ n2896 ^ n1371 ;
  assign n26147 = n23421 ^ n1421 ^ n380 ;
  assign n26148 = n15015 ^ n5032 ^ 1'b0 ;
  assign n26149 = n7488 & n26148 ;
  assign n26150 = n6038 | n25046 ;
  assign n26151 = n25046 & ~n26150 ;
  assign n26152 = n26151 ^ n4213 ^ n3653 ;
  assign n26153 = n1477 | n26152 ;
  assign n26154 = n26153 ^ n11579 ^ 1'b0 ;
  assign n26155 = n26154 ^ n5081 ^ 1'b0 ;
  assign n26156 = n2772 & n26155 ;
  assign n26157 = ~n1959 & n26156 ;
  assign n26158 = n4156 & ~n4410 ;
  assign n26159 = ~n1680 & n25965 ;
  assign n26160 = n22179 ^ n271 ^ 1'b0 ;
  assign n26161 = n18240 ^ n4039 ^ 1'b0 ;
  assign n26162 = n2579 | n8905 ;
  assign n26163 = n2007 | n26162 ;
  assign n26164 = n6571 ^ n3545 ^ 1'b0 ;
  assign n26165 = n1660 | n26164 ;
  assign n26166 = n26165 ^ n13795 ^ 1'b0 ;
  assign n26167 = n25163 ^ n14815 ^ 1'b0 ;
  assign n26168 = n5474 & ~n22774 ;
  assign n26169 = n23352 ^ n19823 ^ 1'b0 ;
  assign n26170 = ~n8208 & n13048 ;
  assign n26171 = n26170 ^ n22784 ^ 1'b0 ;
  assign n26172 = n21503 & ~n23440 ;
  assign n26173 = ( n9002 & ~n26171 ) | ( n9002 & n26172 ) | ( ~n26171 & n26172 ) ;
  assign n26174 = n937 | n10442 ;
  assign n26175 = n26174 ^ n5958 ^ 1'b0 ;
  assign n26176 = ( n10491 & n21173 ) | ( n10491 & ~n26175 ) | ( n21173 & ~n26175 ) ;
  assign n26177 = n4686 & n6333 ;
  assign n26178 = ~n10109 & n26177 ;
  assign n26179 = n26178 ^ n25713 ^ n1610 ;
  assign n26180 = n18721 ^ n697 ^ 1'b0 ;
  assign n26181 = n138 & n14613 ;
  assign n26182 = n10293 & ~n20427 ;
  assign n26183 = n15882 & ~n26182 ;
  assign n26184 = n20064 ^ n13912 ^ 1'b0 ;
  assign n26185 = ~n12667 & n26184 ;
  assign n26186 = ( n2087 & n15050 ) | ( n2087 & n17292 ) | ( n15050 & n17292 ) ;
  assign n26187 = n9327 | n18615 ;
  assign n26188 = n26187 ^ n6687 ^ 1'b0 ;
  assign n26189 = ~n5257 & n26188 ;
  assign n26190 = ( n10259 & n15900 ) | ( n10259 & n19015 ) | ( n15900 & n19015 ) ;
  assign n26191 = ( n4291 & n26189 ) | ( n4291 & n26190 ) | ( n26189 & n26190 ) ;
  assign n26192 = n1082 | n13803 ;
  assign n26193 = n26192 ^ n14404 ^ n13252 ;
  assign n26194 = n18123 ^ n319 ^ 1'b0 ;
  assign n26195 = n19638 ^ n4354 ^ 1'b0 ;
  assign n26196 = n801 & ~n26195 ;
  assign n26197 = ~n3476 & n8002 ;
  assign n26198 = n15582 ^ n12291 ^ 1'b0 ;
  assign n26199 = n26197 & n26198 ;
  assign n26200 = n21088 & n24481 ;
  assign n26201 = n26200 ^ n9304 ^ 1'b0 ;
  assign n26202 = n18984 ^ n10094 ^ n5629 ;
  assign n26203 = n26202 ^ n3752 ^ 1'b0 ;
  assign n26204 = n13892 ^ n9663 ^ n2706 ;
  assign n26205 = n26204 ^ n13085 ^ 1'b0 ;
  assign n26206 = ( ~n3874 & n9800 ) | ( ~n3874 & n21730 ) | ( n9800 & n21730 ) ;
  assign n26207 = n11706 | n16214 ;
  assign n26208 = n26207 ^ n1467 ^ 1'b0 ;
  assign n26209 = n413 & ~n24273 ;
  assign n26210 = n8343 ^ n3756 ^ 1'b0 ;
  assign n26211 = n22269 & ~n26210 ;
  assign n26212 = n26211 ^ n16590 ^ 1'b0 ;
  assign n26213 = n5630 & ~n8135 ;
  assign n26214 = n2146 & n26213 ;
  assign n26215 = n1601 | n16415 ;
  assign n26216 = n26215 ^ n21986 ^ 1'b0 ;
  assign n26217 = n26214 | n26216 ;
  assign n26218 = ( n19452 & n23232 ) | ( n19452 & ~n26050 ) | ( n23232 & ~n26050 ) ;
  assign n26219 = n23334 ^ n21599 ^ n3247 ;
  assign n26220 = n6786 ^ n2335 ^ 1'b0 ;
  assign n26221 = ( ~n7117 & n10569 ) | ( ~n7117 & n26220 ) | ( n10569 & n26220 ) ;
  assign n26222 = ~n5070 & n20377 ;
  assign n26223 = ~n478 & n24032 ;
  assign n26224 = n26223 ^ n2355 ^ 1'b0 ;
  assign n26225 = n2162 | n7311 ;
  assign n26226 = ~n1632 & n5004 ;
  assign n26227 = n17504 | n26226 ;
  assign n26228 = ~n605 & n25678 ;
  assign n26229 = ~n14504 & n26228 ;
  assign n26230 = n9960 ^ n4853 ^ 1'b0 ;
  assign n26231 = ( n1243 & ~n10563 ) | ( n1243 & n26230 ) | ( ~n10563 & n26230 ) ;
  assign n26232 = n6093 & n26231 ;
  assign n26233 = n26232 ^ n14322 ^ 1'b0 ;
  assign n26234 = n26233 ^ n2550 ^ 1'b0 ;
  assign n26235 = n3185 & n5198 ;
  assign n26236 = n2064 | n8584 ;
  assign n26237 = ~n7979 & n24911 ;
  assign n26238 = ( n1521 & n26236 ) | ( n1521 & ~n26237 ) | ( n26236 & ~n26237 ) ;
  assign n26239 = n654 & ~n26238 ;
  assign n26240 = n25794 ^ n14346 ^ 1'b0 ;
  assign n26241 = ~n10057 & n26240 ;
  assign n26242 = n2747 ^ n393 ^ 1'b0 ;
  assign n26243 = n7488 & n26242 ;
  assign n26244 = n26243 ^ n11362 ^ 1'b0 ;
  assign n26245 = n1034 & ~n6050 ;
  assign n26246 = n6050 & n26245 ;
  assign n26247 = ~n265 & n26246 ;
  assign n26248 = n26247 ^ n19558 ^ 1'b0 ;
  assign n26249 = n26248 ^ n24362 ^ n11101 ;
  assign n26250 = x110 & ~n26249 ;
  assign n26251 = n20559 ^ n6038 ^ 1'b0 ;
  assign n26252 = n10868 | n26251 ;
  assign n26253 = n19345 ^ n2152 ^ 1'b0 ;
  assign n26254 = n26252 | n26253 ;
  assign n26255 = n7970 ^ n336 ^ 1'b0 ;
  assign n26256 = ~n24106 & n26255 ;
  assign n26257 = n26256 ^ n8420 ^ 1'b0 ;
  assign n26258 = n12092 & ~n14345 ;
  assign n26259 = n26258 ^ n21335 ^ 1'b0 ;
  assign n26260 = n16274 ^ n14331 ^ 1'b0 ;
  assign n26261 = n26260 ^ n14639 ^ n10693 ;
  assign n26262 = n11812 & n22190 ;
  assign n26264 = n3519 | n11304 ;
  assign n26263 = x113 & ~n15769 ;
  assign n26265 = n26264 ^ n26263 ^ 1'b0 ;
  assign n26266 = n10860 ^ n1413 ^ n805 ;
  assign n26267 = ( ~n11310 & n21038 ) | ( ~n11310 & n26266 ) | ( n21038 & n26266 ) ;
  assign n26268 = ( ~n1689 & n14322 ) | ( ~n1689 & n26267 ) | ( n14322 & n26267 ) ;
  assign n26269 = n26268 ^ n4363 ^ 1'b0 ;
  assign n26270 = n8887 ^ n7663 ^ n5736 ;
  assign n26271 = n26270 ^ n10833 ^ 1'b0 ;
  assign n26272 = n1156 | n8260 ;
  assign n26273 = n26272 ^ n7764 ^ 1'b0 ;
  assign n26274 = n16421 ^ n4893 ^ 1'b0 ;
  assign n26275 = n16524 | n26274 ;
  assign n26276 = n17181 & ~n26275 ;
  assign n26277 = n4017 ^ n802 ^ 1'b0 ;
  assign n26278 = n7189 ^ n2742 ^ 1'b0 ;
  assign n26279 = n26277 & n26278 ;
  assign n26280 = n6426 ^ n169 ^ 1'b0 ;
  assign n26281 = n26230 ^ n21263 ^ n6386 ;
  assign n26282 = ( n1826 & ~n1995 ) | ( n1826 & n26281 ) | ( ~n1995 & n26281 ) ;
  assign n26283 = n26282 ^ n319 ^ 1'b0 ;
  assign n26284 = n11713 & ~n22912 ;
  assign n26285 = x97 & ~n26284 ;
  assign n26286 = n14826 ^ n8038 ^ n5248 ;
  assign n26287 = n11435 ^ n6197 ^ 1'b0 ;
  assign n26288 = n1860 | n26287 ;
  assign n26289 = ( n1072 & n3714 ) | ( n1072 & ~n26288 ) | ( n3714 & ~n26288 ) ;
  assign n26290 = n26115 ^ n18572 ^ 1'b0 ;
  assign n26291 = ~n1413 & n16253 ;
  assign n26292 = n4358 & ~n26291 ;
  assign n26293 = n26292 ^ n11468 ^ 1'b0 ;
  assign n26294 = n4273 | n9448 ;
  assign n26295 = n26293 & ~n26294 ;
  assign n26297 = ~n14504 & n17834 ;
  assign n26296 = ~n12081 & n16246 ;
  assign n26298 = n26297 ^ n26296 ^ 1'b0 ;
  assign n26299 = n22374 | n25614 ;
  assign n26300 = n26299 ^ n16202 ^ 1'b0 ;
  assign n26301 = n849 | n15584 ;
  assign n26302 = n26301 ^ n6888 ^ 1'b0 ;
  assign n26303 = n13859 & n24179 ;
  assign n26304 = ~n3959 & n26303 ;
  assign n26305 = n1684 ^ n632 ^ 1'b0 ;
  assign n26306 = n18446 ^ n13321 ^ n6782 ;
  assign n26307 = ( n6063 & n10682 ) | ( n6063 & ~n26306 ) | ( n10682 & ~n26306 ) ;
  assign n26308 = ( n2918 & n6102 ) | ( n2918 & ~n13246 ) | ( n6102 & ~n13246 ) ;
  assign n26309 = n25787 ^ n18029 ^ n13429 ;
  assign n26310 = ( ~n2200 & n6128 ) | ( ~n2200 & n7094 ) | ( n6128 & n7094 ) ;
  assign n26311 = n25442 & n26310 ;
  assign n26312 = n8491 | n9471 ;
  assign n26313 = n593 & n9630 ;
  assign n26314 = n5928 | n25927 ;
  assign n26315 = n21386 & n23285 ;
  assign n26316 = n22574 | n25614 ;
  assign n26317 = n26316 ^ n6939 ^ 1'b0 ;
  assign n26318 = ( n561 & n4085 ) | ( n561 & n6597 ) | ( n4085 & n6597 ) ;
  assign n26319 = n26318 ^ n22635 ^ n16245 ;
  assign n26320 = n17063 | n26319 ;
  assign n26321 = n26320 ^ n730 ^ 1'b0 ;
  assign n26322 = ~n15616 & n24082 ;
  assign n26323 = n10173 ^ n8276 ^ 1'b0 ;
  assign n26324 = n23294 ^ n10194 ^ 1'b0 ;
  assign n26325 = n7345 | n26324 ;
  assign n26326 = ~n4044 & n4353 ;
  assign n26327 = n26325 | n26326 ;
  assign n26328 = n5085 & n22852 ;
  assign n26329 = n26328 ^ n9432 ^ 1'b0 ;
  assign n26330 = n12037 | n15507 ;
  assign n26331 = n8509 | n26330 ;
  assign n26332 = ~n9728 & n22700 ;
  assign n26333 = n26332 ^ n348 ^ 1'b0 ;
  assign n26334 = ~n5871 & n24967 ;
  assign n26335 = n10388 ^ n10028 ^ 1'b0 ;
  assign n26336 = n3589 | n26335 ;
  assign n26337 = n10373 | n13886 ;
  assign n26338 = n26337 ^ n11300 ^ 1'b0 ;
  assign n26339 = ( n7681 & n12344 ) | ( n7681 & ~n22787 ) | ( n12344 & ~n22787 ) ;
  assign n26340 = ( n352 & n1366 ) | ( n352 & ~n23865 ) | ( n1366 & ~n23865 ) ;
  assign n26341 = n6061 & ~n24648 ;
  assign n26342 = n16674 | n20336 ;
  assign n26343 = n6707 & ~n26342 ;
  assign n26344 = n4822 & n12709 ;
  assign n26345 = n26343 & n26344 ;
  assign n26346 = n26345 ^ n23913 ^ 1'b0 ;
  assign n26347 = n26341 | n26346 ;
  assign n26348 = n4768 & ~n18628 ;
  assign n26349 = n26348 ^ n5347 ^ 1'b0 ;
  assign n26350 = n265 & n5557 ;
  assign n26351 = n3975 & ~n26350 ;
  assign n26352 = ~n8007 & n8568 ;
  assign n26353 = n13501 & n26352 ;
  assign n26354 = n14320 | n26353 ;
  assign n26355 = n14640 & ~n26354 ;
  assign n26356 = n8788 ^ n7476 ^ n415 ;
  assign n26357 = n14354 & n15768 ;
  assign n26358 = n1513 & n9237 ;
  assign n26359 = n14895 & n26358 ;
  assign n26360 = ~n1013 & n26359 ;
  assign n26361 = ( n5141 & n10902 ) | ( n5141 & n26360 ) | ( n10902 & n26360 ) ;
  assign n26362 = n11556 ^ n1022 ^ 1'b0 ;
  assign n26363 = n6977 & ~n26362 ;
  assign n26364 = n26363 ^ n8609 ^ 1'b0 ;
  assign n26366 = n8903 ^ n7850 ^ 1'b0 ;
  assign n26365 = n3125 & ~n16645 ;
  assign n26367 = n26366 ^ n26365 ^ 1'b0 ;
  assign n26368 = n950 & n23875 ;
  assign n26369 = n26368 ^ n3471 ^ 1'b0 ;
  assign n26371 = n18050 ^ n1740 ^ 1'b0 ;
  assign n26372 = n9798 & n26371 ;
  assign n26370 = n7558 & ~n9898 ;
  assign n26373 = n26372 ^ n26370 ^ 1'b0 ;
  assign n26374 = n14432 | n18765 ;
  assign n26375 = n17067 ^ n4090 ^ n2268 ;
  assign n26376 = n4721 & ~n10799 ;
  assign n26377 = ~n26375 & n26376 ;
  assign n26378 = n6456 & ~n23096 ;
  assign n26379 = n17337 ^ n13454 ^ 1'b0 ;
  assign n26380 = n26378 & ~n26379 ;
  assign n26381 = n3015 & n26380 ;
  assign n26382 = n21538 ^ n17910 ^ 1'b0 ;
  assign n26383 = n975 | n17067 ;
  assign n26384 = n1064 & ~n26383 ;
  assign n26385 = n4500 & ~n14729 ;
  assign n26386 = n26385 ^ n7193 ^ 1'b0 ;
  assign n26387 = ~n11172 & n26386 ;
  assign n26388 = ~n8840 & n26387 ;
  assign n26389 = n1972 ^ x56 ^ 1'b0 ;
  assign n26390 = ~n7471 & n26389 ;
  assign n26391 = n9008 ^ n4932 ^ n4038 ;
  assign n26392 = ~n7298 & n17020 ;
  assign n26393 = n26392 ^ n15432 ^ 1'b0 ;
  assign n26394 = n26393 ^ n20711 ^ 1'b0 ;
  assign n26395 = ( n7185 & ~n7218 ) | ( n7185 & n8778 ) | ( ~n7218 & n8778 ) ;
  assign n26396 = n26395 ^ n1553 ^ 1'b0 ;
  assign n26397 = ( n3979 & n5989 ) | ( n3979 & ~n7604 ) | ( n5989 & ~n7604 ) ;
  assign n26398 = n26397 ^ n4893 ^ 1'b0 ;
  assign n26399 = n19574 ^ n13747 ^ 1'b0 ;
  assign n26400 = ~n11344 & n26399 ;
  assign n26401 = n26400 ^ n4023 ^ 1'b0 ;
  assign n26402 = n8824 & n26401 ;
  assign n26403 = n7813 ^ n4382 ^ 1'b0 ;
  assign n26404 = n473 & ~n2842 ;
  assign n26405 = n26404 ^ n23871 ^ 1'b0 ;
  assign n26406 = n3547 | n26405 ;
  assign n26407 = n13687 & ~n20291 ;
  assign n26408 = ( n4027 & n4936 ) | ( n4027 & n23210 ) | ( n4936 & n23210 ) ;
  assign n26409 = n17882 ^ n4283 ^ 1'b0 ;
  assign n26410 = n7471 & n26409 ;
  assign n26411 = n22287 ^ n9974 ^ n3285 ;
  assign n26412 = ~n3073 & n20330 ;
  assign n26413 = n10347 & n26412 ;
  assign n26414 = n14808 ^ n11281 ^ x6 ;
  assign n26415 = n17739 | n26414 ;
  assign n26416 = n1983 & ~n2817 ;
  assign n26417 = ~n17239 & n26416 ;
  assign n26418 = n6856 & ~n26417 ;
  assign n26419 = n26418 ^ n23558 ^ 1'b0 ;
  assign n26420 = n26419 ^ n3815 ^ 1'b0 ;
  assign n26421 = ( n1034 & ~n5989 ) | ( n1034 & n10439 ) | ( ~n5989 & n10439 ) ;
  assign n26422 = ( ~n4863 & n19661 ) | ( ~n4863 & n26421 ) | ( n19661 & n26421 ) ;
  assign n26423 = n26422 ^ n14957 ^ 1'b0 ;
  assign n26424 = ( n706 & ~n3723 ) | ( n706 & n8091 ) | ( ~n3723 & n8091 ) ;
  assign n26425 = n14233 & n26424 ;
  assign n26426 = ~n1454 & n26425 ;
  assign n26428 = n1962 & ~n8481 ;
  assign n26429 = n26428 ^ n2786 ^ 1'b0 ;
  assign n26427 = ( n593 & n10747 ) | ( n593 & n19045 ) | ( n10747 & n19045 ) ;
  assign n26430 = n26429 ^ n26427 ^ n7819 ;
  assign n26431 = n6948 | n17805 ;
  assign n26432 = n1423 & ~n26431 ;
  assign n26433 = ~n17089 & n26432 ;
  assign n26434 = n12309 ^ n10048 ^ 1'b0 ;
  assign n26435 = n1017 & ~n11691 ;
  assign n26436 = ~n4432 & n26435 ;
  assign n26437 = n10414 | n26436 ;
  assign n26438 = n4169 ^ n3181 ^ n2087 ;
  assign n26439 = n23273 ^ n10366 ^ 1'b0 ;
  assign n26440 = n17759 ^ n5911 ^ 1'b0 ;
  assign n26441 = ~n26439 & n26440 ;
  assign n26442 = n21885 ^ n7503 ^ n1930 ;
  assign n26443 = n929 & ~n7786 ;
  assign n26444 = n26443 ^ n17261 ^ 1'b0 ;
  assign n26445 = n16485 ^ n8563 ^ 1'b0 ;
  assign n26446 = n26444 | n26445 ;
  assign n26447 = ( n166 & n26442 ) | ( n166 & n26446 ) | ( n26442 & n26446 ) ;
  assign n26448 = n14666 ^ n11863 ^ 1'b0 ;
  assign n26449 = ~n26447 & n26448 ;
  assign n26450 = n925 & n8306 ;
  assign n26451 = ~n2266 & n13135 ;
  assign n26452 = n26450 & n26451 ;
  assign n26453 = ( n1297 & n15356 ) | ( n1297 & ~n26452 ) | ( n15356 & ~n26452 ) ;
  assign n26454 = n10738 ^ n740 ^ 1'b0 ;
  assign n26455 = n5883 ^ n3994 ^ 1'b0 ;
  assign n26456 = n7579 & n11941 ;
  assign n26457 = n26456 ^ n23871 ^ 1'b0 ;
  assign n26458 = n6511 & ~n15440 ;
  assign n26459 = n26458 ^ n9511 ^ n3881 ;
  assign n26460 = n6753 | n15580 ;
  assign n26461 = n14719 & ~n26460 ;
  assign n26462 = n4252 & n20713 ;
  assign n26463 = n6870 & n26462 ;
  assign n26464 = n7994 & n26463 ;
  assign n26465 = n4219 & n4893 ;
  assign n26466 = n26465 ^ n1680 ^ 1'b0 ;
  assign n26467 = n4847 & n26466 ;
  assign n26468 = ( n26461 & n26464 ) | ( n26461 & ~n26467 ) | ( n26464 & ~n26467 ) ;
  assign n26469 = ~n12691 & n26468 ;
  assign n26470 = ~n4972 & n26469 ;
  assign n26471 = n26470 ^ n17315 ^ 1'b0 ;
  assign n26472 = n26459 | n26471 ;
  assign n26473 = n21401 ^ n14458 ^ 1'b0 ;
  assign n26475 = n1277 | n2701 ;
  assign n26476 = n26475 ^ n2346 ^ 1'b0 ;
  assign n26477 = ~n3073 & n24125 ;
  assign n26478 = ~n15524 & n26477 ;
  assign n26479 = n21552 | n26478 ;
  assign n26480 = n26479 ^ n6265 ^ 1'b0 ;
  assign n26481 = ( ~n8537 & n26476 ) | ( ~n8537 & n26480 ) | ( n26476 & n26480 ) ;
  assign n26482 = n788 & n26481 ;
  assign n26483 = n26482 ^ n938 ^ 1'b0 ;
  assign n26474 = n5531 ^ n1484 ^ 1'b0 ;
  assign n26484 = n26483 ^ n26474 ^ 1'b0 ;
  assign n26485 = n15424 ^ n6330 ^ 1'b0 ;
  assign n26486 = ~n12932 & n26485 ;
  assign n26488 = n4623 & n25673 ;
  assign n26489 = n26488 ^ n8655 ^ 1'b0 ;
  assign n26490 = ~n1918 & n7104 ;
  assign n26491 = n26489 & n26490 ;
  assign n26487 = n398 & ~n763 ;
  assign n26492 = n26491 ^ n26487 ^ 1'b0 ;
  assign n26493 = n14965 ^ n8751 ^ 1'b0 ;
  assign n26494 = n2873 & n26493 ;
  assign n26495 = ~n1452 & n10016 ;
  assign n26496 = n1507 | n25339 ;
  assign n26497 = n4406 & ~n25196 ;
  assign n26498 = n26497 ^ n1724 ^ 1'b0 ;
  assign n26499 = ~n11731 & n26498 ;
  assign n26500 = n16679 & n17146 ;
  assign n26501 = ~n3076 & n20267 ;
  assign n26502 = n19161 ^ n15719 ^ 1'b0 ;
  assign n26504 = n20775 ^ n8892 ^ n893 ;
  assign n26503 = n6007 & n17139 ;
  assign n26505 = n26504 ^ n26503 ^ 1'b0 ;
  assign n26506 = n1248 | n26505 ;
  assign n26507 = n6049 | n16857 ;
  assign n26508 = n3982 & ~n26507 ;
  assign n26509 = n26508 ^ n11663 ^ 1'b0 ;
  assign n26510 = n10876 ^ n5594 ^ 1'b0 ;
  assign n26511 = n2190 | n26510 ;
  assign n26512 = n4836 & n9798 ;
  assign n26513 = n26512 ^ n21992 ^ 1'b0 ;
  assign n26514 = n12969 ^ n2929 ^ 1'b0 ;
  assign n26515 = ~n8479 & n26514 ;
  assign n26516 = n26513 | n26515 ;
  assign n26517 = ( x78 & n5456 ) | ( x78 & n6448 ) | ( n5456 & n6448 ) ;
  assign n26518 = n17394 ^ n5778 ^ 1'b0 ;
  assign n26519 = n897 & ~n26518 ;
  assign n26520 = n26519 ^ n5398 ^ 1'b0 ;
  assign n26521 = n26517 & ~n26520 ;
  assign n26523 = n16686 ^ n871 ^ 1'b0 ;
  assign n26524 = ( n3315 & ~n20807 ) | ( n3315 & n26523 ) | ( ~n20807 & n26523 ) ;
  assign n26522 = n16034 ^ n9442 ^ n4308 ;
  assign n26525 = n26524 ^ n26522 ^ 1'b0 ;
  assign n26526 = ( n14314 & n25744 ) | ( n14314 & ~n26525 ) | ( n25744 & ~n26525 ) ;
  assign n26527 = n21181 ^ n18934 ^ n245 ;
  assign n26528 = n7824 & ~n11149 ;
  assign n26529 = n141 & n26528 ;
  assign n26530 = n16643 & n26529 ;
  assign n26531 = n24204 ^ n21876 ^ 1'b0 ;
  assign n26532 = n419 & ~n26531 ;
  assign n26533 = n12055 ^ n10751 ^ 1'b0 ;
  assign n26534 = n15453 ^ n4880 ^ n1607 ;
  assign n26535 = n6336 & ~n26534 ;
  assign n26536 = n25446 ^ n1089 ^ n505 ;
  assign n26537 = n4112 & n26536 ;
  assign n26539 = n19507 | n25429 ;
  assign n26538 = n3286 & n25938 ;
  assign n26540 = n26539 ^ n26538 ^ 1'b0 ;
  assign n26541 = n668 & n819 ;
  assign n26542 = n26541 ^ n11778 ^ 1'b0 ;
  assign n26543 = n26542 ^ n23703 ^ n9840 ;
  assign n26544 = n16662 ^ n16099 ^ 1'b0 ;
  assign n26545 = ~n8341 & n9225 ;
  assign n26546 = n26545 ^ n2272 ^ 1'b0 ;
  assign n26547 = n26546 ^ n13302 ^ 1'b0 ;
  assign n26548 = n20370 | n26547 ;
  assign n26549 = ~n2020 & n9007 ;
  assign n26550 = n10871 & n26549 ;
  assign n26552 = n9518 ^ n4964 ^ 1'b0 ;
  assign n26551 = n8347 | n17002 ;
  assign n26553 = n26552 ^ n26551 ^ 1'b0 ;
  assign n26554 = n2552 & ~n5223 ;
  assign n26555 = n26554 ^ n10709 ^ 1'b0 ;
  assign n26556 = n1175 | n26555 ;
  assign n26557 = n26556 ^ n16508 ^ n4654 ;
  assign n26558 = n20836 ^ n11819 ^ n3428 ;
  assign n26559 = n15554 ^ n5261 ^ n1758 ;
  assign n26560 = n2999 | n7197 ;
  assign n26561 = n654 | n26560 ;
  assign n26562 = n18398 ^ n11241 ^ 1'b0 ;
  assign n26563 = n2942 ^ n381 ^ 1'b0 ;
  assign n26564 = n21168 ^ n17305 ^ 1'b0 ;
  assign n26565 = n14360 & n26564 ;
  assign n26566 = n26565 ^ n2120 ^ 1'b0 ;
  assign n26567 = n25786 ^ n11607 ^ 1'b0 ;
  assign n26568 = n4745 | n9516 ;
  assign n26569 = n25029 ^ n9686 ^ 1'b0 ;
  assign n26570 = n15100 ^ n2602 ^ 1'b0 ;
  assign n26571 = n26569 & ~n26570 ;
  assign n26572 = n4100 & n8697 ;
  assign n26573 = n26571 & ~n26572 ;
  assign n26577 = n8136 ^ n4576 ^ 1'b0 ;
  assign n26578 = n1022 | n26577 ;
  assign n26574 = ( n1393 & n2782 ) | ( n1393 & ~n6367 ) | ( n2782 & ~n6367 ) ;
  assign n26575 = ~n22318 & n26574 ;
  assign n26576 = ~n4557 & n26575 ;
  assign n26579 = n26578 ^ n26576 ^ 1'b0 ;
  assign n26585 = n26404 ^ n1842 ^ 1'b0 ;
  assign n26586 = n19084 ^ n12534 ^ 1'b0 ;
  assign n26587 = n26585 & n26586 ;
  assign n26580 = n2552 & ~n16415 ;
  assign n26581 = n26580 ^ n17315 ^ 1'b0 ;
  assign n26582 = n2016 & n8828 ;
  assign n26583 = n26582 ^ n21867 ^ 1'b0 ;
  assign n26584 = ( n5850 & ~n26581 ) | ( n5850 & n26583 ) | ( ~n26581 & n26583 ) ;
  assign n26588 = n26587 ^ n26584 ^ 1'b0 ;
  assign n26589 = ( n2063 & n2717 ) | ( n2063 & n23334 ) | ( n2717 & n23334 ) ;
  assign n26590 = n14937 & n26589 ;
  assign n26591 = n7294 & n22616 ;
  assign n26592 = n10317 & n26591 ;
  assign n26593 = n10435 ^ n8054 ^ 1'b0 ;
  assign n26594 = n11755 ^ n6378 ^ 1'b0 ;
  assign n26595 = n25455 ^ n7680 ^ n521 ;
  assign n26596 = n14238 & n26595 ;
  assign n26597 = ~n9216 & n26596 ;
  assign n26598 = n26594 | n26597 ;
  assign n26599 = n939 | n7625 ;
  assign n26600 = n26599 ^ n11739 ^ 1'b0 ;
  assign n26601 = n15640 ^ n13819 ^ 1'b0 ;
  assign n26602 = ~n4235 & n26601 ;
  assign n26603 = n24017 ^ n17311 ^ 1'b0 ;
  assign n26604 = n19935 | n26603 ;
  assign n26605 = n4361 ^ n2701 ^ 1'b0 ;
  assign n26606 = n16454 & n26605 ;
  assign n26607 = ( n5712 & n14433 ) | ( n5712 & ~n25092 ) | ( n14433 & ~n25092 ) ;
  assign n26608 = n3966 ^ n3415 ^ 1'b0 ;
  assign n26609 = ~n2049 & n5185 ;
  assign n26610 = n26609 ^ n5186 ^ 1'b0 ;
  assign n26611 = n26610 ^ n13947 ^ 1'b0 ;
  assign n26612 = ( ~n21144 & n26608 ) | ( ~n21144 & n26611 ) | ( n26608 & n26611 ) ;
  assign n26613 = n14889 ^ n3783 ^ 1'b0 ;
  assign n26614 = n7286 | n13207 ;
  assign n26615 = ~n12823 & n23245 ;
  assign n26616 = ~n20066 & n26615 ;
  assign n26617 = ~n886 & n11094 ;
  assign n26618 = n19751 | n26617 ;
  assign n26619 = n9779 | n26618 ;
  assign n26620 = n5359 ^ n1309 ^ 1'b0 ;
  assign n26621 = n26620 ^ n16742 ^ n11900 ;
  assign n26622 = n332 & n26621 ;
  assign n26623 = n21988 & ~n26622 ;
  assign n26624 = n4410 & n12282 ;
  assign n26625 = n8424 | n15157 ;
  assign n26628 = n1677 ^ n1350 ^ 1'b0 ;
  assign n26629 = n2112 | n26628 ;
  assign n26626 = n16706 ^ n5548 ^ 1'b0 ;
  assign n26627 = n8826 & n26626 ;
  assign n26630 = n26629 ^ n26627 ^ n13810 ;
  assign n26631 = n26380 ^ n5618 ^ n884 ;
  assign n26632 = ( ~x24 & n19830 ) | ( ~x24 & n26631 ) | ( n19830 & n26631 ) ;
  assign n26633 = ~n10910 & n11262 ;
  assign n26634 = n26633 ^ n1171 ^ 1'b0 ;
  assign n26635 = n17858 ^ n3475 ^ 1'b0 ;
  assign n26636 = ~n26634 & n26635 ;
  assign n26637 = n9013 ^ n4208 ^ 1'b0 ;
  assign n26638 = n14686 ^ n314 ^ 1'b0 ;
  assign n26639 = n893 & n24447 ;
  assign n26640 = n7161 ^ n6204 ^ 1'b0 ;
  assign n26641 = ~n17799 & n26640 ;
  assign n26642 = ~n11378 & n14569 ;
  assign n26643 = x23 & n6829 ;
  assign n26644 = n26643 ^ x9 ^ 1'b0 ;
  assign n26645 = ( n6700 & n20668 ) | ( n6700 & ~n26644 ) | ( n20668 & ~n26644 ) ;
  assign n26646 = n4498 & n26645 ;
  assign n26647 = n1520 & n1792 ;
  assign n26648 = ~n1792 & n26647 ;
  assign n26649 = n11569 & ~n14280 ;
  assign n26650 = n22494 & n26649 ;
  assign n26651 = n26650 ^ n4016 ^ 1'b0 ;
  assign n26652 = ~n26648 & n26651 ;
  assign n26653 = n21668 ^ n15598 ^ 1'b0 ;
  assign n26654 = n6241 | n26653 ;
  assign n26655 = n8302 ^ n1714 ^ 1'b0 ;
  assign n26656 = n19064 | n24731 ;
  assign n26657 = n26470 ^ n3589 ^ 1'b0 ;
  assign n26658 = n15111 ^ n2814 ^ 1'b0 ;
  assign n26659 = n18663 | n26658 ;
  assign n26660 = ~n8936 & n19460 ;
  assign n26661 = n26660 ^ n20837 ^ 1'b0 ;
  assign n26662 = n26659 & ~n26661 ;
  assign n26663 = n10788 & n26662 ;
  assign n26664 = n12863 ^ n12420 ^ n12169 ;
  assign n26665 = n4654 & ~n26664 ;
  assign n26666 = n26665 ^ n3788 ^ 1'b0 ;
  assign n26667 = n3585 & ~n10783 ;
  assign n26668 = n26667 ^ n8536 ^ 1'b0 ;
  assign n26669 = n1118 & n19051 ;
  assign n26670 = n5092 & n26669 ;
  assign n26671 = ( x84 & ~n1958 ) | ( x84 & n4362 ) | ( ~n1958 & n4362 ) ;
  assign n26672 = n15696 | n26671 ;
  assign n26673 = n12281 | n26672 ;
  assign n26674 = n1683 | n21031 ;
  assign n26675 = n26673 | n26674 ;
  assign n26677 = n10071 ^ n3079 ^ 1'b0 ;
  assign n26678 = n25961 & ~n26677 ;
  assign n26676 = ( ~n2765 & n10066 ) | ( ~n2765 & n26510 ) | ( n10066 & n26510 ) ;
  assign n26679 = n26678 ^ n26676 ^ n5012 ;
  assign n26680 = n17279 ^ n3576 ^ 1'b0 ;
  assign n26681 = n1161 & ~n26680 ;
  assign n26682 = ( n18685 & n24716 ) | ( n18685 & ~n26681 ) | ( n24716 & ~n26681 ) ;
  assign n26683 = ~n17701 & n23308 ;
  assign n26684 = n8512 ^ n2335 ^ 1'b0 ;
  assign n26685 = n7101 ^ n2983 ^ 1'b0 ;
  assign n26686 = ~n22594 & n26685 ;
  assign n26687 = n11536 & ~n26686 ;
  assign n26688 = n7093 & ~n7370 ;
  assign n26689 = n18163 ^ n2404 ^ 1'b0 ;
  assign n26690 = n26688 | n26689 ;
  assign n26691 = ( n5314 & n19938 ) | ( n5314 & n26690 ) | ( n19938 & n26690 ) ;
  assign n26693 = ( ~n3482 & n8455 ) | ( ~n3482 & n16467 ) | ( n8455 & n16467 ) ;
  assign n26692 = n7758 ^ n2619 ^ 1'b0 ;
  assign n26694 = n26693 ^ n26692 ^ n26595 ;
  assign n26695 = ~n5018 & n22156 ;
  assign n26696 = ~n2496 & n17842 ;
  assign n26697 = n4906 ^ n3355 ^ 1'b0 ;
  assign n26698 = n18530 & ~n26697 ;
  assign n26699 = n9226 & ~n23994 ;
  assign n26700 = n2999 | n13274 ;
  assign n26701 = n671 | n26700 ;
  assign n26702 = n22053 & n26701 ;
  assign n26703 = ~n26699 & n26702 ;
  assign n26704 = n26703 ^ x93 ^ 1'b0 ;
  assign n26705 = n26704 ^ n20397 ^ 1'b0 ;
  assign n26706 = n26698 & n26705 ;
  assign n26707 = n25825 ^ n17603 ^ 1'b0 ;
  assign n26708 = n1858 & ~n6482 ;
  assign n26709 = n15725 & n26708 ;
  assign n26710 = n1521 & ~n26709 ;
  assign n26711 = n3012 | n10099 ;
  assign n26712 = n26711 ^ n2929 ^ 1'b0 ;
  assign n26713 = n26712 ^ n6138 ^ 1'b0 ;
  assign n26714 = n1623 & ~n26713 ;
  assign n26715 = n26714 ^ n8152 ^ 1'b0 ;
  assign n26716 = n7444 ^ n6049 ^ 1'b0 ;
  assign n26717 = n1624 & n26716 ;
  assign n26718 = n26717 ^ n9064 ^ 1'b0 ;
  assign n26719 = ~n14287 & n26718 ;
  assign n26720 = n13356 ^ n10054 ^ 1'b0 ;
  assign n26721 = ~n10677 & n14723 ;
  assign n26722 = n22657 ^ n2005 ^ n1761 ;
  assign n26723 = n632 & n20793 ;
  assign n26724 = n8638 ^ n5077 ^ 1'b0 ;
  assign n26725 = n19946 & ~n26724 ;
  assign n26726 = n6998 ^ n3020 ^ 1'b0 ;
  assign n26727 = n196 & n26726 ;
  assign n26728 = n597 & ~n7740 ;
  assign n26729 = n26728 ^ n8994 ^ 1'b0 ;
  assign n26730 = n10451 & ~n26729 ;
  assign n26731 = n3440 & n26730 ;
  assign n26732 = ~n6899 & n16987 ;
  assign n26733 = ~n23474 & n26732 ;
  assign n26736 = n3206 | n5656 ;
  assign n26737 = n18663 & ~n26736 ;
  assign n26735 = ~n12279 & n23173 ;
  assign n26738 = n26737 ^ n26735 ^ 1'b0 ;
  assign n26734 = n9639 & ~n13756 ;
  assign n26739 = n26738 ^ n26734 ^ 1'b0 ;
  assign n26740 = ( ~n15013 & n26733 ) | ( ~n15013 & n26739 ) | ( n26733 & n26739 ) ;
  assign n26741 = n673 & ~n4938 ;
  assign n26742 = n26741 ^ n22819 ^ 1'b0 ;
  assign n26743 = n5303 ^ n3972 ^ 1'b0 ;
  assign n26744 = n2606 ^ n2289 ^ 1'b0 ;
  assign n26745 = n1307 | n13248 ;
  assign n26746 = n26745 ^ n18062 ^ n4084 ;
  assign n26747 = ~n7627 & n12004 ;
  assign n26748 = ~n26746 & n26747 ;
  assign n26749 = n1072 & n8038 ;
  assign n26750 = n5002 | n9747 ;
  assign n26751 = ( n17799 & n21776 ) | ( n17799 & ~n26750 ) | ( n21776 & ~n26750 ) ;
  assign n26752 = n11402 ^ n6496 ^ 1'b0 ;
  assign n26753 = n7587 & ~n8536 ;
  assign n26754 = n26753 ^ n12864 ^ n2839 ;
  assign n26755 = n23209 & n26754 ;
  assign n26756 = n7909 ^ n692 ^ 1'b0 ;
  assign n26757 = ~n21357 & n26756 ;
  assign n26758 = n17818 ^ n3340 ^ 1'b0 ;
  assign n26759 = n10002 ^ n2987 ^ 1'b0 ;
  assign n26760 = n26758 & ~n26759 ;
  assign n26761 = n20127 ^ n6261 ^ n1888 ;
  assign n26762 = n10788 & n26761 ;
  assign n26763 = n26762 ^ n3321 ^ 1'b0 ;
  assign n26764 = ~n11921 & n23442 ;
  assign n26765 = n11203 ^ n7785 ^ n3149 ;
  assign n26766 = n4006 & ~n26765 ;
  assign n26767 = n9063 | n9571 ;
  assign n26768 = n15812 | n26767 ;
  assign n26769 = n1476 & n26768 ;
  assign n26770 = ~n26766 & n26769 ;
  assign n26771 = n26770 ^ n20639 ^ n18464 ;
  assign n26772 = n11010 ^ n9496 ^ n9037 ;
  assign n26773 = ~n2642 & n20437 ;
  assign n26774 = ~n14439 & n26773 ;
  assign n26775 = x38 & n490 ;
  assign n26776 = ~n6984 & n26775 ;
  assign n26777 = n7196 ^ n1808 ^ 1'b0 ;
  assign n26778 = x74 & n26777 ;
  assign n26779 = ~n12566 & n26778 ;
  assign n26780 = n13307 & n26779 ;
  assign n26781 = n6487 & ~n18698 ;
  assign n26782 = n12362 | n26755 ;
  assign n26783 = n26782 ^ n8786 ^ 1'b0 ;
  assign n26784 = n4957 | n5659 ;
  assign n26785 = n12588 | n26784 ;
  assign n26786 = ~n8890 & n26785 ;
  assign n26787 = n22594 & n26786 ;
  assign n26788 = n8586 ^ n7967 ^ n7575 ;
  assign n26789 = n6117 ^ n1860 ^ 1'b0 ;
  assign n26790 = ~n4684 & n26789 ;
  assign n26791 = n3181 | n26790 ;
  assign n26792 = ( ~n1967 & n2350 ) | ( ~n1967 & n19187 ) | ( n2350 & n19187 ) ;
  assign n26793 = n11792 & ~n26664 ;
  assign n26794 = n26793 ^ n9448 ^ 1'b0 ;
  assign n26795 = n5061 & ~n22112 ;
  assign n26796 = ~n26794 & n26795 ;
  assign n26797 = ~n8481 & n16295 ;
  assign n26798 = n26797 ^ n906 ^ 1'b0 ;
  assign n26799 = n24138 & ~n25188 ;
  assign n26800 = ~n24312 & n26799 ;
  assign n26801 = n26798 & n26800 ;
  assign n26802 = n18266 ^ n8354 ^ 1'b0 ;
  assign n26803 = n19097 & n26802 ;
  assign n26804 = n12927 | n13111 ;
  assign n26805 = n26804 ^ n6076 ^ 1'b0 ;
  assign n26806 = n722 & n1684 ;
  assign n26807 = n13903 ^ n8345 ^ 1'b0 ;
  assign n26808 = n26806 & n26807 ;
  assign n26809 = n26808 ^ n13229 ^ 1'b0 ;
  assign n26810 = n21962 ^ n14601 ^ 1'b0 ;
  assign n26811 = ~n2583 & n24536 ;
  assign n26812 = ( n14312 & n26810 ) | ( n14312 & n26811 ) | ( n26810 & n26811 ) ;
  assign n26813 = n17577 ^ n3315 ^ n2750 ;
  assign n26814 = ~n2341 & n3831 ;
  assign n26815 = n26814 ^ n14267 ^ 1'b0 ;
  assign n26816 = n577 & n5901 ;
  assign n26817 = ~n26815 & n26816 ;
  assign n26818 = n4433 & ~n17365 ;
  assign n26819 = n26818 ^ n9598 ^ 1'b0 ;
  assign n26823 = n3030 | n15540 ;
  assign n26824 = n26823 ^ n3447 ^ 1'b0 ;
  assign n26825 = n17795 & ~n26824 ;
  assign n26826 = ~n1892 & n26825 ;
  assign n26820 = n15500 ^ n8278 ^ 1'b0 ;
  assign n26821 = n10817 & ~n26820 ;
  assign n26822 = ~n24318 & n26821 ;
  assign n26827 = n26826 ^ n26822 ^ 1'b0 ;
  assign n26828 = ~n5292 & n10188 ;
  assign n26829 = n26828 ^ n7714 ^ 1'b0 ;
  assign n26830 = n22457 ^ n15847 ^ n5381 ;
  assign n26831 = n1592 | n21453 ;
  assign n26832 = n5824 | n26831 ;
  assign n26833 = n7029 & n12921 ;
  assign n26834 = n26833 ^ n25236 ^ 1'b0 ;
  assign y0 = x0 ;
  assign y1 = x1 ;
  assign y2 = x15 ;
  assign y3 = x17 ;
  assign y4 = x22 ;
  assign y5 = x27 ;
  assign y6 = x30 ;
  assign y7 = x32 ;
  assign y8 = x44 ;
  assign y9 = x52 ;
  assign y10 = x53 ;
  assign y11 = x66 ;
  assign y12 = x73 ;
  assign y13 = x77 ;
  assign y14 = x79 ;
  assign y15 = x90 ;
  assign y16 = x96 ;
  assign y17 = x104 ;
  assign y18 = x111 ;
  assign y19 = x113 ;
  assign y20 = x124 ;
  assign y21 = x125 ;
  assign y22 = x127 ;
  assign y23 = n129 ;
  assign y24 = n130 ;
  assign y25 = ~1'b0 ;
  assign y26 = n132 ;
  assign y27 = ~1'b0 ;
  assign y28 = n134 ;
  assign y29 = n138 ;
  assign y30 = ~n142 ;
  assign y31 = n143 ;
  assign y32 = n145 ;
  assign y33 = n146 ;
  assign y34 = ~n148 ;
  assign y35 = ~n149 ;
  assign y36 = ~1'b0 ;
  assign y37 = ~1'b0 ;
  assign y38 = ~n155 ;
  assign y39 = n156 ;
  assign y40 = ~n158 ;
  assign y41 = ~n165 ;
  assign y42 = ~n169 ;
  assign y43 = n173 ;
  assign y44 = ~n174 ;
  assign y45 = n175 ;
  assign y46 = ~n177 ;
  assign y47 = ~n179 ;
  assign y48 = n183 ;
  assign y49 = ~n186 ;
  assign y50 = ~n189 ;
  assign y51 = n194 ;
  assign y52 = 1'b0 ;
  assign y53 = n197 ;
  assign y54 = ~n199 ;
  assign y55 = ~1'b0 ;
  assign y56 = ~n202 ;
  assign y57 = ~1'b0 ;
  assign y58 = n210 ;
  assign y59 = ~n212 ;
  assign y60 = ~n215 ;
  assign y61 = n216 ;
  assign y62 = ~n217 ;
  assign y63 = n218 ;
  assign y64 = n223 ;
  assign y65 = ~n225 ;
  assign y66 = ~n231 ;
  assign y67 = ~n240 ;
  assign y68 = n241 ;
  assign y69 = ~n243 ;
  assign y70 = n245 ;
  assign y71 = n252 ;
  assign y72 = ~n254 ;
  assign y73 = n257 ;
  assign y74 = ~n259 ;
  assign y75 = ~n260 ;
  assign y76 = n261 ;
  assign y77 = n262 ;
  assign y78 = ~n267 ;
  assign y79 = ~n275 ;
  assign y80 = n279 ;
  assign y81 = n280 ;
  assign y82 = ~1'b0 ;
  assign y83 = n282 ;
  assign y84 = ~n290 ;
  assign y85 = ~n301 ;
  assign y86 = n309 ;
  assign y87 = ~1'b0 ;
  assign y88 = ~x110 ;
  assign y89 = ~n310 ;
  assign y90 = n312 ;
  assign y91 = ~n316 ;
  assign y92 = n325 ;
  assign y93 = n335 ;
  assign y94 = ~n340 ;
  assign y95 = ~n348 ;
  assign y96 = ~n349 ;
  assign y97 = ~n350 ;
  assign y98 = ~n357 ;
  assign y99 = ~n361 ;
  assign y100 = n362 ;
  assign y101 = ~n363 ;
  assign y102 = ~1'b0 ;
  assign y103 = ~1'b0 ;
  assign y104 = n367 ;
  assign y105 = n371 ;
  assign y106 = ~1'b0 ;
  assign y107 = ~n372 ;
  assign y108 = ~1'b0 ;
  assign y109 = ~1'b0 ;
  assign y110 = ~1'b0 ;
  assign y111 = ~1'b0 ;
  assign y112 = n376 ;
  assign y113 = n380 ;
  assign y114 = ~n381 ;
  assign y115 = n386 ;
  assign y116 = n387 ;
  assign y117 = ~1'b0 ;
  assign y118 = ~1'b0 ;
  assign y119 = n390 ;
  assign y120 = n391 ;
  assign y121 = ~n396 ;
  assign y122 = ~n399 ;
  assign y123 = n401 ;
  assign y124 = ~1'b0 ;
  assign y125 = ~1'b0 ;
  assign y126 = n406 ;
  assign y127 = ~n409 ;
  assign y128 = n410 ;
  assign y129 = ~1'b0 ;
  assign y130 = ~n411 ;
  assign y131 = n419 ;
  assign y132 = n422 ;
  assign y133 = n424 ;
  assign y134 = n429 ;
  assign y135 = ~n438 ;
  assign y136 = n210 ;
  assign y137 = ~n443 ;
  assign y138 = ~n449 ;
  assign y139 = ~1'b0 ;
  assign y140 = n337 ;
  assign y141 = n451 ;
  assign y142 = ~1'b0 ;
  assign y143 = ~n456 ;
  assign y144 = n462 ;
  assign y145 = n463 ;
  assign y146 = ~n467 ;
  assign y147 = n470 ;
  assign y148 = ~n471 ;
  assign y149 = n380 ;
  assign y150 = ~n475 ;
  assign y151 = n478 ;
  assign y152 = ~n479 ;
  assign y153 = n484 ;
  assign y154 = ~1'b0 ;
  assign y155 = ~n485 ;
  assign y156 = ~n486 ;
  assign y157 = n490 ;
  assign y158 = n493 ;
  assign y159 = n497 ;
  assign y160 = ~n498 ;
  assign y161 = ~1'b0 ;
  assign y162 = ~n503 ;
  assign y163 = n507 ;
  assign y164 = n509 ;
  assign y165 = ~n515 ;
  assign y166 = n521 ;
  assign y167 = ~n523 ;
  assign y168 = ~1'b0 ;
  assign y169 = ~n526 ;
  assign y170 = ~1'b0 ;
  assign y171 = n530 ;
  assign y172 = ~n533 ;
  assign y173 = n538 ;
  assign y174 = n539 ;
  assign y175 = ~n541 ;
  assign y176 = n549 ;
  assign y177 = ~n555 ;
  assign y178 = n566 ;
  assign y179 = ~1'b0 ;
  assign y180 = ~1'b0 ;
  assign y181 = n577 ;
  assign y182 = ~n578 ;
  assign y183 = ~n579 ;
  assign y184 = n582 ;
  assign y185 = ~n590 ;
  assign y186 = ~1'b0 ;
  assign y187 = n593 ;
  assign y188 = ~n599 ;
  assign y189 = ~1'b0 ;
  assign y190 = ~n601 ;
  assign y191 = n603 ;
  assign y192 = ~1'b0 ;
  assign y193 = ~n606 ;
  assign y194 = ~1'b0 ;
  assign y195 = ~1'b0 ;
  assign y196 = 1'b0 ;
  assign y197 = n612 ;
  assign y198 = ~n616 ;
  assign y199 = n619 ;
  assign y200 = ~1'b0 ;
  assign y201 = n621 ;
  assign y202 = ~n632 ;
  assign y203 = ~n633 ;
  assign y204 = n636 ;
  assign y205 = n643 ;
  assign y206 = ~1'b0 ;
  assign y207 = ~1'b0 ;
  assign y208 = n644 ;
  assign y209 = ~n645 ;
  assign y210 = n646 ;
  assign y211 = ~n650 ;
  assign y212 = ~n654 ;
  assign y213 = n655 ;
  assign y214 = 1'b0 ;
  assign y215 = ~n664 ;
  assign y216 = ~n665 ;
  assign y217 = ~n667 ;
  assign y218 = n671 ;
  assign y219 = ~1'b0 ;
  assign y220 = n672 ;
  assign y221 = ~n677 ;
  assign y222 = n678 ;
  assign y223 = n681 ;
  assign y224 = ~1'b0 ;
  assign y225 = ~n688 ;
  assign y226 = n690 ;
  assign y227 = ~n694 ;
  assign y228 = ~1'b0 ;
  assign y229 = ~n697 ;
  assign y230 = n702 ;
  assign y231 = ~1'b0 ;
  assign y232 = n713 ;
  assign y233 = n719 ;
  assign y234 = ~n725 ;
  assign y235 = n726 ;
  assign y236 = ~n729 ;
  assign y237 = ~n731 ;
  assign y238 = ~n738 ;
  assign y239 = n422 ;
  assign y240 = ~1'b0 ;
  assign y241 = n739 ;
  assign y242 = ~n745 ;
  assign y243 = n758 ;
  assign y244 = ~n760 ;
  assign y245 = ~n763 ;
  assign y246 = n767 ;
  assign y247 = n777 ;
  assign y248 = ~n786 ;
  assign y249 = n788 ;
  assign y250 = ~n790 ;
  assign y251 = ~n798 ;
  assign y252 = n799 ;
  assign y253 = n802 ;
  assign y254 = n804 ;
  assign y255 = ~n808 ;
  assign y256 = ~n811 ;
  assign y257 = ~1'b0 ;
  assign y258 = n817 ;
  assign y259 = ~n821 ;
  assign y260 = ~1'b0 ;
  assign y261 = ~n824 ;
  assign y262 = ~1'b0 ;
  assign y263 = ~1'b0 ;
  assign y264 = n138 ;
  assign y265 = n826 ;
  assign y266 = n829 ;
  assign y267 = ~1'b0 ;
  assign y268 = ~1'b0 ;
  assign y269 = ~n830 ;
  assign y270 = n831 ;
  assign y271 = ~n832 ;
  assign y272 = ~1'b0 ;
  assign y273 = n836 ;
  assign y274 = ~n837 ;
  assign y275 = ~1'b0 ;
  assign y276 = ~1'b0 ;
  assign y277 = 1'b0 ;
  assign y278 = n840 ;
  assign y279 = ~n842 ;
  assign y280 = n844 ;
  assign y281 = ~n859 ;
  assign y282 = n867 ;
  assign y283 = n869 ;
  assign y284 = ~1'b0 ;
  assign y285 = ~n876 ;
  assign y286 = ~n877 ;
  assign y287 = ~n881 ;
  assign y288 = n882 ;
  assign y289 = n888 ;
  assign y290 = n890 ;
  assign y291 = ~1'b0 ;
  assign y292 = ~1'b0 ;
  assign y293 = n895 ;
  assign y294 = n897 ;
  assign y295 = n901 ;
  assign y296 = ~1'b0 ;
  assign y297 = n906 ;
  assign y298 = n907 ;
  assign y299 = ~n910 ;
  assign y300 = n914 ;
  assign y301 = n925 ;
  assign y302 = ~1'b0 ;
  assign y303 = n927 ;
  assign y304 = ~n928 ;
  assign y305 = ~n937 ;
  assign y306 = ~1'b0 ;
  assign y307 = n939 ;
  assign y308 = ~n942 ;
  assign y309 = ~1'b0 ;
  assign y310 = ~n943 ;
  assign y311 = ~n945 ;
  assign y312 = n950 ;
  assign y313 = ~1'b0 ;
  assign y314 = ~n953 ;
  assign y315 = n955 ;
  assign y316 = ~1'b0 ;
  assign y317 = ~n956 ;
  assign y318 = ~n740 ;
  assign y319 = n957 ;
  assign y320 = ~n959 ;
  assign y321 = n962 ;
  assign y322 = n671 ;
  assign y323 = n964 ;
  assign y324 = ~n967 ;
  assign y325 = ~n972 ;
  assign y326 = ~n975 ;
  assign y327 = ~n570 ;
  assign y328 = ~n977 ;
  assign y329 = ~1'b0 ;
  assign y330 = ~n982 ;
  assign y331 = ~1'b0 ;
  assign y332 = ~n983 ;
  assign y333 = ~n988 ;
  assign y334 = 1'b0 ;
  assign y335 = ~n990 ;
  assign y336 = n664 ;
  assign y337 = ~n997 ;
  assign y338 = ~n998 ;
  assign y339 = n1001 ;
  assign y340 = ~n1004 ;
  assign y341 = ~n282 ;
  assign y342 = n1009 ;
  assign y343 = n1010 ;
  assign y344 = ~n1013 ;
  assign y345 = ~1'b0 ;
  assign y346 = n1017 ;
  assign y347 = n1025 ;
  assign y348 = ~1'b0 ;
  assign y349 = n1026 ;
  assign y350 = ~n1027 ;
  assign y351 = n1030 ;
  assign y352 = ~n1031 ;
  assign y353 = n1036 ;
  assign y354 = ~n1044 ;
  assign y355 = n1050 ;
  assign y356 = ~n1051 ;
  assign y357 = ~n581 ;
  assign y358 = n1053 ;
  assign y359 = ~n1054 ;
  assign y360 = ~1'b0 ;
  assign y361 = n1057 ;
  assign y362 = ~n1065 ;
  assign y363 = n1070 ;
  assign y364 = n1074 ;
  assign y365 = n1075 ;
  assign y366 = n1085 ;
  assign y367 = ~1'b0 ;
  assign y368 = n1089 ;
  assign y369 = ~n1092 ;
  assign y370 = ~n1094 ;
  assign y371 = x3 ;
  assign y372 = n1100 ;
  assign y373 = ~n1101 ;
  assign y374 = n1103 ;
  assign y375 = n1104 ;
  assign y376 = ~1'b0 ;
  assign y377 = ~1'b0 ;
  assign y378 = ~1'b0 ;
  assign y379 = ~n1113 ;
  assign y380 = ~1'b0 ;
  assign y381 = ~1'b0 ;
  assign y382 = ~1'b0 ;
  assign y383 = n1117 ;
  assign y384 = ~1'b0 ;
  assign y385 = ~n1124 ;
  assign y386 = ~1'b0 ;
  assign y387 = ~1'b0 ;
  assign y388 = n1134 ;
  assign y389 = ~n1138 ;
  assign y390 = n1139 ;
  assign y391 = ~1'b0 ;
  assign y392 = ~1'b0 ;
  assign y393 = n1140 ;
  assign y394 = n1141 ;
  assign y395 = ~n1145 ;
  assign y396 = n1147 ;
  assign y397 = n1153 ;
  assign y398 = n1154 ;
  assign y399 = n1159 ;
  assign y400 = ~n1160 ;
  assign y401 = ~1'b0 ;
  assign y402 = ~1'b0 ;
  assign y403 = n1162 ;
  assign y404 = 1'b0 ;
  assign y405 = 1'b0 ;
  assign y406 = n1165 ;
  assign y407 = n1168 ;
  assign y408 = ~n1171 ;
  assign y409 = ~n1181 ;
  assign y410 = ~n1182 ;
  assign y411 = ~n1185 ;
  assign y412 = n1186 ;
  assign y413 = ~1'b0 ;
  assign y414 = ~1'b0 ;
  assign y415 = n516 ;
  assign y416 = ~n1188 ;
  assign y417 = ~n1196 ;
  assign y418 = ~n1197 ;
  assign y419 = ~n1202 ;
  assign y420 = ~n1208 ;
  assign y421 = ~1'b0 ;
  assign y422 = ~n1219 ;
  assign y423 = ~n1224 ;
  assign y424 = ~n1226 ;
  assign y425 = n1231 ;
  assign y426 = ~n1234 ;
  assign y427 = n1235 ;
  assign y428 = n1236 ;
  assign y429 = ~1'b0 ;
  assign y430 = ~1'b0 ;
  assign y431 = ~n1240 ;
  assign y432 = ~n1245 ;
  assign y433 = n1246 ;
  assign y434 = n1251 ;
  assign y435 = n1253 ;
  assign y436 = ~n1256 ;
  assign y437 = ~n1258 ;
  assign y438 = ~n1260 ;
  assign y439 = ~1'b0 ;
  assign y440 = n1263 ;
  assign y441 = n1265 ;
  assign y442 = ~n1269 ;
  assign y443 = n1271 ;
  assign y444 = n582 ;
  assign y445 = ~1'b0 ;
  assign y446 = ~n1273 ;
  assign y447 = n1276 ;
  assign y448 = ~n1278 ;
  assign y449 = n1279 ;
  assign y450 = n1281 ;
  assign y451 = n1283 ;
  assign y452 = n1293 ;
  assign y453 = ~n1300 ;
  assign y454 = ~n1302 ;
  assign y455 = n1311 ;
  assign y456 = n1313 ;
  assign y457 = n1319 ;
  assign y458 = n1320 ;
  assign y459 = n1321 ;
  assign y460 = ~n1323 ;
  assign y461 = ~n1329 ;
  assign y462 = n1330 ;
  assign y463 = ~n1337 ;
  assign y464 = ~1'b0 ;
  assign y465 = ~1'b0 ;
  assign y466 = ~1'b0 ;
  assign y467 = ~1'b0 ;
  assign y468 = n1338 ;
  assign y469 = n1339 ;
  assign y470 = n1342 ;
  assign y471 = 1'b0 ;
  assign y472 = ~1'b0 ;
  assign y473 = ~n1347 ;
  assign y474 = n1348 ;
  assign y475 = ~n1350 ;
  assign y476 = n1352 ;
  assign y477 = ~n1354 ;
  assign y478 = ~n1360 ;
  assign y479 = ~n1365 ;
  assign y480 = ~n1368 ;
  assign y481 = ~1'b0 ;
  assign y482 = ~n1370 ;
  assign y483 = ~n1375 ;
  assign y484 = ~1'b0 ;
  assign y485 = ~n1376 ;
  assign y486 = ~n1382 ;
  assign y487 = n1387 ;
  assign y488 = n1388 ;
  assign y489 = ~n1392 ;
  assign y490 = n1394 ;
  assign y491 = n1397 ;
  assign y492 = ~1'b0 ;
  assign y493 = ~n1401 ;
  assign y494 = ~1'b0 ;
  assign y495 = ~n1403 ;
  assign y496 = ~1'b0 ;
  assign y497 = ~1'b0 ;
  assign y498 = ~n1405 ;
  assign y499 = ~1'b0 ;
  assign y500 = n1406 ;
  assign y501 = ~n1411 ;
  assign y502 = n1415 ;
  assign y503 = ~n1418 ;
  assign y504 = n1422 ;
  assign y505 = ~n1423 ;
  assign y506 = n1424 ;
  assign y507 = ~n1425 ;
  assign y508 = n1428 ;
  assign y509 = ~1'b0 ;
  assign y510 = ~n1430 ;
  assign y511 = ~n1433 ;
  assign y512 = ~1'b0 ;
  assign y513 = n1434 ;
  assign y514 = ~n1438 ;
  assign y515 = ~1'b0 ;
  assign y516 = ~n1439 ;
  assign y517 = ~n1446 ;
  assign y518 = ~n1451 ;
  assign y519 = ~n1461 ;
  assign y520 = ~1'b0 ;
  assign y521 = n1463 ;
  assign y522 = n1471 ;
  assign y523 = n1472 ;
  assign y524 = ~n1475 ;
  assign y525 = n1476 ;
  assign y526 = ~n1477 ;
  assign y527 = n1481 ;
  assign y528 = n1484 ;
  assign y529 = ~n1486 ;
  assign y530 = ~n1490 ;
  assign y531 = n1500 ;
  assign y532 = ~1'b0 ;
  assign y533 = n1501 ;
  assign y534 = n671 ;
  assign y535 = n1503 ;
  assign y536 = n706 ;
  assign y537 = ~1'b0 ;
  assign y538 = ~n1504 ;
  assign y539 = ~n1507 ;
  assign y540 = n1513 ;
  assign y541 = n1516 ;
  assign y542 = ~1'b0 ;
  assign y543 = ~n1519 ;
  assign y544 = n1522 ;
  assign y545 = ~n1526 ;
  assign y546 = n1527 ;
  assign y547 = ~1'b0 ;
  assign y548 = ~1'b0 ;
  assign y549 = ~1'b0 ;
  assign y550 = n1528 ;
  assign y551 = n1532 ;
  assign y552 = n1534 ;
  assign y553 = ~1'b0 ;
  assign y554 = ~n1535 ;
  assign y555 = n1537 ;
  assign y556 = ~1'b0 ;
  assign y557 = ~n1540 ;
  assign y558 = ~1'b0 ;
  assign y559 = ~n1547 ;
  assign y560 = n1552 ;
  assign y561 = n1555 ;
  assign y562 = n1561 ;
  assign y563 = n1562 ;
  assign y564 = n1565 ;
  assign y565 = 1'b0 ;
  assign y566 = ~n1570 ;
  assign y567 = n1575 ;
  assign y568 = ~1'b0 ;
  assign y569 = ~1'b0 ;
  assign y570 = ~n1582 ;
  assign y571 = n1586 ;
  assign y572 = ~n1588 ;
  assign y573 = ~1'b0 ;
  assign y574 = n1590 ;
  assign y575 = ~n1597 ;
  assign y576 = ~n1601 ;
  assign y577 = n1609 ;
  assign y578 = ~n1610 ;
  assign y579 = ~n1613 ;
  assign y580 = n1614 ;
  assign y581 = ~n1617 ;
  assign y582 = n1623 ;
  assign y583 = ~1'b0 ;
  assign y584 = n1628 ;
  assign y585 = n1630 ;
  assign y586 = n1631 ;
  assign y587 = ~n1632 ;
  assign y588 = ~n1634 ;
  assign y589 = ~n1639 ;
  assign y590 = n1644 ;
  assign y591 = ~n1646 ;
  assign y592 = ~1'b0 ;
  assign y593 = n1650 ;
  assign y594 = n1652 ;
  assign y595 = ~n1654 ;
  assign y596 = ~1'b0 ;
  assign y597 = n1655 ;
  assign y598 = ~n1656 ;
  assign y599 = ~n1660 ;
  assign y600 = ~n1661 ;
  assign y601 = ~x3 ;
  assign y602 = ~1'b0 ;
  assign y603 = n1666 ;
  assign y604 = ~n1667 ;
  assign y605 = n1670 ;
  assign y606 = ~1'b0 ;
  assign y607 = n1079 ;
  assign y608 = n1673 ;
  assign y609 = n1679 ;
  assign y610 = n1682 ;
  assign y611 = ~n1684 ;
  assign y612 = ~1'b0 ;
  assign y613 = 1'b0 ;
  assign y614 = ~n1687 ;
  assign y615 = ~1'b0 ;
  assign y616 = 1'b0 ;
  assign y617 = ~n1692 ;
  assign y618 = ~n1695 ;
  assign y619 = ~n1705 ;
  assign y620 = n1708 ;
  assign y621 = n1710 ;
  assign y622 = ~n1713 ;
  assign y623 = n370 ;
  assign y624 = n1714 ;
  assign y625 = ~n1716 ;
  assign y626 = ~n1718 ;
  assign y627 = ~1'b0 ;
  assign y628 = ~n1721 ;
  assign y629 = n1722 ;
  assign y630 = ~1'b0 ;
  assign y631 = ~1'b0 ;
  assign y632 = n1726 ;
  assign y633 = n1732 ;
  assign y634 = n1734 ;
  assign y635 = n1736 ;
  assign y636 = n1374 ;
  assign y637 = n1739 ;
  assign y638 = n1741 ;
  assign y639 = n1745 ;
  assign y640 = ~n1747 ;
  assign y641 = n1749 ;
  assign y642 = n1752 ;
  assign y643 = ~n1753 ;
  assign y644 = n1760 ;
  assign y645 = n1762 ;
  assign y646 = ~n1769 ;
  assign y647 = ~1'b0 ;
  assign y648 = ~1'b0 ;
  assign y649 = ~n1772 ;
  assign y650 = ~n1774 ;
  assign y651 = ~1'b0 ;
  assign y652 = n1776 ;
  assign y653 = ~1'b0 ;
  assign y654 = ~n1777 ;
  assign y655 = ~n1781 ;
  assign y656 = ~1'b0 ;
  assign y657 = ~n1785 ;
  assign y658 = ~n1786 ;
  assign y659 = ~1'b0 ;
  assign y660 = n1788 ;
  assign y661 = ~n1236 ;
  assign y662 = n886 ;
  assign y663 = n1791 ;
  assign y664 = n1798 ;
  assign y665 = ~n1799 ;
  assign y666 = ~n1808 ;
  assign y667 = ~n1811 ;
  assign y668 = ~1'b0 ;
  assign y669 = ~1'b0 ;
  assign y670 = ~n1813 ;
  assign y671 = ~n1817 ;
  assign y672 = ~n1818 ;
  assign y673 = n234 ;
  assign y674 = n1821 ;
  assign y675 = ~n1823 ;
  assign y676 = ~1'b0 ;
  assign y677 = n1265 ;
  assign y678 = n1826 ;
  assign y679 = ~1'b0 ;
  assign y680 = ~n909 ;
  assign y681 = n1828 ;
  assign y682 = ~n1835 ;
  assign y683 = n1839 ;
  assign y684 = n1847 ;
  assign y685 = n1851 ;
  assign y686 = n1853 ;
  assign y687 = ~n1855 ;
  assign y688 = ~1'b0 ;
  assign y689 = ~1'b0 ;
  assign y690 = n1861 ;
  assign y691 = n1864 ;
  assign y692 = ~1'b0 ;
  assign y693 = ~n1866 ;
  assign y694 = n1870 ;
  assign y695 = ~1'b0 ;
  assign y696 = n1871 ;
  assign y697 = ~1'b0 ;
  assign y698 = ~n1872 ;
  assign y699 = ~n1879 ;
  assign y700 = ~n1880 ;
  assign y701 = n1884 ;
  assign y702 = ~n1885 ;
  assign y703 = ~n1886 ;
  assign y704 = n1887 ;
  assign y705 = ~1'b0 ;
  assign y706 = ~1'b0 ;
  assign y707 = ~n1899 ;
  assign y708 = ~n1901 ;
  assign y709 = ~n1907 ;
  assign y710 = n161 ;
  assign y711 = ~1'b0 ;
  assign y712 = n1909 ;
  assign y713 = ~1'b0 ;
  assign y714 = n1912 ;
  assign y715 = ~1'b0 ;
  assign y716 = ~n1917 ;
  assign y717 = ~1'b0 ;
  assign y718 = ~1'b0 ;
  assign y719 = ~1'b0 ;
  assign y720 = ~n1924 ;
  assign y721 = ~n1925 ;
  assign y722 = n1931 ;
  assign y723 = ~n1935 ;
  assign y724 = n1938 ;
  assign y725 = n1939 ;
  assign y726 = n1941 ;
  assign y727 = ~1'b0 ;
  assign y728 = ~n612 ;
  assign y729 = ~1'b0 ;
  assign y730 = n1943 ;
  assign y731 = n1944 ;
  assign y732 = n1946 ;
  assign y733 = n1948 ;
  assign y734 = n1958 ;
  assign y735 = ~n1963 ;
  assign y736 = ~n1970 ;
  assign y737 = ~n1971 ;
  assign y738 = n1972 ;
  assign y739 = n1977 ;
  assign y740 = n1981 ;
  assign y741 = ~n1982 ;
  assign y742 = ~1'b0 ;
  assign y743 = n1983 ;
  assign y744 = ~n1989 ;
  assign y745 = ~1'b0 ;
  assign y746 = ~n1585 ;
  assign y747 = ~n1990 ;
  assign y748 = n1992 ;
  assign y749 = n1997 ;
  assign y750 = n1999 ;
  assign y751 = ~1'b0 ;
  assign y752 = ~1'b0 ;
  assign y753 = ~1'b0 ;
  assign y754 = ~1'b0 ;
  assign y755 = ~n2003 ;
  assign y756 = ~n2006 ;
  assign y757 = ~1'b0 ;
  assign y758 = ~1'b0 ;
  assign y759 = ~1'b0 ;
  assign y760 = ~n2007 ;
  assign y761 = n2008 ;
  assign y762 = ~n2011 ;
  assign y763 = ~1'b0 ;
  assign y764 = n2014 ;
  assign y765 = ~1'b0 ;
  assign y766 = ~n2015 ;
  assign y767 = n2019 ;
  assign y768 = ~1'b0 ;
  assign y769 = ~1'b0 ;
  assign y770 = ~n2021 ;
  assign y771 = ~1'b0 ;
  assign y772 = ~n2022 ;
  assign y773 = ~1'b0 ;
  assign y774 = n2023 ;
  assign y775 = ~1'b0 ;
  assign y776 = ~1'b0 ;
  assign y777 = ~1'b0 ;
  assign y778 = 1'b0 ;
  assign y779 = ~1'b0 ;
  assign y780 = ~1'b0 ;
  assign y781 = n336 ;
  assign y782 = n2026 ;
  assign y783 = ~n2027 ;
  assign y784 = n2028 ;
  assign y785 = n2035 ;
  assign y786 = ~n2036 ;
  assign y787 = ~n2039 ;
  assign y788 = ~1'b0 ;
  assign y789 = n2040 ;
  assign y790 = ~1'b0 ;
  assign y791 = ~1'b0 ;
  assign y792 = ~n2045 ;
  assign y793 = ~1'b0 ;
  assign y794 = n2048 ;
  assign y795 = n2049 ;
  assign y796 = ~n2062 ;
  assign y797 = ~n2063 ;
  assign y798 = n2065 ;
  assign y799 = ~1'b0 ;
  assign y800 = ~n2066 ;
  assign y801 = n2069 ;
  assign y802 = ~1'b0 ;
  assign y803 = n2076 ;
  assign y804 = ~n2090 ;
  assign y805 = ~1'b0 ;
  assign y806 = ~1'b0 ;
  assign y807 = ~n933 ;
  assign y808 = n2098 ;
  assign y809 = ~1'b0 ;
  assign y810 = n2103 ;
  assign y811 = n2105 ;
  assign y812 = n2108 ;
  assign y813 = n2109 ;
  assign y814 = ~1'b0 ;
  assign y815 = ~n2111 ;
  assign y816 = ~n2113 ;
  assign y817 = n2063 ;
  assign y818 = ~1'b0 ;
  assign y819 = ~n2117 ;
  assign y820 = ~1'b0 ;
  assign y821 = ~1'b0 ;
  assign y822 = ~1'b0 ;
  assign y823 = ~n2119 ;
  assign y824 = ~n2122 ;
  assign y825 = ~n1597 ;
  assign y826 = ~n2126 ;
  assign y827 = ~1'b0 ;
  assign y828 = ~n2132 ;
  assign y829 = ~n2133 ;
  assign y830 = ~n584 ;
  assign y831 = ~n2137 ;
  assign y832 = n2138 ;
  assign y833 = n2142 ;
  assign y834 = ~1'b0 ;
  assign y835 = ~n2146 ;
  assign y836 = ~1'b0 ;
  assign y837 = 1'b0 ;
  assign y838 = ~n2147 ;
  assign y839 = n395 ;
  assign y840 = ~n2148 ;
  assign y841 = n2151 ;
  assign y842 = n2152 ;
  assign y843 = n2155 ;
  assign y844 = ~n2157 ;
  assign y845 = ~1'b0 ;
  assign y846 = ~n2160 ;
  assign y847 = n2162 ;
  assign y848 = ~n2164 ;
  assign y849 = n2166 ;
  assign y850 = ~n2170 ;
  assign y851 = n2180 ;
  assign y852 = ~1'b0 ;
  assign y853 = ~n2184 ;
  assign y854 = ~n2187 ;
  assign y855 = ~n2194 ;
  assign y856 = ~n2199 ;
  assign y857 = n612 ;
  assign y858 = n2204 ;
  assign y859 = n2205 ;
  assign y860 = n2207 ;
  assign y861 = ~n2217 ;
  assign y862 = ~n2218 ;
  assign y863 = ~1'b0 ;
  assign y864 = ~n1135 ;
  assign y865 = ~1'b0 ;
  assign y866 = ~1'b0 ;
  assign y867 = ~n2219 ;
  assign y868 = ~1'b0 ;
  assign y869 = n2220 ;
  assign y870 = n2221 ;
  assign y871 = ~1'b0 ;
  assign y872 = ~1'b0 ;
  assign y873 = n2244 ;
  assign y874 = ~1'b0 ;
  assign y875 = ~1'b0 ;
  assign y876 = 1'b0 ;
  assign y877 = n2249 ;
  assign y878 = n1506 ;
  assign y879 = ~1'b0 ;
  assign y880 = n2250 ;
  assign y881 = ~1'b0 ;
  assign y882 = n2252 ;
  assign y883 = ~n2254 ;
  assign y884 = ~1'b0 ;
  assign y885 = ~n2259 ;
  assign y886 = n2260 ;
  assign y887 = ~n2266 ;
  assign y888 = n2271 ;
  assign y889 = ~n2272 ;
  assign y890 = ~1'b0 ;
  assign y891 = n2278 ;
  assign y892 = ~1'b0 ;
  assign y893 = ~1'b0 ;
  assign y894 = n2282 ;
  assign y895 = ~n2292 ;
  assign y896 = ~1'b0 ;
  assign y897 = n2293 ;
  assign y898 = ~n2297 ;
  assign y899 = n2300 ;
  assign y900 = n2302 ;
  assign y901 = n2304 ;
  assign y902 = ~1'b0 ;
  assign y903 = ~n2306 ;
  assign y904 = n2309 ;
  assign y905 = n2312 ;
  assign y906 = n2313 ;
  assign y907 = n2315 ;
  assign y908 = ~1'b0 ;
  assign y909 = ~1'b0 ;
  assign y910 = ~n2317 ;
  assign y911 = n2325 ;
  assign y912 = n2326 ;
  assign y913 = ~n2330 ;
  assign y914 = n2334 ;
  assign y915 = n373 ;
  assign y916 = n2335 ;
  assign y917 = ~n2339 ;
  assign y918 = ~n2341 ;
  assign y919 = n2342 ;
  assign y920 = ~n2345 ;
  assign y921 = ~n2346 ;
  assign y922 = n2351 ;
  assign y923 = n2357 ;
  assign y924 = ~1'b0 ;
  assign y925 = ~1'b0 ;
  assign y926 = n2359 ;
  assign y927 = ~n2361 ;
  assign y928 = ~n2362 ;
  assign y929 = ~n1106 ;
  assign y930 = ~1'b0 ;
  assign y931 = n2364 ;
  assign y932 = ~1'b0 ;
  assign y933 = n2365 ;
  assign y934 = ~1'b0 ;
  assign y935 = n2368 ;
  assign y936 = ~n2379 ;
  assign y937 = ~1'b0 ;
  assign y938 = ~1'b0 ;
  assign y939 = n386 ;
  assign y940 = ~n2383 ;
  assign y941 = ~n2386 ;
  assign y942 = ~n2389 ;
  assign y943 = ~1'b0 ;
  assign y944 = n2393 ;
  assign y945 = ~n1971 ;
  assign y946 = ~n2395 ;
  assign y947 = ~n2397 ;
  assign y948 = n2401 ;
  assign y949 = n2404 ;
  assign y950 = n2409 ;
  assign y951 = ~n2413 ;
  assign y952 = n2421 ;
  assign y953 = ~n2423 ;
  assign y954 = ~1'b0 ;
  assign y955 = ~n2428 ;
  assign y956 = ~n1573 ;
  assign y957 = ~1'b0 ;
  assign y958 = n2432 ;
  assign y959 = n2433 ;
  assign y960 = ~n2435 ;
  assign y961 = ~n2438 ;
  assign y962 = n2443 ;
  assign y963 = ~n2445 ;
  assign y964 = ~n2453 ;
  assign y965 = n2456 ;
  assign y966 = n2457 ;
  assign y967 = ~n2459 ;
  assign y968 = ~n2466 ;
  assign y969 = ~1'b0 ;
  assign y970 = ~n2471 ;
  assign y971 = ~1'b0 ;
  assign y972 = ~n2473 ;
  assign y973 = n2474 ;
  assign y974 = ~n2484 ;
  assign y975 = ~1'b0 ;
  assign y976 = ~n2493 ;
  assign y977 = ~1'b0 ;
  assign y978 = n2496 ;
  assign y979 = ~n2498 ;
  assign y980 = ~1'b0 ;
  assign y981 = n2500 ;
  assign y982 = ~1'b0 ;
  assign y983 = ~n2501 ;
  assign y984 = n2505 ;
  assign y985 = ~n2506 ;
  assign y986 = ~n2507 ;
  assign y987 = ~n2509 ;
  assign y988 = ~n2513 ;
  assign y989 = ~n2517 ;
  assign y990 = n2519 ;
  assign y991 = ~n2521 ;
  assign y992 = n2525 ;
  assign y993 = n2528 ;
  assign y994 = ~n2529 ;
  assign y995 = ~n2531 ;
  assign y996 = ~n2532 ;
  assign y997 = ~n2537 ;
  assign y998 = ~1'b0 ;
  assign y999 = n2538 ;
  assign y1000 = ~1'b0 ;
  assign y1001 = ~n2550 ;
  assign y1002 = ~1'b0 ;
  assign y1003 = ~n2554 ;
  assign y1004 = ~n2556 ;
  assign y1005 = ~1'b0 ;
  assign y1006 = ~1'b0 ;
  assign y1007 = 1'b0 ;
  assign y1008 = ~1'b0 ;
  assign y1009 = n2566 ;
  assign y1010 = ~n2569 ;
  assign y1011 = ~1'b0 ;
  assign y1012 = ~1'b0 ;
  assign y1013 = n2570 ;
  assign y1014 = ~n2571 ;
  assign y1015 = ~n2575 ;
  assign y1016 = n2577 ;
  assign y1017 = ~1'b0 ;
  assign y1018 = ~1'b0 ;
  assign y1019 = ~n2579 ;
  assign y1020 = n2582 ;
  assign y1021 = n2585 ;
  assign y1022 = n383 ;
  assign y1023 = n2586 ;
  assign y1024 = n2590 ;
  assign y1025 = ~1'b0 ;
  assign y1026 = ~n2194 ;
  assign y1027 = 1'b0 ;
  assign y1028 = ~n2591 ;
  assign y1029 = n2594 ;
  assign y1030 = n2595 ;
  assign y1031 = n1162 ;
  assign y1032 = ~n2596 ;
  assign y1033 = ~1'b0 ;
  assign y1034 = ~1'b0 ;
  assign y1035 = ~n2597 ;
  assign y1036 = n2599 ;
  assign y1037 = n2600 ;
  assign y1038 = n2605 ;
  assign y1039 = n2606 ;
  assign y1040 = ~n2607 ;
  assign y1041 = n2609 ;
  assign y1042 = ~n2611 ;
  assign y1043 = n2617 ;
  assign y1044 = ~n1713 ;
  assign y1045 = ~n2618 ;
  assign y1046 = n2619 ;
  assign y1047 = n2620 ;
  assign y1048 = n2621 ;
  assign y1049 = ~n2629 ;
  assign y1050 = ~1'b0 ;
  assign y1051 = ~n1272 ;
  assign y1052 = ~n2642 ;
  assign y1053 = ~n1139 ;
  assign y1054 = n2649 ;
  assign y1055 = ~n2652 ;
  assign y1056 = ~n2654 ;
  assign y1057 = ~n2656 ;
  assign y1058 = ~1'b0 ;
  assign y1059 = ~1'b0 ;
  assign y1060 = ~n2662 ;
  assign y1061 = n2666 ;
  assign y1062 = n2667 ;
  assign y1063 = n1115 ;
  assign y1064 = ~n2670 ;
  assign y1065 = ~n2671 ;
  assign y1066 = ~1'b0 ;
  assign y1067 = n2676 ;
  assign y1068 = ~n2692 ;
  assign y1069 = ~n2693 ;
  assign y1070 = ~n2694 ;
  assign y1071 = n2695 ;
  assign y1072 = ~n2699 ;
  assign y1073 = ~n2701 ;
  assign y1074 = n2703 ;
  assign y1075 = ~n2708 ;
  assign y1076 = ~1'b0 ;
  assign y1077 = n2710 ;
  assign y1078 = ~n2717 ;
  assign y1079 = n2723 ;
  assign y1080 = ~n2726 ;
  assign y1081 = ~1'b0 ;
  assign y1082 = ~1'b0 ;
  assign y1083 = n2728 ;
  assign y1084 = n2737 ;
  assign y1085 = n2740 ;
  assign y1086 = ~n2741 ;
  assign y1087 = ~n2744 ;
  assign y1088 = n2746 ;
  assign y1089 = ~n2749 ;
  assign y1090 = ~n854 ;
  assign y1091 = ~n2751 ;
  assign y1092 = ~n2752 ;
  assign y1093 = n2758 ;
  assign y1094 = n2759 ;
  assign y1095 = ~1'b0 ;
  assign y1096 = n2760 ;
  assign y1097 = n2761 ;
  assign y1098 = ~1'b0 ;
  assign y1099 = ~n2767 ;
  assign y1100 = ~n2770 ;
  assign y1101 = ~1'b0 ;
  assign y1102 = n2772 ;
  assign y1103 = ~n2780 ;
  assign y1104 = ~n2785 ;
  assign y1105 = ~1'b0 ;
  assign y1106 = ~n1716 ;
  assign y1107 = n2786 ;
  assign y1108 = n2787 ;
  assign y1109 = ~n2788 ;
  assign y1110 = n1684 ;
  assign y1111 = ~n2793 ;
  assign y1112 = ~1'b0 ;
  assign y1113 = ~n2801 ;
  assign y1114 = n2804 ;
  assign y1115 = ~n2805 ;
  assign y1116 = n2806 ;
  assign y1117 = n2809 ;
  assign y1118 = n2811 ;
  assign y1119 = n2815 ;
  assign y1120 = ~1'b0 ;
  assign y1121 = ~n2821 ;
  assign y1122 = n2824 ;
  assign y1123 = n2830 ;
  assign y1124 = ~n2831 ;
  assign y1125 = ~n2837 ;
  assign y1126 = ~n2840 ;
  assign y1127 = n1578 ;
  assign y1128 = ~1'b0 ;
  assign y1129 = n2841 ;
  assign y1130 = ~1'b0 ;
  assign y1131 = ~1'b0 ;
  assign y1132 = ~n2845 ;
  assign y1133 = n2849 ;
  assign y1134 = n2852 ;
  assign y1135 = ~n2855 ;
  assign y1136 = n2858 ;
  assign y1137 = ~1'b0 ;
  assign y1138 = ~1'b0 ;
  assign y1139 = ~n2860 ;
  assign y1140 = ~n2864 ;
  assign y1141 = n2866 ;
  assign y1142 = ~n2868 ;
  assign y1143 = n2870 ;
  assign y1144 = ~n2355 ;
  assign y1145 = n2871 ;
  assign y1146 = n2875 ;
  assign y1147 = ~1'b0 ;
  assign y1148 = ~n2880 ;
  assign y1149 = ~1'b0 ;
  assign y1150 = ~n2882 ;
  assign y1151 = ~n2883 ;
  assign y1152 = n2885 ;
  assign y1153 = ~1'b0 ;
  assign y1154 = n2892 ;
  assign y1155 = ~1'b0 ;
  assign y1156 = n2894 ;
  assign y1157 = ~1'b0 ;
  assign y1158 = ~n2903 ;
  assign y1159 = n2907 ;
  assign y1160 = ~n2909 ;
  assign y1161 = ~n1639 ;
  assign y1162 = n2914 ;
  assign y1163 = ~n1784 ;
  assign y1164 = n2915 ;
  assign y1165 = ~1'b0 ;
  assign y1166 = ~n2921 ;
  assign y1167 = ~n2922 ;
  assign y1168 = ~1'b0 ;
  assign y1169 = ~n2923 ;
  assign y1170 = n2924 ;
  assign y1171 = ~n2925 ;
  assign y1172 = ~1'b0 ;
  assign y1173 = n2926 ;
  assign y1174 = n2928 ;
  assign y1175 = ~n2929 ;
  assign y1176 = ~n2930 ;
  assign y1177 = n2934 ;
  assign y1178 = ~n2935 ;
  assign y1179 = ~1'b0 ;
  assign y1180 = n2940 ;
  assign y1181 = ~n2944 ;
  assign y1182 = 1'b0 ;
  assign y1183 = ~n337 ;
  assign y1184 = ~1'b0 ;
  assign y1185 = n2947 ;
  assign y1186 = ~n2949 ;
  assign y1187 = n2951 ;
  assign y1188 = n2952 ;
  assign y1189 = ~n2954 ;
  assign y1190 = ~n2961 ;
  assign y1191 = ~n2968 ;
  assign y1192 = ~n2969 ;
  assign y1193 = ~n2976 ;
  assign y1194 = ~1'b0 ;
  assign y1195 = ~n975 ;
  assign y1196 = n2979 ;
  assign y1197 = ~n2988 ;
  assign y1198 = ~n2997 ;
  assign y1199 = ~n2999 ;
  assign y1200 = n3005 ;
  assign y1201 = ~n3009 ;
  assign y1202 = ~1'b0 ;
  assign y1203 = ~n3011 ;
  assign y1204 = ~n3014 ;
  assign y1205 = ~n3017 ;
  assign y1206 = n3019 ;
  assign y1207 = ~1'b0 ;
  assign y1208 = n3024 ;
  assign y1209 = ~n3026 ;
  assign y1210 = ~n1827 ;
  assign y1211 = ~n3027 ;
  assign y1212 = ~n3031 ;
  assign y1213 = ~n3033 ;
  assign y1214 = n3035 ;
  assign y1215 = ~1'b0 ;
  assign y1216 = ~1'b0 ;
  assign y1217 = ~1'b0 ;
  assign y1218 = n3041 ;
  assign y1219 = n3046 ;
  assign y1220 = ~n3050 ;
  assign y1221 = ~n3051 ;
  assign y1222 = ~n3055 ;
  assign y1223 = n3056 ;
  assign y1224 = ~n3057 ;
  assign y1225 = n3061 ;
  assign y1226 = n3062 ;
  assign y1227 = ~n3070 ;
  assign y1228 = n3071 ;
  assign y1229 = ~n3073 ;
  assign y1230 = ~1'b0 ;
  assign y1231 = n3077 ;
  assign y1232 = n3079 ;
  assign y1233 = n3080 ;
  assign y1234 = n3083 ;
  assign y1235 = ~n3084 ;
  assign y1236 = n3096 ;
  assign y1237 = ~n3100 ;
  assign y1238 = n3103 ;
  assign y1239 = ~1'b0 ;
  assign y1240 = ~1'b0 ;
  assign y1241 = ~n1581 ;
  assign y1242 = ~1'b0 ;
  assign y1243 = ~n3105 ;
  assign y1244 = ~n3107 ;
  assign y1245 = ~1'b0 ;
  assign y1246 = ~n3109 ;
  assign y1247 = ~1'b0 ;
  assign y1248 = ~1'b0 ;
  assign y1249 = ~1'b0 ;
  assign y1250 = n3114 ;
  assign y1251 = ~n3116 ;
  assign y1252 = ~n3117 ;
  assign y1253 = ~n3119 ;
  assign y1254 = ~n3126 ;
  assign y1255 = ~1'b0 ;
  assign y1256 = n2489 ;
  assign y1257 = ~1'b0 ;
  assign y1258 = n3130 ;
  assign y1259 = ~n3132 ;
  assign y1260 = n3135 ;
  assign y1261 = n3140 ;
  assign y1262 = ~n3143 ;
  assign y1263 = ~1'b0 ;
  assign y1264 = ~1'b0 ;
  assign y1265 = ~1'b0 ;
  assign y1266 = ~n3147 ;
  assign y1267 = ~1'b0 ;
  assign y1268 = ~n3152 ;
  assign y1269 = ~n3157 ;
  assign y1270 = n2980 ;
  assign y1271 = n3161 ;
  assign y1272 = ~n3163 ;
  assign y1273 = ~n3165 ;
  assign y1274 = ~n3166 ;
  assign y1275 = ~n3169 ;
  assign y1276 = ~n3171 ;
  assign y1277 = ~n3172 ;
  assign y1278 = n3173 ;
  assign y1279 = ~n3175 ;
  assign y1280 = ~1'b0 ;
  assign y1281 = ~n3176 ;
  assign y1282 = n3179 ;
  assign y1283 = n3181 ;
  assign y1284 = ~n3188 ;
  assign y1285 = ~n3191 ;
  assign y1286 = ~n3198 ;
  assign y1287 = ~n3202 ;
  assign y1288 = ~n3204 ;
  assign y1289 = n1627 ;
  assign y1290 = ~n3206 ;
  assign y1291 = n3210 ;
  assign y1292 = ~n3211 ;
  assign y1293 = n3213 ;
  assign y1294 = n3216 ;
  assign y1295 = ~n3217 ;
  assign y1296 = n3221 ;
  assign y1297 = ~1'b0 ;
  assign y1298 = ~n3228 ;
  assign y1299 = ~1'b0 ;
  assign y1300 = ~n3232 ;
  assign y1301 = ~n3239 ;
  assign y1302 = n3243 ;
  assign y1303 = ~1'b0 ;
  assign y1304 = n3245 ;
  assign y1305 = ~1'b0 ;
  assign y1306 = ~1'b0 ;
  assign y1307 = ~n3252 ;
  assign y1308 = ~1'b0 ;
  assign y1309 = ~1'b0 ;
  assign y1310 = n3253 ;
  assign y1311 = ~n3255 ;
  assign y1312 = ~n3258 ;
  assign y1313 = ~1'b0 ;
  assign y1314 = ~n3265 ;
  assign y1315 = ~n3266 ;
  assign y1316 = n3267 ;
  assign y1317 = ~n3268 ;
  assign y1318 = n3270 ;
  assign y1319 = n3274 ;
  assign y1320 = n3275 ;
  assign y1321 = n3279 ;
  assign y1322 = ~n403 ;
  assign y1323 = ~1'b0 ;
  assign y1324 = n3286 ;
  assign y1325 = n3287 ;
  assign y1326 = n3288 ;
  assign y1327 = ~n3289 ;
  assign y1328 = ~n3294 ;
  assign y1329 = n3298 ;
  assign y1330 = n3302 ;
  assign y1331 = ~n3304 ;
  assign y1332 = ~n3307 ;
  assign y1333 = ~n3310 ;
  assign y1334 = ~1'b0 ;
  assign y1335 = n3312 ;
  assign y1336 = ~n3317 ;
  assign y1337 = ~n3319 ;
  assign y1338 = ~n3320 ;
  assign y1339 = ~1'b0 ;
  assign y1340 = x84 ;
  assign y1341 = ~n3325 ;
  assign y1342 = ~1'b0 ;
  assign y1343 = ~n3329 ;
  assign y1344 = n3330 ;
  assign y1345 = ~1'b0 ;
  assign y1346 = ~1'b0 ;
  assign y1347 = n3334 ;
  assign y1348 = n3335 ;
  assign y1349 = n3336 ;
  assign y1350 = ~n3344 ;
  assign y1351 = ~n3347 ;
  assign y1352 = ~1'b0 ;
  assign y1353 = ~n3348 ;
  assign y1354 = n3353 ;
  assign y1355 = n3355 ;
  assign y1356 = n3358 ;
  assign y1357 = ~n3366 ;
  assign y1358 = ~n372 ;
  assign y1359 = n3367 ;
  assign y1360 = n3372 ;
  assign y1361 = n3377 ;
  assign y1362 = n3380 ;
  assign y1363 = ~1'b0 ;
  assign y1364 = ~n3382 ;
  assign y1365 = n3383 ;
  assign y1366 = ~1'b0 ;
  assign y1367 = ~n3384 ;
  assign y1368 = ~1'b0 ;
  assign y1369 = ~1'b0 ;
  assign y1370 = n3385 ;
  assign y1371 = ~n3391 ;
  assign y1372 = ~n3393 ;
  assign y1373 = n3395 ;
  assign y1374 = ~n3401 ;
  assign y1375 = ~n3402 ;
  assign y1376 = ~1'b0 ;
  assign y1377 = ~n3404 ;
  assign y1378 = n3408 ;
  assign y1379 = ~n3409 ;
  assign y1380 = n3417 ;
  assign y1381 = n3418 ;
  assign y1382 = ~1'b0 ;
  assign y1383 = n3424 ;
  assign y1384 = ~n3431 ;
  assign y1385 = ~n3432 ;
  assign y1386 = ~n3435 ;
  assign y1387 = n2485 ;
  assign y1388 = n3436 ;
  assign y1389 = n3437 ;
  assign y1390 = ~n3438 ;
  assign y1391 = ~n3439 ;
  assign y1392 = ~1'b0 ;
  assign y1393 = ~n3442 ;
  assign y1394 = ~n3444 ;
  assign y1395 = ~n3446 ;
  assign y1396 = ~n2622 ;
  assign y1397 = ~1'b0 ;
  assign y1398 = n3450 ;
  assign y1399 = ~n3461 ;
  assign y1400 = n3464 ;
  assign y1401 = ~n3466 ;
  assign y1402 = ~n3467 ;
  assign y1403 = n2032 ;
  assign y1404 = n3475 ;
  assign y1405 = ~n3478 ;
  assign y1406 = n3480 ;
  assign y1407 = n3484 ;
  assign y1408 = ~1'b0 ;
  assign y1409 = ~1'b0 ;
  assign y1410 = ~1'b0 ;
  assign y1411 = n3307 ;
  assign y1412 = ~1'b0 ;
  assign y1413 = ~1'b0 ;
  assign y1414 = ~n3491 ;
  assign y1415 = n3496 ;
  assign y1416 = ~n3512 ;
  assign y1417 = 1'b0 ;
  assign y1418 = ~n3515 ;
  assign y1419 = ~n3519 ;
  assign y1420 = n3521 ;
  assign y1421 = ~n3523 ;
  assign y1422 = ~n3524 ;
  assign y1423 = ~1'b0 ;
  assign y1424 = n3526 ;
  assign y1425 = ~1'b0 ;
  assign y1426 = ~n3531 ;
  assign y1427 = ~n3532 ;
  assign y1428 = n3536 ;
  assign y1429 = ~n3544 ;
  assign y1430 = n530 ;
  assign y1431 = ~n3546 ;
  assign y1432 = ~n3553 ;
  assign y1433 = ~n3559 ;
  assign y1434 = n3564 ;
  assign y1435 = ~1'b0 ;
  assign y1436 = ~1'b0 ;
  assign y1437 = ~1'b0 ;
  assign y1438 = n3565 ;
  assign y1439 = n3567 ;
  assign y1440 = 1'b0 ;
  assign y1441 = ~n3571 ;
  assign y1442 = n1479 ;
  assign y1443 = ~1'b0 ;
  assign y1444 = ~n3575 ;
  assign y1445 = ~n3581 ;
  assign y1446 = ~n3584 ;
  assign y1447 = n3585 ;
  assign y1448 = ~n691 ;
  assign y1449 = n3594 ;
  assign y1450 = n3596 ;
  assign y1451 = n2430 ;
  assign y1452 = n3600 ;
  assign y1453 = ~n3604 ;
  assign y1454 = ~1'b0 ;
  assign y1455 = ~n3618 ;
  assign y1456 = ~1'b0 ;
  assign y1457 = ~1'b0 ;
  assign y1458 = n3619 ;
  assign y1459 = ~n3622 ;
  assign y1460 = ~n3624 ;
  assign y1461 = ~n3625 ;
  assign y1462 = ~n3628 ;
  assign y1463 = ~n3630 ;
  assign y1464 = n3635 ;
  assign y1465 = n1637 ;
  assign y1466 = ~n3636 ;
  assign y1467 = ~1'b0 ;
  assign y1468 = n3637 ;
  assign y1469 = ~n3638 ;
  assign y1470 = n3639 ;
  assign y1471 = ~n3641 ;
  assign y1472 = ~n3646 ;
  assign y1473 = n3651 ;
  assign y1474 = ~n3652 ;
  assign y1475 = ~1'b0 ;
  assign y1476 = ~n3653 ;
  assign y1477 = ~n3655 ;
  assign y1478 = ~n3656 ;
  assign y1479 = ~n3663 ;
  assign y1480 = ~n3669 ;
  assign y1481 = n3670 ;
  assign y1482 = ~n3672 ;
  assign y1483 = ~1'b0 ;
  assign y1484 = ~1'b0 ;
  assign y1485 = ~n3674 ;
  assign y1486 = n3675 ;
  assign y1487 = n3676 ;
  assign y1488 = n3681 ;
  assign y1489 = ~n3686 ;
  assign y1490 = ~n3687 ;
  assign y1491 = ~n3693 ;
  assign y1492 = ~1'b0 ;
  assign y1493 = ~n3697 ;
  assign y1494 = ~1'b0 ;
  assign y1495 = ~n3699 ;
  assign y1496 = n3702 ;
  assign y1497 = n3708 ;
  assign y1498 = ~n3709 ;
  assign y1499 = n3717 ;
  assign y1500 = ~n3719 ;
  assign y1501 = ~n3723 ;
  assign y1502 = ~1'b0 ;
  assign y1503 = ~n3724 ;
  assign y1504 = n3727 ;
  assign y1505 = n910 ;
  assign y1506 = n3728 ;
  assign y1507 = n3731 ;
  assign y1508 = ~1'b0 ;
  assign y1509 = ~n3739 ;
  assign y1510 = ~n3740 ;
  assign y1511 = ~n3741 ;
  assign y1512 = n3744 ;
  assign y1513 = ~n3749 ;
  assign y1514 = n3753 ;
  assign y1515 = n3754 ;
  assign y1516 = ~1'b0 ;
  assign y1517 = ~1'b0 ;
  assign y1518 = ~1'b0 ;
  assign y1519 = ~n2549 ;
  assign y1520 = ~n3758 ;
  assign y1521 = n3760 ;
  assign y1522 = ~1'b0 ;
  assign y1523 = n3761 ;
  assign y1524 = ~1'b0 ;
  assign y1525 = n3768 ;
  assign y1526 = ~n3776 ;
  assign y1527 = ~1'b0 ;
  assign y1528 = ~n3781 ;
  assign y1529 = ~1'b0 ;
  assign y1530 = ~n3786 ;
  assign y1531 = ~1'b0 ;
  assign y1532 = n3789 ;
  assign y1533 = ~n2608 ;
  assign y1534 = ~1'b0 ;
  assign y1535 = n3791 ;
  assign y1536 = n3793 ;
  assign y1537 = ~n3800 ;
  assign y1538 = ~1'b0 ;
  assign y1539 = n3802 ;
  assign y1540 = n3807 ;
  assign y1541 = n3808 ;
  assign y1542 = n3811 ;
  assign y1543 = ~1'b0 ;
  assign y1544 = n3812 ;
  assign y1545 = ~n3815 ;
  assign y1546 = ~1'b0 ;
  assign y1547 = ~n3818 ;
  assign y1548 = ~n3820 ;
  assign y1549 = ~1'b0 ;
  assign y1550 = n3821 ;
  assign y1551 = n3826 ;
  assign y1552 = ~n3828 ;
  assign y1553 = n3831 ;
  assign y1554 = ~n3832 ;
  assign y1555 = ~1'b0 ;
  assign y1556 = n1101 ;
  assign y1557 = n3835 ;
  assign y1558 = ~n3836 ;
  assign y1559 = ~n3842 ;
  assign y1560 = ~n3844 ;
  assign y1561 = ~1'b0 ;
  assign y1562 = ~n3856 ;
  assign y1563 = n3858 ;
  assign y1564 = n3860 ;
  assign y1565 = ~1'b0 ;
  assign y1566 = ~1'b0 ;
  assign y1567 = ~1'b0 ;
  assign y1568 = n3866 ;
  assign y1569 = ~n3868 ;
  assign y1570 = ~1'b0 ;
  assign y1571 = ~n3872 ;
  assign y1572 = ~1'b0 ;
  assign y1573 = ~1'b0 ;
  assign y1574 = n3881 ;
  assign y1575 = ~1'b0 ;
  assign y1576 = ~1'b0 ;
  assign y1577 = 1'b0 ;
  assign y1578 = ~n3882 ;
  assign y1579 = ~n3906 ;
  assign y1580 = ~1'b0 ;
  assign y1581 = n2953 ;
  assign y1582 = n3910 ;
  assign y1583 = ~n3911 ;
  assign y1584 = ~n3916 ;
  assign y1585 = n3922 ;
  assign y1586 = n341 ;
  assign y1587 = n3924 ;
  assign y1588 = n3927 ;
  assign y1589 = n3931 ;
  assign y1590 = ~1'b0 ;
  assign y1591 = ~1'b0 ;
  assign y1592 = ~n3934 ;
  assign y1593 = ~n3937 ;
  assign y1594 = n3940 ;
  assign y1595 = n3946 ;
  assign y1596 = n3948 ;
  assign y1597 = ~n3952 ;
  assign y1598 = ~n3956 ;
  assign y1599 = n3957 ;
  assign y1600 = ~n3958 ;
  assign y1601 = n3960 ;
  assign y1602 = n3961 ;
  assign y1603 = ~1'b0 ;
  assign y1604 = ~n3962 ;
  assign y1605 = ~n3974 ;
  assign y1606 = n3151 ;
  assign y1607 = n3975 ;
  assign y1608 = n3977 ;
  assign y1609 = n3979 ;
  assign y1610 = ~n3980 ;
  assign y1611 = ~n3981 ;
  assign y1612 = ~1'b0 ;
  assign y1613 = ~n3982 ;
  assign y1614 = n3984 ;
  assign y1615 = ~1'b0 ;
  assign y1616 = ~n3986 ;
  assign y1617 = n3989 ;
  assign y1618 = ~n3991 ;
  assign y1619 = ~n3993 ;
  assign y1620 = n3994 ;
  assign y1621 = ~1'b0 ;
  assign y1622 = ~1'b0 ;
  assign y1623 = ~1'b0 ;
  assign y1624 = ~n1860 ;
  assign y1625 = ~1'b0 ;
  assign y1626 = ~n3997 ;
  assign y1627 = ~1'b0 ;
  assign y1628 = ~n3998 ;
  assign y1629 = n4000 ;
  assign y1630 = ~n4002 ;
  assign y1631 = ~1'b0 ;
  assign y1632 = ~n4008 ;
  assign y1633 = n4010 ;
  assign y1634 = n4011 ;
  assign y1635 = ~1'b0 ;
  assign y1636 = ~n4012 ;
  assign y1637 = ~n4016 ;
  assign y1638 = ~n4018 ;
  assign y1639 = n4023 ;
  assign y1640 = n4024 ;
  assign y1641 = n431 ;
  assign y1642 = n4028 ;
  assign y1643 = n4030 ;
  assign y1644 = n4032 ;
  assign y1645 = ~n4037 ;
  assign y1646 = ~1'b0 ;
  assign y1647 = n4038 ;
  assign y1648 = n2694 ;
  assign y1649 = ~1'b0 ;
  assign y1650 = n4041 ;
  assign y1651 = n4043 ;
  assign y1652 = ~n4050 ;
  assign y1653 = ~n4053 ;
  assign y1654 = ~1'b0 ;
  assign y1655 = ~n306 ;
  assign y1656 = ~n4055 ;
  assign y1657 = n4057 ;
  assign y1658 = n4058 ;
  assign y1659 = ~1'b0 ;
  assign y1660 = n4075 ;
  assign y1661 = n4076 ;
  assign y1662 = n4081 ;
  assign y1663 = n4082 ;
  assign y1664 = n4090 ;
  assign y1665 = n4092 ;
  assign y1666 = ~n4096 ;
  assign y1667 = n4097 ;
  assign y1668 = n4099 ;
  assign y1669 = n4104 ;
  assign y1670 = ~1'b0 ;
  assign y1671 = ~n4105 ;
  assign y1672 = ~n4106 ;
  assign y1673 = ~1'b0 ;
  assign y1674 = ~n4113 ;
  assign y1675 = n4118 ;
  assign y1676 = ~n4120 ;
  assign y1677 = ~n4122 ;
  assign y1678 = ~1'b0 ;
  assign y1679 = ~n4123 ;
  assign y1680 = n283 ;
  assign y1681 = ~n4129 ;
  assign y1682 = ~n4130 ;
  assign y1683 = ~1'b0 ;
  assign y1684 = ~1'b0 ;
  assign y1685 = ~n1492 ;
  assign y1686 = ~n4131 ;
  assign y1687 = ~1'b0 ;
  assign y1688 = ~n4133 ;
  assign y1689 = ~n4135 ;
  assign y1690 = n4136 ;
  assign y1691 = ~n4140 ;
  assign y1692 = ~n4143 ;
  assign y1693 = n4144 ;
  assign y1694 = n4147 ;
  assign y1695 = ~n4149 ;
  assign y1696 = ~n4151 ;
  assign y1697 = ~n764 ;
  assign y1698 = ~n4153 ;
  assign y1699 = ~n4154 ;
  assign y1700 = ~1'b0 ;
  assign y1701 = n4156 ;
  assign y1702 = ~1'b0 ;
  assign y1703 = ~n4161 ;
  assign y1704 = n4171 ;
  assign y1705 = ~n4174 ;
  assign y1706 = ~n4178 ;
  assign y1707 = ~n3681 ;
  assign y1708 = ~n4183 ;
  assign y1709 = n4184 ;
  assign y1710 = n4188 ;
  assign y1711 = ~n4192 ;
  assign y1712 = 1'b0 ;
  assign y1713 = ~n4195 ;
  assign y1714 = ~1'b0 ;
  assign y1715 = n4197 ;
  assign y1716 = ~n4208 ;
  assign y1717 = n4213 ;
  assign y1718 = n4214 ;
  assign y1719 = ~n4216 ;
  assign y1720 = ~n4220 ;
  assign y1721 = ~n4222 ;
  assign y1722 = ~1'b0 ;
  assign y1723 = n4223 ;
  assign y1724 = n4227 ;
  assign y1725 = ~n4229 ;
  assign y1726 = n4231 ;
  assign y1727 = n4232 ;
  assign y1728 = x58 ;
  assign y1729 = ~n4233 ;
  assign y1730 = ~n4238 ;
  assign y1731 = ~n4241 ;
  assign y1732 = ~1'b0 ;
  assign y1733 = n4249 ;
  assign y1734 = ~n4250 ;
  assign y1735 = ~1'b0 ;
  assign y1736 = n3192 ;
  assign y1737 = ~n4253 ;
  assign y1738 = ~n2190 ;
  assign y1739 = ~n4254 ;
  assign y1740 = ~n4262 ;
  assign y1741 = n4264 ;
  assign y1742 = n4275 ;
  assign y1743 = n4277 ;
  assign y1744 = ~1'b0 ;
  assign y1745 = ~1'b0 ;
  assign y1746 = n4280 ;
  assign y1747 = ~1'b0 ;
  assign y1748 = ~1'b0 ;
  assign y1749 = ~n4281 ;
  assign y1750 = n4286 ;
  assign y1751 = n4289 ;
  assign y1752 = n4292 ;
  assign y1753 = ~1'b0 ;
  assign y1754 = n4295 ;
  assign y1755 = ~1'b0 ;
  assign y1756 = ~1'b0 ;
  assign y1757 = ~n4301 ;
  assign y1758 = ~1'b0 ;
  assign y1759 = n4305 ;
  assign y1760 = ~1'b0 ;
  assign y1761 = n4306 ;
  assign y1762 = ~n4307 ;
  assign y1763 = ~n4308 ;
  assign y1764 = ~1'b0 ;
  assign y1765 = ~n4311 ;
  assign y1766 = n4312 ;
  assign y1767 = ~1'b0 ;
  assign y1768 = ~1'b0 ;
  assign y1769 = ~n4314 ;
  assign y1770 = ~n4319 ;
  assign y1771 = ~1'b0 ;
  assign y1772 = ~1'b0 ;
  assign y1773 = n4323 ;
  assign y1774 = ~n4327 ;
  assign y1775 = ~1'b0 ;
  assign y1776 = ~n4333 ;
  assign y1777 = ~n4336 ;
  assign y1778 = ~1'b0 ;
  assign y1779 = n4343 ;
  assign y1780 = ~1'b0 ;
  assign y1781 = ~n4344 ;
  assign y1782 = ~n4348 ;
  assign y1783 = ~n4355 ;
  assign y1784 = ~1'b0 ;
  assign y1785 = ~1'b0 ;
  assign y1786 = n4357 ;
  assign y1787 = ~1'b0 ;
  assign y1788 = n4358 ;
  assign y1789 = ~n4359 ;
  assign y1790 = n4363 ;
  assign y1791 = ~n4364 ;
  assign y1792 = ~n4366 ;
  assign y1793 = ~n4371 ;
  assign y1794 = ~n4374 ;
  assign y1795 = ~1'b0 ;
  assign y1796 = ~n4378 ;
  assign y1797 = ~n642 ;
  assign y1798 = ~1'b0 ;
  assign y1799 = ~n4379 ;
  assign y1800 = n4390 ;
  assign y1801 = ~1'b0 ;
  assign y1802 = n4392 ;
  assign y1803 = ~n4393 ;
  assign y1804 = 1'b0 ;
  assign y1805 = ~1'b0 ;
  assign y1806 = ~n4397 ;
  assign y1807 = ~n4398 ;
  assign y1808 = ~n4407 ;
  assign y1809 = 1'b0 ;
  assign y1810 = ~n4410 ;
  assign y1811 = ~n4424 ;
  assign y1812 = ~n4426 ;
  assign y1813 = 1'b0 ;
  assign y1814 = ~1'b0 ;
  assign y1815 = n4436 ;
  assign y1816 = ~n4441 ;
  assign y1817 = n4446 ;
  assign y1818 = ~n4447 ;
  assign y1819 = ~1'b0 ;
  assign y1820 = n4448 ;
  assign y1821 = n4450 ;
  assign y1822 = n4452 ;
  assign y1823 = ~n4453 ;
  assign y1824 = n4454 ;
  assign y1825 = ~1'b0 ;
  assign y1826 = n4456 ;
  assign y1827 = ~n4457 ;
  assign y1828 = n4459 ;
  assign y1829 = n4460 ;
  assign y1830 = ~1'b0 ;
  assign y1831 = n4464 ;
  assign y1832 = n4465 ;
  assign y1833 = 1'b0 ;
  assign y1834 = n4470 ;
  assign y1835 = ~1'b0 ;
  assign y1836 = n4471 ;
  assign y1837 = ~n4474 ;
  assign y1838 = ~n4475 ;
  assign y1839 = n306 ;
  assign y1840 = n4477 ;
  assign y1841 = n4478 ;
  assign y1842 = n4479 ;
  assign y1843 = ~n1861 ;
  assign y1844 = ~n4481 ;
  assign y1845 = ~n4485 ;
  assign y1846 = n4490 ;
  assign y1847 = n4500 ;
  assign y1848 = ~n4503 ;
  assign y1849 = ~n4508 ;
  assign y1850 = ~1'b0 ;
  assign y1851 = ~n4512 ;
  assign y1852 = ~1'b0 ;
  assign y1853 = ~n4514 ;
  assign y1854 = n4515 ;
  assign y1855 = n4516 ;
  assign y1856 = n1529 ;
  assign y1857 = ~n4520 ;
  assign y1858 = ~n4524 ;
  assign y1859 = ~n4526 ;
  assign y1860 = n4529 ;
  assign y1861 = ~1'b0 ;
  assign y1862 = n4535 ;
  assign y1863 = n4538 ;
  assign y1864 = ~n4539 ;
  assign y1865 = ~n1044 ;
  assign y1866 = ~1'b0 ;
  assign y1867 = ~n4543 ;
  assign y1868 = ~n4548 ;
  assign y1869 = n4553 ;
  assign y1870 = ~1'b0 ;
  assign y1871 = n4555 ;
  assign y1872 = n4562 ;
  assign y1873 = n4564 ;
  assign y1874 = ~n4566 ;
  assign y1875 = ~n4570 ;
  assign y1876 = ~n4573 ;
  assign y1877 = n4575 ;
  assign y1878 = ~1'b0 ;
  assign y1879 = n4578 ;
  assign y1880 = ~1'b0 ;
  assign y1881 = ~1'b0 ;
  assign y1882 = ~1'b0 ;
  assign y1883 = ~n4579 ;
  assign y1884 = ~n4580 ;
  assign y1885 = ~1'b0 ;
  assign y1886 = ~n4585 ;
  assign y1887 = n4591 ;
  assign y1888 = ~n4594 ;
  assign y1889 = ~n4600 ;
  assign y1890 = ~n4602 ;
  assign y1891 = ~n4605 ;
  assign y1892 = n4610 ;
  assign y1893 = ~n4612 ;
  assign y1894 = n4613 ;
  assign y1895 = ~n4616 ;
  assign y1896 = n4622 ;
  assign y1897 = ~1'b0 ;
  assign y1898 = n4625 ;
  assign y1899 = ~1'b0 ;
  assign y1900 = n4626 ;
  assign y1901 = ~n4631 ;
  assign y1902 = ~n4632 ;
  assign y1903 = ~1'b0 ;
  assign y1904 = ~n4634 ;
  assign y1905 = ~1'b0 ;
  assign y1906 = n4636 ;
  assign y1907 = ~n4637 ;
  assign y1908 = n4640 ;
  assign y1909 = n4642 ;
  assign y1910 = ~n4645 ;
  assign y1911 = ~1'b0 ;
  assign y1912 = ~n4648 ;
  assign y1913 = n4654 ;
  assign y1914 = ~1'b0 ;
  assign y1915 = ~n4655 ;
  assign y1916 = ~n4658 ;
  assign y1917 = n4660 ;
  assign y1918 = n4665 ;
  assign y1919 = ~n4672 ;
  assign y1920 = n4674 ;
  assign y1921 = ~n4678 ;
  assign y1922 = 1'b0 ;
  assign y1923 = ~n4679 ;
  assign y1924 = ~n4681 ;
  assign y1925 = n4683 ;
  assign y1926 = x110 ;
  assign y1927 = ~x65 ;
  assign y1928 = ~n4684 ;
  assign y1929 = ~n3550 ;
  assign y1930 = ~1'b0 ;
  assign y1931 = n4685 ;
  assign y1932 = ~1'b0 ;
  assign y1933 = n4693 ;
  assign y1934 = n4695 ;
  assign y1935 = n4697 ;
  assign y1936 = n4698 ;
  assign y1937 = ~1'b0 ;
  assign y1938 = n4700 ;
  assign y1939 = n4380 ;
  assign y1940 = ~n4701 ;
  assign y1941 = ~n4702 ;
  assign y1942 = n4703 ;
  assign y1943 = n4705 ;
  assign y1944 = n4708 ;
  assign y1945 = n4713 ;
  assign y1946 = n4714 ;
  assign y1947 = ~n4715 ;
  assign y1948 = ~n4717 ;
  assign y1949 = ~n4718 ;
  assign y1950 = ~n4722 ;
  assign y1951 = n4729 ;
  assign y1952 = ~n4739 ;
  assign y1953 = n4742 ;
  assign y1954 = ~n4743 ;
  assign y1955 = ~n4745 ;
  assign y1956 = ~1'b0 ;
  assign y1957 = ~n4746 ;
  assign y1958 = n4748 ;
  assign y1959 = n4750 ;
  assign y1960 = ~n4754 ;
  assign y1961 = n4757 ;
  assign y1962 = n4758 ;
  assign y1963 = ~1'b0 ;
  assign y1964 = ~n4759 ;
  assign y1965 = n4760 ;
  assign y1966 = n4761 ;
  assign y1967 = n4764 ;
  assign y1968 = ~1'b0 ;
  assign y1969 = n4768 ;
  assign y1970 = n4772 ;
  assign y1971 = n4775 ;
  assign y1972 = ~1'b0 ;
  assign y1973 = n4776 ;
  assign y1974 = n4779 ;
  assign y1975 = n4780 ;
  assign y1976 = ~n4782 ;
  assign y1977 = n4783 ;
  assign y1978 = ~n4785 ;
  assign y1979 = ~n4787 ;
  assign y1980 = ~n4788 ;
  assign y1981 = ~n4793 ;
  assign y1982 = n4797 ;
  assign y1983 = n4802 ;
  assign y1984 = ~n4805 ;
  assign y1985 = ~n4808 ;
  assign y1986 = ~1'b0 ;
  assign y1987 = n4811 ;
  assign y1988 = ~n4812 ;
  assign y1989 = ~n4821 ;
  assign y1990 = ~1'b0 ;
  assign y1991 = n4829 ;
  assign y1992 = ~1'b0 ;
  assign y1993 = ~n4837 ;
  assign y1994 = ~n4842 ;
  assign y1995 = ~n4845 ;
  assign y1996 = n4846 ;
  assign y1997 = ~n4847 ;
  assign y1998 = n2104 ;
  assign y1999 = ~n4848 ;
  assign y2000 = ~1'b0 ;
  assign y2001 = ~n4857 ;
  assign y2002 = ~1'b0 ;
  assign y2003 = n4859 ;
  assign y2004 = ~1'b0 ;
  assign y2005 = ~n4860 ;
  assign y2006 = ~n4864 ;
  assign y2007 = ~n4867 ;
  assign y2008 = ~n4868 ;
  assign y2009 = ~n4874 ;
  assign y2010 = ~n4883 ;
  assign y2011 = ~n4884 ;
  assign y2012 = ~1'b0 ;
  assign y2013 = ~n4886 ;
  assign y2014 = ~1'b0 ;
  assign y2015 = ~n4887 ;
  assign y2016 = ~1'b0 ;
  assign y2017 = ~1'b0 ;
  assign y2018 = n4891 ;
  assign y2019 = n4893 ;
  assign y2020 = n4896 ;
  assign y2021 = ~n4897 ;
  assign y2022 = n4898 ;
  assign y2023 = ~n1815 ;
  assign y2024 = ~n4900 ;
  assign y2025 = ~1'b0 ;
  assign y2026 = ~n4907 ;
  assign y2027 = n4909 ;
  assign y2028 = n4915 ;
  assign y2029 = ~1'b0 ;
  assign y2030 = ~n4917 ;
  assign y2031 = n4929 ;
  assign y2032 = ~1'b0 ;
  assign y2033 = n4930 ;
  assign y2034 = n4931 ;
  assign y2035 = n4933 ;
  assign y2036 = ~1'b0 ;
  assign y2037 = n4938 ;
  assign y2038 = n4945 ;
  assign y2039 = ~1'b0 ;
  assign y2040 = ~n4952 ;
  assign y2041 = ~n4954 ;
  assign y2042 = n4955 ;
  assign y2043 = ~1'b0 ;
  assign y2044 = ~n4957 ;
  assign y2045 = ~n4961 ;
  assign y2046 = 1'b0 ;
  assign y2047 = ~1'b0 ;
  assign y2048 = ~1'b0 ;
  assign y2049 = n4963 ;
  assign y2050 = ~1'b0 ;
  assign y2051 = ~n4964 ;
  assign y2052 = n804 ;
  assign y2053 = ~n4966 ;
  assign y2054 = n4974 ;
  assign y2055 = ~n4977 ;
  assign y2056 = n4984 ;
  assign y2057 = 1'b0 ;
  assign y2058 = ~n4987 ;
  assign y2059 = ~n1108 ;
  assign y2060 = ~n4991 ;
  assign y2061 = ~n4995 ;
  assign y2062 = ~n4996 ;
  assign y2063 = ~n5001 ;
  assign y2064 = n5002 ;
  assign y2065 = ~n5003 ;
  assign y2066 = n5008 ;
  assign y2067 = ~1'b0 ;
  assign y2068 = n4749 ;
  assign y2069 = ~n5013 ;
  assign y2070 = n1599 ;
  assign y2071 = ~n5014 ;
  assign y2072 = ~1'b0 ;
  assign y2073 = n5016 ;
  assign y2074 = ~n5017 ;
  assign y2075 = n5020 ;
  assign y2076 = n5021 ;
  assign y2077 = ~n5025 ;
  assign y2078 = ~n5029 ;
  assign y2079 = ~1'b0 ;
  assign y2080 = ~n5032 ;
  assign y2081 = ~1'b0 ;
  assign y2082 = ~1'b0 ;
  assign y2083 = ~n5036 ;
  assign y2084 = ~n5039 ;
  assign y2085 = ~1'b0 ;
  assign y2086 = ~n5045 ;
  assign y2087 = n5046 ;
  assign y2088 = n5048 ;
  assign y2089 = ~1'b0 ;
  assign y2090 = ~1'b0 ;
  assign y2091 = n5051 ;
  assign y2092 = n5053 ;
  assign y2093 = ~n5058 ;
  assign y2094 = n5061 ;
  assign y2095 = ~n5069 ;
  assign y2096 = ~n5072 ;
  assign y2097 = ~n5079 ;
  assign y2098 = n5083 ;
  assign y2099 = n5085 ;
  assign y2100 = n3995 ;
  assign y2101 = n5090 ;
  assign y2102 = n5094 ;
  assign y2103 = n5097 ;
  assign y2104 = ~n5098 ;
  assign y2105 = ~1'b0 ;
  assign y2106 = ~n5099 ;
  assign y2107 = ~n5102 ;
  assign y2108 = ~n5105 ;
  assign y2109 = n5106 ;
  assign y2110 = ~n5107 ;
  assign y2111 = ~n5112 ;
  assign y2112 = n5114 ;
  assign y2113 = ~1'b0 ;
  assign y2114 = ~n5118 ;
  assign y2115 = n5119 ;
  assign y2116 = n5121 ;
  assign y2117 = n5122 ;
  assign y2118 = n5127 ;
  assign y2119 = n5130 ;
  assign y2120 = ~1'b0 ;
  assign y2121 = n5133 ;
  assign y2122 = n5138 ;
  assign y2123 = n5142 ;
  assign y2124 = ~n5149 ;
  assign y2125 = ~n5150 ;
  assign y2126 = n2654 ;
  assign y2127 = n5152 ;
  assign y2128 = n5156 ;
  assign y2129 = ~1'b0 ;
  assign y2130 = n5160 ;
  assign y2131 = ~1'b0 ;
  assign y2132 = n5161 ;
  assign y2133 = ~n5168 ;
  assign y2134 = ~1'b0 ;
  assign y2135 = ~1'b0 ;
  assign y2136 = ~n5169 ;
  assign y2137 = n5173 ;
  assign y2138 = n5176 ;
  assign y2139 = 1'b0 ;
  assign y2140 = n5181 ;
  assign y2141 = n5185 ;
  assign y2142 = n5191 ;
  assign y2143 = n5194 ;
  assign y2144 = ~n5196 ;
  assign y2145 = ~n5199 ;
  assign y2146 = ~n5203 ;
  assign y2147 = n5204 ;
  assign y2148 = ~n5206 ;
  assign y2149 = ~n5212 ;
  assign y2150 = ~1'b0 ;
  assign y2151 = ~1'b0 ;
  assign y2152 = ~1'b0 ;
  assign y2153 = n5216 ;
  assign y2154 = n5218 ;
  assign y2155 = ~n5219 ;
  assign y2156 = ~n5221 ;
  assign y2157 = ~n5222 ;
  assign y2158 = n5223 ;
  assign y2159 = n5224 ;
  assign y2160 = ~n5225 ;
  assign y2161 = ~n5227 ;
  assign y2162 = ~1'b0 ;
  assign y2163 = ~n5229 ;
  assign y2164 = n5231 ;
  assign y2165 = ~1'b0 ;
  assign y2166 = ~1'b0 ;
  assign y2167 = n5235 ;
  assign y2168 = n4909 ;
  assign y2169 = n5236 ;
  assign y2170 = n5237 ;
  assign y2171 = ~n5240 ;
  assign y2172 = ~n5242 ;
  assign y2173 = ~n5243 ;
  assign y2174 = ~n5246 ;
  assign y2175 = n4827 ;
  assign y2176 = ~1'b0 ;
  assign y2177 = ~n5247 ;
  assign y2178 = n5251 ;
  assign y2179 = n5253 ;
  assign y2180 = ~n5255 ;
  assign y2181 = 1'b0 ;
  assign y2182 = ~1'b0 ;
  assign y2183 = 1'b0 ;
  assign y2184 = n5258 ;
  assign y2185 = ~n5262 ;
  assign y2186 = ~n5264 ;
  assign y2187 = n5265 ;
  assign y2188 = ~n5266 ;
  assign y2189 = ~n5269 ;
  assign y2190 = ~n5273 ;
  assign y2191 = ~1'b0 ;
  assign y2192 = ~n5275 ;
  assign y2193 = ~n5278 ;
  assign y2194 = ~1'b0 ;
  assign y2195 = ~1'b0 ;
  assign y2196 = ~n5279 ;
  assign y2197 = ~1'b0 ;
  assign y2198 = n5282 ;
  assign y2199 = ~n5284 ;
  assign y2200 = ~1'b0 ;
  assign y2201 = ~1'b0 ;
  assign y2202 = n5285 ;
  assign y2203 = n5286 ;
  assign y2204 = ~n5292 ;
  assign y2205 = n5295 ;
  assign y2206 = ~n5297 ;
  assign y2207 = ~1'b0 ;
  assign y2208 = ~n5298 ;
  assign y2209 = ~n5300 ;
  assign y2210 = ~n5205 ;
  assign y2211 = ~n5306 ;
  assign y2212 = ~n5308 ;
  assign y2213 = ~n5310 ;
  assign y2214 = n5312 ;
  assign y2215 = ~1'b0 ;
  assign y2216 = ~n5316 ;
  assign y2217 = ~1'b0 ;
  assign y2218 = n5320 ;
  assign y2219 = ~1'b0 ;
  assign y2220 = n5321 ;
  assign y2221 = ~1'b0 ;
  assign y2222 = n5331 ;
  assign y2223 = ~1'b0 ;
  assign y2224 = n5333 ;
  assign y2225 = n5340 ;
  assign y2226 = ~n5344 ;
  assign y2227 = ~1'b0 ;
  assign y2228 = n5353 ;
  assign y2229 = ~n5355 ;
  assign y2230 = ~n5360 ;
  assign y2231 = ~1'b0 ;
  assign y2232 = ~1'b0 ;
  assign y2233 = ~n5365 ;
  assign y2234 = n5367 ;
  assign y2235 = n5371 ;
  assign y2236 = n5376 ;
  assign y2237 = ~n5378 ;
  assign y2238 = ~1'b0 ;
  assign y2239 = ~n5385 ;
  assign y2240 = ~n5387 ;
  assign y2241 = n5392 ;
  assign y2242 = ~n5397 ;
  assign y2243 = ~n5398 ;
  assign y2244 = ~1'b0 ;
  assign y2245 = ~n5404 ;
  assign y2246 = n5409 ;
  assign y2247 = n5410 ;
  assign y2248 = ~1'b0 ;
  assign y2249 = n5412 ;
  assign y2250 = ~n5414 ;
  assign y2251 = ~n5415 ;
  assign y2252 = ~n5416 ;
  assign y2253 = n5419 ;
  assign y2254 = ~1'b0 ;
  assign y2255 = ~n5421 ;
  assign y2256 = ~n5423 ;
  assign y2257 = ~n5429 ;
  assign y2258 = n5434 ;
  assign y2259 = ~n5437 ;
  assign y2260 = ~1'b0 ;
  assign y2261 = ~n5441 ;
  assign y2262 = ~n5446 ;
  assign y2263 = ~n5449 ;
  assign y2264 = ~n5454 ;
  assign y2265 = n5456 ;
  assign y2266 = n5458 ;
  assign y2267 = ~1'b0 ;
  assign y2268 = ~n5466 ;
  assign y2269 = n5472 ;
  assign y2270 = ~n5473 ;
  assign y2271 = ~1'b0 ;
  assign y2272 = ~1'b0 ;
  assign y2273 = ~1'b0 ;
  assign y2274 = ~n5475 ;
  assign y2275 = ~1'b0 ;
  assign y2276 = ~1'b0 ;
  assign y2277 = ~1'b0 ;
  assign y2278 = n5477 ;
  assign y2279 = ~n5479 ;
  assign y2280 = ~n5482 ;
  assign y2281 = ~1'b0 ;
  assign y2282 = n5483 ;
  assign y2283 = ~n5488 ;
  assign y2284 = 1'b0 ;
  assign y2285 = ~n5491 ;
  assign y2286 = ~1'b0 ;
  assign y2287 = ~n5493 ;
  assign y2288 = ~1'b0 ;
  assign y2289 = n5497 ;
  assign y2290 = ~n5499 ;
  assign y2291 = ~1'b0 ;
  assign y2292 = ~n5511 ;
  assign y2293 = ~1'b0 ;
  assign y2294 = n5515 ;
  assign y2295 = n5524 ;
  assign y2296 = ~n5533 ;
  assign y2297 = ~1'b0 ;
  assign y2298 = ~n5542 ;
  assign y2299 = ~n5545 ;
  assign y2300 = x71 ;
  assign y2301 = n5547 ;
  assign y2302 = ~1'b0 ;
  assign y2303 = ~n5548 ;
  assign y2304 = ~1'b0 ;
  assign y2305 = n5549 ;
  assign y2306 = ~1'b0 ;
  assign y2307 = n5553 ;
  assign y2308 = n5556 ;
  assign y2309 = ~n5559 ;
  assign y2310 = ~n5562 ;
  assign y2311 = ~n5565 ;
  assign y2312 = n5567 ;
  assign y2313 = ~n5571 ;
  assign y2314 = n5572 ;
  assign y2315 = ~n5145 ;
  assign y2316 = ~n5577 ;
  assign y2317 = 1'b0 ;
  assign y2318 = ~n5580 ;
  assign y2319 = ~1'b0 ;
  assign y2320 = n5587 ;
  assign y2321 = ~1'b0 ;
  assign y2322 = ~1'b0 ;
  assign y2323 = n5588 ;
  assign y2324 = n5596 ;
  assign y2325 = n5597 ;
  assign y2326 = ~n5604 ;
  assign y2327 = n5606 ;
  assign y2328 = ~n5610 ;
  assign y2329 = ~1'b0 ;
  assign y2330 = ~1'b0 ;
  assign y2331 = n5611 ;
  assign y2332 = ~n5612 ;
  assign y2333 = ~1'b0 ;
  assign y2334 = ~n5616 ;
  assign y2335 = ~1'b0 ;
  assign y2336 = ~1'b0 ;
  assign y2337 = n5620 ;
  assign y2338 = ~1'b0 ;
  assign y2339 = n2958 ;
  assign y2340 = ~1'b0 ;
  assign y2341 = ~1'b0 ;
  assign y2342 = ~n5631 ;
  assign y2343 = ~n5632 ;
  assign y2344 = ~n5635 ;
  assign y2345 = n5637 ;
  assign y2346 = ~1'b0 ;
  assign y2347 = ~n4845 ;
  assign y2348 = ~n5640 ;
  assign y2349 = ~n5650 ;
  assign y2350 = n5654 ;
  assign y2351 = n5655 ;
  assign y2352 = ~n5656 ;
  assign y2353 = ~n5662 ;
  assign y2354 = ~n5664 ;
  assign y2355 = n5669 ;
  assign y2356 = n5675 ;
  assign y2357 = ~1'b0 ;
  assign y2358 = ~n391 ;
  assign y2359 = ~1'b0 ;
  assign y2360 = n5681 ;
  assign y2361 = ~1'b0 ;
  assign y2362 = ~n5691 ;
  assign y2363 = ~n5692 ;
  assign y2364 = n5696 ;
  assign y2365 = ~n5699 ;
  assign y2366 = ~1'b0 ;
  assign y2367 = n5702 ;
  assign y2368 = n5703 ;
  assign y2369 = n5708 ;
  assign y2370 = ~1'b0 ;
  assign y2371 = ~1'b0 ;
  assign y2372 = ~1'b0 ;
  assign y2373 = n5711 ;
  assign y2374 = n5715 ;
  assign y2375 = ~1'b0 ;
  assign y2376 = ~n5717 ;
  assign y2377 = ~n5721 ;
  assign y2378 = ~n5722 ;
  assign y2379 = ~n5724 ;
  assign y2380 = ~1'b0 ;
  assign y2381 = ~n1397 ;
  assign y2382 = ~n5725 ;
  assign y2383 = n5726 ;
  assign y2384 = ~1'b0 ;
  assign y2385 = ~n5728 ;
  assign y2386 = ~n5734 ;
  assign y2387 = ~n2064 ;
  assign y2388 = n5736 ;
  assign y2389 = ~n5739 ;
  assign y2390 = ~n5741 ;
  assign y2391 = n5742 ;
  assign y2392 = ~n5756 ;
  assign y2393 = ~n5760 ;
  assign y2394 = ~n5761 ;
  assign y2395 = ~1'b0 ;
  assign y2396 = n5763 ;
  assign y2397 = ~1'b0 ;
  assign y2398 = ~1'b0 ;
  assign y2399 = ~n5765 ;
  assign y2400 = n5770 ;
  assign y2401 = ~n5772 ;
  assign y2402 = ~n5773 ;
  assign y2403 = n5776 ;
  assign y2404 = n5780 ;
  assign y2405 = n5783 ;
  assign y2406 = n5784 ;
  assign y2407 = n5792 ;
  assign y2408 = ~1'b0 ;
  assign y2409 = ~n5794 ;
  assign y2410 = n5796 ;
  assign y2411 = n1966 ;
  assign y2412 = ~n2928 ;
  assign y2413 = ~n5802 ;
  assign y2414 = ~n5805 ;
  assign y2415 = n5811 ;
  assign y2416 = ~n5812 ;
  assign y2417 = ~n5814 ;
  assign y2418 = ~n5815 ;
  assign y2419 = ~1'b0 ;
  assign y2420 = ~n5816 ;
  assign y2421 = n5822 ;
  assign y2422 = n5823 ;
  assign y2423 = ~n5826 ;
  assign y2424 = ~n5827 ;
  assign y2425 = ~n5829 ;
  assign y2426 = ~n5831 ;
  assign y2427 = ~1'b0 ;
  assign y2428 = n5833 ;
  assign y2429 = n5845 ;
  assign y2430 = ~1'b0 ;
  assign y2431 = n5846 ;
  assign y2432 = ~n5854 ;
  assign y2433 = ~n5858 ;
  assign y2434 = ~n5861 ;
  assign y2435 = ~1'b0 ;
  assign y2436 = n5866 ;
  assign y2437 = n5872 ;
  assign y2438 = ~1'b0 ;
  assign y2439 = n5874 ;
  assign y2440 = n5876 ;
  assign y2441 = ~n4169 ;
  assign y2442 = n5886 ;
  assign y2443 = ~1'b0 ;
  assign y2444 = ~1'b0 ;
  assign y2445 = ~n5887 ;
  assign y2446 = n5888 ;
  assign y2447 = ~n5889 ;
  assign y2448 = ~n5890 ;
  assign y2449 = ~n5891 ;
  assign y2450 = ~n5892 ;
  assign y2451 = ~n5896 ;
  assign y2452 = ~1'b0 ;
  assign y2453 = ~n5897 ;
  assign y2454 = ~n5899 ;
  assign y2455 = n2102 ;
  assign y2456 = ~n5906 ;
  assign y2457 = ~1'b0 ;
  assign y2458 = ~1'b0 ;
  assign y2459 = ~n5908 ;
  assign y2460 = n5909 ;
  assign y2461 = ~1'b0 ;
  assign y2462 = ~n5911 ;
  assign y2463 = n5913 ;
  assign y2464 = ~n5915 ;
  assign y2465 = ~n5922 ;
  assign y2466 = ~n5924 ;
  assign y2467 = ~n5929 ;
  assign y2468 = ~1'b0 ;
  assign y2469 = n5940 ;
  assign y2470 = n5944 ;
  assign y2471 = ~n5945 ;
  assign y2472 = n5946 ;
  assign y2473 = ~n5950 ;
  assign y2474 = ~n5955 ;
  assign y2475 = ~n5957 ;
  assign y2476 = n5101 ;
  assign y2477 = n5959 ;
  assign y2478 = ~n5962 ;
  assign y2479 = ~1'b0 ;
  assign y2480 = ~n5963 ;
  assign y2481 = n425 ;
  assign y2482 = ~1'b0 ;
  assign y2483 = ~n5964 ;
  assign y2484 = ~1'b0 ;
  assign y2485 = ~n5970 ;
  assign y2486 = ~n5972 ;
  assign y2487 = ~1'b0 ;
  assign y2488 = ~1'b0 ;
  assign y2489 = n5977 ;
  assign y2490 = ~1'b0 ;
  assign y2491 = n5985 ;
  assign y2492 = ~n5986 ;
  assign y2493 = ~1'b0 ;
  assign y2494 = ~n5988 ;
  assign y2495 = n5990 ;
  assign y2496 = n5994 ;
  assign y2497 = 1'b0 ;
  assign y2498 = n6000 ;
  assign y2499 = n6004 ;
  assign y2500 = ~n6005 ;
  assign y2501 = ~n6010 ;
  assign y2502 = 1'b0 ;
  assign y2503 = ~1'b0 ;
  assign y2504 = n6013 ;
  assign y2505 = ~n6014 ;
  assign y2506 = n6016 ;
  assign y2507 = ~n6020 ;
  assign y2508 = ~n6022 ;
  assign y2509 = ~1'b0 ;
  assign y2510 = ~1'b0 ;
  assign y2511 = ~n6028 ;
  assign y2512 = n6029 ;
  assign y2513 = n6030 ;
  assign y2514 = ~n6034 ;
  assign y2515 = n6035 ;
  assign y2516 = n6039 ;
  assign y2517 = ~n6046 ;
  assign y2518 = ~1'b0 ;
  assign y2519 = n6047 ;
  assign y2520 = ~n6053 ;
  assign y2521 = ~1'b0 ;
  assign y2522 = n6055 ;
  assign y2523 = ~1'b0 ;
  assign y2524 = ~1'b0 ;
  assign y2525 = ~n6056 ;
  assign y2526 = ~n6060 ;
  assign y2527 = n6061 ;
  assign y2528 = ~n6066 ;
  assign y2529 = ~n6067 ;
  assign y2530 = n6078 ;
  assign y2531 = n6081 ;
  assign y2532 = ~1'b0 ;
  assign y2533 = n6087 ;
  assign y2534 = ~n6088 ;
  assign y2535 = n6093 ;
  assign y2536 = ~n6099 ;
  assign y2537 = n4391 ;
  assign y2538 = ~n6101 ;
  assign y2539 = ~n6106 ;
  assign y2540 = n3556 ;
  assign y2541 = ~1'b0 ;
  assign y2542 = n6107 ;
  assign y2543 = n6111 ;
  assign y2544 = ~n6112 ;
  assign y2545 = n6116 ;
  assign y2546 = ~n6117 ;
  assign y2547 = n6126 ;
  assign y2548 = ~1'b0 ;
  assign y2549 = ~1'b0 ;
  assign y2550 = ~n6130 ;
  assign y2551 = ~1'b0 ;
  assign y2552 = n6131 ;
  assign y2553 = ~n1582 ;
  assign y2554 = ~1'b0 ;
  assign y2555 = ~1'b0 ;
  assign y2556 = ~n6132 ;
  assign y2557 = n6136 ;
  assign y2558 = ~1'b0 ;
  assign y2559 = ~n6143 ;
  assign y2560 = n2333 ;
  assign y2561 = ~1'b0 ;
  assign y2562 = ~n6144 ;
  assign y2563 = ~n6146 ;
  assign y2564 = ~n6151 ;
  assign y2565 = n6155 ;
  assign y2566 = ~1'b0 ;
  assign y2567 = ~1'b0 ;
  assign y2568 = n6162 ;
  assign y2569 = n6164 ;
  assign y2570 = ~n6168 ;
  assign y2571 = ~n6171 ;
  assign y2572 = ~n6172 ;
  assign y2573 = n6176 ;
  assign y2574 = ~n1175 ;
  assign y2575 = ~n770 ;
  assign y2576 = ~n6182 ;
  assign y2577 = n5117 ;
  assign y2578 = n6191 ;
  assign y2579 = ~1'b0 ;
  assign y2580 = n6193 ;
  assign y2581 = ~n3067 ;
  assign y2582 = ~1'b0 ;
  assign y2583 = 1'b0 ;
  assign y2584 = n6197 ;
  assign y2585 = ~n6204 ;
  assign y2586 = ~n6205 ;
  assign y2587 = n6212 ;
  assign y2588 = ~1'b0 ;
  assign y2589 = ~n6217 ;
  assign y2590 = n6220 ;
  assign y2591 = n6221 ;
  assign y2592 = ~n6227 ;
  assign y2593 = ~n6230 ;
  assign y2594 = ~n6231 ;
  assign y2595 = n6232 ;
  assign y2596 = ~n1918 ;
  assign y2597 = n6235 ;
  assign y2598 = ~n6236 ;
  assign y2599 = ~1'b0 ;
  assign y2600 = ~n6238 ;
  assign y2601 = 1'b0 ;
  assign y2602 = ~n6239 ;
  assign y2603 = n6243 ;
  assign y2604 = n6251 ;
  assign y2605 = ~n6255 ;
  assign y2606 = ~1'b0 ;
  assign y2607 = ~n6261 ;
  assign y2608 = ~n6266 ;
  assign y2609 = n6268 ;
  assign y2610 = ~n6269 ;
  assign y2611 = n6271 ;
  assign y2612 = n1040 ;
  assign y2613 = ~1'b0 ;
  assign y2614 = ~1'b0 ;
  assign y2615 = ~1'b0 ;
  assign y2616 = n6273 ;
  assign y2617 = ~n6277 ;
  assign y2618 = ~n6280 ;
  assign y2619 = ~n6284 ;
  assign y2620 = ~n6285 ;
  assign y2621 = ~1'b0 ;
  assign y2622 = ~1'b0 ;
  assign y2623 = ~1'b0 ;
  assign y2624 = n6287 ;
  assign y2625 = ~n6288 ;
  assign y2626 = n6289 ;
  assign y2627 = n6290 ;
  assign y2628 = ~n6295 ;
  assign y2629 = n6296 ;
  assign y2630 = ~n6299 ;
  assign y2631 = ~n6306 ;
  assign y2632 = ~n6307 ;
  assign y2633 = ~1'b0 ;
  assign y2634 = ~1'b0 ;
  assign y2635 = n6310 ;
  assign y2636 = ~n6314 ;
  assign y2637 = n6315 ;
  assign y2638 = n6319 ;
  assign y2639 = ~1'b0 ;
  assign y2640 = ~n6320 ;
  assign y2641 = n6322 ;
  assign y2642 = n6323 ;
  assign y2643 = ~n6327 ;
  assign y2644 = n6329 ;
  assign y2645 = ~n6336 ;
  assign y2646 = ~n6341 ;
  assign y2647 = ~1'b0 ;
  assign y2648 = ~n6343 ;
  assign y2649 = ~n6344 ;
  assign y2650 = ~n6346 ;
  assign y2651 = ~1'b0 ;
  assign y2652 = ~n6348 ;
  assign y2653 = ~n4760 ;
  assign y2654 = ~n6351 ;
  assign y2655 = ~1'b0 ;
  assign y2656 = n6360 ;
  assign y2657 = n6362 ;
  assign y2658 = ~1'b0 ;
  assign y2659 = ~n6364 ;
  assign y2660 = ~n6369 ;
  assign y2661 = 1'b0 ;
  assign y2662 = n6371 ;
  assign y2663 = n6376 ;
  assign y2664 = ~n6378 ;
  assign y2665 = ~1'b0 ;
  assign y2666 = ~n6379 ;
  assign y2667 = ~n6380 ;
  assign y2668 = ~n6381 ;
  assign y2669 = ~n6383 ;
  assign y2670 = ~n6385 ;
  assign y2671 = n6390 ;
  assign y2672 = n6391 ;
  assign y2673 = n1915 ;
  assign y2674 = n6394 ;
  assign y2675 = n6398 ;
  assign y2676 = ~n6400 ;
  assign y2677 = ~1'b0 ;
  assign y2678 = n6401 ;
  assign y2679 = ~n6408 ;
  assign y2680 = n6410 ;
  assign y2681 = n6412 ;
  assign y2682 = n892 ;
  assign y2683 = ~n6413 ;
  assign y2684 = ~1'b0 ;
  assign y2685 = n6419 ;
  assign y2686 = n6424 ;
  assign y2687 = n5916 ;
  assign y2688 = ~n6430 ;
  assign y2689 = ~n6434 ;
  assign y2690 = n625 ;
  assign y2691 = ~n6435 ;
  assign y2692 = ~1'b0 ;
  assign y2693 = n6436 ;
  assign y2694 = ~n6438 ;
  assign y2695 = ~n6439 ;
  assign y2696 = ~n6441 ;
  assign y2697 = n6446 ;
  assign y2698 = ~1'b0 ;
  assign y2699 = ~1'b0 ;
  assign y2700 = n6453 ;
  assign y2701 = n6459 ;
  assign y2702 = ~n6461 ;
  assign y2703 = n6466 ;
  assign y2704 = ~1'b0 ;
  assign y2705 = n6468 ;
  assign y2706 = ~n6470 ;
  assign y2707 = ~1'b0 ;
  assign y2708 = ~n6472 ;
  assign y2709 = n6473 ;
  assign y2710 = n6476 ;
  assign y2711 = ~1'b0 ;
  assign y2712 = n6479 ;
  assign y2713 = ~1'b0 ;
  assign y2714 = n6481 ;
  assign y2715 = ~n6483 ;
  assign y2716 = ~n3336 ;
  assign y2717 = ~n6489 ;
  assign y2718 = ~n6493 ;
  assign y2719 = ~n6494 ;
  assign y2720 = ~n6498 ;
  assign y2721 = ~n6499 ;
  assign y2722 = n6501 ;
  assign y2723 = ~n6504 ;
  assign y2724 = n6509 ;
  assign y2725 = n6515 ;
  assign y2726 = n6516 ;
  assign y2727 = n6517 ;
  assign y2728 = ~n6532 ;
  assign y2729 = n6536 ;
  assign y2730 = ~n6537 ;
  assign y2731 = n6545 ;
  assign y2732 = ~1'b0 ;
  assign y2733 = n1669 ;
  assign y2734 = n6548 ;
  assign y2735 = ~n6549 ;
  assign y2736 = ~1'b0 ;
  assign y2737 = ~1'b0 ;
  assign y2738 = n6550 ;
  assign y2739 = ~n6552 ;
  assign y2740 = ~1'b0 ;
  assign y2741 = n6553 ;
  assign y2742 = ~n6374 ;
  assign y2743 = n6555 ;
  assign y2744 = n6560 ;
  assign y2745 = ~n6567 ;
  assign y2746 = ~n6570 ;
  assign y2747 = ~n6573 ;
  assign y2748 = ~1'b0 ;
  assign y2749 = ~1'b0 ;
  assign y2750 = n6575 ;
  assign y2751 = n6579 ;
  assign y2752 = 1'b0 ;
  assign y2753 = n6580 ;
  assign y2754 = ~1'b0 ;
  assign y2755 = n6591 ;
  assign y2756 = ~1'b0 ;
  assign y2757 = ~1'b0 ;
  assign y2758 = ~n6593 ;
  assign y2759 = ~n6600 ;
  assign y2760 = ~n6605 ;
  assign y2761 = ~1'b0 ;
  assign y2762 = ~1'b0 ;
  assign y2763 = ~n6611 ;
  assign y2764 = ~n6617 ;
  assign y2765 = n6171 ;
  assign y2766 = n6621 ;
  assign y2767 = ~n6622 ;
  assign y2768 = n190 ;
  assign y2769 = ~n6624 ;
  assign y2770 = ~n6634 ;
  assign y2771 = ~n6636 ;
  assign y2772 = ~n6639 ;
  assign y2773 = ~n6641 ;
  assign y2774 = ~1'b0 ;
  assign y2775 = ~n6642 ;
  assign y2776 = ~n6643 ;
  assign y2777 = ~1'b0 ;
  assign y2778 = n6646 ;
  assign y2779 = ~1'b0 ;
  assign y2780 = ~n6647 ;
  assign y2781 = ~n6651 ;
  assign y2782 = n6655 ;
  assign y2783 = 1'b0 ;
  assign y2784 = n6656 ;
  assign y2785 = n6658 ;
  assign y2786 = n6660 ;
  assign y2787 = ~n6662 ;
  assign y2788 = ~n6663 ;
  assign y2789 = ~1'b0 ;
  assign y2790 = ~n6669 ;
  assign y2791 = ~n6671 ;
  assign y2792 = ~n6674 ;
  assign y2793 = n1765 ;
  assign y2794 = ~n6678 ;
  assign y2795 = ~1'b0 ;
  assign y2796 = ~1'b0 ;
  assign y2797 = ~1'b0 ;
  assign y2798 = n3633 ;
  assign y2799 = ~1'b0 ;
  assign y2800 = n6680 ;
  assign y2801 = n6681 ;
  assign y2802 = n6682 ;
  assign y2803 = ~n6683 ;
  assign y2804 = x2 ;
  assign y2805 = n6688 ;
  assign y2806 = n6691 ;
  assign y2807 = ~n6694 ;
  assign y2808 = n6696 ;
  assign y2809 = ~1'b0 ;
  assign y2810 = n6702 ;
  assign y2811 = ~n6706 ;
  assign y2812 = ~n6707 ;
  assign y2813 = n6708 ;
  assign y2814 = n6714 ;
  assign y2815 = ~1'b0 ;
  assign y2816 = ~n6716 ;
  assign y2817 = ~n6721 ;
  assign y2818 = n6726 ;
  assign y2819 = ~1'b0 ;
  assign y2820 = n6729 ;
  assign y2821 = n6736 ;
  assign y2822 = n6739 ;
  assign y2823 = ~1'b0 ;
  assign y2824 = ~n6742 ;
  assign y2825 = ~1'b0 ;
  assign y2826 = ~1'b0 ;
  assign y2827 = n6743 ;
  assign y2828 = ~1'b0 ;
  assign y2829 = n6745 ;
  assign y2830 = ~n6746 ;
  assign y2831 = ~n6750 ;
  assign y2832 = n6751 ;
  assign y2833 = n6755 ;
  assign y2834 = ~1'b0 ;
  assign y2835 = n6327 ;
  assign y2836 = ~1'b0 ;
  assign y2837 = ~n6758 ;
  assign y2838 = ~n6759 ;
  assign y2839 = n6761 ;
  assign y2840 = n6767 ;
  assign y2841 = n6768 ;
  assign y2842 = ~1'b0 ;
  assign y2843 = n6773 ;
  assign y2844 = ~n6778 ;
  assign y2845 = ~1'b0 ;
  assign y2846 = n6781 ;
  assign y2847 = ~n6784 ;
  assign y2848 = n1256 ;
  assign y2849 = ~n6785 ;
  assign y2850 = ~1'b0 ;
  assign y2851 = n6789 ;
  assign y2852 = ~1'b0 ;
  assign y2853 = ~1'b0 ;
  assign y2854 = ~n5043 ;
  assign y2855 = n6790 ;
  assign y2856 = ~n6795 ;
  assign y2857 = n6801 ;
  assign y2858 = ~n6802 ;
  assign y2859 = ~n6805 ;
  assign y2860 = ~1'b0 ;
  assign y2861 = ~n6809 ;
  assign y2862 = ~n6811 ;
  assign y2863 = ~n6812 ;
  assign y2864 = n6817 ;
  assign y2865 = ~1'b0 ;
  assign y2866 = ~n6818 ;
  assign y2867 = n6819 ;
  assign y2868 = n6825 ;
  assign y2869 = n6828 ;
  assign y2870 = ~1'b0 ;
  assign y2871 = ~1'b0 ;
  assign y2872 = ~n6835 ;
  assign y2873 = n6841 ;
  assign y2874 = ~1'b0 ;
  assign y2875 = n6842 ;
  assign y2876 = n6845 ;
  assign y2877 = ~n6848 ;
  assign y2878 = ~1'b0 ;
  assign y2879 = ~n6850 ;
  assign y2880 = ~n6852 ;
  assign y2881 = ~1'b0 ;
  assign y2882 = n1679 ;
  assign y2883 = n6856 ;
  assign y2884 = ~1'b0 ;
  assign y2885 = ~n6858 ;
  assign y2886 = ~1'b0 ;
  assign y2887 = n6859 ;
  assign y2888 = ~1'b0 ;
  assign y2889 = n3831 ;
  assign y2890 = ~n6862 ;
  assign y2891 = ~n6866 ;
  assign y2892 = ~1'b0 ;
  assign y2893 = ~1'b0 ;
  assign y2894 = ~n6870 ;
  assign y2895 = n6875 ;
  assign y2896 = ~1'b0 ;
  assign y2897 = ~n6880 ;
  assign y2898 = n6882 ;
  assign y2899 = n6885 ;
  assign y2900 = ~n6886 ;
  assign y2901 = ~1'b0 ;
  assign y2902 = ~1'b0 ;
  assign y2903 = ~n6893 ;
  assign y2904 = ~n6896 ;
  assign y2905 = ~1'b0 ;
  assign y2906 = ~1'b0 ;
  assign y2907 = n6897 ;
  assign y2908 = ~n6901 ;
  assign y2909 = ~n6912 ;
  assign y2910 = n6914 ;
  assign y2911 = n6916 ;
  assign y2912 = n6919 ;
  assign y2913 = ~1'b0 ;
  assign y2914 = ~n6925 ;
  assign y2915 = ~1'b0 ;
  assign y2916 = n6926 ;
  assign y2917 = ~n6928 ;
  assign y2918 = ~n6930 ;
  assign y2919 = n6931 ;
  assign y2920 = n6943 ;
  assign y2921 = ~n6948 ;
  assign y2922 = n2355 ;
  assign y2923 = ~1'b0 ;
  assign y2924 = ~n6951 ;
  assign y2925 = n4214 ;
  assign y2926 = ~n6954 ;
  assign y2927 = n6955 ;
  assign y2928 = n6964 ;
  assign y2929 = ~1'b0 ;
  assign y2930 = ~n6969 ;
  assign y2931 = ~n6975 ;
  assign y2932 = ~1'b0 ;
  assign y2933 = ~n6978 ;
  assign y2934 = n6983 ;
  assign y2935 = n6987 ;
  assign y2936 = ~n6988 ;
  assign y2937 = ~n6990 ;
  assign y2938 = n6999 ;
  assign y2939 = ~1'b0 ;
  assign y2940 = ~1'b0 ;
  assign y2941 = ~n7003 ;
  assign y2942 = ~1'b0 ;
  assign y2943 = n7008 ;
  assign y2944 = n7015 ;
  assign y2945 = ~1'b0 ;
  assign y2946 = ~n7025 ;
  assign y2947 = ~n7032 ;
  assign y2948 = n2841 ;
  assign y2949 = ~n7038 ;
  assign y2950 = ~1'b0 ;
  assign y2951 = n7040 ;
  assign y2952 = ~n7044 ;
  assign y2953 = ~n7047 ;
  assign y2954 = n7055 ;
  assign y2955 = ~n7057 ;
  assign y2956 = ~n984 ;
  assign y2957 = ~1'b0 ;
  assign y2958 = ~n7059 ;
  assign y2959 = ~n7062 ;
  assign y2960 = ~1'b0 ;
  assign y2961 = ~n7065 ;
  assign y2962 = n7068 ;
  assign y2963 = n7069 ;
  assign y2964 = n7071 ;
  assign y2965 = ~n7078 ;
  assign y2966 = ~n7081 ;
  assign y2967 = n7084 ;
  assign y2968 = ~n7086 ;
  assign y2969 = ~1'b0 ;
  assign y2970 = ~n654 ;
  assign y2971 = ~1'b0 ;
  assign y2972 = ~n7088 ;
  assign y2973 = ~1'b0 ;
  assign y2974 = ~1'b0 ;
  assign y2975 = ~n7089 ;
  assign y2976 = ~1'b0 ;
  assign y2977 = n7091 ;
  assign y2978 = ~1'b0 ;
  assign y2979 = ~n7099 ;
  assign y2980 = ~n7101 ;
  assign y2981 = n7106 ;
  assign y2982 = n7112 ;
  assign y2983 = n7114 ;
  assign y2984 = ~n4564 ;
  assign y2985 = n7119 ;
  assign y2986 = ~1'b0 ;
  assign y2987 = ~1'b0 ;
  assign y2988 = n7121 ;
  assign y2989 = ~n7126 ;
  assign y2990 = ~1'b0 ;
  assign y2991 = n7128 ;
  assign y2992 = n7130 ;
  assign y2993 = ~1'b0 ;
  assign y2994 = ~1'b0 ;
  assign y2995 = ~1'b0 ;
  assign y2996 = ~n7133 ;
  assign y2997 = ~n7135 ;
  assign y2998 = ~1'b0 ;
  assign y2999 = ~1'b0 ;
  assign y3000 = n7138 ;
  assign y3001 = ~1'b0 ;
  assign y3002 = ~n7143 ;
  assign y3003 = ~n7145 ;
  assign y3004 = n7146 ;
  assign y3005 = ~n7153 ;
  assign y3006 = n7154 ;
  assign y3007 = ~n7166 ;
  assign y3008 = n7169 ;
  assign y3009 = ~n7170 ;
  assign y3010 = ~n7171 ;
  assign y3011 = ~n7172 ;
  assign y3012 = ~1'b0 ;
  assign y3013 = n7173 ;
  assign y3014 = ~n7187 ;
  assign y3015 = n7190 ;
  assign y3016 = ~n7193 ;
  assign y3017 = n7197 ;
  assign y3018 = ~1'b0 ;
  assign y3019 = ~1'b0 ;
  assign y3020 = ~n7203 ;
  assign y3021 = 1'b0 ;
  assign y3022 = n7204 ;
  assign y3023 = n7208 ;
  assign y3024 = ~1'b0 ;
  assign y3025 = ~n7210 ;
  assign y3026 = 1'b0 ;
  assign y3027 = ~1'b0 ;
  assign y3028 = n7212 ;
  assign y3029 = n7215 ;
  assign y3030 = n7218 ;
  assign y3031 = ~n7220 ;
  assign y3032 = ~1'b0 ;
  assign y3033 = ~n7225 ;
  assign y3034 = n4330 ;
  assign y3035 = ~n7226 ;
  assign y3036 = ~1'b0 ;
  assign y3037 = ~n7227 ;
  assign y3038 = n7233 ;
  assign y3039 = ~1'b0 ;
  assign y3040 = n6815 ;
  assign y3041 = ~n7235 ;
  assign y3042 = ~n7236 ;
  assign y3043 = ~1'b0 ;
  assign y3044 = ~1'b0 ;
  assign y3045 = n7238 ;
  assign y3046 = ~n7239 ;
  assign y3047 = ~n7240 ;
  assign y3048 = ~1'b0 ;
  assign y3049 = ~1'b0 ;
  assign y3050 = ~n7241 ;
  assign y3051 = 1'b0 ;
  assign y3052 = ~n7242 ;
  assign y3053 = ~n7245 ;
  assign y3054 = ~1'b0 ;
  assign y3055 = ~1'b0 ;
  assign y3056 = n7249 ;
  assign y3057 = ~n7254 ;
  assign y3058 = ~1'b0 ;
  assign y3059 = ~n7255 ;
  assign y3060 = n4107 ;
  assign y3061 = ~1'b0 ;
  assign y3062 = n7259 ;
  assign y3063 = n7260 ;
  assign y3064 = ~n7262 ;
  assign y3065 = ~n7263 ;
  assign y3066 = ~n7268 ;
  assign y3067 = ~n7279 ;
  assign y3068 = ~1'b0 ;
  assign y3069 = ~1'b0 ;
  assign y3070 = ~n7286 ;
  assign y3071 = ~n7287 ;
  assign y3072 = ~1'b0 ;
  assign y3073 = ~1'b0 ;
  assign y3074 = ~n7288 ;
  assign y3075 = ~1'b0 ;
  assign y3076 = n7289 ;
  assign y3077 = ~n7290 ;
  assign y3078 = n1821 ;
  assign y3079 = n7294 ;
  assign y3080 = n7296 ;
  assign y3081 = n7297 ;
  assign y3082 = ~n7298 ;
  assign y3083 = n7303 ;
  assign y3084 = n7304 ;
  assign y3085 = n7306 ;
  assign y3086 = ~1'b0 ;
  assign y3087 = ~1'b0 ;
  assign y3088 = ~n7308 ;
  assign y3089 = ~n7309 ;
  assign y3090 = n7313 ;
  assign y3091 = n7316 ;
  assign y3092 = n7320 ;
  assign y3093 = n7321 ;
  assign y3094 = ~n4650 ;
  assign y3095 = ~1'b0 ;
  assign y3096 = ~1'b0 ;
  assign y3097 = ~1'b0 ;
  assign y3098 = ~n7324 ;
  assign y3099 = ~n7325 ;
  assign y3100 = ~n7326 ;
  assign y3101 = ~1'b0 ;
  assign y3102 = n7329 ;
  assign y3103 = ~n7330 ;
  assign y3104 = n7338 ;
  assign y3105 = n7339 ;
  assign y3106 = ~1'b0 ;
  assign y3107 = n7340 ;
  assign y3108 = n7341 ;
  assign y3109 = ~n7351 ;
  assign y3110 = ~n7352 ;
  assign y3111 = ~n7357 ;
  assign y3112 = 1'b0 ;
  assign y3113 = ~n7365 ;
  assign y3114 = ~1'b0 ;
  assign y3115 = ~n7367 ;
  assign y3116 = n7372 ;
  assign y3117 = ~n7374 ;
  assign y3118 = n7380 ;
  assign y3119 = n7382 ;
  assign y3120 = ~1'b0 ;
  assign y3121 = n7383 ;
  assign y3122 = n7384 ;
  assign y3123 = ~n7386 ;
  assign y3124 = n4219 ;
  assign y3125 = ~1'b0 ;
  assign y3126 = ~1'b0 ;
  assign y3127 = n7389 ;
  assign y3128 = ~1'b0 ;
  assign y3129 = ~n7390 ;
  assign y3130 = ~n7393 ;
  assign y3131 = ~1'b0 ;
  assign y3132 = ~n7399 ;
  assign y3133 = ~1'b0 ;
  assign y3134 = ~1'b0 ;
  assign y3135 = n7400 ;
  assign y3136 = ~n7407 ;
  assign y3137 = n7413 ;
  assign y3138 = n7418 ;
  assign y3139 = ~1'b0 ;
  assign y3140 = n7421 ;
  assign y3141 = ~1'b0 ;
  assign y3142 = ~n7422 ;
  assign y3143 = ~1'b0 ;
  assign y3144 = ~1'b0 ;
  assign y3145 = ~n7424 ;
  assign y3146 = ~n7428 ;
  assign y3147 = ~1'b0 ;
  assign y3148 = ~n7432 ;
  assign y3149 = ~1'b0 ;
  assign y3150 = ~1'b0 ;
  assign y3151 = ~1'b0 ;
  assign y3152 = ~n7438 ;
  assign y3153 = n7442 ;
  assign y3154 = ~1'b0 ;
  assign y3155 = n7448 ;
  assign y3156 = ~n7449 ;
  assign y3157 = ~1'b0 ;
  assign y3158 = ~n7451 ;
  assign y3159 = 1'b0 ;
  assign y3160 = n4369 ;
  assign y3161 = ~1'b0 ;
  assign y3162 = n4097 ;
  assign y3163 = n7453 ;
  assign y3164 = ~1'b0 ;
  assign y3165 = ~1'b0 ;
  assign y3166 = n7455 ;
  assign y3167 = ~n7457 ;
  assign y3168 = n7460 ;
  assign y3169 = ~1'b0 ;
  assign y3170 = ~1'b0 ;
  assign y3171 = n7463 ;
  assign y3172 = ~1'b0 ;
  assign y3173 = ~1'b0 ;
  assign y3174 = ~1'b0 ;
  assign y3175 = n2365 ;
  assign y3176 = n7465 ;
  assign y3177 = 1'b0 ;
  assign y3178 = ~n7478 ;
  assign y3179 = n7479 ;
  assign y3180 = ~1'b0 ;
  assign y3181 = n7482 ;
  assign y3182 = ~n7485 ;
  assign y3183 = n7488 ;
  assign y3184 = n7491 ;
  assign y3185 = ~n7496 ;
  assign y3186 = ~n7502 ;
  assign y3187 = n7511 ;
  assign y3188 = ~1'b0 ;
  assign y3189 = n7514 ;
  assign y3190 = ~n7516 ;
  assign y3191 = ~n7524 ;
  assign y3192 = ~n7525 ;
  assign y3193 = ~1'b0 ;
  assign y3194 = ~n7526 ;
  assign y3195 = ~1'b0 ;
  assign y3196 = ~n7527 ;
  assign y3197 = ~n7536 ;
  assign y3198 = 1'b0 ;
  assign y3199 = ~1'b0 ;
  assign y3200 = n7539 ;
  assign y3201 = n7545 ;
  assign y3202 = ~n7547 ;
  assign y3203 = n4504 ;
  assign y3204 = ~1'b0 ;
  assign y3205 = n7557 ;
  assign y3206 = n7559 ;
  assign y3207 = ~1'b0 ;
  assign y3208 = ~n7560 ;
  assign y3209 = n7562 ;
  assign y3210 = ~n3981 ;
  assign y3211 = ~1'b0 ;
  assign y3212 = n7567 ;
  assign y3213 = ~n7570 ;
  assign y3214 = n7573 ;
  assign y3215 = ~n7576 ;
  assign y3216 = ~1'b0 ;
  assign y3217 = ~1'b0 ;
  assign y3218 = n4394 ;
  assign y3219 = ~n7580 ;
  assign y3220 = n7583 ;
  assign y3221 = n7587 ;
  assign y3222 = ~n7594 ;
  assign y3223 = n7595 ;
  assign y3224 = ~n7604 ;
  assign y3225 = n7608 ;
  assign y3226 = n7609 ;
  assign y3227 = n7614 ;
  assign y3228 = ~1'b0 ;
  assign y3229 = ~n7616 ;
  assign y3230 = ~1'b0 ;
  assign y3231 = ~n7618 ;
  assign y3232 = ~1'b0 ;
  assign y3233 = n7619 ;
  assign y3234 = ~1'b0 ;
  assign y3235 = n7622 ;
  assign y3236 = ~n7623 ;
  assign y3237 = ~n7625 ;
  assign y3238 = ~1'b0 ;
  assign y3239 = ~1'b0 ;
  assign y3240 = ~1'b0 ;
  assign y3241 = ~n7630 ;
  assign y3242 = ~n7631 ;
  assign y3243 = ~n7635 ;
  assign y3244 = n7638 ;
  assign y3245 = 1'b0 ;
  assign y3246 = ~1'b0 ;
  assign y3247 = ~1'b0 ;
  assign y3248 = n7641 ;
  assign y3249 = ~n6097 ;
  assign y3250 = ~n7648 ;
  assign y3251 = ~n7649 ;
  assign y3252 = n7660 ;
  assign y3253 = n7666 ;
  assign y3254 = ~n7667 ;
  assign y3255 = ~n7672 ;
  assign y3256 = ~1'b0 ;
  assign y3257 = n7673 ;
  assign y3258 = ~1'b0 ;
  assign y3259 = n7682 ;
  assign y3260 = n7683 ;
  assign y3261 = n7685 ;
  assign y3262 = ~n2958 ;
  assign y3263 = n7687 ;
  assign y3264 = ~1'b0 ;
  assign y3265 = ~n7689 ;
  assign y3266 = ~n7692 ;
  assign y3267 = n5076 ;
  assign y3268 = ~1'b0 ;
  assign y3269 = ~n7695 ;
  assign y3270 = ~n7698 ;
  assign y3271 = ~n3528 ;
  assign y3272 = ~n7700 ;
  assign y3273 = ~n7703 ;
  assign y3274 = ~n7713 ;
  assign y3275 = ~n7715 ;
  assign y3276 = n7720 ;
  assign y3277 = ~n7721 ;
  assign y3278 = ~1'b0 ;
  assign y3279 = n7723 ;
  assign y3280 = n3710 ;
  assign y3281 = ~n7724 ;
  assign y3282 = n7729 ;
  assign y3283 = n7735 ;
  assign y3284 = n7737 ;
  assign y3285 = n7739 ;
  assign y3286 = ~n7740 ;
  assign y3287 = ~n7746 ;
  assign y3288 = ~n7748 ;
  assign y3289 = n7752 ;
  assign y3290 = n7756 ;
  assign y3291 = ~n7757 ;
  assign y3292 = n7003 ;
  assign y3293 = n7759 ;
  assign y3294 = ~n7771 ;
  assign y3295 = ~1'b0 ;
  assign y3296 = ~1'b0 ;
  assign y3297 = ~1'b0 ;
  assign y3298 = n7773 ;
  assign y3299 = ~n7774 ;
  assign y3300 = ~n7776 ;
  assign y3301 = ~n7780 ;
  assign y3302 = ~1'b0 ;
  assign y3303 = n7785 ;
  assign y3304 = ~n7790 ;
  assign y3305 = n7791 ;
  assign y3306 = ~1'b0 ;
  assign y3307 = ~n7792 ;
  assign y3308 = ~1'b0 ;
  assign y3309 = ~n7577 ;
  assign y3310 = n7794 ;
  assign y3311 = ~n7797 ;
  assign y3312 = ~1'b0 ;
  assign y3313 = ~1'b0 ;
  assign y3314 = ~n7798 ;
  assign y3315 = n7800 ;
  assign y3316 = ~n1739 ;
  assign y3317 = n7802 ;
  assign y3318 = ~n7803 ;
  assign y3319 = n7812 ;
  assign y3320 = ~n7813 ;
  assign y3321 = ~n7816 ;
  assign y3322 = ~n7820 ;
  assign y3323 = ~n7825 ;
  assign y3324 = ~n7828 ;
  assign y3325 = n7835 ;
  assign y3326 = ~n7837 ;
  assign y3327 = n7839 ;
  assign y3328 = ~1'b0 ;
  assign y3329 = ~1'b0 ;
  assign y3330 = ~1'b0 ;
  assign y3331 = ~n7840 ;
  assign y3332 = ~n7841 ;
  assign y3333 = ~n7848 ;
  assign y3334 = ~n7857 ;
  assign y3335 = ~n7858 ;
  assign y3336 = ~n7859 ;
  assign y3337 = ~n7861 ;
  assign y3338 = ~1'b0 ;
  assign y3339 = ~1'b0 ;
  assign y3340 = ~n7864 ;
  assign y3341 = n7865 ;
  assign y3342 = ~n7867 ;
  assign y3343 = n7868 ;
  assign y3344 = ~1'b0 ;
  assign y3345 = ~n7871 ;
  assign y3346 = ~1'b0 ;
  assign y3347 = ~n7872 ;
  assign y3348 = n7873 ;
  assign y3349 = n7878 ;
  assign y3350 = n7882 ;
  assign y3351 = ~n7885 ;
  assign y3352 = n7888 ;
  assign y3353 = n7891 ;
  assign y3354 = ~1'b0 ;
  assign y3355 = ~1'b0 ;
  assign y3356 = n7896 ;
  assign y3357 = ~1'b0 ;
  assign y3358 = n7897 ;
  assign y3359 = ~1'b0 ;
  assign y3360 = ~n7909 ;
  assign y3361 = ~n7911 ;
  assign y3362 = ~n4157 ;
  assign y3363 = ~n7913 ;
  assign y3364 = ~n7922 ;
  assign y3365 = ~1'b0 ;
  assign y3366 = ~n7927 ;
  assign y3367 = ~n7933 ;
  assign y3368 = ~n7934 ;
  assign y3369 = ~1'b0 ;
  assign y3370 = ~n7935 ;
  assign y3371 = n7943 ;
  assign y3372 = n3994 ;
  assign y3373 = ~1'b0 ;
  assign y3374 = ~1'b0 ;
  assign y3375 = ~n7944 ;
  assign y3376 = ~1'b0 ;
  assign y3377 = ~1'b0 ;
  assign y3378 = n7946 ;
  assign y3379 = ~1'b0 ;
  assign y3380 = ~1'b0 ;
  assign y3381 = ~n7947 ;
  assign y3382 = 1'b0 ;
  assign y3383 = n7951 ;
  assign y3384 = n7954 ;
  assign y3385 = ~1'b0 ;
  assign y3386 = n7957 ;
  assign y3387 = n2649 ;
  assign y3388 = ~1'b0 ;
  assign y3389 = n7958 ;
  assign y3390 = n7962 ;
  assign y3391 = ~1'b0 ;
  assign y3392 = ~1'b0 ;
  assign y3393 = ~n7963 ;
  assign y3394 = ~n7964 ;
  assign y3395 = ~n7968 ;
  assign y3396 = n7969 ;
  assign y3397 = ~n7973 ;
  assign y3398 = ~1'b0 ;
  assign y3399 = ~1'b0 ;
  assign y3400 = n7983 ;
  assign y3401 = ~1'b0 ;
  assign y3402 = ~n7986 ;
  assign y3403 = ~n7987 ;
  assign y3404 = ~n7989 ;
  assign y3405 = n7990 ;
  assign y3406 = n7991 ;
  assign y3407 = ~n7992 ;
  assign y3408 = ~1'b0 ;
  assign y3409 = ~1'b0 ;
  assign y3410 = ~1'b0 ;
  assign y3411 = ~1'b0 ;
  assign y3412 = ~1'b0 ;
  assign y3413 = n7993 ;
  assign y3414 = ~n7995 ;
  assign y3415 = n8001 ;
  assign y3416 = n8004 ;
  assign y3417 = n8005 ;
  assign y3418 = n8008 ;
  assign y3419 = ~1'b0 ;
  assign y3420 = ~n8009 ;
  assign y3421 = n8015 ;
  assign y3422 = ~1'b0 ;
  assign y3423 = ~1'b0 ;
  assign y3424 = ~1'b0 ;
  assign y3425 = ~n8029 ;
  assign y3426 = ~n8030 ;
  assign y3427 = n8038 ;
  assign y3428 = ~n4050 ;
  assign y3429 = ~n8040 ;
  assign y3430 = ~1'b0 ;
  assign y3431 = ~1'b0 ;
  assign y3432 = n8046 ;
  assign y3433 = ~n8055 ;
  assign y3434 = n8056 ;
  assign y3435 = n8061 ;
  assign y3436 = ~1'b0 ;
  assign y3437 = n8062 ;
  assign y3438 = ~n8063 ;
  assign y3439 = ~n8071 ;
  assign y3440 = ~n6138 ;
  assign y3441 = ~n8078 ;
  assign y3442 = n8079 ;
  assign y3443 = ~n8082 ;
  assign y3444 = ~1'b0 ;
  assign y3445 = n2632 ;
  assign y3446 = ~1'b0 ;
  assign y3447 = n8083 ;
  assign y3448 = n8086 ;
  assign y3449 = ~1'b0 ;
  assign y3450 = ~n8087 ;
  assign y3451 = ~n8091 ;
  assign y3452 = ~n8093 ;
  assign y3453 = n8094 ;
  assign y3454 = n8097 ;
  assign y3455 = n8100 ;
  assign y3456 = n8103 ;
  assign y3457 = n8107 ;
  assign y3458 = ~n8113 ;
  assign y3459 = n8114 ;
  assign y3460 = ~1'b0 ;
  assign y3461 = ~n8115 ;
  assign y3462 = ~1'b0 ;
  assign y3463 = n8116 ;
  assign y3464 = ~1'b0 ;
  assign y3465 = n8118 ;
  assign y3466 = ~n8120 ;
  assign y3467 = ~n3193 ;
  assign y3468 = ~n8121 ;
  assign y3469 = ~n8123 ;
  assign y3470 = n8126 ;
  assign y3471 = ~n895 ;
  assign y3472 = ~n8127 ;
  assign y3473 = ~n8128 ;
  assign y3474 = ~n1452 ;
  assign y3475 = n8134 ;
  assign y3476 = ~1'b0 ;
  assign y3477 = ~n8135 ;
  assign y3478 = ~1'b0 ;
  assign y3479 = ~n8136 ;
  assign y3480 = ~1'b0 ;
  assign y3481 = ~n8137 ;
  assign y3482 = n8140 ;
  assign y3483 = n8141 ;
  assign y3484 = ~n8145 ;
  assign y3485 = n8146 ;
  assign y3486 = n8147 ;
  assign y3487 = ~n8154 ;
  assign y3488 = ~n8162 ;
  assign y3489 = ~n8165 ;
  assign y3490 = ~n8166 ;
  assign y3491 = ~n8167 ;
  assign y3492 = ~n8170 ;
  assign y3493 = ~1'b0 ;
  assign y3494 = n8171 ;
  assign y3495 = n8172 ;
  assign y3496 = n8180 ;
  assign y3497 = n8182 ;
  assign y3498 = n8183 ;
  assign y3499 = ~1'b0 ;
  assign y3500 = ~n8189 ;
  assign y3501 = ~1'b0 ;
  assign y3502 = ~n8193 ;
  assign y3503 = n1382 ;
  assign y3504 = ~1'b0 ;
  assign y3505 = ~n8195 ;
  assign y3506 = ~n8197 ;
  assign y3507 = ~1'b0 ;
  assign y3508 = ~1'b0 ;
  assign y3509 = n8199 ;
  assign y3510 = ~n8200 ;
  assign y3511 = ~1'b0 ;
  assign y3512 = ~n8204 ;
  assign y3513 = ~1'b0 ;
  assign y3514 = n8206 ;
  assign y3515 = ~1'b0 ;
  assign y3516 = ~n8208 ;
  assign y3517 = n8210 ;
  assign y3518 = ~1'b0 ;
  assign y3519 = n8213 ;
  assign y3520 = ~1'b0 ;
  assign y3521 = ~1'b0 ;
  assign y3522 = ~1'b0 ;
  assign y3523 = ~n8214 ;
  assign y3524 = n8220 ;
  assign y3525 = n8222 ;
  assign y3526 = ~1'b0 ;
  assign y3527 = ~1'b0 ;
  assign y3528 = ~n8227 ;
  assign y3529 = ~1'b0 ;
  assign y3530 = ~1'b0 ;
  assign y3531 = n8229 ;
  assign y3532 = n8232 ;
  assign y3533 = n8245 ;
  assign y3534 = ~n8248 ;
  assign y3535 = ~1'b0 ;
  assign y3536 = ~n8250 ;
  assign y3537 = ~n8252 ;
  assign y3538 = ~1'b0 ;
  assign y3539 = ~n8256 ;
  assign y3540 = ~n8260 ;
  assign y3541 = ~n8262 ;
  assign y3542 = 1'b0 ;
  assign y3543 = n8264 ;
  assign y3544 = ~1'b0 ;
  assign y3545 = ~n8269 ;
  assign y3546 = ~n8272 ;
  assign y3547 = ~n8275 ;
  assign y3548 = ~1'b0 ;
  assign y3549 = ~n8277 ;
  assign y3550 = ~n5752 ;
  assign y3551 = n8278 ;
  assign y3552 = ~n8282 ;
  assign y3553 = n8286 ;
  assign y3554 = ~1'b0 ;
  assign y3555 = ~n8288 ;
  assign y3556 = ~1'b0 ;
  assign y3557 = n8293 ;
  assign y3558 = ~n8296 ;
  assign y3559 = ~n8302 ;
  assign y3560 = ~n8303 ;
  assign y3561 = ~n8305 ;
  assign y3562 = ~n8306 ;
  assign y3563 = ~n8315 ;
  assign y3564 = ~n8322 ;
  assign y3565 = ~1'b0 ;
  assign y3566 = n8324 ;
  assign y3567 = ~n8326 ;
  assign y3568 = ~1'b0 ;
  assign y3569 = ~n8328 ;
  assign y3570 = ~1'b0 ;
  assign y3571 = ~n8329 ;
  assign y3572 = ~n8332 ;
  assign y3573 = 1'b0 ;
  assign y3574 = n8340 ;
  assign y3575 = n8342 ;
  assign y3576 = ~n8344 ;
  assign y3577 = ~1'b0 ;
  assign y3578 = n8345 ;
  assign y3579 = ~n8349 ;
  assign y3580 = ~1'b0 ;
  assign y3581 = ~n8351 ;
  assign y3582 = n8354 ;
  assign y3583 = n8356 ;
  assign y3584 = n8366 ;
  assign y3585 = 1'b0 ;
  assign y3586 = ~n8367 ;
  assign y3587 = n4064 ;
  assign y3588 = ~1'b0 ;
  assign y3589 = n8368 ;
  assign y3590 = ~n8369 ;
  assign y3591 = ~1'b0 ;
  assign y3592 = ~n1578 ;
  assign y3593 = ~n8374 ;
  assign y3594 = ~n8380 ;
  assign y3595 = n4512 ;
  assign y3596 = ~n8381 ;
  assign y3597 = n8382 ;
  assign y3598 = ~1'b0 ;
  assign y3599 = n8384 ;
  assign y3600 = n8385 ;
  assign y3601 = n8387 ;
  assign y3602 = ~1'b0 ;
  assign y3603 = n8393 ;
  assign y3604 = ~n8399 ;
  assign y3605 = n8404 ;
  assign y3606 = ~n8415 ;
  assign y3607 = n8424 ;
  assign y3608 = n8426 ;
  assign y3609 = ~n8428 ;
  assign y3610 = ~n8429 ;
  assign y3611 = n8434 ;
  assign y3612 = ~n8436 ;
  assign y3613 = n2877 ;
  assign y3614 = ~n8441 ;
  assign y3615 = n8449 ;
  assign y3616 = n8452 ;
  assign y3617 = ~1'b0 ;
  assign y3618 = ~n8453 ;
  assign y3619 = ~n8454 ;
  assign y3620 = n8459 ;
  assign y3621 = ~1'b0 ;
  assign y3622 = ~1'b0 ;
  assign y3623 = n8461 ;
  assign y3624 = n8462 ;
  assign y3625 = ~n5063 ;
  assign y3626 = ~n8464 ;
  assign y3627 = n8467 ;
  assign y3628 = ~n8469 ;
  assign y3629 = n8470 ;
  assign y3630 = n8471 ;
  assign y3631 = ~1'b0 ;
  assign y3632 = ~1'b0 ;
  assign y3633 = ~n8476 ;
  assign y3634 = ~n8478 ;
  assign y3635 = ~1'b0 ;
  assign y3636 = n8480 ;
  assign y3637 = ~n8484 ;
  assign y3638 = ~n8486 ;
  assign y3639 = n8490 ;
  assign y3640 = ~n8493 ;
  assign y3641 = n8496 ;
  assign y3642 = ~1'b0 ;
  assign y3643 = n8499 ;
  assign y3644 = ~n8500 ;
  assign y3645 = n8503 ;
  assign y3646 = n8504 ;
  assign y3647 = n8505 ;
  assign y3648 = n8507 ;
  assign y3649 = n8510 ;
  assign y3650 = ~n8514 ;
  assign y3651 = ~n8515 ;
  assign y3652 = n8516 ;
  assign y3653 = ~n8522 ;
  assign y3654 = ~1'b0 ;
  assign y3655 = n8526 ;
  assign y3656 = ~n8534 ;
  assign y3657 = n8544 ;
  assign y3658 = ~n8548 ;
  assign y3659 = n8550 ;
  assign y3660 = n6558 ;
  assign y3661 = ~n8553 ;
  assign y3662 = ~1'b0 ;
  assign y3663 = n8556 ;
  assign y3664 = ~1'b0 ;
  assign y3665 = ~n8558 ;
  assign y3666 = ~n8559 ;
  assign y3667 = ~n8560 ;
  assign y3668 = n8561 ;
  assign y3669 = n8563 ;
  assign y3670 = ~n8566 ;
  assign y3671 = n8568 ;
  assign y3672 = ~1'b0 ;
  assign y3673 = n8570 ;
  assign y3674 = ~1'b0 ;
  assign y3675 = n8573 ;
  assign y3676 = 1'b0 ;
  assign y3677 = n8574 ;
  assign y3678 = n8577 ;
  assign y3679 = ~1'b0 ;
  assign y3680 = ~1'b0 ;
  assign y3681 = n8579 ;
  assign y3682 = n8581 ;
  assign y3683 = ~1'b0 ;
  assign y3684 = ~n8590 ;
  assign y3685 = n8592 ;
  assign y3686 = n8596 ;
  assign y3687 = ~n8597 ;
  assign y3688 = ~1'b0 ;
  assign y3689 = ~1'b0 ;
  assign y3690 = ~n8598 ;
  assign y3691 = ~n8600 ;
  assign y3692 = ~n8602 ;
  assign y3693 = n8611 ;
  assign y3694 = n8613 ;
  assign y3695 = ~n8615 ;
  assign y3696 = ~1'b0 ;
  assign y3697 = ~x63 ;
  assign y3698 = n8621 ;
  assign y3699 = ~n8626 ;
  assign y3700 = ~1'b0 ;
  assign y3701 = n8630 ;
  assign y3702 = n8634 ;
  assign y3703 = n8636 ;
  assign y3704 = n8638 ;
  assign y3705 = n8649 ;
  assign y3706 = ~n8652 ;
  assign y3707 = n8653 ;
  assign y3708 = n8655 ;
  assign y3709 = ~n8657 ;
  assign y3710 = n8659 ;
  assign y3711 = ~n8660 ;
  assign y3712 = ~1'b0 ;
  assign y3713 = n8663 ;
  assign y3714 = n8664 ;
  assign y3715 = n8665 ;
  assign y3716 = n8666 ;
  assign y3717 = n8669 ;
  assign y3718 = ~n8671 ;
  assign y3719 = n8674 ;
  assign y3720 = n8678 ;
  assign y3721 = ~n8682 ;
  assign y3722 = n8684 ;
  assign y3723 = ~n8692 ;
  assign y3724 = ~n8700 ;
  assign y3725 = ~1'b0 ;
  assign y3726 = ~1'b0 ;
  assign y3727 = ~n8703 ;
  assign y3728 = n8705 ;
  assign y3729 = ~n8707 ;
  assign y3730 = ~n8712 ;
  assign y3731 = ~1'b0 ;
  assign y3732 = ~n997 ;
  assign y3733 = 1'b0 ;
  assign y3734 = ~n8715 ;
  assign y3735 = ~1'b0 ;
  assign y3736 = n5389 ;
  assign y3737 = ~1'b0 ;
  assign y3738 = ~n8716 ;
  assign y3739 = ~n8717 ;
  assign y3740 = ~n8718 ;
  assign y3741 = ~n8722 ;
  assign y3742 = n8723 ;
  assign y3743 = ~1'b0 ;
  assign y3744 = ~n8725 ;
  assign y3745 = n7169 ;
  assign y3746 = ~1'b0 ;
  assign y3747 = ~n8729 ;
  assign y3748 = n8730 ;
  assign y3749 = ~n8732 ;
  assign y3750 = n8733 ;
  assign y3751 = ~n8734 ;
  assign y3752 = ~1'b0 ;
  assign y3753 = ~n8740 ;
  assign y3754 = ~n8742 ;
  assign y3755 = ~1'b0 ;
  assign y3756 = ~n8743 ;
  assign y3757 = ~1'b0 ;
  assign y3758 = ~1'b0 ;
  assign y3759 = n8747 ;
  assign y3760 = ~n8749 ;
  assign y3761 = 1'b0 ;
  assign y3762 = n8753 ;
  assign y3763 = ~1'b0 ;
  assign y3764 = ~n8756 ;
  assign y3765 = n8758 ;
  assign y3766 = n3076 ;
  assign y3767 = n8764 ;
  assign y3768 = ~n8773 ;
  assign y3769 = ~1'b0 ;
  assign y3770 = ~1'b0 ;
  assign y3771 = ~n8775 ;
  assign y3772 = ~1'b0 ;
  assign y3773 = ~1'b0 ;
  assign y3774 = ~1'b0 ;
  assign y3775 = ~n8777 ;
  assign y3776 = ~1'b0 ;
  assign y3777 = ~1'b0 ;
  assign y3778 = n8779 ;
  assign y3779 = n8787 ;
  assign y3780 = ~n8794 ;
  assign y3781 = n2053 ;
  assign y3782 = n8798 ;
  assign y3783 = ~1'b0 ;
  assign y3784 = n8801 ;
  assign y3785 = n8803 ;
  assign y3786 = ~1'b0 ;
  assign y3787 = ~1'b0 ;
  assign y3788 = n8807 ;
  assign y3789 = n8809 ;
  assign y3790 = n8811 ;
  assign y3791 = n8813 ;
  assign y3792 = ~1'b0 ;
  assign y3793 = n8817 ;
  assign y3794 = ~n8820 ;
  assign y3795 = ~1'b0 ;
  assign y3796 = n8821 ;
  assign y3797 = ~1'b0 ;
  assign y3798 = ~1'b0 ;
  assign y3799 = n8828 ;
  assign y3800 = n8831 ;
  assign y3801 = ~1'b0 ;
  assign y3802 = ~1'b0 ;
  assign y3803 = n8841 ;
  assign y3804 = n8842 ;
  assign y3805 = ~n8845 ;
  assign y3806 = n7872 ;
  assign y3807 = ~n6742 ;
  assign y3808 = ~1'b0 ;
  assign y3809 = ~1'b0 ;
  assign y3810 = n8847 ;
  assign y3811 = n8849 ;
  assign y3812 = ~n8852 ;
  assign y3813 = ~1'b0 ;
  assign y3814 = ~n8857 ;
  assign y3815 = ~n8867 ;
  assign y3816 = n8869 ;
  assign y3817 = n4084 ;
  assign y3818 = ~n8873 ;
  assign y3819 = n8874 ;
  assign y3820 = ~1'b0 ;
  assign y3821 = ~n196 ;
  assign y3822 = ~n5036 ;
  assign y3823 = ~n8878 ;
  assign y3824 = n8880 ;
  assign y3825 = n8884 ;
  assign y3826 = ~1'b0 ;
  assign y3827 = ~n8886 ;
  assign y3828 = n4981 ;
  assign y3829 = ~n8890 ;
  assign y3830 = n8894 ;
  assign y3831 = ~n5723 ;
  assign y3832 = n8896 ;
  assign y3833 = ~1'b0 ;
  assign y3834 = ~n8902 ;
  assign y3835 = n8909 ;
  assign y3836 = n8913 ;
  assign y3837 = ~n8922 ;
  assign y3838 = ~n8928 ;
  assign y3839 = ~1'b0 ;
  assign y3840 = ~n8936 ;
  assign y3841 = n8937 ;
  assign y3842 = n8940 ;
  assign y3843 = ~n8944 ;
  assign y3844 = n8945 ;
  assign y3845 = ~n8952 ;
  assign y3846 = ~n8955 ;
  assign y3847 = ~n8957 ;
  assign y3848 = ~n8958 ;
  assign y3849 = ~n8959 ;
  assign y3850 = n8963 ;
  assign y3851 = ~n8967 ;
  assign y3852 = ~n8969 ;
  assign y3853 = n8971 ;
  assign y3854 = n8972 ;
  assign y3855 = ~n8980 ;
  assign y3856 = ~1'b0 ;
  assign y3857 = ~1'b0 ;
  assign y3858 = n8989 ;
  assign y3859 = ~1'b0 ;
  assign y3860 = ~n8993 ;
  assign y3861 = ~n8998 ;
  assign y3862 = ~n8999 ;
  assign y3863 = n9003 ;
  assign y3864 = n9005 ;
  assign y3865 = ~1'b0 ;
  assign y3866 = n9015 ;
  assign y3867 = n9022 ;
  assign y3868 = n9024 ;
  assign y3869 = n2850 ;
  assign y3870 = n9033 ;
  assign y3871 = ~n9035 ;
  assign y3872 = ~n9048 ;
  assign y3873 = n9054 ;
  assign y3874 = n9055 ;
  assign y3875 = ~n9061 ;
  assign y3876 = n9062 ;
  assign y3877 = n9064 ;
  assign y3878 = ~n9066 ;
  assign y3879 = n9071 ;
  assign y3880 = ~n9075 ;
  assign y3881 = n9077 ;
  assign y3882 = 1'b0 ;
  assign y3883 = ~n9079 ;
  assign y3884 = n9083 ;
  assign y3885 = n9088 ;
  assign y3886 = ~1'b0 ;
  assign y3887 = ~n9096 ;
  assign y3888 = ~n8081 ;
  assign y3889 = ~n9129 ;
  assign y3890 = ~n9130 ;
  assign y3891 = ~n9131 ;
  assign y3892 = n9135 ;
  assign y3893 = ~1'b0 ;
  assign y3894 = ~n9138 ;
  assign y3895 = 1'b0 ;
  assign y3896 = n9140 ;
  assign y3897 = ~1'b0 ;
  assign y3898 = n9143 ;
  assign y3899 = n9150 ;
  assign y3900 = ~1'b0 ;
  assign y3901 = n9152 ;
  assign y3902 = ~1'b0 ;
  assign y3903 = 1'b0 ;
  assign y3904 = ~n9156 ;
  assign y3905 = ~n9163 ;
  assign y3906 = ~n9166 ;
  assign y3907 = ~1'b0 ;
  assign y3908 = ~n9172 ;
  assign y3909 = n9177 ;
  assign y3910 = n9179 ;
  assign y3911 = ~1'b0 ;
  assign y3912 = ~1'b0 ;
  assign y3913 = ~1'b0 ;
  assign y3914 = ~n9186 ;
  assign y3915 = n9187 ;
  assign y3916 = n9193 ;
  assign y3917 = n9194 ;
  assign y3918 = ~n9196 ;
  assign y3919 = n9197 ;
  assign y3920 = n9201 ;
  assign y3921 = ~n9206 ;
  assign y3922 = ~n9208 ;
  assign y3923 = ~n9211 ;
  assign y3924 = ~1'b0 ;
  assign y3925 = ~n2049 ;
  assign y3926 = n9215 ;
  assign y3927 = n9218 ;
  assign y3928 = ~1'b0 ;
  assign y3929 = ~1'b0 ;
  assign y3930 = ~n2847 ;
  assign y3931 = ~1'b0 ;
  assign y3932 = n9220 ;
  assign y3933 = ~n9226 ;
  assign y3934 = ~n9227 ;
  assign y3935 = ~1'b0 ;
  assign y3936 = ~n9228 ;
  assign y3937 = ~n9229 ;
  assign y3938 = n9236 ;
  assign y3939 = n3497 ;
  assign y3940 = n9237 ;
  assign y3941 = ~n9240 ;
  assign y3942 = n9245 ;
  assign y3943 = ~1'b0 ;
  assign y3944 = n9249 ;
  assign y3945 = n9253 ;
  assign y3946 = ~1'b0 ;
  assign y3947 = n9257 ;
  assign y3948 = n9258 ;
  assign y3949 = n9260 ;
  assign y3950 = ~n9262 ;
  assign y3951 = ~n9263 ;
  assign y3952 = ~1'b0 ;
  assign y3953 = n9267 ;
  assign y3954 = n4562 ;
  assign y3955 = ~n9271 ;
  assign y3956 = n9274 ;
  assign y3957 = ~n9280 ;
  assign y3958 = ~n9284 ;
  assign y3959 = n9287 ;
  assign y3960 = ~n9291 ;
  assign y3961 = ~1'b0 ;
  assign y3962 = ~n9296 ;
  assign y3963 = ~n9299 ;
  assign y3964 = n9300 ;
  assign y3965 = ~n9305 ;
  assign y3966 = ~n9308 ;
  assign y3967 = ~1'b0 ;
  assign y3968 = ~1'b0 ;
  assign y3969 = ~n9312 ;
  assign y3970 = ~1'b0 ;
  assign y3971 = n9314 ;
  assign y3972 = ~n9315 ;
  assign y3973 = ~n9317 ;
  assign y3974 = ~n9318 ;
  assign y3975 = n7558 ;
  assign y3976 = ~1'b0 ;
  assign y3977 = n9322 ;
  assign y3978 = ~n9325 ;
  assign y3979 = ~n9334 ;
  assign y3980 = ~1'b0 ;
  assign y3981 = n9335 ;
  assign y3982 = ~n9337 ;
  assign y3983 = n9344 ;
  assign y3984 = n9346 ;
  assign y3985 = ~n9352 ;
  assign y3986 = n9357 ;
  assign y3987 = ~n9362 ;
  assign y3988 = ~1'b0 ;
  assign y3989 = n9363 ;
  assign y3990 = ~n9368 ;
  assign y3991 = n9371 ;
  assign y3992 = n1649 ;
  assign y3993 = n9375 ;
  assign y3994 = ~n9379 ;
  assign y3995 = ~n9384 ;
  assign y3996 = n9385 ;
  assign y3997 = ~1'b0 ;
  assign y3998 = ~n9387 ;
  assign y3999 = ~n9390 ;
  assign y4000 = ~n9393 ;
  assign y4001 = n9395 ;
  assign y4002 = n9399 ;
  assign y4003 = ~1'b0 ;
  assign y4004 = ~n9405 ;
  assign y4005 = ~n9407 ;
  assign y4006 = ~1'b0 ;
  assign y4007 = ~n9411 ;
  assign y4008 = n9415 ;
  assign y4009 = 1'b0 ;
  assign y4010 = n9420 ;
  assign y4011 = ~n9422 ;
  assign y4012 = ~n9424 ;
  assign y4013 = ~n9427 ;
  assign y4014 = ~n9428 ;
  assign y4015 = n9430 ;
  assign y4016 = ~1'b0 ;
  assign y4017 = ~1'b0 ;
  assign y4018 = n9431 ;
  assign y4019 = ~n9434 ;
  assign y4020 = n9441 ;
  assign y4021 = ~1'b0 ;
  assign y4022 = ~n9444 ;
  assign y4023 = ~n3979 ;
  assign y4024 = ~1'b0 ;
  assign y4025 = ~n9448 ;
  assign y4026 = ~1'b0 ;
  assign y4027 = ~1'b0 ;
  assign y4028 = ~1'b0 ;
  assign y4029 = n9449 ;
  assign y4030 = ~1'b0 ;
  assign y4031 = n9460 ;
  assign y4032 = ~n9463 ;
  assign y4033 = n1347 ;
  assign y4034 = ~1'b0 ;
  assign y4035 = ~n9467 ;
  assign y4036 = n9472 ;
  assign y4037 = ~1'b0 ;
  assign y4038 = ~1'b0 ;
  assign y4039 = ~n9475 ;
  assign y4040 = ~n9478 ;
  assign y4041 = n9483 ;
  assign y4042 = ~n5724 ;
  assign y4043 = ~1'b0 ;
  assign y4044 = ~1'b0 ;
  assign y4045 = n9487 ;
  assign y4046 = ~n9491 ;
  assign y4047 = ~1'b0 ;
  assign y4048 = n9492 ;
  assign y4049 = ~1'b0 ;
  assign y4050 = ~1'b0 ;
  assign y4051 = ~n9493 ;
  assign y4052 = ~n9495 ;
  assign y4053 = n9497 ;
  assign y4054 = ~n9499 ;
  assign y4055 = ~n9501 ;
  assign y4056 = n9502 ;
  assign y4057 = n9503 ;
  assign y4058 = ~n9505 ;
  assign y4059 = ~n9509 ;
  assign y4060 = ~1'b0 ;
  assign y4061 = ~n9514 ;
  assign y4062 = ~n9516 ;
  assign y4063 = ~n5662 ;
  assign y4064 = ~1'b0 ;
  assign y4065 = ~n9518 ;
  assign y4066 = ~n9520 ;
  assign y4067 = ~n9521 ;
  assign y4068 = ~n2182 ;
  assign y4069 = ~1'b0 ;
  assign y4070 = ~1'b0 ;
  assign y4071 = ~n9529 ;
  assign y4072 = ~n9530 ;
  assign y4073 = n9156 ;
  assign y4074 = ~n9534 ;
  assign y4075 = n9535 ;
  assign y4076 = ~n9536 ;
  assign y4077 = ~1'b0 ;
  assign y4078 = ~n9538 ;
  assign y4079 = ~n9541 ;
  assign y4080 = n9542 ;
  assign y4081 = 1'b0 ;
  assign y4082 = n4116 ;
  assign y4083 = ~1'b0 ;
  assign y4084 = ~1'b0 ;
  assign y4085 = ~1'b0 ;
  assign y4086 = ~n9544 ;
  assign y4087 = n9546 ;
  assign y4088 = n9549 ;
  assign y4089 = n9551 ;
  assign y4090 = ~n9552 ;
  assign y4091 = ~n9555 ;
  assign y4092 = ~n9557 ;
  assign y4093 = n9560 ;
  assign y4094 = ~1'b0 ;
  assign y4095 = n9564 ;
  assign y4096 = ~n9565 ;
  assign y4097 = ~n9566 ;
  assign y4098 = ~n9567 ;
  assign y4099 = ~1'b0 ;
  assign y4100 = ~n9569 ;
  assign y4101 = n9570 ;
  assign y4102 = ~n9572 ;
  assign y4103 = n9573 ;
  assign y4104 = n5267 ;
  assign y4105 = ~n9582 ;
  assign y4106 = n9586 ;
  assign y4107 = n9589 ;
  assign y4108 = ~n9592 ;
  assign y4109 = n9595 ;
  assign y4110 = n9598 ;
  assign y4111 = n9603 ;
  assign y4112 = n9604 ;
  assign y4113 = ~n9606 ;
  assign y4114 = ~n9608 ;
  assign y4115 = ~n9611 ;
  assign y4116 = ~n9612 ;
  assign y4117 = ~n9613 ;
  assign y4118 = ~1'b0 ;
  assign y4119 = ~n9615 ;
  assign y4120 = ~n9616 ;
  assign y4121 = n9619 ;
  assign y4122 = ~n9623 ;
  assign y4123 = n9624 ;
  assign y4124 = n9628 ;
  assign y4125 = n9634 ;
  assign y4126 = ~1'b0 ;
  assign y4127 = ~n9635 ;
  assign y4128 = ~n9642 ;
  assign y4129 = ~n9648 ;
  assign y4130 = ~n9651 ;
  assign y4131 = n9658 ;
  assign y4132 = ~n9661 ;
  assign y4133 = ~1'b0 ;
  assign y4134 = ~1'b0 ;
  assign y4135 = ~1'b0 ;
  assign y4136 = ~n7076 ;
  assign y4137 = n9662 ;
  assign y4138 = ~n9666 ;
  assign y4139 = n9669 ;
  assign y4140 = n9676 ;
  assign y4141 = n9679 ;
  assign y4142 = 1'b0 ;
  assign y4143 = n9681 ;
  assign y4144 = ~1'b0 ;
  assign y4145 = ~n9682 ;
  assign y4146 = ~1'b0 ;
  assign y4147 = ~n9691 ;
  assign y4148 = ~n9692 ;
  assign y4149 = ~n9693 ;
  assign y4150 = ~n9696 ;
  assign y4151 = ~1'b0 ;
  assign y4152 = 1'b0 ;
  assign y4153 = ~n9700 ;
  assign y4154 = ~n9704 ;
  assign y4155 = ~n9706 ;
  assign y4156 = ~n9707 ;
  assign y4157 = n9710 ;
  assign y4158 = n9711 ;
  assign y4159 = ~n9713 ;
  assign y4160 = 1'b0 ;
  assign y4161 = ~n9714 ;
  assign y4162 = ~n9715 ;
  assign y4163 = n9720 ;
  assign y4164 = ~n9728 ;
  assign y4165 = n9730 ;
  assign y4166 = 1'b0 ;
  assign y4167 = ~n9731 ;
  assign y4168 = n9735 ;
  assign y4169 = n9736 ;
  assign y4170 = ~n9739 ;
  assign y4171 = ~n9741 ;
  assign y4172 = ~1'b0 ;
  assign y4173 = ~n9744 ;
  assign y4174 = ~1'b0 ;
  assign y4175 = n9748 ;
  assign y4176 = ~1'b0 ;
  assign y4177 = n9749 ;
  assign y4178 = ~1'b0 ;
  assign y4179 = ~1'b0 ;
  assign y4180 = ~n9752 ;
  assign y4181 = ~n9759 ;
  assign y4182 = ~1'b0 ;
  assign y4183 = ~n9763 ;
  assign y4184 = n9764 ;
  assign y4185 = n4897 ;
  assign y4186 = ~1'b0 ;
  assign y4187 = n9765 ;
  assign y4188 = ~n9775 ;
  assign y4189 = ~n9776 ;
  assign y4190 = ~1'b0 ;
  assign y4191 = ~1'b0 ;
  assign y4192 = ~n9779 ;
  assign y4193 = ~1'b0 ;
  assign y4194 = ~1'b0 ;
  assign y4195 = ~n9781 ;
  assign y4196 = ~n9783 ;
  assign y4197 = ~1'b0 ;
  assign y4198 = n9785 ;
  assign y4199 = ~n6067 ;
  assign y4200 = ~1'b0 ;
  assign y4201 = n9788 ;
  assign y4202 = ~n9791 ;
  assign y4203 = ~1'b0 ;
  assign y4204 = ~n9793 ;
  assign y4205 = ~1'b0 ;
  assign y4206 = n9796 ;
  assign y4207 = ~1'b0 ;
  assign y4208 = ~1'b0 ;
  assign y4209 = ~n9797 ;
  assign y4210 = ~1'b0 ;
  assign y4211 = ~1'b0 ;
  assign y4212 = ~1'b0 ;
  assign y4213 = ~n9802 ;
  assign y4214 = ~1'b0 ;
  assign y4215 = ~1'b0 ;
  assign y4216 = ~n9805 ;
  assign y4217 = ~n9807 ;
  assign y4218 = ~n9809 ;
  assign y4219 = ~1'b0 ;
  assign y4220 = ~n9813 ;
  assign y4221 = ~n9814 ;
  assign y4222 = ~n9817 ;
  assign y4223 = n9818 ;
  assign y4224 = ~1'b0 ;
  assign y4225 = ~1'b0 ;
  assign y4226 = ~n9827 ;
  assign y4227 = ~n9834 ;
  assign y4228 = ~1'b0 ;
  assign y4229 = ~n9836 ;
  assign y4230 = n9838 ;
  assign y4231 = n9843 ;
  assign y4232 = n9858 ;
  assign y4233 = ~n4315 ;
  assign y4234 = ~n9859 ;
  assign y4235 = n9865 ;
  assign y4236 = ~n9867 ;
  assign y4237 = ~n9870 ;
  assign y4238 = ~n9873 ;
  assign y4239 = ~1'b0 ;
  assign y4240 = n9881 ;
  assign y4241 = n9883 ;
  assign y4242 = n9885 ;
  assign y4243 = n9888 ;
  assign y4244 = n9892 ;
  assign y4245 = ~1'b0 ;
  assign y4246 = ~n9896 ;
  assign y4247 = ~n9897 ;
  assign y4248 = ~n9898 ;
  assign y4249 = ~n9901 ;
  assign y4250 = n9902 ;
  assign y4251 = n9903 ;
  assign y4252 = ~n9906 ;
  assign y4253 = ~n9912 ;
  assign y4254 = ~1'b0 ;
  assign y4255 = n9914 ;
  assign y4256 = n8311 ;
  assign y4257 = n9915 ;
  assign y4258 = ~1'b0 ;
  assign y4259 = ~n9918 ;
  assign y4260 = n9922 ;
  assign y4261 = ~1'b0 ;
  assign y4262 = ~1'b0 ;
  assign y4263 = ~n9937 ;
  assign y4264 = n9942 ;
  assign y4265 = ~1'b0 ;
  assign y4266 = ~n9943 ;
  assign y4267 = ~1'b0 ;
  assign y4268 = n9946 ;
  assign y4269 = n9948 ;
  assign y4270 = n9954 ;
  assign y4271 = ~1'b0 ;
  assign y4272 = ~1'b0 ;
  assign y4273 = ~1'b0 ;
  assign y4274 = n9958 ;
  assign y4275 = n9968 ;
  assign y4276 = n9969 ;
  assign y4277 = ~n9974 ;
  assign y4278 = ~n9982 ;
  assign y4279 = n9983 ;
  assign y4280 = n9986 ;
  assign y4281 = ~n9991 ;
  assign y4282 = ~n9992 ;
  assign y4283 = n9995 ;
  assign y4284 = ~1'b0 ;
  assign y4285 = n10002 ;
  assign y4286 = ~1'b0 ;
  assign y4287 = ~n10003 ;
  assign y4288 = ~1'b0 ;
  assign y4289 = 1'b0 ;
  assign y4290 = n10005 ;
  assign y4291 = n10006 ;
  assign y4292 = n10011 ;
  assign y4293 = ~1'b0 ;
  assign y4294 = ~n10013 ;
  assign y4295 = ~n10015 ;
  assign y4296 = ~1'b0 ;
  assign y4297 = n10016 ;
  assign y4298 = ~1'b0 ;
  assign y4299 = ~n10020 ;
  assign y4300 = ~n10022 ;
  assign y4301 = ~1'b0 ;
  assign y4302 = n10023 ;
  assign y4303 = n10033 ;
  assign y4304 = ~1'b0 ;
  assign y4305 = n10034 ;
  assign y4306 = n10036 ;
  assign y4307 = n10039 ;
  assign y4308 = ~1'b0 ;
  assign y4309 = ~n10040 ;
  assign y4310 = ~n10046 ;
  assign y4311 = ~1'b0 ;
  assign y4312 = n10050 ;
  assign y4313 = ~n10055 ;
  assign y4314 = ~n10059 ;
  assign y4315 = n10062 ;
  assign y4316 = n10064 ;
  assign y4317 = n10067 ;
  assign y4318 = ~n10069 ;
  assign y4319 = ~n10072 ;
  assign y4320 = n10074 ;
  assign y4321 = ~n10076 ;
  assign y4322 = ~n10077 ;
  assign y4323 = ~n10078 ;
  assign y4324 = 1'b0 ;
  assign y4325 = ~1'b0 ;
  assign y4326 = ~1'b0 ;
  assign y4327 = ~n10080 ;
  assign y4328 = ~n7567 ;
  assign y4329 = n10082 ;
  assign y4330 = ~n10087 ;
  assign y4331 = n10088 ;
  assign y4332 = n10092 ;
  assign y4333 = n10100 ;
  assign y4334 = ~1'b0 ;
  assign y4335 = ~n2143 ;
  assign y4336 = ~1'b0 ;
  assign y4337 = ~1'b0 ;
  assign y4338 = ~n10101 ;
  assign y4339 = n10108 ;
  assign y4340 = ~n10110 ;
  assign y4341 = ~1'b0 ;
  assign y4342 = ~n10114 ;
  assign y4343 = ~n10120 ;
  assign y4344 = n10123 ;
  assign y4345 = ~1'b0 ;
  assign y4346 = n10125 ;
  assign y4347 = ~n10127 ;
  assign y4348 = ~1'b0 ;
  assign y4349 = ~n10129 ;
  assign y4350 = ~n10131 ;
  assign y4351 = ~1'b0 ;
  assign y4352 = n10132 ;
  assign y4353 = ~n10137 ;
  assign y4354 = n10139 ;
  assign y4355 = n10142 ;
  assign y4356 = ~n10145 ;
  assign y4357 = ~n10148 ;
  assign y4358 = n10152 ;
  assign y4359 = n10154 ;
  assign y4360 = ~n10162 ;
  assign y4361 = ~1'b0 ;
  assign y4362 = ~1'b0 ;
  assign y4363 = ~n10164 ;
  assign y4364 = ~1'b0 ;
  assign y4365 = 1'b0 ;
  assign y4366 = n10166 ;
  assign y4367 = ~1'b0 ;
  assign y4368 = n10168 ;
  assign y4369 = n10172 ;
  assign y4370 = n10176 ;
  assign y4371 = n10178 ;
  assign y4372 = ~n10179 ;
  assign y4373 = n10180 ;
  assign y4374 = n10184 ;
  assign y4375 = ~n10192 ;
  assign y4376 = n10196 ;
  assign y4377 = n10199 ;
  assign y4378 = 1'b0 ;
  assign y4379 = n10204 ;
  assign y4380 = n7240 ;
  assign y4381 = n10205 ;
  assign y4382 = ~1'b0 ;
  assign y4383 = ~n10206 ;
  assign y4384 = ~n10209 ;
  assign y4385 = n10212 ;
  assign y4386 = ~n10214 ;
  assign y4387 = ~n10215 ;
  assign y4388 = ~n10217 ;
  assign y4389 = ~n10218 ;
  assign y4390 = n10223 ;
  assign y4391 = n10225 ;
  assign y4392 = n10231 ;
  assign y4393 = ~n10232 ;
  assign y4394 = ~1'b0 ;
  assign y4395 = n10234 ;
  assign y4396 = ~n10236 ;
  assign y4397 = ~n10239 ;
  assign y4398 = ~n10240 ;
  assign y4399 = ~n10242 ;
  assign y4400 = ~1'b0 ;
  assign y4401 = ~n10245 ;
  assign y4402 = n10250 ;
  assign y4403 = n10253 ;
  assign y4404 = ~n10255 ;
  assign y4405 = 1'b0 ;
  assign y4406 = ~n7850 ;
  assign y4407 = ~n10261 ;
  assign y4408 = ~1'b0 ;
  assign y4409 = ~1'b0 ;
  assign y4410 = ~n10263 ;
  assign y4411 = ~n10267 ;
  assign y4412 = ~1'b0 ;
  assign y4413 = ~n10268 ;
  assign y4414 = ~n10270 ;
  assign y4415 = n10271 ;
  assign y4416 = ~1'b0 ;
  assign y4417 = n10275 ;
  assign y4418 = ~n10286 ;
  assign y4419 = ~1'b0 ;
  assign y4420 = ~n10289 ;
  assign y4421 = ~n10294 ;
  assign y4422 = n10297 ;
  assign y4423 = n10301 ;
  assign y4424 = n10308 ;
  assign y4425 = ~1'b0 ;
  assign y4426 = ~n10309 ;
  assign y4427 = ~1'b0 ;
  assign y4428 = ~1'b0 ;
  assign y4429 = n10311 ;
  assign y4430 = n10313 ;
  assign y4431 = n10320 ;
  assign y4432 = ~1'b0 ;
  assign y4433 = ~n10321 ;
  assign y4434 = ~n399 ;
  assign y4435 = ~1'b0 ;
  assign y4436 = ~1'b0 ;
  assign y4437 = ~n362 ;
  assign y4438 = n10323 ;
  assign y4439 = ~1'b0 ;
  assign y4440 = ~1'b0 ;
  assign y4441 = n10325 ;
  assign y4442 = n10326 ;
  assign y4443 = n10327 ;
  assign y4444 = ~1'b0 ;
  assign y4445 = ~n10330 ;
  assign y4446 = ~1'b0 ;
  assign y4447 = n10336 ;
  assign y4448 = ~n10337 ;
  assign y4449 = ~n1973 ;
  assign y4450 = n10341 ;
  assign y4451 = ~1'b0 ;
  assign y4452 = ~n10343 ;
  assign y4453 = n10350 ;
  assign y4454 = ~n10352 ;
  assign y4455 = ~n10361 ;
  assign y4456 = ~n10366 ;
  assign y4457 = ~1'b0 ;
  assign y4458 = ~1'b0 ;
  assign y4459 = ~n10372 ;
  assign y4460 = n10126 ;
  assign y4461 = ~1'b0 ;
  assign y4462 = ~1'b0 ;
  assign y4463 = n10373 ;
  assign y4464 = ~1'b0 ;
  assign y4465 = ~n10376 ;
  assign y4466 = ~n10379 ;
  assign y4467 = ~1'b0 ;
  assign y4468 = ~1'b0 ;
  assign y4469 = ~n10383 ;
  assign y4470 = ~1'b0 ;
  assign y4471 = n10385 ;
  assign y4472 = n10388 ;
  assign y4473 = n10389 ;
  assign y4474 = ~n10390 ;
  assign y4475 = n1813 ;
  assign y4476 = ~1'b0 ;
  assign y4477 = ~n10392 ;
  assign y4478 = ~n10393 ;
  assign y4479 = ~1'b0 ;
  assign y4480 = n10394 ;
  assign y4481 = ~n10400 ;
  assign y4482 = ~1'b0 ;
  assign y4483 = n10401 ;
  assign y4484 = 1'b0 ;
  assign y4485 = ~n10402 ;
  assign y4486 = ~n10404 ;
  assign y4487 = n10413 ;
  assign y4488 = ~n10414 ;
  assign y4489 = n10415 ;
  assign y4490 = ~n10416 ;
  assign y4491 = n10419 ;
  assign y4492 = ~n10420 ;
  assign y4493 = n10421 ;
  assign y4494 = n10432 ;
  assign y4495 = ~n10435 ;
  assign y4496 = n10436 ;
  assign y4497 = n10440 ;
  assign y4498 = ~1'b0 ;
  assign y4499 = ~1'b0 ;
  assign y4500 = n10444 ;
  assign y4501 = n10449 ;
  assign y4502 = ~1'b0 ;
  assign y4503 = n10451 ;
  assign y4504 = n10453 ;
  assign y4505 = n10455 ;
  assign y4506 = ~n10459 ;
  assign y4507 = ~n10463 ;
  assign y4508 = ~n10464 ;
  assign y4509 = ~n10467 ;
  assign y4510 = ~n4294 ;
  assign y4511 = ~n10468 ;
  assign y4512 = n10470 ;
  assign y4513 = ~n10475 ;
  assign y4514 = ~1'b0 ;
  assign y4515 = n10479 ;
  assign y4516 = ~n10483 ;
  assign y4517 = n10486 ;
  assign y4518 = n10487 ;
  assign y4519 = ~1'b0 ;
  assign y4520 = n10488 ;
  assign y4521 = n10490 ;
  assign y4522 = ~n10493 ;
  assign y4523 = ~n10497 ;
  assign y4524 = ~n10501 ;
  assign y4525 = ~n4559 ;
  assign y4526 = n10502 ;
  assign y4527 = ~1'b0 ;
  assign y4528 = ~n10506 ;
  assign y4529 = n10507 ;
  assign y4530 = n10508 ;
  assign y4531 = ~1'b0 ;
  assign y4532 = ~1'b0 ;
  assign y4533 = n10509 ;
  assign y4534 = ~n10511 ;
  assign y4535 = ~n10515 ;
  assign y4536 = ~1'b0 ;
  assign y4537 = n9323 ;
  assign y4538 = n10519 ;
  assign y4539 = ~n10521 ;
  assign y4540 = n10523 ;
  assign y4541 = ~n10524 ;
  assign y4542 = n10531 ;
  assign y4543 = ~n10533 ;
  assign y4544 = ~n4664 ;
  assign y4545 = ~1'b0 ;
  assign y4546 = n10535 ;
  assign y4547 = ~n10537 ;
  assign y4548 = ~n10538 ;
  assign y4549 = n673 ;
  assign y4550 = ~n10540 ;
  assign y4551 = ~1'b0 ;
  assign y4552 = n10544 ;
  assign y4553 = n10546 ;
  assign y4554 = n10551 ;
  assign y4555 = n4927 ;
  assign y4556 = ~n10553 ;
  assign y4557 = ~1'b0 ;
  assign y4558 = n10555 ;
  assign y4559 = n10558 ;
  assign y4560 = n10560 ;
  assign y4561 = ~n10564 ;
  assign y4562 = n10565 ;
  assign y4563 = n10566 ;
  assign y4564 = n10574 ;
  assign y4565 = n10577 ;
  assign y4566 = ~n9138 ;
  assign y4567 = ~n10579 ;
  assign y4568 = ~n10582 ;
  assign y4569 = ~n10584 ;
  assign y4570 = ~1'b0 ;
  assign y4571 = ~n10590 ;
  assign y4572 = ~1'b0 ;
  assign y4573 = ~n10592 ;
  assign y4574 = ~1'b0 ;
  assign y4575 = n10593 ;
  assign y4576 = n10595 ;
  assign y4577 = n10600 ;
  assign y4578 = n10602 ;
  assign y4579 = n10605 ;
  assign y4580 = ~n10611 ;
  assign y4581 = ~n6457 ;
  assign y4582 = n10615 ;
  assign y4583 = ~n10618 ;
  assign y4584 = ~n10621 ;
  assign y4585 = ~n10622 ;
  assign y4586 = n10623 ;
  assign y4587 = n10624 ;
  assign y4588 = n10627 ;
  assign y4589 = ~1'b0 ;
  assign y4590 = ~1'b0 ;
  assign y4591 = ~1'b0 ;
  assign y4592 = n10628 ;
  assign y4593 = ~1'b0 ;
  assign y4594 = ~n10631 ;
  assign y4595 = n10638 ;
  assign y4596 = ~n10642 ;
  assign y4597 = n10643 ;
  assign y4598 = ~n10644 ;
  assign y4599 = ~n305 ;
  assign y4600 = n10645 ;
  assign y4601 = n10650 ;
  assign y4602 = n10653 ;
  assign y4603 = n8038 ;
  assign y4604 = ~1'b0 ;
  assign y4605 = ~1'b0 ;
  assign y4606 = ~1'b0 ;
  assign y4607 = n10657 ;
  assign y4608 = ~n10658 ;
  assign y4609 = ~1'b0 ;
  assign y4610 = n10660 ;
  assign y4611 = ~1'b0 ;
  assign y4612 = ~1'b0 ;
  assign y4613 = n1758 ;
  assign y4614 = n10666 ;
  assign y4615 = 1'b0 ;
  assign y4616 = ~n10670 ;
  assign y4617 = ~n10672 ;
  assign y4618 = ~1'b0 ;
  assign y4619 = n10679 ;
  assign y4620 = ~n10681 ;
  assign y4621 = ~1'b0 ;
  assign y4622 = ~n10688 ;
  assign y4623 = ~1'b0 ;
  assign y4624 = ~n10689 ;
  assign y4625 = ~1'b0 ;
  assign y4626 = n10691 ;
  assign y4627 = ~n10695 ;
  assign y4628 = ~n10698 ;
  assign y4629 = ~1'b0 ;
  assign y4630 = ~1'b0 ;
  assign y4631 = n10700 ;
  assign y4632 = ~n10702 ;
  assign y4633 = n10703 ;
  assign y4634 = ~n10705 ;
  assign y4635 = n10712 ;
  assign y4636 = n10714 ;
  assign y4637 = n10718 ;
  assign y4638 = ~1'b0 ;
  assign y4639 = ~n10721 ;
  assign y4640 = ~n10722 ;
  assign y4641 = ~n10724 ;
  assign y4642 = ~1'b0 ;
  assign y4643 = ~n10730 ;
  assign y4644 = ~n10731 ;
  assign y4645 = n10736 ;
  assign y4646 = ~n10737 ;
  assign y4647 = 1'b0 ;
  assign y4648 = n1183 ;
  assign y4649 = n10740 ;
  assign y4650 = n10746 ;
  assign y4651 = ~n10754 ;
  assign y4652 = ~1'b0 ;
  assign y4653 = ~n10756 ;
  assign y4654 = ~n10757 ;
  assign y4655 = ~1'b0 ;
  assign y4656 = n10761 ;
  assign y4657 = ~n10763 ;
  assign y4658 = ~n10766 ;
  assign y4659 = n10779 ;
  assign y4660 = ~n10780 ;
  assign y4661 = n10784 ;
  assign y4662 = n10788 ;
  assign y4663 = ~1'b0 ;
  assign y4664 = n10789 ;
  assign y4665 = ~n10793 ;
  assign y4666 = n10796 ;
  assign y4667 = ~n8403 ;
  assign y4668 = ~n10799 ;
  assign y4669 = 1'b0 ;
  assign y4670 = n10804 ;
  assign y4671 = ~n10806 ;
  assign y4672 = ~1'b0 ;
  assign y4673 = ~1'b0 ;
  assign y4674 = ~n10810 ;
  assign y4675 = ~1'b0 ;
  assign y4676 = n10812 ;
  assign y4677 = ~n10815 ;
  assign y4678 = ~n10820 ;
  assign y4679 = 1'b0 ;
  assign y4680 = n10821 ;
  assign y4681 = ~1'b0 ;
  assign y4682 = ~n10822 ;
  assign y4683 = ~n10823 ;
  assign y4684 = ~1'b0 ;
  assign y4685 = n10825 ;
  assign y4686 = ~n10831 ;
  assign y4687 = ~1'b0 ;
  assign y4688 = ~n10832 ;
  assign y4689 = n10842 ;
  assign y4690 = ~n10845 ;
  assign y4691 = ~1'b0 ;
  assign y4692 = n10851 ;
  assign y4693 = ~1'b0 ;
  assign y4694 = ~n10854 ;
  assign y4695 = ~n10855 ;
  assign y4696 = ~1'b0 ;
  assign y4697 = ~n10856 ;
  assign y4698 = ~n10865 ;
  assign y4699 = ~n10867 ;
  assign y4700 = n10869 ;
  assign y4701 = ~1'b0 ;
  assign y4702 = n10870 ;
  assign y4703 = n10871 ;
  assign y4704 = n10874 ;
  assign y4705 = ~1'b0 ;
  assign y4706 = ~n10877 ;
  assign y4707 = n9090 ;
  assign y4708 = n10889 ;
  assign y4709 = ~n10891 ;
  assign y4710 = n10893 ;
  assign y4711 = n10896 ;
  assign y4712 = n10897 ;
  assign y4713 = ~n10898 ;
  assign y4714 = ~1'b0 ;
  assign y4715 = ~n10900 ;
  assign y4716 = ~n10903 ;
  assign y4717 = n10907 ;
  assign y4718 = ~1'b0 ;
  assign y4719 = ~1'b0 ;
  assign y4720 = x3 ;
  assign y4721 = ~n10908 ;
  assign y4722 = ~1'b0 ;
  assign y4723 = n8605 ;
  assign y4724 = ~n10912 ;
  assign y4725 = n10923 ;
  assign y4726 = ~1'b0 ;
  assign y4727 = ~n10924 ;
  assign y4728 = n10925 ;
  assign y4729 = ~n10930 ;
  assign y4730 = n10931 ;
  assign y4731 = n10933 ;
  assign y4732 = ~1'b0 ;
  assign y4733 = n10934 ;
  assign y4734 = n10938 ;
  assign y4735 = n10943 ;
  assign y4736 = n10944 ;
  assign y4737 = ~n10946 ;
  assign y4738 = ~1'b0 ;
  assign y4739 = n10947 ;
  assign y4740 = n10948 ;
  assign y4741 = n10953 ;
  assign y4742 = n9657 ;
  assign y4743 = n10957 ;
  assign y4744 = n10959 ;
  assign y4745 = ~n10964 ;
  assign y4746 = ~n10968 ;
  assign y4747 = ~n10969 ;
  assign y4748 = n10971 ;
  assign y4749 = ~n10974 ;
  assign y4750 = ~1'b0 ;
  assign y4751 = n10988 ;
  assign y4752 = n10993 ;
  assign y4753 = n10994 ;
  assign y4754 = ~n10995 ;
  assign y4755 = ~n10999 ;
  assign y4756 = n11000 ;
  assign y4757 = ~n11001 ;
  assign y4758 = n11003 ;
  assign y4759 = n11012 ;
  assign y4760 = n193 ;
  assign y4761 = n11014 ;
  assign y4762 = ~1'b0 ;
  assign y4763 = ~n11021 ;
  assign y4764 = ~1'b0 ;
  assign y4765 = n11022 ;
  assign y4766 = ~n11028 ;
  assign y4767 = ~n11029 ;
  assign y4768 = ~n11031 ;
  assign y4769 = ~n11032 ;
  assign y4770 = ~n11033 ;
  assign y4771 = ~n11034 ;
  assign y4772 = ~1'b0 ;
  assign y4773 = ~1'b0 ;
  assign y4774 = n11035 ;
  assign y4775 = ~1'b0 ;
  assign y4776 = ~n11036 ;
  assign y4777 = ~1'b0 ;
  assign y4778 = ~n11037 ;
  assign y4779 = n11038 ;
  assign y4780 = ~n11040 ;
  assign y4781 = ~1'b0 ;
  assign y4782 = n11050 ;
  assign y4783 = ~n11051 ;
  assign y4784 = n11059 ;
  assign y4785 = ~n11064 ;
  assign y4786 = n11070 ;
  assign y4787 = n11073 ;
  assign y4788 = ~n11076 ;
  assign y4789 = n11078 ;
  assign y4790 = ~1'b0 ;
  assign y4791 = n11081 ;
  assign y4792 = ~1'b0 ;
  assign y4793 = n11082 ;
  assign y4794 = ~n11084 ;
  assign y4795 = ~n11087 ;
  assign y4796 = ~n11090 ;
  assign y4797 = ~n11091 ;
  assign y4798 = ~n11097 ;
  assign y4799 = ~1'b0 ;
  assign y4800 = ~n11098 ;
  assign y4801 = ~n11104 ;
  assign y4802 = n11107 ;
  assign y4803 = ~n11110 ;
  assign y4804 = n11112 ;
  assign y4805 = ~n11118 ;
  assign y4806 = ~n11126 ;
  assign y4807 = ~1'b0 ;
  assign y4808 = n11129 ;
  assign y4809 = n11131 ;
  assign y4810 = n11132 ;
  assign y4811 = ~1'b0 ;
  assign y4812 = ~n196 ;
  assign y4813 = ~1'b0 ;
  assign y4814 = n11152 ;
  assign y4815 = ~x78 ;
  assign y4816 = ~1'b0 ;
  assign y4817 = n11153 ;
  assign y4818 = ~1'b0 ;
  assign y4819 = ~n11155 ;
  assign y4820 = n11160 ;
  assign y4821 = n11162 ;
  assign y4822 = ~n11167 ;
  assign y4823 = n11168 ;
  assign y4824 = ~n11170 ;
  assign y4825 = ~1'b0 ;
  assign y4826 = ~1'b0 ;
  assign y4827 = ~n11172 ;
  assign y4828 = n11177 ;
  assign y4829 = ~1'b0 ;
  assign y4830 = ~1'b0 ;
  assign y4831 = ~n11182 ;
  assign y4832 = n11189 ;
  assign y4833 = ~1'b0 ;
  assign y4834 = ~1'b0 ;
  assign y4835 = ~n11192 ;
  assign y4836 = ~n11193 ;
  assign y4837 = 1'b0 ;
  assign y4838 = ~n11208 ;
  assign y4839 = ~1'b0 ;
  assign y4840 = n11210 ;
  assign y4841 = n11215 ;
  assign y4842 = ~n11221 ;
  assign y4843 = ~1'b0 ;
  assign y4844 = ~n11222 ;
  assign y4845 = ~n11223 ;
  assign y4846 = ~n11224 ;
  assign y4847 = ~1'b0 ;
  assign y4848 = n11226 ;
  assign y4849 = ~n11229 ;
  assign y4850 = ~n11235 ;
  assign y4851 = ~n11236 ;
  assign y4852 = ~n11238 ;
  assign y4853 = ~1'b0 ;
  assign y4854 = n11239 ;
  assign y4855 = n11242 ;
  assign y4856 = ~n11250 ;
  assign y4857 = ~n11251 ;
  assign y4858 = n11253 ;
  assign y4859 = ~n11254 ;
  assign y4860 = ~n11255 ;
  assign y4861 = ~1'b0 ;
  assign y4862 = n11256 ;
  assign y4863 = ~n11258 ;
  assign y4864 = n11260 ;
  assign y4865 = ~n1578 ;
  assign y4866 = ~1'b0 ;
  assign y4867 = n11262 ;
  assign y4868 = ~n11265 ;
  assign y4869 = ~1'b0 ;
  assign y4870 = n11268 ;
  assign y4871 = n11276 ;
  assign y4872 = ~1'b0 ;
  assign y4873 = n11277 ;
  assign y4874 = ~1'b0 ;
  assign y4875 = ~1'b0 ;
  assign y4876 = ~1'b0 ;
  assign y4877 = ~n11278 ;
  assign y4878 = n11279 ;
  assign y4879 = n11282 ;
  assign y4880 = ~n11283 ;
  assign y4881 = n11284 ;
  assign y4882 = n9592 ;
  assign y4883 = ~n11290 ;
  assign y4884 = n11291 ;
  assign y4885 = ~1'b0 ;
  assign y4886 = ~n11293 ;
  assign y4887 = ~n11295 ;
  assign y4888 = n11297 ;
  assign y4889 = n11299 ;
  assign y4890 = n11302 ;
  assign y4891 = ~n11303 ;
  assign y4892 = ~n11305 ;
  assign y4893 = ~n11309 ;
  assign y4894 = ~n11314 ;
  assign y4895 = n11318 ;
  assign y4896 = ~n11322 ;
  assign y4897 = ~n11326 ;
  assign y4898 = n11332 ;
  assign y4899 = ~n11334 ;
  assign y4900 = ~1'b0 ;
  assign y4901 = ~1'b0 ;
  assign y4902 = n11336 ;
  assign y4903 = ~n11345 ;
  assign y4904 = n11346 ;
  assign y4905 = n11350 ;
  assign y4906 = ~n11354 ;
  assign y4907 = ~n10100 ;
  assign y4908 = ~n11358 ;
  assign y4909 = n11360 ;
  assign y4910 = ~n11363 ;
  assign y4911 = ~n11365 ;
  assign y4912 = ~1'b0 ;
  assign y4913 = n11372 ;
  assign y4914 = n11374 ;
  assign y4915 = ~n11380 ;
  assign y4916 = n11382 ;
  assign y4917 = ~n11383 ;
  assign y4918 = n11385 ;
  assign y4919 = ~1'b0 ;
  assign y4920 = ~1'b0 ;
  assign y4921 = n11386 ;
  assign y4922 = ~1'b0 ;
  assign y4923 = ~1'b0 ;
  assign y4924 = ~1'b0 ;
  assign y4925 = ~1'b0 ;
  assign y4926 = ~n11397 ;
  assign y4927 = ~n11398 ;
  assign y4928 = ~1'b0 ;
  assign y4929 = ~1'b0 ;
  assign y4930 = n11401 ;
  assign y4931 = n11405 ;
  assign y4932 = n11410 ;
  assign y4933 = ~n10741 ;
  assign y4934 = ~1'b0 ;
  assign y4935 = ~n11412 ;
  assign y4936 = ~1'b0 ;
  assign y4937 = ~n11424 ;
  assign y4938 = ~n11425 ;
  assign y4939 = ~1'b0 ;
  assign y4940 = ~1'b0 ;
  assign y4941 = ~1'b0 ;
  assign y4942 = ~1'b0 ;
  assign y4943 = ~n11428 ;
  assign y4944 = n11434 ;
  assign y4945 = ~n11436 ;
  assign y4946 = n11438 ;
  assign y4947 = ~n11441 ;
  assign y4948 = ~1'b0 ;
  assign y4949 = ~1'b0 ;
  assign y4950 = n11443 ;
  assign y4951 = ~1'b0 ;
  assign y4952 = n11445 ;
  assign y4953 = ~1'b0 ;
  assign y4954 = n11448 ;
  assign y4955 = n11450 ;
  assign y4956 = ~n11452 ;
  assign y4957 = ~n11455 ;
  assign y4958 = n11461 ;
  assign y4959 = ~n11464 ;
  assign y4960 = ~n4342 ;
  assign y4961 = ~n11481 ;
  assign y4962 = ~n11485 ;
  assign y4963 = ~n11488 ;
  assign y4964 = ~n11489 ;
  assign y4965 = ~n11491 ;
  assign y4966 = ~n11492 ;
  assign y4967 = n11495 ;
  assign y4968 = ~n11497 ;
  assign y4969 = n910 ;
  assign y4970 = ~1'b0 ;
  assign y4971 = ~n11500 ;
  assign y4972 = n11501 ;
  assign y4973 = ~1'b0 ;
  assign y4974 = n11506 ;
  assign y4975 = n11509 ;
  assign y4976 = ~1'b0 ;
  assign y4977 = 1'b0 ;
  assign y4978 = ~n11511 ;
  assign y4979 = n11514 ;
  assign y4980 = ~n11515 ;
  assign y4981 = ~1'b0 ;
  assign y4982 = ~1'b0 ;
  assign y4983 = ~n11517 ;
  assign y4984 = n11521 ;
  assign y4985 = ~n11522 ;
  assign y4986 = ~n11525 ;
  assign y4987 = ~n11526 ;
  assign y4988 = ~n11529 ;
  assign y4989 = ~n11533 ;
  assign y4990 = n11536 ;
  assign y4991 = ~n11542 ;
  assign y4992 = ~n11546 ;
  assign y4993 = ~n11548 ;
  assign y4994 = n11555 ;
  assign y4995 = n11561 ;
  assign y4996 = ~1'b0 ;
  assign y4997 = n5152 ;
  assign y4998 = ~n11564 ;
  assign y4999 = ~1'b0 ;
  assign y5000 = n11565 ;
  assign y5001 = n11570 ;
  assign y5002 = ~1'b0 ;
  assign y5003 = ~n11572 ;
  assign y5004 = n11576 ;
  assign y5005 = n11582 ;
  assign y5006 = ~1'b0 ;
  assign y5007 = n11585 ;
  assign y5008 = ~n11591 ;
  assign y5009 = ~n11594 ;
  assign y5010 = n11595 ;
  assign y5011 = n11600 ;
  assign y5012 = ~n11602 ;
  assign y5013 = ~1'b0 ;
  assign y5014 = n11605 ;
  assign y5015 = n11606 ;
  assign y5016 = ~1'b0 ;
  assign y5017 = ~1'b0 ;
  assign y5018 = n11609 ;
  assign y5019 = ~n11612 ;
  assign y5020 = n11617 ;
  assign y5021 = ~n11624 ;
  assign y5022 = ~n11629 ;
  assign y5023 = ~n11635 ;
  assign y5024 = n11636 ;
  assign y5025 = ~n11641 ;
  assign y5026 = n11643 ;
  assign y5027 = ~n11644 ;
  assign y5028 = ~1'b0 ;
  assign y5029 = n11649 ;
  assign y5030 = ~1'b0 ;
  assign y5031 = n11651 ;
  assign y5032 = ~n11655 ;
  assign y5033 = ~1'b0 ;
  assign y5034 = ~1'b0 ;
  assign y5035 = ~1'b0 ;
  assign y5036 = ~n11658 ;
  assign y5037 = n11659 ;
  assign y5038 = n6855 ;
  assign y5039 = ~1'b0 ;
  assign y5040 = ~n11663 ;
  assign y5041 = ~n11665 ;
  assign y5042 = ~n11666 ;
  assign y5043 = ~n11667 ;
  assign y5044 = 1'b0 ;
  assign y5045 = n11671 ;
  assign y5046 = n11673 ;
  assign y5047 = ~1'b0 ;
  assign y5048 = n11677 ;
  assign y5049 = ~n11680 ;
  assign y5050 = n11681 ;
  assign y5051 = n11683 ;
  assign y5052 = n11685 ;
  assign y5053 = ~n11688 ;
  assign y5054 = n11694 ;
  assign y5055 = n11700 ;
  assign y5056 = ~n11701 ;
  assign y5057 = n11704 ;
  assign y5058 = n5574 ;
  assign y5059 = ~n11707 ;
  assign y5060 = n8826 ;
  assign y5061 = ~1'b0 ;
  assign y5062 = n11716 ;
  assign y5063 = n4836 ;
  assign y5064 = ~1'b0 ;
  assign y5065 = ~1'b0 ;
  assign y5066 = ~n11718 ;
  assign y5067 = n11719 ;
  assign y5068 = ~n11721 ;
  assign y5069 = ~n11725 ;
  assign y5070 = ~1'b0 ;
  assign y5071 = ~1'b0 ;
  assign y5072 = n11735 ;
  assign y5073 = n11741 ;
  assign y5074 = ~n11743 ;
  assign y5075 = ~1'b0 ;
  assign y5076 = n11746 ;
  assign y5077 = n11747 ;
  assign y5078 = ~n11748 ;
  assign y5079 = ~1'b0 ;
  assign y5080 = n11749 ;
  assign y5081 = n11751 ;
  assign y5082 = ~n11753 ;
  assign y5083 = ~1'b0 ;
  assign y5084 = ~1'b0 ;
  assign y5085 = ~n11756 ;
  assign y5086 = n11758 ;
  assign y5087 = ~n11759 ;
  assign y5088 = ~n11760 ;
  assign y5089 = n11761 ;
  assign y5090 = ~n11765 ;
  assign y5091 = ~1'b0 ;
  assign y5092 = ~n11771 ;
  assign y5093 = ~n11772 ;
  assign y5094 = ~1'b0 ;
  assign y5095 = ~1'b0 ;
  assign y5096 = ~1'b0 ;
  assign y5097 = ~n11774 ;
  assign y5098 = n11785 ;
  assign y5099 = n11789 ;
  assign y5100 = ~n11791 ;
  assign y5101 = n11792 ;
  assign y5102 = n11798 ;
  assign y5103 = n11802 ;
  assign y5104 = ~1'b0 ;
  assign y5105 = ~n11803 ;
  assign y5106 = ~1'b0 ;
  assign y5107 = ~1'b0 ;
  assign y5108 = ~n11807 ;
  assign y5109 = n11814 ;
  assign y5110 = ~n11815 ;
  assign y5111 = ~n11817 ;
  assign y5112 = n11818 ;
  assign y5113 = ~n11821 ;
  assign y5114 = ~1'b0 ;
  assign y5115 = n1118 ;
  assign y5116 = ~n11823 ;
  assign y5117 = n11827 ;
  assign y5118 = n11828 ;
  assign y5119 = ~n11829 ;
  assign y5120 = n11835 ;
  assign y5121 = 1'b0 ;
  assign y5122 = n11838 ;
  assign y5123 = ~1'b0 ;
  assign y5124 = n11840 ;
  assign y5125 = ~n11842 ;
  assign y5126 = ~n11843 ;
  assign y5127 = ~1'b0 ;
  assign y5128 = n11238 ;
  assign y5129 = n11844 ;
  assign y5130 = ~1'b0 ;
  assign y5131 = ~n11849 ;
  assign y5132 = ~1'b0 ;
  assign y5133 = ~1'b0 ;
  assign y5134 = n11851 ;
  assign y5135 = ~n11856 ;
  assign y5136 = n11872 ;
  assign y5137 = n11874 ;
  assign y5138 = n11875 ;
  assign y5139 = ~n11877 ;
  assign y5140 = ~1'b0 ;
  assign y5141 = ~n11880 ;
  assign y5142 = n11885 ;
  assign y5143 = n11886 ;
  assign y5144 = n11890 ;
  assign y5145 = ~1'b0 ;
  assign y5146 = n11894 ;
  assign y5147 = n11896 ;
  assign y5148 = n11902 ;
  assign y5149 = ~1'b0 ;
  assign y5150 = ~1'b0 ;
  assign y5151 = n11912 ;
  assign y5152 = n11915 ;
  assign y5153 = n11917 ;
  assign y5154 = ~1'b0 ;
  assign y5155 = n11920 ;
  assign y5156 = ~1'b0 ;
  assign y5157 = ~n11922 ;
  assign y5158 = ~1'b0 ;
  assign y5159 = ~n11924 ;
  assign y5160 = n11925 ;
  assign y5161 = n7416 ;
  assign y5162 = ~1'b0 ;
  assign y5163 = ~n11937 ;
  assign y5164 = ~1'b0 ;
  assign y5165 = ~n11940 ;
  assign y5166 = n11941 ;
  assign y5167 = n11942 ;
  assign y5168 = n11950 ;
  assign y5169 = ~1'b0 ;
  assign y5170 = ~n11951 ;
  assign y5171 = n11955 ;
  assign y5172 = ~n11959 ;
  assign y5173 = ~1'b0 ;
  assign y5174 = ~1'b0 ;
  assign y5175 = n11960 ;
  assign y5176 = ~n11961 ;
  assign y5177 = n11964 ;
  assign y5178 = ~n11967 ;
  assign y5179 = n11970 ;
  assign y5180 = ~n11972 ;
  assign y5181 = ~1'b0 ;
  assign y5182 = ~1'b0 ;
  assign y5183 = ~1'b0 ;
  assign y5184 = ~n11975 ;
  assign y5185 = ~1'b0 ;
  assign y5186 = ~n11976 ;
  assign y5187 = ~1'b0 ;
  assign y5188 = n11977 ;
  assign y5189 = ~n11981 ;
  assign y5190 = ~n11982 ;
  assign y5191 = n8618 ;
  assign y5192 = n11987 ;
  assign y5193 = 1'b0 ;
  assign y5194 = ~n11988 ;
  assign y5195 = ~1'b0 ;
  assign y5196 = n11990 ;
  assign y5197 = ~n11992 ;
  assign y5198 = ~n11998 ;
  assign y5199 = 1'b0 ;
  assign y5200 = ~1'b0 ;
  assign y5201 = ~1'b0 ;
  assign y5202 = n12002 ;
  assign y5203 = n12003 ;
  assign y5204 = n12004 ;
  assign y5205 = n12008 ;
  assign y5206 = ~n12009 ;
  assign y5207 = ~1'b0 ;
  assign y5208 = ~n12013 ;
  assign y5209 = ~1'b0 ;
  assign y5210 = n12014 ;
  assign y5211 = ~n12016 ;
  assign y5212 = n12017 ;
  assign y5213 = n12018 ;
  assign y5214 = ~n12022 ;
  assign y5215 = ~1'b0 ;
  assign y5216 = ~1'b0 ;
  assign y5217 = ~n12023 ;
  assign y5218 = n12024 ;
  assign y5219 = ~1'b0 ;
  assign y5220 = ~n12029 ;
  assign y5221 = ~1'b0 ;
  assign y5222 = ~n12035 ;
  assign y5223 = ~n12036 ;
  assign y5224 = 1'b0 ;
  assign y5225 = ~1'b0 ;
  assign y5226 = ~n12044 ;
  assign y5227 = ~1'b0 ;
  assign y5228 = ~1'b0 ;
  assign y5229 = ~n12045 ;
  assign y5230 = n12046 ;
  assign y5231 = ~1'b0 ;
  assign y5232 = n12049 ;
  assign y5233 = ~n4875 ;
  assign y5234 = n12051 ;
  assign y5235 = n12060 ;
  assign y5236 = ~1'b0 ;
  assign y5237 = n12061 ;
  assign y5238 = n12063 ;
  assign y5239 = n12065 ;
  assign y5240 = n12067 ;
  assign y5241 = n12070 ;
  assign y5242 = n12071 ;
  assign y5243 = n12076 ;
  assign y5244 = n12077 ;
  assign y5245 = ~n12079 ;
  assign y5246 = ~1'b0 ;
  assign y5247 = ~n12083 ;
  assign y5248 = ~n12084 ;
  assign y5249 = ~n12085 ;
  assign y5250 = n12089 ;
  assign y5251 = ~n12096 ;
  assign y5252 = ~n12097 ;
  assign y5253 = ~n12099 ;
  assign y5254 = ~n12101 ;
  assign y5255 = n12107 ;
  assign y5256 = ~1'b0 ;
  assign y5257 = ~1'b0 ;
  assign y5258 = n6075 ;
  assign y5259 = n12110 ;
  assign y5260 = n12112 ;
  assign y5261 = ~1'b0 ;
  assign y5262 = n12113 ;
  assign y5263 = n12115 ;
  assign y5264 = n12119 ;
  assign y5265 = ~n12120 ;
  assign y5266 = ~1'b0 ;
  assign y5267 = ~n12121 ;
  assign y5268 = ~n12122 ;
  assign y5269 = n12124 ;
  assign y5270 = ~n12125 ;
  assign y5271 = n12126 ;
  assign y5272 = ~n12129 ;
  assign y5273 = ~n12130 ;
  assign y5274 = ~n12132 ;
  assign y5275 = n12135 ;
  assign y5276 = ~1'b0 ;
  assign y5277 = n12136 ;
  assign y5278 = ~n12137 ;
  assign y5279 = n12140 ;
  assign y5280 = ~1'b0 ;
  assign y5281 = ~1'b0 ;
  assign y5282 = n12141 ;
  assign y5283 = ~n12145 ;
  assign y5284 = n12152 ;
  assign y5285 = n12164 ;
  assign y5286 = n12165 ;
  assign y5287 = n12167 ;
  assign y5288 = ~n12168 ;
  assign y5289 = n12173 ;
  assign y5290 = ~1'b0 ;
  assign y5291 = ~n10439 ;
  assign y5292 = ~n12180 ;
  assign y5293 = n12184 ;
  assign y5294 = n1583 ;
  assign y5295 = n12187 ;
  assign y5296 = ~1'b0 ;
  assign y5297 = ~n12192 ;
  assign y5298 = n12194 ;
  assign y5299 = ~1'b0 ;
  assign y5300 = ~1'b0 ;
  assign y5301 = ~n12195 ;
  assign y5302 = n12198 ;
  assign y5303 = ~1'b0 ;
  assign y5304 = n12199 ;
  assign y5305 = ~n12201 ;
  assign y5306 = ~n12204 ;
  assign y5307 = ~n12206 ;
  assign y5308 = ~1'b0 ;
  assign y5309 = ~1'b0 ;
  assign y5310 = ~n12216 ;
  assign y5311 = ~n12218 ;
  assign y5312 = ~1'b0 ;
  assign y5313 = n12219 ;
  assign y5314 = ~1'b0 ;
  assign y5315 = ~1'b0 ;
  assign y5316 = n12220 ;
  assign y5317 = ~n12229 ;
  assign y5318 = ~1'b0 ;
  assign y5319 = ~1'b0 ;
  assign y5320 = ~n12230 ;
  assign y5321 = ~n12231 ;
  assign y5322 = ~n12235 ;
  assign y5323 = ~n12239 ;
  assign y5324 = ~n12241 ;
  assign y5325 = ~n12242 ;
  assign y5326 = n12244 ;
  assign y5327 = ~n12248 ;
  assign y5328 = ~1'b0 ;
  assign y5329 = ~1'b0 ;
  assign y5330 = n12251 ;
  assign y5331 = n12253 ;
  assign y5332 = ~n12263 ;
  assign y5333 = ~n12264 ;
  assign y5334 = ~1'b0 ;
  assign y5335 = n12266 ;
  assign y5336 = n12267 ;
  assign y5337 = ~n12269 ;
  assign y5338 = ~1'b0 ;
  assign y5339 = n12273 ;
  assign y5340 = n12275 ;
  assign y5341 = ~1'b0 ;
  assign y5342 = ~n12282 ;
  assign y5343 = ~n12286 ;
  assign y5344 = ~n12289 ;
  assign y5345 = ~n12291 ;
  assign y5346 = ~n12303 ;
  assign y5347 = 1'b0 ;
  assign y5348 = ~1'b0 ;
  assign y5349 = ~n12309 ;
  assign y5350 = ~n12310 ;
  assign y5351 = ~1'b0 ;
  assign y5352 = ~n12316 ;
  assign y5353 = ~1'b0 ;
  assign y5354 = ~n12317 ;
  assign y5355 = ~n12318 ;
  assign y5356 = ~1'b0 ;
  assign y5357 = ~1'b0 ;
  assign y5358 = ~n3896 ;
  assign y5359 = ~n12319 ;
  assign y5360 = n7075 ;
  assign y5361 = 1'b0 ;
  assign y5362 = n12320 ;
  assign y5363 = n12322 ;
  assign y5364 = ~n3861 ;
  assign y5365 = ~n12323 ;
  assign y5366 = ~n2594 ;
  assign y5367 = ~n12326 ;
  assign y5368 = n12329 ;
  assign y5369 = n12333 ;
  assign y5370 = ~1'b0 ;
  assign y5371 = ~n12334 ;
  assign y5372 = ~n12336 ;
  assign y5373 = n12341 ;
  assign y5374 = ~1'b0 ;
  assign y5375 = ~n12343 ;
  assign y5376 = ~1'b0 ;
  assign y5377 = ~n12348 ;
  assign y5378 = n12351 ;
  assign y5379 = n12355 ;
  assign y5380 = ~1'b0 ;
  assign y5381 = ~n12357 ;
  assign y5382 = n12358 ;
  assign y5383 = ~1'b0 ;
  assign y5384 = ~1'b0 ;
  assign y5385 = ~1'b0 ;
  assign y5386 = ~n12361 ;
  assign y5387 = n12364 ;
  assign y5388 = n12366 ;
  assign y5389 = ~n12369 ;
  assign y5390 = ~1'b0 ;
  assign y5391 = n12373 ;
  assign y5392 = ~n12374 ;
  assign y5393 = ~n12376 ;
  assign y5394 = ~n12378 ;
  assign y5395 = ~n12380 ;
  assign y5396 = n12384 ;
  assign y5397 = ~1'b0 ;
  assign y5398 = ~n12385 ;
  assign y5399 = n4827 ;
  assign y5400 = ~1'b0 ;
  assign y5401 = ~n5412 ;
  assign y5402 = n12387 ;
  assign y5403 = ~n12390 ;
  assign y5404 = ~1'b0 ;
  assign y5405 = ~1'b0 ;
  assign y5406 = n12391 ;
  assign y5407 = n12397 ;
  assign y5408 = ~1'b0 ;
  assign y5409 = n12402 ;
  assign y5410 = ~n12404 ;
  assign y5411 = ~n12415 ;
  assign y5412 = n12416 ;
  assign y5413 = ~1'b0 ;
  assign y5414 = ~n6603 ;
  assign y5415 = n12417 ;
  assign y5416 = n12418 ;
  assign y5417 = ~n12419 ;
  assign y5418 = n12420 ;
  assign y5419 = ~1'b0 ;
  assign y5420 = ~1'b0 ;
  assign y5421 = n12423 ;
  assign y5422 = ~n12425 ;
  assign y5423 = ~1'b0 ;
  assign y5424 = ~n12426 ;
  assign y5425 = n12430 ;
  assign y5426 = n12432 ;
  assign y5427 = ~n12433 ;
  assign y5428 = ~n12438 ;
  assign y5429 = n12441 ;
  assign y5430 = ~1'b0 ;
  assign y5431 = ~1'b0 ;
  assign y5432 = ~n12447 ;
  assign y5433 = n12453 ;
  assign y5434 = ~1'b0 ;
  assign y5435 = ~n12456 ;
  assign y5436 = n12459 ;
  assign y5437 = ~1'b0 ;
  assign y5438 = ~1'b0 ;
  assign y5439 = n12463 ;
  assign y5440 = n12465 ;
  assign y5441 = n12466 ;
  assign y5442 = ~n12471 ;
  assign y5443 = ~1'b0 ;
  assign y5444 = n12474 ;
  assign y5445 = ~n12475 ;
  assign y5446 = ~n12480 ;
  assign y5447 = ~n12486 ;
  assign y5448 = n12492 ;
  assign y5449 = ~1'b0 ;
  assign y5450 = ~n12493 ;
  assign y5451 = ~n12495 ;
  assign y5452 = 1'b0 ;
  assign y5453 = ~1'b0 ;
  assign y5454 = n12497 ;
  assign y5455 = ~1'b0 ;
  assign y5456 = n12498 ;
  assign y5457 = ~n12499 ;
  assign y5458 = ~1'b0 ;
  assign y5459 = n12503 ;
  assign y5460 = ~1'b0 ;
  assign y5461 = ~n12504 ;
  assign y5462 = ~n12506 ;
  assign y5463 = n12508 ;
  assign y5464 = ~n12509 ;
  assign y5465 = ~1'b0 ;
  assign y5466 = ~n12510 ;
  assign y5467 = ~n6197 ;
  assign y5468 = ~1'b0 ;
  assign y5469 = n12514 ;
  assign y5470 = ~1'b0 ;
  assign y5471 = n12515 ;
  assign y5472 = ~n12516 ;
  assign y5473 = n12521 ;
  assign y5474 = ~1'b0 ;
  assign y5475 = ~1'b0 ;
  assign y5476 = ~1'b0 ;
  assign y5477 = ~n12522 ;
  assign y5478 = n12523 ;
  assign y5479 = ~1'b0 ;
  assign y5480 = ~n12524 ;
  assign y5481 = ~n11101 ;
  assign y5482 = ~n12528 ;
  assign y5483 = n6124 ;
  assign y5484 = n12534 ;
  assign y5485 = n12537 ;
  assign y5486 = ~1'b0 ;
  assign y5487 = ~1'b0 ;
  assign y5488 = n12540 ;
  assign y5489 = ~n12541 ;
  assign y5490 = 1'b0 ;
  assign y5491 = n12544 ;
  assign y5492 = n12550 ;
  assign y5493 = ~n12552 ;
  assign y5494 = ~n12554 ;
  assign y5495 = ~n12556 ;
  assign y5496 = ~1'b0 ;
  assign y5497 = n12561 ;
  assign y5498 = ~n5324 ;
  assign y5499 = ~n12566 ;
  assign y5500 = ~n12568 ;
  assign y5501 = ~n12570 ;
  assign y5502 = ~n12572 ;
  assign y5503 = ~n12573 ;
  assign y5504 = ~n12575 ;
  assign y5505 = ~1'b0 ;
  assign y5506 = ~n12580 ;
  assign y5507 = ~1'b0 ;
  assign y5508 = ~1'b0 ;
  assign y5509 = ~n12582 ;
  assign y5510 = ~n12585 ;
  assign y5511 = ~n12586 ;
  assign y5512 = n12587 ;
  assign y5513 = n12589 ;
  assign y5514 = ~1'b0 ;
  assign y5515 = ~n12591 ;
  assign y5516 = ~1'b0 ;
  assign y5517 = ~1'b0 ;
  assign y5518 = ~n12593 ;
  assign y5519 = ~n12594 ;
  assign y5520 = ~n12595 ;
  assign y5521 = n12596 ;
  assign y5522 = n12598 ;
  assign y5523 = ~1'b0 ;
  assign y5524 = ~n12600 ;
  assign y5525 = ~n12601 ;
  assign y5526 = n510 ;
  assign y5527 = n12603 ;
  assign y5528 = ~n3858 ;
  assign y5529 = ~1'b0 ;
  assign y5530 = ~n12608 ;
  assign y5531 = n12611 ;
  assign y5532 = n12616 ;
  assign y5533 = n12618 ;
  assign y5534 = n12619 ;
  assign y5535 = ~n12620 ;
  assign y5536 = n12623 ;
  assign y5537 = n12628 ;
  assign y5538 = ~n5117 ;
  assign y5539 = ~n12629 ;
  assign y5540 = ~1'b0 ;
  assign y5541 = ~n12630 ;
  assign y5542 = n6119 ;
  assign y5543 = ~n12633 ;
  assign y5544 = ~n12635 ;
  assign y5545 = ~1'b0 ;
  assign y5546 = n12636 ;
  assign y5547 = ~n12638 ;
  assign y5548 = n12639 ;
  assign y5549 = ~n12640 ;
  assign y5550 = ~1'b0 ;
  assign y5551 = ~1'b0 ;
  assign y5552 = n12641 ;
  assign y5553 = ~n12642 ;
  assign y5554 = ~n12644 ;
  assign y5555 = n7837 ;
  assign y5556 = ~n12645 ;
  assign y5557 = n12648 ;
  assign y5558 = n12657 ;
  assign y5559 = n12658 ;
  assign y5560 = ~1'b0 ;
  assign y5561 = n12663 ;
  assign y5562 = n12672 ;
  assign y5563 = ~n12673 ;
  assign y5564 = ~n12674 ;
  assign y5565 = ~n12677 ;
  assign y5566 = ~n12678 ;
  assign y5567 = n12679 ;
  assign y5568 = n12685 ;
  assign y5569 = n12687 ;
  assign y5570 = ~1'b0 ;
  assign y5571 = ~n12691 ;
  assign y5572 = n12692 ;
  assign y5573 = ~n12695 ;
  assign y5574 = ~n12697 ;
  assign y5575 = n12702 ;
  assign y5576 = ~1'b0 ;
  assign y5577 = ~n12703 ;
  assign y5578 = n12704 ;
  assign y5579 = ~n12706 ;
  assign y5580 = n12709 ;
  assign y5581 = n12712 ;
  assign y5582 = n12713 ;
  assign y5583 = n6312 ;
  assign y5584 = ~1'b0 ;
  assign y5585 = ~1'b0 ;
  assign y5586 = ~1'b0 ;
  assign y5587 = ~n12714 ;
  assign y5588 = ~n12718 ;
  assign y5589 = n12719 ;
  assign y5590 = 1'b0 ;
  assign y5591 = n12722 ;
  assign y5592 = ~n12723 ;
  assign y5593 = ~1'b0 ;
  assign y5594 = ~1'b0 ;
  assign y5595 = ~1'b0 ;
  assign y5596 = n12725 ;
  assign y5597 = ~n12726 ;
  assign y5598 = n12731 ;
  assign y5599 = ~n12732 ;
  assign y5600 = ~n12736 ;
  assign y5601 = n8996 ;
  assign y5602 = ~1'b0 ;
  assign y5603 = n12741 ;
  assign y5604 = ~n12748 ;
  assign y5605 = n12753 ;
  assign y5606 = n12757 ;
  assign y5607 = ~n12763 ;
  assign y5608 = ~n12766 ;
  assign y5609 = ~n12769 ;
  assign y5610 = ~n12773 ;
  assign y5611 = n12777 ;
  assign y5612 = ~n12782 ;
  assign y5613 = n12787 ;
  assign y5614 = ~n12790 ;
  assign y5615 = ~n12799 ;
  assign y5616 = n12801 ;
  assign y5617 = ~1'b0 ;
  assign y5618 = ~1'b0 ;
  assign y5619 = ~n12802 ;
  assign y5620 = n12803 ;
  assign y5621 = ~1'b0 ;
  assign y5622 = n12805 ;
  assign y5623 = n12807 ;
  assign y5624 = n12810 ;
  assign y5625 = ~1'b0 ;
  assign y5626 = ~n12821 ;
  assign y5627 = ~n12823 ;
  assign y5628 = ~n12825 ;
  assign y5629 = n12826 ;
  assign y5630 = n12829 ;
  assign y5631 = ~n12833 ;
  assign y5632 = ~1'b0 ;
  assign y5633 = n12836 ;
  assign y5634 = ~n12838 ;
  assign y5635 = n12845 ;
  assign y5636 = n12854 ;
  assign y5637 = ~n12856 ;
  assign y5638 = ~n12862 ;
  assign y5639 = n12865 ;
  assign y5640 = ~n12866 ;
  assign y5641 = ~1'b0 ;
  assign y5642 = ~1'b0 ;
  assign y5643 = n12868 ;
  assign y5644 = n12875 ;
  assign y5645 = ~n12887 ;
  assign y5646 = ~1'b0 ;
  assign y5647 = ~n12889 ;
  assign y5648 = ~n12891 ;
  assign y5649 = n12894 ;
  assign y5650 = ~n12898 ;
  assign y5651 = ~n12908 ;
  assign y5652 = n12911 ;
  assign y5653 = ~n12913 ;
  assign y5654 = n12917 ;
  assign y5655 = n12918 ;
  assign y5656 = n12921 ;
  assign y5657 = ~n12922 ;
  assign y5658 = ~n12927 ;
  assign y5659 = n12931 ;
  assign y5660 = ~n12935 ;
  assign y5661 = ~n12936 ;
  assign y5662 = ~n12937 ;
  assign y5663 = n12940 ;
  assign y5664 = n12943 ;
  assign y5665 = ~n12961 ;
  assign y5666 = ~1'b0 ;
  assign y5667 = n12962 ;
  assign y5668 = n12965 ;
  assign y5669 = ~1'b0 ;
  assign y5670 = ~n12966 ;
  assign y5671 = ~n12969 ;
  assign y5672 = n12970 ;
  assign y5673 = ~n12974 ;
  assign y5674 = n12975 ;
  assign y5675 = ~1'b0 ;
  assign y5676 = ~1'b0 ;
  assign y5677 = ~1'b0 ;
  assign y5678 = ~n12976 ;
  assign y5679 = ~n12978 ;
  assign y5680 = ~n12981 ;
  assign y5681 = n12987 ;
  assign y5682 = ~1'b0 ;
  assign y5683 = ~n12991 ;
  assign y5684 = ~1'b0 ;
  assign y5685 = n12993 ;
  assign y5686 = ~1'b0 ;
  assign y5687 = ~1'b0 ;
  assign y5688 = n12367 ;
  assign y5689 = ~n12802 ;
  assign y5690 = ~n12995 ;
  assign y5691 = ~1'b0 ;
  assign y5692 = n12996 ;
  assign y5693 = ~1'b0 ;
  assign y5694 = n12997 ;
  assign y5695 = ~n13000 ;
  assign y5696 = n13004 ;
  assign y5697 = 1'b0 ;
  assign y5698 = ~n13005 ;
  assign y5699 = ~n13011 ;
  assign y5700 = ~n13014 ;
  assign y5701 = ~1'b0 ;
  assign y5702 = ~1'b0 ;
  assign y5703 = ~n13016 ;
  assign y5704 = n2882 ;
  assign y5705 = ~1'b0 ;
  assign y5706 = n4432 ;
  assign y5707 = ~n13017 ;
  assign y5708 = ~n13024 ;
  assign y5709 = n13029 ;
  assign y5710 = ~1'b0 ;
  assign y5711 = ~n13031 ;
  assign y5712 = n13032 ;
  assign y5713 = ~1'b0 ;
  assign y5714 = n13035 ;
  assign y5715 = ~n13037 ;
  assign y5716 = n13039 ;
  assign y5717 = ~1'b0 ;
  assign y5718 = ~1'b0 ;
  assign y5719 = n13041 ;
  assign y5720 = n13044 ;
  assign y5721 = n13046 ;
  assign y5722 = ~n13049 ;
  assign y5723 = ~n13056 ;
  assign y5724 = n13061 ;
  assign y5725 = n13067 ;
  assign y5726 = n13072 ;
  assign y5727 = n326 ;
  assign y5728 = ~n13075 ;
  assign y5729 = n13077 ;
  assign y5730 = ~n13079 ;
  assign y5731 = n13086 ;
  assign y5732 = ~n13088 ;
  assign y5733 = ~1'b0 ;
  assign y5734 = ~1'b0 ;
  assign y5735 = ~1'b0 ;
  assign y5736 = ~1'b0 ;
  assign y5737 = ~n13092 ;
  assign y5738 = ~n13094 ;
  assign y5739 = n13098 ;
  assign y5740 = ~n13100 ;
  assign y5741 = 1'b0 ;
  assign y5742 = n13101 ;
  assign y5743 = ~n13103 ;
  assign y5744 = ~n13105 ;
  assign y5745 = ~n13109 ;
  assign y5746 = ~1'b0 ;
  assign y5747 = ~n13116 ;
  assign y5748 = ~n13130 ;
  assign y5749 = n13132 ;
  assign y5750 = ~1'b0 ;
  assign y5751 = ~n13136 ;
  assign y5752 = ~n13137 ;
  assign y5753 = ~n13138 ;
  assign y5754 = ~1'b0 ;
  assign y5755 = n13141 ;
  assign y5756 = n13145 ;
  assign y5757 = ~n13147 ;
  assign y5758 = ~n13151 ;
  assign y5759 = ~n13156 ;
  assign y5760 = ~n13158 ;
  assign y5761 = ~n13160 ;
  assign y5762 = n13162 ;
  assign y5763 = ~n13168 ;
  assign y5764 = n13169 ;
  assign y5765 = n13170 ;
  assign y5766 = n13173 ;
  assign y5767 = ~1'b0 ;
  assign y5768 = ~1'b0 ;
  assign y5769 = n13174 ;
  assign y5770 = n13176 ;
  assign y5771 = ~1'b0 ;
  assign y5772 = n13178 ;
  assign y5773 = n13189 ;
  assign y5774 = ~1'b0 ;
  assign y5775 = n13193 ;
  assign y5776 = n13202 ;
  assign y5777 = n13204 ;
  assign y5778 = ~1'b0 ;
  assign y5779 = ~n13210 ;
  assign y5780 = 1'b0 ;
  assign y5781 = n1305 ;
  assign y5782 = ~1'b0 ;
  assign y5783 = ~1'b0 ;
  assign y5784 = n5911 ;
  assign y5785 = n13213 ;
  assign y5786 = n13216 ;
  assign y5787 = 1'b0 ;
  assign y5788 = n13217 ;
  assign y5789 = ~1'b0 ;
  assign y5790 = ~1'b0 ;
  assign y5791 = ~n13224 ;
  assign y5792 = ~n13234 ;
  assign y5793 = n13241 ;
  assign y5794 = ~n13243 ;
  assign y5795 = ~n13250 ;
  assign y5796 = n1268 ;
  assign y5797 = n13253 ;
  assign y5798 = ~n13255 ;
  assign y5799 = n13256 ;
  assign y5800 = ~1'b0 ;
  assign y5801 = n13257 ;
  assign y5802 = ~n12500 ;
  assign y5803 = ~1'b0 ;
  assign y5804 = ~n13258 ;
  assign y5805 = ~n13259 ;
  assign y5806 = ~n13267 ;
  assign y5807 = ~n13272 ;
  assign y5808 = ~n13277 ;
  assign y5809 = ~1'b0 ;
  assign y5810 = ~1'b0 ;
  assign y5811 = n13279 ;
  assign y5812 = ~n13280 ;
  assign y5813 = n13282 ;
  assign y5814 = n13283 ;
  assign y5815 = ~1'b0 ;
  assign y5816 = ~n13284 ;
  assign y5817 = ~1'b0 ;
  assign y5818 = ~1'b0 ;
  assign y5819 = ~n13285 ;
  assign y5820 = ~1'b0 ;
  assign y5821 = n13291 ;
  assign y5822 = ~1'b0 ;
  assign y5823 = ~1'b0 ;
  assign y5824 = n13292 ;
  assign y5825 = ~n13293 ;
  assign y5826 = ~1'b0 ;
  assign y5827 = ~n13294 ;
  assign y5828 = n3178 ;
  assign y5829 = ~n13301 ;
  assign y5830 = ~n13305 ;
  assign y5831 = n13309 ;
  assign y5832 = n13312 ;
  assign y5833 = ~1'b0 ;
  assign y5834 = ~1'b0 ;
  assign y5835 = ~1'b0 ;
  assign y5836 = n13314 ;
  assign y5837 = n13315 ;
  assign y5838 = ~1'b0 ;
  assign y5839 = ~1'b0 ;
  assign y5840 = ~n13318 ;
  assign y5841 = ~n13321 ;
  assign y5842 = n13322 ;
  assign y5843 = ~n13323 ;
  assign y5844 = ~n13325 ;
  assign y5845 = ~n13326 ;
  assign y5846 = ~n13327 ;
  assign y5847 = n13331 ;
  assign y5848 = ~1'b0 ;
  assign y5849 = ~n10959 ;
  assign y5850 = ~n13333 ;
  assign y5851 = n13334 ;
  assign y5852 = ~n13337 ;
  assign y5853 = ~1'b0 ;
  assign y5854 = n2441 ;
  assign y5855 = n13338 ;
  assign y5856 = ~n13344 ;
  assign y5857 = n13348 ;
  assign y5858 = ~1'b0 ;
  assign y5859 = n13350 ;
  assign y5860 = ~n13353 ;
  assign y5861 = n13358 ;
  assign y5862 = ~1'b0 ;
  assign y5863 = ~1'b0 ;
  assign y5864 = ~1'b0 ;
  assign y5865 = ~n13364 ;
  assign y5866 = ~1'b0 ;
  assign y5867 = ~n13367 ;
  assign y5868 = n13369 ;
  assign y5869 = ~n13375 ;
  assign y5870 = ~n13376 ;
  assign y5871 = n13378 ;
  assign y5872 = ~n13380 ;
  assign y5873 = n13382 ;
  assign y5874 = ~1'b0 ;
  assign y5875 = n13385 ;
  assign y5876 = ~n13387 ;
  assign y5877 = n13388 ;
  assign y5878 = n13389 ;
  assign y5879 = ~1'b0 ;
  assign y5880 = n13391 ;
  assign y5881 = n13392 ;
  assign y5882 = n13395 ;
  assign y5883 = n13402 ;
  assign y5884 = ~1'b0 ;
  assign y5885 = ~1'b0 ;
  assign y5886 = ~1'b0 ;
  assign y5887 = ~n13405 ;
  assign y5888 = ~1'b0 ;
  assign y5889 = ~n13406 ;
  assign y5890 = n6524 ;
  assign y5891 = n13408 ;
  assign y5892 = ~1'b0 ;
  assign y5893 = n13409 ;
  assign y5894 = ~n13413 ;
  assign y5895 = n13415 ;
  assign y5896 = ~n13417 ;
  assign y5897 = ~n13421 ;
  assign y5898 = ~1'b0 ;
  assign y5899 = n13422 ;
  assign y5900 = n13427 ;
  assign y5901 = ~n13430 ;
  assign y5902 = n13431 ;
  assign y5903 = n4806 ;
  assign y5904 = ~n13434 ;
  assign y5905 = ~1'b0 ;
  assign y5906 = ~1'b0 ;
  assign y5907 = ~1'b0 ;
  assign y5908 = ~1'b0 ;
  assign y5909 = ~n13435 ;
  assign y5910 = ~n13441 ;
  assign y5911 = n13447 ;
  assign y5912 = n13452 ;
  assign y5913 = ~n13455 ;
  assign y5914 = n13458 ;
  assign y5915 = n13465 ;
  assign y5916 = ~n13469 ;
  assign y5917 = ~n13472 ;
  assign y5918 = n13473 ;
  assign y5919 = ~1'b0 ;
  assign y5920 = n13489 ;
  assign y5921 = ~1'b0 ;
  assign y5922 = ~1'b0 ;
  assign y5923 = ~n13501 ;
  assign y5924 = n13505 ;
  assign y5925 = ~1'b0 ;
  assign y5926 = ~n13506 ;
  assign y5927 = ~n13508 ;
  assign y5928 = ~n13509 ;
  assign y5929 = n13510 ;
  assign y5930 = ~1'b0 ;
  assign y5931 = ~n13514 ;
  assign y5932 = ~1'b0 ;
  assign y5933 = n13516 ;
  assign y5934 = ~1'b0 ;
  assign y5935 = n13518 ;
  assign y5936 = ~n13522 ;
  assign y5937 = ~1'b0 ;
  assign y5938 = ~1'b0 ;
  assign y5939 = n13524 ;
  assign y5940 = n13525 ;
  assign y5941 = ~1'b0 ;
  assign y5942 = n13526 ;
  assign y5943 = ~n13529 ;
  assign y5944 = ~1'b0 ;
  assign y5945 = n13540 ;
  assign y5946 = ~n13542 ;
  assign y5947 = ~n13544 ;
  assign y5948 = ~1'b0 ;
  assign y5949 = ~1'b0 ;
  assign y5950 = ~n13552 ;
  assign y5951 = ~n13553 ;
  assign y5952 = n13556 ;
  assign y5953 = n13558 ;
  assign y5954 = ~1'b0 ;
  assign y5955 = ~1'b0 ;
  assign y5956 = ~n13563 ;
  assign y5957 = ~1'b0 ;
  assign y5958 = n13564 ;
  assign y5959 = ~1'b0 ;
  assign y5960 = ~n13566 ;
  assign y5961 = ~1'b0 ;
  assign y5962 = n13568 ;
  assign y5963 = ~n13572 ;
  assign y5964 = ~n13573 ;
  assign y5965 = ~1'b0 ;
  assign y5966 = n13581 ;
  assign y5967 = n13583 ;
  assign y5968 = ~n11440 ;
  assign y5969 = n13585 ;
  assign y5970 = n13587 ;
  assign y5971 = ~n13592 ;
  assign y5972 = ~1'b0 ;
  assign y5973 = n13594 ;
  assign y5974 = ~n13595 ;
  assign y5975 = n13596 ;
  assign y5976 = ~n13599 ;
  assign y5977 = ~n8500 ;
  assign y5978 = ~n13601 ;
  assign y5979 = n13602 ;
  assign y5980 = n13608 ;
  assign y5981 = 1'b0 ;
  assign y5982 = ~n13610 ;
  assign y5983 = n13614 ;
  assign y5984 = ~1'b0 ;
  assign y5985 = ~1'b0 ;
  assign y5986 = n13616 ;
  assign y5987 = ~n13617 ;
  assign y5988 = ~n13624 ;
  assign y5989 = n13628 ;
  assign y5990 = n13629 ;
  assign y5991 = n13637 ;
  assign y5992 = n13639 ;
  assign y5993 = n13641 ;
  assign y5994 = ~n13643 ;
  assign y5995 = ~n13646 ;
  assign y5996 = n13652 ;
  assign y5997 = n6133 ;
  assign y5998 = ~n13656 ;
  assign y5999 = ~1'b0 ;
  assign y6000 = n13658 ;
  assign y6001 = n13659 ;
  assign y6002 = n13660 ;
  assign y6003 = n13663 ;
  assign y6004 = n13669 ;
  assign y6005 = ~n13670 ;
  assign y6006 = ~1'b0 ;
  assign y6007 = ~1'b0 ;
  assign y6008 = ~1'b0 ;
  assign y6009 = ~1'b0 ;
  assign y6010 = ~n13672 ;
  assign y6011 = n13673 ;
  assign y6012 = ~1'b0 ;
  assign y6013 = ~n13675 ;
  assign y6014 = ~n13676 ;
  assign y6015 = ~n13679 ;
  assign y6016 = ~n13681 ;
  assign y6017 = n13685 ;
  assign y6018 = n13693 ;
  assign y6019 = ~1'b0 ;
  assign y6020 = n10843 ;
  assign y6021 = n13694 ;
  assign y6022 = ~1'b0 ;
  assign y6023 = ~1'b0 ;
  assign y6024 = n13695 ;
  assign y6025 = n13704 ;
  assign y6026 = n13707 ;
  assign y6027 = ~1'b0 ;
  assign y6028 = n13708 ;
  assign y6029 = n13710 ;
  assign y6030 = n13715 ;
  assign y6031 = n13717 ;
  assign y6032 = ~1'b0 ;
  assign y6033 = ~1'b0 ;
  assign y6034 = ~1'b0 ;
  assign y6035 = n13718 ;
  assign y6036 = n13723 ;
  assign y6037 = n13725 ;
  assign y6038 = ~n13726 ;
  assign y6039 = n13728 ;
  assign y6040 = ~n13729 ;
  assign y6041 = ~n13735 ;
  assign y6042 = ~n13737 ;
  assign y6043 = 1'b0 ;
  assign y6044 = ~n13739 ;
  assign y6045 = ~n13741 ;
  assign y6046 = ~1'b0 ;
  assign y6047 = n13746 ;
  assign y6048 = ~n13753 ;
  assign y6049 = ~n13755 ;
  assign y6050 = ~n13756 ;
  assign y6051 = n13759 ;
  assign y6052 = ~1'b0 ;
  assign y6053 = n13762 ;
  assign y6054 = n13771 ;
  assign y6055 = n13773 ;
  assign y6056 = n13774 ;
  assign y6057 = ~1'b0 ;
  assign y6058 = ~n13777 ;
  assign y6059 = ~1'b0 ;
  assign y6060 = ~n13781 ;
  assign y6061 = n13785 ;
  assign y6062 = ~n13789 ;
  assign y6063 = n13797 ;
  assign y6064 = n13805 ;
  assign y6065 = ~1'b0 ;
  assign y6066 = ~n13816 ;
  assign y6067 = ~1'b0 ;
  assign y6068 = ~1'b0 ;
  assign y6069 = n13817 ;
  assign y6070 = n13818 ;
  assign y6071 = n13819 ;
  assign y6072 = ~1'b0 ;
  assign y6073 = ~n13822 ;
  assign y6074 = ~n13825 ;
  assign y6075 = ~n13830 ;
  assign y6076 = n13832 ;
  assign y6077 = ~1'b0 ;
  assign y6078 = ~1'b0 ;
  assign y6079 = ~n13835 ;
  assign y6080 = ~n13836 ;
  assign y6081 = ~1'b0 ;
  assign y6082 = ~1'b0 ;
  assign y6083 = ~n13837 ;
  assign y6084 = n13839 ;
  assign y6085 = n13840 ;
  assign y6086 = ~n13844 ;
  assign y6087 = ~n13845 ;
  assign y6088 = ~n13848 ;
  assign y6089 = n13851 ;
  assign y6090 = ~1'b0 ;
  assign y6091 = ~n13853 ;
  assign y6092 = n13856 ;
  assign y6093 = ~n13858 ;
  assign y6094 = ~1'b0 ;
  assign y6095 = n13859 ;
  assign y6096 = ~n13862 ;
  assign y6097 = ~n13875 ;
  assign y6098 = ~n13877 ;
  assign y6099 = ~1'b0 ;
  assign y6100 = n13880 ;
  assign y6101 = ~n13887 ;
  assign y6102 = ~n13888 ;
  assign y6103 = n13890 ;
  assign y6104 = ~1'b0 ;
  assign y6105 = n13891 ;
  assign y6106 = n13896 ;
  assign y6107 = ~n13897 ;
  assign y6108 = ~n13898 ;
  assign y6109 = ~n10435 ;
  assign y6110 = n13900 ;
  assign y6111 = n13904 ;
  assign y6112 = ~1'b0 ;
  assign y6113 = n13905 ;
  assign y6114 = ~n13907 ;
  assign y6115 = n13910 ;
  assign y6116 = ~1'b0 ;
  assign y6117 = ~1'b0 ;
  assign y6118 = n13917 ;
  assign y6119 = n13924 ;
  assign y6120 = n3465 ;
  assign y6121 = ~1'b0 ;
  assign y6122 = ~n13933 ;
  assign y6123 = n13934 ;
  assign y6124 = n13935 ;
  assign y6125 = ~1'b0 ;
  assign y6126 = n13939 ;
  assign y6127 = ~1'b0 ;
  assign y6128 = n13945 ;
  assign y6129 = n13953 ;
  assign y6130 = ~n13957 ;
  assign y6131 = ~1'b0 ;
  assign y6132 = ~n12132 ;
  assign y6133 = ~n13962 ;
  assign y6134 = n13963 ;
  assign y6135 = ~1'b0 ;
  assign y6136 = ~1'b0 ;
  assign y6137 = ~n13965 ;
  assign y6138 = n13967 ;
  assign y6139 = n13971 ;
  assign y6140 = ~n13972 ;
  assign y6141 = ~n13977 ;
  assign y6142 = ~1'b0 ;
  assign y6143 = ~1'b0 ;
  assign y6144 = n13984 ;
  assign y6145 = ~n13853 ;
  assign y6146 = ~n13985 ;
  assign y6147 = ~n13986 ;
  assign y6148 = ~1'b0 ;
  assign y6149 = ~1'b0 ;
  assign y6150 = ~1'b0 ;
  assign y6151 = n13990 ;
  assign y6152 = ~1'b0 ;
  assign y6153 = n13998 ;
  assign y6154 = ~1'b0 ;
  assign y6155 = n14000 ;
  assign y6156 = n14004 ;
  assign y6157 = ~1'b0 ;
  assign y6158 = ~n14009 ;
  assign y6159 = ~1'b0 ;
  assign y6160 = ~n14011 ;
  assign y6161 = ~n14013 ;
  assign y6162 = ~n14018 ;
  assign y6163 = ~n14021 ;
  assign y6164 = ~n14022 ;
  assign y6165 = ~n14024 ;
  assign y6166 = ~n14026 ;
  assign y6167 = n14027 ;
  assign y6168 = ~n14029 ;
  assign y6169 = n11100 ;
  assign y6170 = n14030 ;
  assign y6171 = ~n8587 ;
  assign y6172 = 1'b0 ;
  assign y6173 = n14034 ;
  assign y6174 = ~n3411 ;
  assign y6175 = ~n14036 ;
  assign y6176 = n14037 ;
  assign y6177 = n14041 ;
  assign y6178 = n14042 ;
  assign y6179 = 1'b0 ;
  assign y6180 = ~n14043 ;
  assign y6181 = ~1'b0 ;
  assign y6182 = n14044 ;
  assign y6183 = ~n14047 ;
  assign y6184 = ~1'b0 ;
  assign y6185 = ~1'b0 ;
  assign y6186 = n14050 ;
  assign y6187 = ~n6468 ;
  assign y6188 = ~n14066 ;
  assign y6189 = ~n14067 ;
  assign y6190 = ~n14068 ;
  assign y6191 = n14078 ;
  assign y6192 = ~1'b0 ;
  assign y6193 = n10284 ;
  assign y6194 = n14079 ;
  assign y6195 = ~n14084 ;
  assign y6196 = ~n14087 ;
  assign y6197 = n14091 ;
  assign y6198 = n14093 ;
  assign y6199 = n14095 ;
  assign y6200 = n14100 ;
  assign y6201 = ~1'b0 ;
  assign y6202 = ~n14101 ;
  assign y6203 = ~1'b0 ;
  assign y6204 = n14110 ;
  assign y6205 = n14111 ;
  assign y6206 = ~n14112 ;
  assign y6207 = ~1'b0 ;
  assign y6208 = ~1'b0 ;
  assign y6209 = n14113 ;
  assign y6210 = n14114 ;
  assign y6211 = ~1'b0 ;
  assign y6212 = ~n14115 ;
  assign y6213 = n14120 ;
  assign y6214 = ~1'b0 ;
  assign y6215 = ~1'b0 ;
  assign y6216 = ~n14121 ;
  assign y6217 = ~n2779 ;
  assign y6218 = n14123 ;
  assign y6219 = ~1'b0 ;
  assign y6220 = n14125 ;
  assign y6221 = ~n14127 ;
  assign y6222 = n14131 ;
  assign y6223 = n14136 ;
  assign y6224 = ~1'b0 ;
  assign y6225 = ~1'b0 ;
  assign y6226 = ~x91 ;
  assign y6227 = n14137 ;
  assign y6228 = ~1'b0 ;
  assign y6229 = n14138 ;
  assign y6230 = ~n14140 ;
  assign y6231 = ~n14141 ;
  assign y6232 = ~1'b0 ;
  assign y6233 = n14149 ;
  assign y6234 = n14150 ;
  assign y6235 = ~n14156 ;
  assign y6236 = ~n14159 ;
  assign y6237 = ~1'b0 ;
  assign y6238 = ~n14162 ;
  assign y6239 = ~n14165 ;
  assign y6240 = n14167 ;
  assign y6241 = n14171 ;
  assign y6242 = ~n14173 ;
  assign y6243 = ~n14174 ;
  assign y6244 = ~n14176 ;
  assign y6245 = n14180 ;
  assign y6246 = n14184 ;
  assign y6247 = n14191 ;
  assign y6248 = ~n14193 ;
  assign y6249 = n14194 ;
  assign y6250 = n14195 ;
  assign y6251 = n14197 ;
  assign y6252 = n14202 ;
  assign y6253 = ~n14205 ;
  assign y6254 = n14208 ;
  assign y6255 = n14210 ;
  assign y6256 = n14211 ;
  assign y6257 = n14213 ;
  assign y6258 = ~1'b0 ;
  assign y6259 = ~n14214 ;
  assign y6260 = n14215 ;
  assign y6261 = n14218 ;
  assign y6262 = ~1'b0 ;
  assign y6263 = ~n14219 ;
  assign y6264 = n14220 ;
  assign y6265 = ~n14224 ;
  assign y6266 = n14227 ;
  assign y6267 = ~1'b0 ;
  assign y6268 = ~n14228 ;
  assign y6269 = ~n12664 ;
  assign y6270 = ~n14230 ;
  assign y6271 = ~n14231 ;
  assign y6272 = n14233 ;
  assign y6273 = ~1'b0 ;
  assign y6274 = 1'b0 ;
  assign y6275 = ~1'b0 ;
  assign y6276 = n14236 ;
  assign y6277 = ~1'b0 ;
  assign y6278 = ~1'b0 ;
  assign y6279 = ~n14243 ;
  assign y6280 = ~1'b0 ;
  assign y6281 = ~n14244 ;
  assign y6282 = n14251 ;
  assign y6283 = ~n14255 ;
  assign y6284 = ~n14258 ;
  assign y6285 = ~1'b0 ;
  assign y6286 = ~n14260 ;
  assign y6287 = ~1'b0 ;
  assign y6288 = ~n14261 ;
  assign y6289 = ~1'b0 ;
  assign y6290 = ~1'b0 ;
  assign y6291 = n14270 ;
  assign y6292 = ~n14271 ;
  assign y6293 = n14275 ;
  assign y6294 = ~n14278 ;
  assign y6295 = n14281 ;
  assign y6296 = ~1'b0 ;
  assign y6297 = n14283 ;
  assign y6298 = ~n12575 ;
  assign y6299 = n14286 ;
  assign y6300 = n14290 ;
  assign y6301 = n14291 ;
  assign y6302 = ~1'b0 ;
  assign y6303 = ~1'b0 ;
  assign y6304 = n14296 ;
  assign y6305 = n14298 ;
  assign y6306 = ~1'b0 ;
  assign y6307 = n14299 ;
  assign y6308 = ~n14300 ;
  assign y6309 = n14302 ;
  assign y6310 = ~1'b0 ;
  assign y6311 = ~n14306 ;
  assign y6312 = ~1'b0 ;
  assign y6313 = n14313 ;
  assign y6314 = ~n14318 ;
  assign y6315 = ~n14319 ;
  assign y6316 = ~n14320 ;
  assign y6317 = ~1'b0 ;
  assign y6318 = ~n14325 ;
  assign y6319 = ~1'b0 ;
  assign y6320 = ~n8040 ;
  assign y6321 = n14327 ;
  assign y6322 = ~n14330 ;
  assign y6323 = ~n14336 ;
  assign y6324 = ~n14345 ;
  assign y6325 = n14346 ;
  assign y6326 = ~n2243 ;
  assign y6327 = ~1'b0 ;
  assign y6328 = n14351 ;
  assign y6329 = n14357 ;
  assign y6330 = n7311 ;
  assign y6331 = n14360 ;
  assign y6332 = n14361 ;
  assign y6333 = ~1'b0 ;
  assign y6334 = ~n14362 ;
  assign y6335 = ~n4084 ;
  assign y6336 = n14364 ;
  assign y6337 = n14366 ;
  assign y6338 = n14367 ;
  assign y6339 = ~1'b0 ;
  assign y6340 = ~1'b0 ;
  assign y6341 = n14369 ;
  assign y6342 = ~1'b0 ;
  assign y6343 = n14370 ;
  assign y6344 = ~n229 ;
  assign y6345 = ~n14379 ;
  assign y6346 = ~n8664 ;
  assign y6347 = ~n14383 ;
  assign y6348 = ~1'b0 ;
  assign y6349 = ~1'b0 ;
  assign y6350 = ~n14389 ;
  assign y6351 = ~1'b0 ;
  assign y6352 = n14392 ;
  assign y6353 = ~n14399 ;
  assign y6354 = n14402 ;
  assign y6355 = ~n14409 ;
  assign y6356 = n14414 ;
  assign y6357 = n14416 ;
  assign y6358 = n14420 ;
  assign y6359 = ~n14421 ;
  assign y6360 = 1'b0 ;
  assign y6361 = n14423 ;
  assign y6362 = n14424 ;
  assign y6363 = ~n14427 ;
  assign y6364 = ~1'b0 ;
  assign y6365 = n14429 ;
  assign y6366 = n14432 ;
  assign y6367 = n14435 ;
  assign y6368 = ~n2623 ;
  assign y6369 = ~1'b0 ;
  assign y6370 = n9821 ;
  assign y6371 = ~1'b0 ;
  assign y6372 = n14442 ;
  assign y6373 = ~n14444 ;
  assign y6374 = ~1'b0 ;
  assign y6375 = n14445 ;
  assign y6376 = n1205 ;
  assign y6377 = ~x40 ;
  assign y6378 = ~1'b0 ;
  assign y6379 = n14449 ;
  assign y6380 = ~1'b0 ;
  assign y6381 = ~1'b0 ;
  assign y6382 = ~n14452 ;
  assign y6383 = n14459 ;
  assign y6384 = ~n14460 ;
  assign y6385 = n14464 ;
  assign y6386 = 1'b0 ;
  assign y6387 = ~n14215 ;
  assign y6388 = n14466 ;
  assign y6389 = n14467 ;
  assign y6390 = ~n14468 ;
  assign y6391 = n14469 ;
  assign y6392 = n14485 ;
  assign y6393 = ~n319 ;
  assign y6394 = ~1'b0 ;
  assign y6395 = n14489 ;
  assign y6396 = ~1'b0 ;
  assign y6397 = ~n14491 ;
  assign y6398 = n14492 ;
  assign y6399 = n14497 ;
  assign y6400 = 1'b0 ;
  assign y6401 = n14499 ;
  assign y6402 = n14500 ;
  assign y6403 = ~1'b0 ;
  assign y6404 = ~n14502 ;
  assign y6405 = n14505 ;
  assign y6406 = n14512 ;
  assign y6407 = 1'b0 ;
  assign y6408 = n14514 ;
  assign y6409 = ~n14516 ;
  assign y6410 = ~1'b0 ;
  assign y6411 = n14518 ;
  assign y6412 = ~n14524 ;
  assign y6413 = ~n14525 ;
  assign y6414 = ~1'b0 ;
  assign y6415 = n14528 ;
  assign y6416 = n14530 ;
  assign y6417 = ~n14531 ;
  assign y6418 = n14539 ;
  assign y6419 = ~1'b0 ;
  assign y6420 = n14540 ;
  assign y6421 = ~n14542 ;
  assign y6422 = ~n8900 ;
  assign y6423 = ~1'b0 ;
  assign y6424 = ~1'b0 ;
  assign y6425 = n14543 ;
  assign y6426 = ~n14544 ;
  assign y6427 = n14545 ;
  assign y6428 = ~1'b0 ;
  assign y6429 = ~1'b0 ;
  assign y6430 = ~n10341 ;
  assign y6431 = n14547 ;
  assign y6432 = ~n14548 ;
  assign y6433 = ~n14554 ;
  assign y6434 = n14555 ;
  assign y6435 = ~n14559 ;
  assign y6436 = ~1'b0 ;
  assign y6437 = ~1'b0 ;
  assign y6438 = ~n14561 ;
  assign y6439 = n14563 ;
  assign y6440 = ~n14564 ;
  assign y6441 = ~n14565 ;
  assign y6442 = ~n14569 ;
  assign y6443 = ~n14570 ;
  assign y6444 = n14574 ;
  assign y6445 = n14576 ;
  assign y6446 = 1'b0 ;
  assign y6447 = n14577 ;
  assign y6448 = ~n14579 ;
  assign y6449 = ~1'b0 ;
  assign y6450 = n14581 ;
  assign y6451 = ~1'b0 ;
  assign y6452 = ~1'b0 ;
  assign y6453 = ~n13659 ;
  assign y6454 = n14583 ;
  assign y6455 = ~n14585 ;
  assign y6456 = ~1'b0 ;
  assign y6457 = n14591 ;
  assign y6458 = ~1'b0 ;
  assign y6459 = n14595 ;
  assign y6460 = n14597 ;
  assign y6461 = ~n14598 ;
  assign y6462 = ~n14599 ;
  assign y6463 = ~n14606 ;
  assign y6464 = ~n14615 ;
  assign y6465 = ~n14617 ;
  assign y6466 = n14620 ;
  assign y6467 = ~n14621 ;
  assign y6468 = n14622 ;
  assign y6469 = ~1'b0 ;
  assign y6470 = ~n14629 ;
  assign y6471 = n14633 ;
  assign y6472 = n14634 ;
  assign y6473 = n14635 ;
  assign y6474 = ~1'b0 ;
  assign y6475 = ~n14644 ;
  assign y6476 = n14645 ;
  assign y6477 = ~n14647 ;
  assign y6478 = ~1'b0 ;
  assign y6479 = ~n14650 ;
  assign y6480 = n14653 ;
  assign y6481 = n14654 ;
  assign y6482 = n14655 ;
  assign y6483 = n14657 ;
  assign y6484 = ~1'b0 ;
  assign y6485 = n14661 ;
  assign y6486 = ~n14662 ;
  assign y6487 = ~n14664 ;
  assign y6488 = ~n14666 ;
  assign y6489 = ~1'b0 ;
  assign y6490 = ~1'b0 ;
  assign y6491 = ~n14667 ;
  assign y6492 = ~n14670 ;
  assign y6493 = ~n14677 ;
  assign y6494 = ~1'b0 ;
  assign y6495 = n14678 ;
  assign y6496 = n14684 ;
  assign y6497 = ~1'b0 ;
  assign y6498 = ~n14686 ;
  assign y6499 = n14688 ;
  assign y6500 = ~1'b0 ;
  assign y6501 = n14689 ;
  assign y6502 = n14691 ;
  assign y6503 = n14692 ;
  assign y6504 = ~1'b0 ;
  assign y6505 = n14693 ;
  assign y6506 = n14694 ;
  assign y6507 = ~n14699 ;
  assign y6508 = n14702 ;
  assign y6509 = ~1'b0 ;
  assign y6510 = ~n14703 ;
  assign y6511 = ~n14706 ;
  assign y6512 = ~n14709 ;
  assign y6513 = ~n14711 ;
  assign y6514 = n14713 ;
  assign y6515 = n14717 ;
  assign y6516 = n14722 ;
  assign y6517 = n14724 ;
  assign y6518 = 1'b0 ;
  assign y6519 = ~1'b0 ;
  assign y6520 = n14730 ;
  assign y6521 = ~1'b0 ;
  assign y6522 = n14731 ;
  assign y6523 = ~n14734 ;
  assign y6524 = ~1'b0 ;
  assign y6525 = ~n14735 ;
  assign y6526 = n1581 ;
  assign y6527 = ~n14736 ;
  assign y6528 = ~n14740 ;
  assign y6529 = ~n14741 ;
  assign y6530 = n14742 ;
  assign y6531 = ~1'b0 ;
  assign y6532 = n14743 ;
  assign y6533 = ~n11940 ;
  assign y6534 = ~1'b0 ;
  assign y6535 = ~1'b0 ;
  assign y6536 = ~n14748 ;
  assign y6537 = ~n14754 ;
  assign y6538 = ~1'b0 ;
  assign y6539 = n14756 ;
  assign y6540 = ~1'b0 ;
  assign y6541 = ~n14757 ;
  assign y6542 = n14759 ;
  assign y6543 = n14760 ;
  assign y6544 = ~n14761 ;
  assign y6545 = ~n14762 ;
  assign y6546 = ~n14764 ;
  assign y6547 = ~1'b0 ;
  assign y6548 = n9413 ;
  assign y6549 = ~n10327 ;
  assign y6550 = n14767 ;
  assign y6551 = n14768 ;
  assign y6552 = n14769 ;
  assign y6553 = ~n14775 ;
  assign y6554 = ~n14778 ;
  assign y6555 = ~1'b0 ;
  assign y6556 = ~1'b0 ;
  assign y6557 = n1506 ;
  assign y6558 = n14779 ;
  assign y6559 = ~n14786 ;
  assign y6560 = ~n14791 ;
  assign y6561 = n14797 ;
  assign y6562 = n14800 ;
  assign y6563 = 1'b0 ;
  assign y6564 = n14803 ;
  assign y6565 = n12631 ;
  assign y6566 = ~1'b0 ;
  assign y6567 = ~n14805 ;
  assign y6568 = ~n14811 ;
  assign y6569 = n14814 ;
  assign y6570 = n14815 ;
  assign y6571 = ~1'b0 ;
  assign y6572 = ~1'b0 ;
  assign y6573 = n14817 ;
  assign y6574 = n14818 ;
  assign y6575 = n14823 ;
  assign y6576 = ~n14825 ;
  assign y6577 = n14830 ;
  assign y6578 = ~n14833 ;
  assign y6579 = ~1'b0 ;
  assign y6580 = ~n8445 ;
  assign y6581 = ~1'b0 ;
  assign y6582 = ~1'b0 ;
  assign y6583 = n14840 ;
  assign y6584 = ~n14843 ;
  assign y6585 = ~n14845 ;
  assign y6586 = ~1'b0 ;
  assign y6587 = n14848 ;
  assign y6588 = n14850 ;
  assign y6589 = ~n14851 ;
  assign y6590 = ~n14854 ;
  assign y6591 = ~n14856 ;
  assign y6592 = ~n14857 ;
  assign y6593 = ~n14858 ;
  assign y6594 = n14859 ;
  assign y6595 = n14860 ;
  assign y6596 = ~n14862 ;
  assign y6597 = ~1'b0 ;
  assign y6598 = n14866 ;
  assign y6599 = ~1'b0 ;
  assign y6600 = ~1'b0 ;
  assign y6601 = n14867 ;
  assign y6602 = ~n14868 ;
  assign y6603 = ~n14869 ;
  assign y6604 = ~1'b0 ;
  assign y6605 = n14871 ;
  assign y6606 = ~1'b0 ;
  assign y6607 = ~n14874 ;
  assign y6608 = n14882 ;
  assign y6609 = ~n14884 ;
  assign y6610 = ~n14887 ;
  assign y6611 = ~1'b0 ;
  assign y6612 = ~n14888 ;
  assign y6613 = n14891 ;
  assign y6614 = ~n6698 ;
  assign y6615 = ~1'b0 ;
  assign y6616 = ~n14893 ;
  assign y6617 = n14898 ;
  assign y6618 = n14903 ;
  assign y6619 = ~1'b0 ;
  assign y6620 = ~1'b0 ;
  assign y6621 = ~1'b0 ;
  assign y6622 = ~1'b0 ;
  assign y6623 = n14905 ;
  assign y6624 = ~n14909 ;
  assign y6625 = ~n14917 ;
  assign y6626 = n14919 ;
  assign y6627 = ~1'b0 ;
  assign y6628 = ~n14922 ;
  assign y6629 = ~n14923 ;
  assign y6630 = ~1'b0 ;
  assign y6631 = n14927 ;
  assign y6632 = n14932 ;
  assign y6633 = ~n14935 ;
  assign y6634 = ~n14938 ;
  assign y6635 = ~1'b0 ;
  assign y6636 = ~n14939 ;
  assign y6637 = n14942 ;
  assign y6638 = ~n14944 ;
  assign y6639 = ~1'b0 ;
  assign y6640 = ~n14948 ;
  assign y6641 = ~n14949 ;
  assign y6642 = ~1'b0 ;
  assign y6643 = ~1'b0 ;
  assign y6644 = n14950 ;
  assign y6645 = ~n14956 ;
  assign y6646 = n14957 ;
  assign y6647 = ~1'b0 ;
  assign y6648 = n14959 ;
  assign y6649 = ~n14962 ;
  assign y6650 = n14963 ;
  assign y6651 = ~n14964 ;
  assign y6652 = n14965 ;
  assign y6653 = n13216 ;
  assign y6654 = ~n14971 ;
  assign y6655 = ~n14974 ;
  assign y6656 = ~n14983 ;
  assign y6657 = n14984 ;
  assign y6658 = ~n6463 ;
  assign y6659 = n14985 ;
  assign y6660 = ~n14986 ;
  assign y6661 = n14988 ;
  assign y6662 = n14991 ;
  assign y6663 = ~n14995 ;
  assign y6664 = ~n14999 ;
  assign y6665 = n15000 ;
  assign y6666 = ~1'b0 ;
  assign y6667 = ~n15004 ;
  assign y6668 = ~1'b0 ;
  assign y6669 = ~1'b0 ;
  assign y6670 = ~1'b0 ;
  assign y6671 = n15005 ;
  assign y6672 = ~n15010 ;
  assign y6673 = ~1'b0 ;
  assign y6674 = n15020 ;
  assign y6675 = ~1'b0 ;
  assign y6676 = ~n15021 ;
  assign y6677 = ~1'b0 ;
  assign y6678 = n918 ;
  assign y6679 = ~n15023 ;
  assign y6680 = ~n9131 ;
  assign y6681 = ~n15028 ;
  assign y6682 = ~1'b0 ;
  assign y6683 = n15032 ;
  assign y6684 = ~n2444 ;
  assign y6685 = ~n15036 ;
  assign y6686 = n15040 ;
  assign y6687 = ~1'b0 ;
  assign y6688 = ~n15046 ;
  assign y6689 = ~n15047 ;
  assign y6690 = ~1'b0 ;
  assign y6691 = ~n15052 ;
  assign y6692 = ~n15053 ;
  assign y6693 = n15054 ;
  assign y6694 = ~n15055 ;
  assign y6695 = ~1'b0 ;
  assign y6696 = ~1'b0 ;
  assign y6697 = ~1'b0 ;
  assign y6698 = ~n15056 ;
  assign y6699 = ~n15057 ;
  assign y6700 = n15060 ;
  assign y6701 = ~n15062 ;
  assign y6702 = ~1'b0 ;
  assign y6703 = n15067 ;
  assign y6704 = ~1'b0 ;
  assign y6705 = n15068 ;
  assign y6706 = ~n15069 ;
  assign y6707 = ~n15073 ;
  assign y6708 = ~1'b0 ;
  assign y6709 = ~n15075 ;
  assign y6710 = ~n15078 ;
  assign y6711 = ~n15085 ;
  assign y6712 = n15087 ;
  assign y6713 = n15088 ;
  assign y6714 = ~n15090 ;
  assign y6715 = ~n15092 ;
  assign y6716 = n15094 ;
  assign y6717 = ~n15097 ;
  assign y6718 = ~1'b0 ;
  assign y6719 = n15098 ;
  assign y6720 = ~1'b0 ;
  assign y6721 = n3497 ;
  assign y6722 = ~1'b0 ;
  assign y6723 = n15100 ;
  assign y6724 = ~n15102 ;
  assign y6725 = ~1'b0 ;
  assign y6726 = ~1'b0 ;
  assign y6727 = n2369 ;
  assign y6728 = n15103 ;
  assign y6729 = n15105 ;
  assign y6730 = ~1'b0 ;
  assign y6731 = ~n15110 ;
  assign y6732 = n15111 ;
  assign y6733 = n15113 ;
  assign y6734 = n15120 ;
  assign y6735 = ~n15122 ;
  assign y6736 = ~n15126 ;
  assign y6737 = ~n15128 ;
  assign y6738 = n15129 ;
  assign y6739 = ~n15130 ;
  assign y6740 = ~n15131 ;
  assign y6741 = ~n15134 ;
  assign y6742 = ~n15136 ;
  assign y6743 = ~1'b0 ;
  assign y6744 = ~n7726 ;
  assign y6745 = ~n15138 ;
  assign y6746 = ~n15140 ;
  assign y6747 = ~1'b0 ;
  assign y6748 = n15141 ;
  assign y6749 = ~1'b0 ;
  assign y6750 = ~1'b0 ;
  assign y6751 = ~n15143 ;
  assign y6752 = ~n6114 ;
  assign y6753 = ~1'b0 ;
  assign y6754 = ~n15145 ;
  assign y6755 = n15146 ;
  assign y6756 = n15147 ;
  assign y6757 = ~n15153 ;
  assign y6758 = ~n15154 ;
  assign y6759 = ~1'b0 ;
  assign y6760 = n15156 ;
  assign y6761 = n15158 ;
  assign y6762 = n15160 ;
  assign y6763 = ~n15161 ;
  assign y6764 = ~n15164 ;
  assign y6765 = n15170 ;
  assign y6766 = ~n262 ;
  assign y6767 = ~1'b0 ;
  assign y6768 = ~1'b0 ;
  assign y6769 = ~n15175 ;
  assign y6770 = n15181 ;
  assign y6771 = ~n15184 ;
  assign y6772 = n15189 ;
  assign y6773 = n15191 ;
  assign y6774 = n15196 ;
  assign y6775 = ~1'b0 ;
  assign y6776 = ~1'b0 ;
  assign y6777 = ~1'b0 ;
  assign y6778 = n15200 ;
  assign y6779 = n15205 ;
  assign y6780 = ~1'b0 ;
  assign y6781 = n15212 ;
  assign y6782 = ~n15220 ;
  assign y6783 = ~n15221 ;
  assign y6784 = ~n15222 ;
  assign y6785 = ~n15223 ;
  assign y6786 = n15225 ;
  assign y6787 = ~1'b0 ;
  assign y6788 = ~n15230 ;
  assign y6789 = ~n15232 ;
  assign y6790 = n15236 ;
  assign y6791 = ~n15239 ;
  assign y6792 = ~n15240 ;
  assign y6793 = n15244 ;
  assign y6794 = ~1'b0 ;
  assign y6795 = ~n15245 ;
  assign y6796 = ~n15246 ;
  assign y6797 = ~n15249 ;
  assign y6798 = ~n15250 ;
  assign y6799 = ~1'b0 ;
  assign y6800 = ~1'b0 ;
  assign y6801 = n15255 ;
  assign y6802 = ~n15257 ;
  assign y6803 = n15264 ;
  assign y6804 = ~n15265 ;
  assign y6805 = n15269 ;
  assign y6806 = ~1'b0 ;
  assign y6807 = n15277 ;
  assign y6808 = n7874 ;
  assign y6809 = ~1'b0 ;
  assign y6810 = ~1'b0 ;
  assign y6811 = n8545 ;
  assign y6812 = ~1'b0 ;
  assign y6813 = ~n15279 ;
  assign y6814 = ~n15280 ;
  assign y6815 = ~n15281 ;
  assign y6816 = n15283 ;
  assign y6817 = ~n15287 ;
  assign y6818 = ~n15291 ;
  assign y6819 = 1'b0 ;
  assign y6820 = ~n13058 ;
  assign y6821 = n15292 ;
  assign y6822 = ~n15294 ;
  assign y6823 = ~n15299 ;
  assign y6824 = ~1'b0 ;
  assign y6825 = ~n15301 ;
  assign y6826 = ~1'b0 ;
  assign y6827 = ~n15305 ;
  assign y6828 = ~1'b0 ;
  assign y6829 = n15307 ;
  assign y6830 = n15308 ;
  assign y6831 = n15309 ;
  assign y6832 = ~n15316 ;
  assign y6833 = n15318 ;
  assign y6834 = ~n15321 ;
  assign y6835 = n15328 ;
  assign y6836 = ~1'b0 ;
  assign y6837 = n15329 ;
  assign y6838 = n15330 ;
  assign y6839 = n15334 ;
  assign y6840 = ~1'b0 ;
  assign y6841 = 1'b0 ;
  assign y6842 = ~n15338 ;
  assign y6843 = ~1'b0 ;
  assign y6844 = ~n15339 ;
  assign y6845 = n15341 ;
  assign y6846 = n15343 ;
  assign y6847 = n15354 ;
  assign y6848 = ~1'b0 ;
  assign y6849 = ~1'b0 ;
  assign y6850 = ~1'b0 ;
  assign y6851 = ~n15355 ;
  assign y6852 = n15357 ;
  assign y6853 = ~n15358 ;
  assign y6854 = ~n15359 ;
  assign y6855 = n15360 ;
  assign y6856 = ~n15366 ;
  assign y6857 = 1'b0 ;
  assign y6858 = ~1'b0 ;
  assign y6859 = n15367 ;
  assign y6860 = ~n14729 ;
  assign y6861 = n15369 ;
  assign y6862 = ~n15372 ;
  assign y6863 = n15376 ;
  assign y6864 = ~1'b0 ;
  assign y6865 = ~1'b0 ;
  assign y6866 = ~n15378 ;
  assign y6867 = ~1'b0 ;
  assign y6868 = ~n3035 ;
  assign y6869 = ~n15379 ;
  assign y6870 = n15383 ;
  assign y6871 = n15388 ;
  assign y6872 = ~n15390 ;
  assign y6873 = n15392 ;
  assign y6874 = n15393 ;
  assign y6875 = n15394 ;
  assign y6876 = n6214 ;
  assign y6877 = ~n15395 ;
  assign y6878 = n15396 ;
  assign y6879 = 1'b0 ;
  assign y6880 = n15399 ;
  assign y6881 = ~n15406 ;
  assign y6882 = n15407 ;
  assign y6883 = ~n15410 ;
  assign y6884 = ~n15412 ;
  assign y6885 = ~1'b0 ;
  assign y6886 = ~n15415 ;
  assign y6887 = n15416 ;
  assign y6888 = ~1'b0 ;
  assign y6889 = n15431 ;
  assign y6890 = n15436 ;
  assign y6891 = n15437 ;
  assign y6892 = ~n15441 ;
  assign y6893 = ~n15444 ;
  assign y6894 = n15446 ;
  assign y6895 = n15332 ;
  assign y6896 = n4285 ;
  assign y6897 = ~n15449 ;
  assign y6898 = ~n9273 ;
  assign y6899 = n15451 ;
  assign y6900 = ~n15457 ;
  assign y6901 = ~n15460 ;
  assign y6902 = n15462 ;
  assign y6903 = n15464 ;
  assign y6904 = n15467 ;
  assign y6905 = n15468 ;
  assign y6906 = ~1'b0 ;
  assign y6907 = ~n15471 ;
  assign y6908 = n15472 ;
  assign y6909 = ~n15473 ;
  assign y6910 = ~1'b0 ;
  assign y6911 = ~1'b0 ;
  assign y6912 = ~n15475 ;
  assign y6913 = n15476 ;
  assign y6914 = ~1'b0 ;
  assign y6915 = ~n15482 ;
  assign y6916 = ~n15484 ;
  assign y6917 = ~1'b0 ;
  assign y6918 = n15485 ;
  assign y6919 = ~1'b0 ;
  assign y6920 = ~n15490 ;
  assign y6921 = ~n15491 ;
  assign y6922 = n15492 ;
  assign y6923 = ~1'b0 ;
  assign y6924 = ~n15496 ;
  assign y6925 = ~n15500 ;
  assign y6926 = n15501 ;
  assign y6927 = n15503 ;
  assign y6928 = ~n15506 ;
  assign y6929 = ~1'b0 ;
  assign y6930 = ~n15507 ;
  assign y6931 = ~n15509 ;
  assign y6932 = n15513 ;
  assign y6933 = n15514 ;
  assign y6934 = n15515 ;
  assign y6935 = n15517 ;
  assign y6936 = ~1'b0 ;
  assign y6937 = ~n15519 ;
  assign y6938 = ~1'b0 ;
  assign y6939 = n15521 ;
  assign y6940 = ~1'b0 ;
  assign y6941 = n15522 ;
  assign y6942 = n15527 ;
  assign y6943 = n15533 ;
  assign y6944 = n15535 ;
  assign y6945 = n15541 ;
  assign y6946 = 1'b0 ;
  assign y6947 = n15542 ;
  assign y6948 = ~n15543 ;
  assign y6949 = n15545 ;
  assign y6950 = ~1'b0 ;
  assign y6951 = ~1'b0 ;
  assign y6952 = n15546 ;
  assign y6953 = n7206 ;
  assign y6954 = ~n15547 ;
  assign y6955 = ~n15552 ;
  assign y6956 = ~n10248 ;
  assign y6957 = ~1'b0 ;
  assign y6958 = ~n15556 ;
  assign y6959 = ~n15558 ;
  assign y6960 = ~n15560 ;
  assign y6961 = ~1'b0 ;
  assign y6962 = n15563 ;
  assign y6963 = ~n15571 ;
  assign y6964 = ~n15572 ;
  assign y6965 = ~n15573 ;
  assign y6966 = ~n15575 ;
  assign y6967 = ~n15576 ;
  assign y6968 = ~1'b0 ;
  assign y6969 = ~1'b0 ;
  assign y6970 = ~n15578 ;
  assign y6971 = ~n15584 ;
  assign y6972 = ~n12265 ;
  assign y6973 = ~1'b0 ;
  assign y6974 = n15589 ;
  assign y6975 = ~n15594 ;
  assign y6976 = ~1'b0 ;
  assign y6977 = ~1'b0 ;
  assign y6978 = ~1'b0 ;
  assign y6979 = ~n15597 ;
  assign y6980 = n15598 ;
  assign y6981 = ~1'b0 ;
  assign y6982 = ~n15602 ;
  assign y6983 = n15607 ;
  assign y6984 = ~1'b0 ;
  assign y6985 = n15613 ;
  assign y6986 = ~1'b0 ;
  assign y6987 = ~n15615 ;
  assign y6988 = n15617 ;
  assign y6989 = n15623 ;
  assign y6990 = ~n15625 ;
  assign y6991 = ~n15627 ;
  assign y6992 = n15628 ;
  assign y6993 = n15630 ;
  assign y6994 = ~n15538 ;
  assign y6995 = ~1'b0 ;
  assign y6996 = ~n15636 ;
  assign y6997 = ~n3304 ;
  assign y6998 = n15639 ;
  assign y6999 = n15641 ;
  assign y7000 = n15643 ;
  assign y7001 = ~1'b0 ;
  assign y7002 = ~1'b0 ;
  assign y7003 = ~1'b0 ;
  assign y7004 = ~n15648 ;
  assign y7005 = ~n15649 ;
  assign y7006 = ~n15657 ;
  assign y7007 = n15660 ;
  assign y7008 = n15661 ;
  assign y7009 = ~1'b0 ;
  assign y7010 = ~1'b0 ;
  assign y7011 = n15662 ;
  assign y7012 = ~n15666 ;
  assign y7013 = ~n15676 ;
  assign y7014 = n15685 ;
  assign y7015 = ~1'b0 ;
  assign y7016 = ~n15686 ;
  assign y7017 = ~1'b0 ;
  assign y7018 = n15687 ;
  assign y7019 = ~1'b0 ;
  assign y7020 = ~1'b0 ;
  assign y7021 = ~1'b0 ;
  assign y7022 = ~1'b0 ;
  assign y7023 = ~n4824 ;
  assign y7024 = ~n15689 ;
  assign y7025 = ~n15691 ;
  assign y7026 = ~n15693 ;
  assign y7027 = ~1'b0 ;
  assign y7028 = ~n15696 ;
  assign y7029 = n15698 ;
  assign y7030 = ~n15700 ;
  assign y7031 = n15702 ;
  assign y7032 = ~n15709 ;
  assign y7033 = n15717 ;
  assign y7034 = n15720 ;
  assign y7035 = n15723 ;
  assign y7036 = n15732 ;
  assign y7037 = n15733 ;
  assign y7038 = ~n15736 ;
  assign y7039 = ~1'b0 ;
  assign y7040 = ~1'b0 ;
  assign y7041 = ~n15738 ;
  assign y7042 = n15749 ;
  assign y7043 = n15750 ;
  assign y7044 = ~n15752 ;
  assign y7045 = n15756 ;
  assign y7046 = ~n15757 ;
  assign y7047 = n15760 ;
  assign y7048 = n15761 ;
  assign y7049 = ~n15763 ;
  assign y7050 = n15764 ;
  assign y7051 = 1'b0 ;
  assign y7052 = ~n15765 ;
  assign y7053 = ~1'b0 ;
  assign y7054 = ~n2419 ;
  assign y7055 = ~1'b0 ;
  assign y7056 = ~n15771 ;
  assign y7057 = n15774 ;
  assign y7058 = n15775 ;
  assign y7059 = ~n15781 ;
  assign y7060 = n15789 ;
  assign y7061 = ~n15790 ;
  assign y7062 = ~n15798 ;
  assign y7063 = ~1'b0 ;
  assign y7064 = n15800 ;
  assign y7065 = ~n15804 ;
  assign y7066 = ~1'b0 ;
  assign y7067 = n15806 ;
  assign y7068 = ~n15808 ;
  assign y7069 = n15810 ;
  assign y7070 = n15814 ;
  assign y7071 = n15818 ;
  assign y7072 = n15819 ;
  assign y7073 = n15821 ;
  assign y7074 = n15823 ;
  assign y7075 = n15830 ;
  assign y7076 = ~1'b0 ;
  assign y7077 = ~n15833 ;
  assign y7078 = ~n15839 ;
  assign y7079 = n5278 ;
  assign y7080 = ~n1660 ;
  assign y7081 = ~n15841 ;
  assign y7082 = ~1'b0 ;
  assign y7083 = n15845 ;
  assign y7084 = ~n15850 ;
  assign y7085 = ~1'b0 ;
  assign y7086 = n15852 ;
  assign y7087 = ~n15858 ;
  assign y7088 = ~n15859 ;
  assign y7089 = ~n15863 ;
  assign y7090 = n15865 ;
  assign y7091 = n15869 ;
  assign y7092 = ~n15870 ;
  assign y7093 = n15872 ;
  assign y7094 = ~n15873 ;
  assign y7095 = ~n15875 ;
  assign y7096 = ~1'b0 ;
  assign y7097 = n11926 ;
  assign y7098 = ~n15878 ;
  assign y7099 = ~n15882 ;
  assign y7100 = ~1'b0 ;
  assign y7101 = ~n15884 ;
  assign y7102 = ~n14034 ;
  assign y7103 = n15885 ;
  assign y7104 = ~n15886 ;
  assign y7105 = n15890 ;
  assign y7106 = n15894 ;
  assign y7107 = n9305 ;
  assign y7108 = ~n15896 ;
  assign y7109 = ~1'b0 ;
  assign y7110 = n6506 ;
  assign y7111 = ~n15902 ;
  assign y7112 = ~1'b0 ;
  assign y7113 = ~1'b0 ;
  assign y7114 = ~n15903 ;
  assign y7115 = n15906 ;
  assign y7116 = ~1'b0 ;
  assign y7117 = n15909 ;
  assign y7118 = n15914 ;
  assign y7119 = n15922 ;
  assign y7120 = ~n15923 ;
  assign y7121 = n15928 ;
  assign y7122 = ~n15931 ;
  assign y7123 = n15933 ;
  assign y7124 = n7446 ;
  assign y7125 = ~n2741 ;
  assign y7126 = ~n15940 ;
  assign y7127 = ~1'b0 ;
  assign y7128 = ~n15941 ;
  assign y7129 = ~n15943 ;
  assign y7130 = n15945 ;
  assign y7131 = ~1'b0 ;
  assign y7132 = ~1'b0 ;
  assign y7133 = n9008 ;
  assign y7134 = ~n15950 ;
  assign y7135 = n15951 ;
  assign y7136 = ~n15957 ;
  assign y7137 = ~n15960 ;
  assign y7138 = ~n13548 ;
  assign y7139 = n15963 ;
  assign y7140 = ~1'b0 ;
  assign y7141 = ~n15966 ;
  assign y7142 = n15971 ;
  assign y7143 = n15974 ;
  assign y7144 = ~1'b0 ;
  assign y7145 = n15975 ;
  assign y7146 = ~n15979 ;
  assign y7147 = ~n15981 ;
  assign y7148 = n15982 ;
  assign y7149 = n15984 ;
  assign y7150 = ~n15986 ;
  assign y7151 = n15996 ;
  assign y7152 = ~n15999 ;
  assign y7153 = n16001 ;
  assign y7154 = n16007 ;
  assign y7155 = n16009 ;
  assign y7156 = n16010 ;
  assign y7157 = ~n16016 ;
  assign y7158 = ~n16018 ;
  assign y7159 = ~n16020 ;
  assign y7160 = n16021 ;
  assign y7161 = ~1'b0 ;
  assign y7162 = n16023 ;
  assign y7163 = n16028 ;
  assign y7164 = n16030 ;
  assign y7165 = n16032 ;
  assign y7166 = ~n16036 ;
  assign y7167 = ~n16037 ;
  assign y7168 = ~n16038 ;
  assign y7169 = ~n16040 ;
  assign y7170 = n16041 ;
  assign y7171 = ~n16044 ;
  assign y7172 = ~n3491 ;
  assign y7173 = ~n16048 ;
  assign y7174 = n16051 ;
  assign y7175 = ~n16059 ;
  assign y7176 = ~1'b0 ;
  assign y7177 = n12109 ;
  assign y7178 = n16061 ;
  assign y7179 = ~1'b0 ;
  assign y7180 = ~n16068 ;
  assign y7181 = ~n15634 ;
  assign y7182 = n16069 ;
  assign y7183 = n16074 ;
  assign y7184 = n16076 ;
  assign y7185 = ~1'b0 ;
  assign y7186 = ~1'b0 ;
  assign y7187 = n16078 ;
  assign y7188 = n16081 ;
  assign y7189 = n4690 ;
  assign y7190 = ~1'b0 ;
  assign y7191 = n16087 ;
  assign y7192 = ~n16089 ;
  assign y7193 = ~1'b0 ;
  assign y7194 = ~n16091 ;
  assign y7195 = n16092 ;
  assign y7196 = ~1'b0 ;
  assign y7197 = ~n16093 ;
  assign y7198 = ~n16094 ;
  assign y7199 = ~n16098 ;
  assign y7200 = ~n16099 ;
  assign y7201 = ~n16100 ;
  assign y7202 = ~n16101 ;
  assign y7203 = n16102 ;
  assign y7204 = ~1'b0 ;
  assign y7205 = n16104 ;
  assign y7206 = n16105 ;
  assign y7207 = ~n16107 ;
  assign y7208 = n16108 ;
  assign y7209 = n16109 ;
  assign y7210 = n16110 ;
  assign y7211 = n16113 ;
  assign y7212 = ~n16118 ;
  assign y7213 = ~1'b0 ;
  assign y7214 = ~n16128 ;
  assign y7215 = ~n10260 ;
  assign y7216 = n16132 ;
  assign y7217 = ~1'b0 ;
  assign y7218 = n16133 ;
  assign y7219 = ~n16136 ;
  assign y7220 = ~n16137 ;
  assign y7221 = n16139 ;
  assign y7222 = n16140 ;
  assign y7223 = ~1'b0 ;
  assign y7224 = n16143 ;
  assign y7225 = ~n16146 ;
  assign y7226 = n16147 ;
  assign y7227 = ~n16152 ;
  assign y7228 = ~1'b0 ;
  assign y7229 = ~n16153 ;
  assign y7230 = ~n16159 ;
  assign y7231 = n16160 ;
  assign y7232 = n16164 ;
  assign y7233 = ~1'b0 ;
  assign y7234 = ~n16166 ;
  assign y7235 = ~1'b0 ;
  assign y7236 = n16167 ;
  assign y7237 = n16168 ;
  assign y7238 = n16172 ;
  assign y7239 = n8608 ;
  assign y7240 = ~n16181 ;
  assign y7241 = ~n7622 ;
  assign y7242 = ~n7243 ;
  assign y7243 = ~n16182 ;
  assign y7244 = n16188 ;
  assign y7245 = ~1'b0 ;
  assign y7246 = n16191 ;
  assign y7247 = n16193 ;
  assign y7248 = ~n16196 ;
  assign y7249 = n16197 ;
  assign y7250 = n16200 ;
  assign y7251 = x91 ;
  assign y7252 = ~1'b0 ;
  assign y7253 = ~n16201 ;
  assign y7254 = ~n16206 ;
  assign y7255 = n16208 ;
  assign y7256 = ~n16209 ;
  assign y7257 = n16212 ;
  assign y7258 = ~n16213 ;
  assign y7259 = ~n16214 ;
  assign y7260 = ~x70 ;
  assign y7261 = ~n16217 ;
  assign y7262 = n16220 ;
  assign y7263 = n16221 ;
  assign y7264 = ~n16224 ;
  assign y7265 = n16227 ;
  assign y7266 = ~n16232 ;
  assign y7267 = ~1'b0 ;
  assign y7268 = ~1'b0 ;
  assign y7269 = ~n16233 ;
  assign y7270 = ~n16239 ;
  assign y7271 = n16240 ;
  assign y7272 = ~n492 ;
  assign y7273 = ~1'b0 ;
  assign y7274 = ~1'b0 ;
  assign y7275 = ~1'b0 ;
  assign y7276 = ~n16242 ;
  assign y7277 = ~n16243 ;
  assign y7278 = n2101 ;
  assign y7279 = ~1'b0 ;
  assign y7280 = ~1'b0 ;
  assign y7281 = ~1'b0 ;
  assign y7282 = n16246 ;
  assign y7283 = ~n16249 ;
  assign y7284 = ~n16250 ;
  assign y7285 = ~1'b0 ;
  assign y7286 = ~n16259 ;
  assign y7287 = ~1'b0 ;
  assign y7288 = ~1'b0 ;
  assign y7289 = ~n16261 ;
  assign y7290 = n16268 ;
  assign y7291 = n16270 ;
  assign y7292 = n16272 ;
  assign y7293 = n16275 ;
  assign y7294 = ~n16277 ;
  assign y7295 = n16279 ;
  assign y7296 = ~n16281 ;
  assign y7297 = n16283 ;
  assign y7298 = ~n16284 ;
  assign y7299 = ~n16287 ;
  assign y7300 = n16293 ;
  assign y7301 = n16294 ;
  assign y7302 = n16295 ;
  assign y7303 = n3254 ;
  assign y7304 = ~1'b0 ;
  assign y7305 = n5651 ;
  assign y7306 = ~1'b0 ;
  assign y7307 = n16297 ;
  assign y7308 = n16298 ;
  assign y7309 = n16299 ;
  assign y7310 = ~n16302 ;
  assign y7311 = ~n16304 ;
  assign y7312 = ~n16305 ;
  assign y7313 = n16306 ;
  assign y7314 = ~n16307 ;
  assign y7315 = n16309 ;
  assign y7316 = n16311 ;
  assign y7317 = ~n16312 ;
  assign y7318 = ~n16315 ;
  assign y7319 = n9274 ;
  assign y7320 = n16318 ;
  assign y7321 = ~1'b0 ;
  assign y7322 = ~1'b0 ;
  assign y7323 = n16319 ;
  assign y7324 = ~n16321 ;
  assign y7325 = 1'b0 ;
  assign y7326 = ~n16325 ;
  assign y7327 = n16326 ;
  assign y7328 = ~n16328 ;
  assign y7329 = n16333 ;
  assign y7330 = n16334 ;
  assign y7331 = ~n16335 ;
  assign y7332 = n16338 ;
  assign y7333 = n16340 ;
  assign y7334 = ~n16341 ;
  assign y7335 = ~1'b0 ;
  assign y7336 = ~n16346 ;
  assign y7337 = n16348 ;
  assign y7338 = n12671 ;
  assign y7339 = ~1'b0 ;
  assign y7340 = ~n4954 ;
  assign y7341 = ~n16354 ;
  assign y7342 = n16356 ;
  assign y7343 = ~n16359 ;
  assign y7344 = ~n16366 ;
  assign y7345 = n16367 ;
  assign y7346 = ~1'b0 ;
  assign y7347 = n16369 ;
  assign y7348 = 1'b0 ;
  assign y7349 = ~n16376 ;
  assign y7350 = ~1'b0 ;
  assign y7351 = ~1'b0 ;
  assign y7352 = ~n16387 ;
  assign y7353 = ~1'b0 ;
  assign y7354 = n16388 ;
  assign y7355 = n16389 ;
  assign y7356 = n362 ;
  assign y7357 = ~n16392 ;
  assign y7358 = ~n16394 ;
  assign y7359 = n5902 ;
  assign y7360 = n16395 ;
  assign y7361 = ~n16396 ;
  assign y7362 = 1'b0 ;
  assign y7363 = n16398 ;
  assign y7364 = ~1'b0 ;
  assign y7365 = ~1'b0 ;
  assign y7366 = ~n2426 ;
  assign y7367 = n16404 ;
  assign y7368 = ~1'b0 ;
  assign y7369 = ~1'b0 ;
  assign y7370 = n1582 ;
  assign y7371 = n16405 ;
  assign y7372 = ~n16406 ;
  assign y7373 = ~n16408 ;
  assign y7374 = n16412 ;
  assign y7375 = ~1'b0 ;
  assign y7376 = ~1'b0 ;
  assign y7377 = ~1'b0 ;
  assign y7378 = n16419 ;
  assign y7379 = n16423 ;
  assign y7380 = n16429 ;
  assign y7381 = ~n16436 ;
  assign y7382 = ~1'b0 ;
  assign y7383 = n16438 ;
  assign y7384 = ~1'b0 ;
  assign y7385 = n16440 ;
  assign y7386 = ~1'b0 ;
  assign y7387 = n16441 ;
  assign y7388 = ~n16445 ;
  assign y7389 = ~1'b0 ;
  assign y7390 = ~n16457 ;
  assign y7391 = ~1'b0 ;
  assign y7392 = n16458 ;
  assign y7393 = ~1'b0 ;
  assign y7394 = n16459 ;
  assign y7395 = ~n16465 ;
  assign y7396 = ~1'b0 ;
  assign y7397 = ~1'b0 ;
  assign y7398 = ~n16470 ;
  assign y7399 = n16474 ;
  assign y7400 = ~1'b0 ;
  assign y7401 = n16475 ;
  assign y7402 = ~n16477 ;
  assign y7403 = ~1'b0 ;
  assign y7404 = ~n16480 ;
  assign y7405 = ~n16482 ;
  assign y7406 = n16483 ;
  assign y7407 = ~n16484 ;
  assign y7408 = n16488 ;
  assign y7409 = n16489 ;
  assign y7410 = n16491 ;
  assign y7411 = n16493 ;
  assign y7412 = n16494 ;
  assign y7413 = ~n16495 ;
  assign y7414 = n16497 ;
  assign y7415 = ~n16502 ;
  assign y7416 = ~n16503 ;
  assign y7417 = ~n16506 ;
  assign y7418 = n16510 ;
  assign y7419 = n16515 ;
  assign y7420 = ~1'b0 ;
  assign y7421 = n16516 ;
  assign y7422 = ~n16518 ;
  assign y7423 = ~n8613 ;
  assign y7424 = 1'b0 ;
  assign y7425 = ~n16524 ;
  assign y7426 = ~1'b0 ;
  assign y7427 = n16526 ;
  assign y7428 = ~n16527 ;
  assign y7429 = ~1'b0 ;
  assign y7430 = n16531 ;
  assign y7431 = ~n16536 ;
  assign y7432 = ~n16539 ;
  assign y7433 = ~1'b0 ;
  assign y7434 = ~n16540 ;
  assign y7435 = ~n16543 ;
  assign y7436 = n16546 ;
  assign y7437 = ~1'b0 ;
  assign y7438 = ~1'b0 ;
  assign y7439 = n16549 ;
  assign y7440 = ~n16551 ;
  assign y7441 = ~n16554 ;
  assign y7442 = ~n16559 ;
  assign y7443 = ~n16560 ;
  assign y7444 = ~1'b0 ;
  assign y7445 = ~1'b0 ;
  assign y7446 = ~1'b0 ;
  assign y7447 = n16562 ;
  assign y7448 = ~n16564 ;
  assign y7449 = ~1'b0 ;
  assign y7450 = ~n16565 ;
  assign y7451 = ~1'b0 ;
  assign y7452 = n16568 ;
  assign y7453 = n16570 ;
  assign y7454 = n16572 ;
  assign y7455 = n16574 ;
  assign y7456 = n16578 ;
  assign y7457 = ~n16579 ;
  assign y7458 = ~n16584 ;
  assign y7459 = ~1'b0 ;
  assign y7460 = ~n16587 ;
  assign y7461 = n16589 ;
  assign y7462 = n16591 ;
  assign y7463 = n16592 ;
  assign y7464 = ~n16603 ;
  assign y7465 = n2535 ;
  assign y7466 = ~n16605 ;
  assign y7467 = n16606 ;
  assign y7468 = ~n16611 ;
  assign y7469 = ~n16615 ;
  assign y7470 = n16617 ;
  assign y7471 = n9192 ;
  assign y7472 = ~n16620 ;
  assign y7473 = ~n16623 ;
  assign y7474 = ~n16624 ;
  assign y7475 = ~1'b0 ;
  assign y7476 = ~1'b0 ;
  assign y7477 = n12349 ;
  assign y7478 = ~n16629 ;
  assign y7479 = n16632 ;
  assign y7480 = n13372 ;
  assign y7481 = n16633 ;
  assign y7482 = n16638 ;
  assign y7483 = ~1'b0 ;
  assign y7484 = ~1'b0 ;
  assign y7485 = ~n5910 ;
  assign y7486 = n922 ;
  assign y7487 = n16639 ;
  assign y7488 = n16640 ;
  assign y7489 = ~n16645 ;
  assign y7490 = n16647 ;
  assign y7491 = ~1'b0 ;
  assign y7492 = ~n16651 ;
  assign y7493 = n16653 ;
  assign y7494 = ~n16655 ;
  assign y7495 = 1'b0 ;
  assign y7496 = n16656 ;
  assign y7497 = ~n16659 ;
  assign y7498 = ~n1309 ;
  assign y7499 = ~n16660 ;
  assign y7500 = ~n16665 ;
  assign y7501 = ~n16669 ;
  assign y7502 = ~n16671 ;
  assign y7503 = ~1'b0 ;
  assign y7504 = n16679 ;
  assign y7505 = n16681 ;
  assign y7506 = n16683 ;
  assign y7507 = ~1'b0 ;
  assign y7508 = ~1'b0 ;
  assign y7509 = ~n16685 ;
  assign y7510 = ~n16688 ;
  assign y7511 = n16691 ;
  assign y7512 = ~n16698 ;
  assign y7513 = ~n5158 ;
  assign y7514 = n16699 ;
  assign y7515 = ~n16701 ;
  assign y7516 = ~n16703 ;
  assign y7517 = ~n16705 ;
  assign y7518 = ~n16708 ;
  assign y7519 = n16712 ;
  assign y7520 = ~1'b0 ;
  assign y7521 = ~n16715 ;
  assign y7522 = n16717 ;
  assign y7523 = ~n16722 ;
  assign y7524 = ~1'b0 ;
  assign y7525 = n16723 ;
  assign y7526 = ~1'b0 ;
  assign y7527 = ~n8182 ;
  assign y7528 = ~n16727 ;
  assign y7529 = n16730 ;
  assign y7530 = n16737 ;
  assign y7531 = n16740 ;
  assign y7532 = n16744 ;
  assign y7533 = ~n16749 ;
  assign y7534 = ~n16750 ;
  assign y7535 = ~n16751 ;
  assign y7536 = ~1'b0 ;
  assign y7537 = ~n16753 ;
  assign y7538 = ~1'b0 ;
  assign y7539 = ~n16761 ;
  assign y7540 = ~n16768 ;
  assign y7541 = ~n16771 ;
  assign y7542 = ~1'b0 ;
  assign y7543 = ~n16782 ;
  assign y7544 = n16783 ;
  assign y7545 = n16784 ;
  assign y7546 = ~n16788 ;
  assign y7547 = n16791 ;
  assign y7548 = ~1'b0 ;
  assign y7549 = ~1'b0 ;
  assign y7550 = n16794 ;
  assign y7551 = n16807 ;
  assign y7552 = n16812 ;
  assign y7553 = ~n16821 ;
  assign y7554 = ~n16822 ;
  assign y7555 = ~n16824 ;
  assign y7556 = n16827 ;
  assign y7557 = ~n16829 ;
  assign y7558 = n16830 ;
  assign y7559 = n4844 ;
  assign y7560 = n16832 ;
  assign y7561 = ~n2835 ;
  assign y7562 = ~n16833 ;
  assign y7563 = n16837 ;
  assign y7564 = ~1'b0 ;
  assign y7565 = n16839 ;
  assign y7566 = ~n16841 ;
  assign y7567 = n16843 ;
  assign y7568 = ~n16851 ;
  assign y7569 = ~n16855 ;
  assign y7570 = n16858 ;
  assign y7571 = ~n16864 ;
  assign y7572 = ~1'b0 ;
  assign y7573 = n12317 ;
  assign y7574 = ~n16866 ;
  assign y7575 = n1846 ;
  assign y7576 = ~1'b0 ;
  assign y7577 = ~n16867 ;
  assign y7578 = 1'b0 ;
  assign y7579 = n16869 ;
  assign y7580 = ~n16877 ;
  assign y7581 = 1'b0 ;
  assign y7582 = ~1'b0 ;
  assign y7583 = ~n16882 ;
  assign y7584 = ~1'b0 ;
  assign y7585 = ~1'b0 ;
  assign y7586 = n8208 ;
  assign y7587 = 1'b0 ;
  assign y7588 = ~n16883 ;
  assign y7589 = ~n16888 ;
  assign y7590 = ~n16890 ;
  assign y7591 = n16891 ;
  assign y7592 = 1'b0 ;
  assign y7593 = ~n16892 ;
  assign y7594 = ~n16894 ;
  assign y7595 = ~n16897 ;
  assign y7596 = n16899 ;
  assign y7597 = ~1'b0 ;
  assign y7598 = n14835 ;
  assign y7599 = ~1'b0 ;
  assign y7600 = n16900 ;
  assign y7601 = ~n16901 ;
  assign y7602 = ~n16902 ;
  assign y7603 = ~1'b0 ;
  assign y7604 = n16912 ;
  assign y7605 = n16915 ;
  assign y7606 = n16916 ;
  assign y7607 = ~n16920 ;
  assign y7608 = n16923 ;
  assign y7609 = n16924 ;
  assign y7610 = ~n16928 ;
  assign y7611 = ~n4863 ;
  assign y7612 = ~n16934 ;
  assign y7613 = n16935 ;
  assign y7614 = n16936 ;
  assign y7615 = ~n16939 ;
  assign y7616 = ~n16942 ;
  assign y7617 = n16946 ;
  assign y7618 = ~1'b0 ;
  assign y7619 = n16948 ;
  assign y7620 = ~1'b0 ;
  assign y7621 = ~1'b0 ;
  assign y7622 = ~n16949 ;
  assign y7623 = ~n16950 ;
  assign y7624 = ~1'b0 ;
  assign y7625 = ~1'b0 ;
  assign y7626 = ~1'b0 ;
  assign y7627 = ~n16952 ;
  assign y7628 = ~n16953 ;
  assign y7629 = ~1'b0 ;
  assign y7630 = n16955 ;
  assign y7631 = n16956 ;
  assign y7632 = ~1'b0 ;
  assign y7633 = n16961 ;
  assign y7634 = n16963 ;
  assign y7635 = ~1'b0 ;
  assign y7636 = n16965 ;
  assign y7637 = n16967 ;
  assign y7638 = n16969 ;
  assign y7639 = n16970 ;
  assign y7640 = n16972 ;
  assign y7641 = ~1'b0 ;
  assign y7642 = ~n16973 ;
  assign y7643 = ~1'b0 ;
  assign y7644 = ~1'b0 ;
  assign y7645 = ~1'b0 ;
  assign y7646 = ~n16975 ;
  assign y7647 = ~n16978 ;
  assign y7648 = n16981 ;
  assign y7649 = ~n16982 ;
  assign y7650 = n16985 ;
  assign y7651 = ~n16986 ;
  assign y7652 = ~1'b0 ;
  assign y7653 = n10263 ;
  assign y7654 = ~1'b0 ;
  assign y7655 = ~n16988 ;
  assign y7656 = ~1'b0 ;
  assign y7657 = n16989 ;
  assign y7658 = ~n16994 ;
  assign y7659 = n16995 ;
  assign y7660 = ~n16999 ;
  assign y7661 = n7605 ;
  assign y7662 = ~n17001 ;
  assign y7663 = ~1'b0 ;
  assign y7664 = ~1'b0 ;
  assign y7665 = ~n17002 ;
  assign y7666 = n17003 ;
  assign y7667 = ~n17007 ;
  assign y7668 = ~n17008 ;
  assign y7669 = ~n16849 ;
  assign y7670 = ~1'b0 ;
  assign y7671 = ~1'b0 ;
  assign y7672 = n6363 ;
  assign y7673 = n17009 ;
  assign y7674 = n17011 ;
  assign y7675 = ~1'b0 ;
  assign y7676 = ~1'b0 ;
  assign y7677 = ~1'b0 ;
  assign y7678 = ~n1046 ;
  assign y7679 = n17012 ;
  assign y7680 = n17013 ;
  assign y7681 = n17015 ;
  assign y7682 = n17023 ;
  assign y7683 = ~n17025 ;
  assign y7684 = ~1'b0 ;
  assign y7685 = ~n17026 ;
  assign y7686 = 1'b0 ;
  assign y7687 = n17028 ;
  assign y7688 = n17032 ;
  assign y7689 = ~n17033 ;
  assign y7690 = n17040 ;
  assign y7691 = ~1'b0 ;
  assign y7692 = n17043 ;
  assign y7693 = ~n17046 ;
  assign y7694 = n17048 ;
  assign y7695 = ~n17049 ;
  assign y7696 = ~1'b0 ;
  assign y7697 = ~n17052 ;
  assign y7698 = n17053 ;
  assign y7699 = n11343 ;
  assign y7700 = n17055 ;
  assign y7701 = ~n17062 ;
  assign y7702 = n17063 ;
  assign y7703 = n17079 ;
  assign y7704 = ~n17081 ;
  assign y7705 = ~n17086 ;
  assign y7706 = n17091 ;
  assign y7707 = ~n17092 ;
  assign y7708 = ~n17093 ;
  assign y7709 = ~1'b0 ;
  assign y7710 = ~1'b0 ;
  assign y7711 = ~n17094 ;
  assign y7712 = n17097 ;
  assign y7713 = n17098 ;
  assign y7714 = ~1'b0 ;
  assign y7715 = n17101 ;
  assign y7716 = ~n17102 ;
  assign y7717 = ~n17107 ;
  assign y7718 = n367 ;
  assign y7719 = ~n17108 ;
  assign y7720 = n17114 ;
  assign y7721 = ~1'b0 ;
  assign y7722 = ~1'b0 ;
  assign y7723 = n17116 ;
  assign y7724 = n6722 ;
  assign y7725 = ~n17118 ;
  assign y7726 = n17120 ;
  assign y7727 = ~n17121 ;
  assign y7728 = n17125 ;
  assign y7729 = n17131 ;
  assign y7730 = ~1'b0 ;
  assign y7731 = ~1'b0 ;
  assign y7732 = ~n14391 ;
  assign y7733 = ~n17132 ;
  assign y7734 = n17139 ;
  assign y7735 = ~n17141 ;
  assign y7736 = ~1'b0 ;
  assign y7737 = ~n17143 ;
  assign y7738 = ~n17144 ;
  assign y7739 = n17147 ;
  assign y7740 = ~n17149 ;
  assign y7741 = n17152 ;
  assign y7742 = ~n17154 ;
  assign y7743 = ~n17157 ;
  assign y7744 = ~1'b0 ;
  assign y7745 = n17161 ;
  assign y7746 = ~n17165 ;
  assign y7747 = ~1'b0 ;
  assign y7748 = n17168 ;
  assign y7749 = 1'b0 ;
  assign y7750 = ~n17169 ;
  assign y7751 = n17175 ;
  assign y7752 = ~n17177 ;
  assign y7753 = ~n17180 ;
  assign y7754 = ~n17190 ;
  assign y7755 = n17192 ;
  assign y7756 = n17193 ;
  assign y7757 = ~n17194 ;
  assign y7758 = ~1'b0 ;
  assign y7759 = ~n17195 ;
  assign y7760 = ~1'b0 ;
  assign y7761 = ~n17196 ;
  assign y7762 = n17197 ;
  assign y7763 = n17198 ;
  assign y7764 = ~n17199 ;
  assign y7765 = ~n17200 ;
  assign y7766 = n13257 ;
  assign y7767 = ~n17201 ;
  assign y7768 = n17203 ;
  assign y7769 = n17204 ;
  assign y7770 = n17205 ;
  assign y7771 = ~n17209 ;
  assign y7772 = n17210 ;
  assign y7773 = ~n17212 ;
  assign y7774 = ~n17214 ;
  assign y7775 = n17218 ;
  assign y7776 = n17221 ;
  assign y7777 = n17223 ;
  assign y7778 = ~n17231 ;
  assign y7779 = n17233 ;
  assign y7780 = n17236 ;
  assign y7781 = n17238 ;
  assign y7782 = n17240 ;
  assign y7783 = n17241 ;
  assign y7784 = ~n17242 ;
  assign y7785 = n17243 ;
  assign y7786 = n17248 ;
  assign y7787 = ~n17250 ;
  assign y7788 = n17251 ;
  assign y7789 = ~n17253 ;
  assign y7790 = ~n17258 ;
  assign y7791 = ~1'b0 ;
  assign y7792 = ~n17264 ;
  assign y7793 = ~1'b0 ;
  assign y7794 = ~n17267 ;
  assign y7795 = ~n17268 ;
  assign y7796 = ~n17271 ;
  assign y7797 = n17272 ;
  assign y7798 = ~n17273 ;
  assign y7799 = ~1'b0 ;
  assign y7800 = n17275 ;
  assign y7801 = ~1'b0 ;
  assign y7802 = ~n17276 ;
  assign y7803 = n17277 ;
  assign y7804 = ~n7853 ;
  assign y7805 = n17281 ;
  assign y7806 = ~n17286 ;
  assign y7807 = ~1'b0 ;
  assign y7808 = ~n17287 ;
  assign y7809 = ~1'b0 ;
  assign y7810 = ~n17288 ;
  assign y7811 = n17291 ;
  assign y7812 = ~n14236 ;
  assign y7813 = ~n17293 ;
  assign y7814 = n16230 ;
  assign y7815 = n17295 ;
  assign y7816 = ~n17298 ;
  assign y7817 = ~n17300 ;
  assign y7818 = ~n17301 ;
  assign y7819 = ~n17308 ;
  assign y7820 = n17309 ;
  assign y7821 = ~n17310 ;
  assign y7822 = ~n17311 ;
  assign y7823 = ~1'b0 ;
  assign y7824 = ~1'b0 ;
  assign y7825 = n17316 ;
  assign y7826 = ~n17317 ;
  assign y7827 = n17320 ;
  assign y7828 = n17325 ;
  assign y7829 = ~n17327 ;
  assign y7830 = ~1'b0 ;
  assign y7831 = n17328 ;
  assign y7832 = ~1'b0 ;
  assign y7833 = ~1'b0 ;
  assign y7834 = n17333 ;
  assign y7835 = n17334 ;
  assign y7836 = ~1'b0 ;
  assign y7837 = n17335 ;
  assign y7838 = n17344 ;
  assign y7839 = ~n17345 ;
  assign y7840 = n17349 ;
  assign y7841 = n17355 ;
  assign y7842 = n17357 ;
  assign y7843 = ~1'b0 ;
  assign y7844 = ~1'b0 ;
  assign y7845 = ~n17362 ;
  assign y7846 = 1'b0 ;
  assign y7847 = ~1'b0 ;
  assign y7848 = n17364 ;
  assign y7849 = ~n17369 ;
  assign y7850 = n17372 ;
  assign y7851 = ~1'b0 ;
  assign y7852 = ~n17379 ;
  assign y7853 = ~n529 ;
  assign y7854 = n17381 ;
  assign y7855 = ~n17385 ;
  assign y7856 = n17386 ;
  assign y7857 = n17387 ;
  assign y7858 = n17389 ;
  assign y7859 = n17393 ;
  assign y7860 = ~n17394 ;
  assign y7861 = n17396 ;
  assign y7862 = ~1'b0 ;
  assign y7863 = n17401 ;
  assign y7864 = n17403 ;
  assign y7865 = ~1'b0 ;
  assign y7866 = n17405 ;
  assign y7867 = ~n2089 ;
  assign y7868 = ~n17407 ;
  assign y7869 = ~1'b0 ;
  assign y7870 = ~n17408 ;
  assign y7871 = n17409 ;
  assign y7872 = ~1'b0 ;
  assign y7873 = ~1'b0 ;
  assign y7874 = ~1'b0 ;
  assign y7875 = ~1'b0 ;
  assign y7876 = ~n17410 ;
  assign y7877 = n17413 ;
  assign y7878 = ~1'b0 ;
  assign y7879 = ~n17419 ;
  assign y7880 = n17422 ;
  assign y7881 = ~n17423 ;
  assign y7882 = ~1'b0 ;
  assign y7883 = ~n17428 ;
  assign y7884 = n17430 ;
  assign y7885 = n17431 ;
  assign y7886 = n3275 ;
  assign y7887 = n17432 ;
  assign y7888 = ~n17433 ;
  assign y7889 = ~n14320 ;
  assign y7890 = n17439 ;
  assign y7891 = n17447 ;
  assign y7892 = ~n17450 ;
  assign y7893 = ~1'b0 ;
  assign y7894 = ~n17451 ;
  assign y7895 = ~1'b0 ;
  assign y7896 = ~n17457 ;
  assign y7897 = n17465 ;
  assign y7898 = n17469 ;
  assign y7899 = n17472 ;
  assign y7900 = n17474 ;
  assign y7901 = n17482 ;
  assign y7902 = n7265 ;
  assign y7903 = ~n17484 ;
  assign y7904 = ~1'b0 ;
  assign y7905 = ~1'b0 ;
  assign y7906 = n17488 ;
  assign y7907 = ~n17491 ;
  assign y7908 = n17493 ;
  assign y7909 = ~n17500 ;
  assign y7910 = ~1'b0 ;
  assign y7911 = ~n17502 ;
  assign y7912 = n17503 ;
  assign y7913 = ~n17504 ;
  assign y7914 = ~n17507 ;
  assign y7915 = ~1'b0 ;
  assign y7916 = n17509 ;
  assign y7917 = n17511 ;
  assign y7918 = ~n17512 ;
  assign y7919 = ~n17515 ;
  assign y7920 = ~n17207 ;
  assign y7921 = n17521 ;
  assign y7922 = ~1'b0 ;
  assign y7923 = ~n17523 ;
  assign y7924 = ~n17524 ;
  assign y7925 = n17527 ;
  assign y7926 = n17529 ;
  assign y7927 = ~n17530 ;
  assign y7928 = ~n17532 ;
  assign y7929 = ~n8740 ;
  assign y7930 = ~n17535 ;
  assign y7931 = n17538 ;
  assign y7932 = ~n17539 ;
  assign y7933 = n17541 ;
  assign y7934 = ~n14246 ;
  assign y7935 = n17542 ;
  assign y7936 = n17543 ;
  assign y7937 = 1'b0 ;
  assign y7938 = ~1'b0 ;
  assign y7939 = ~n17553 ;
  assign y7940 = ~n17557 ;
  assign y7941 = ~1'b0 ;
  assign y7942 = ~n17562 ;
  assign y7943 = n17568 ;
  assign y7944 = n6582 ;
  assign y7945 = ~n17569 ;
  assign y7946 = n7359 ;
  assign y7947 = ~n17571 ;
  assign y7948 = n17583 ;
  assign y7949 = ~1'b0 ;
  assign y7950 = ~n17586 ;
  assign y7951 = n13343 ;
  assign y7952 = ~n17592 ;
  assign y7953 = ~n17594 ;
  assign y7954 = ~n17595 ;
  assign y7955 = ~n17599 ;
  assign y7956 = ~1'b0 ;
  assign y7957 = ~n17603 ;
  assign y7958 = ~n17604 ;
  assign y7959 = n5443 ;
  assign y7960 = ~n17606 ;
  assign y7961 = ~n17610 ;
  assign y7962 = n712 ;
  assign y7963 = ~n17612 ;
  assign y7964 = n17620 ;
  assign y7965 = ~n17622 ;
  assign y7966 = 1'b0 ;
  assign y7967 = ~1'b0 ;
  assign y7968 = n17627 ;
  assign y7969 = ~1'b0 ;
  assign y7970 = n17630 ;
  assign y7971 = ~n17632 ;
  assign y7972 = ~n17635 ;
  assign y7973 = n17636 ;
  assign y7974 = ~1'b0 ;
  assign y7975 = 1'b0 ;
  assign y7976 = n17637 ;
  assign y7977 = ~n17427 ;
  assign y7978 = ~1'b0 ;
  assign y7979 = ~1'b0 ;
  assign y7980 = ~n130 ;
  assign y7981 = ~1'b0 ;
  assign y7982 = ~n17639 ;
  assign y7983 = n4366 ;
  assign y7984 = ~n17642 ;
  assign y7985 = n17647 ;
  assign y7986 = ~n17651 ;
  assign y7987 = ~1'b0 ;
  assign y7988 = n17652 ;
  assign y7989 = ~n17655 ;
  assign y7990 = ~n17659 ;
  assign y7991 = ~n17664 ;
  assign y7992 = 1'b0 ;
  assign y7993 = n17667 ;
  assign y7994 = ~n17674 ;
  assign y7995 = n17675 ;
  assign y7996 = ~1'b0 ;
  assign y7997 = ~n17684 ;
  assign y7998 = ~n17689 ;
  assign y7999 = n12712 ;
  assign y8000 = n17693 ;
  assign y8001 = ~1'b0 ;
  assign y8002 = ~n17694 ;
  assign y8003 = ~n17698 ;
  assign y8004 = n17706 ;
  assign y8005 = ~1'b0 ;
  assign y8006 = ~1'b0 ;
  assign y8007 = ~n10266 ;
  assign y8008 = n17714 ;
  assign y8009 = n16048 ;
  assign y8010 = ~n17716 ;
  assign y8011 = n17717 ;
  assign y8012 = n17718 ;
  assign y8013 = ~1'b0 ;
  assign y8014 = 1'b0 ;
  assign y8015 = n17719 ;
  assign y8016 = ~1'b0 ;
  assign y8017 = ~n17720 ;
  assign y8018 = n17721 ;
  assign y8019 = ~n17722 ;
  assign y8020 = ~1'b0 ;
  assign y8021 = ~n17727 ;
  assign y8022 = ~n17738 ;
  assign y8023 = ~1'b0 ;
  assign y8024 = ~n17739 ;
  assign y8025 = n17742 ;
  assign y8026 = n17743 ;
  assign y8027 = ~1'b0 ;
  assign y8028 = ~1'b0 ;
  assign y8029 = n17746 ;
  assign y8030 = ~n17748 ;
  assign y8031 = ~n17750 ;
  assign y8032 = ~1'b0 ;
  assign y8033 = ~n17751 ;
  assign y8034 = n17752 ;
  assign y8035 = ~n17757 ;
  assign y8036 = n17760 ;
  assign y8037 = ~1'b0 ;
  assign y8038 = ~n17763 ;
  assign y8039 = ~1'b0 ;
  assign y8040 = ~n17764 ;
  assign y8041 = ~n17766 ;
  assign y8042 = ~n8260 ;
  assign y8043 = n17769 ;
  assign y8044 = ~n17770 ;
  assign y8045 = n17773 ;
  assign y8046 = n17774 ;
  assign y8047 = ~n17775 ;
  assign y8048 = ~n17776 ;
  assign y8049 = ~n17778 ;
  assign y8050 = ~n17792 ;
  assign y8051 = n17794 ;
  assign y8052 = ~1'b0 ;
  assign y8053 = ~n17797 ;
  assign y8054 = ~n17798 ;
  assign y8055 = ~n17801 ;
  assign y8056 = ~n17803 ;
  assign y8057 = ~1'b0 ;
  assign y8058 = n17809 ;
  assign y8059 = ~n17811 ;
  assign y8060 = ~n17812 ;
  assign y8061 = ~n17816 ;
  assign y8062 = n17825 ;
  assign y8063 = n17828 ;
  assign y8064 = ~n17829 ;
  assign y8065 = n17833 ;
  assign y8066 = ~n17838 ;
  assign y8067 = ~n17839 ;
  assign y8068 = n17840 ;
  assign y8069 = n17845 ;
  assign y8070 = ~n17847 ;
  assign y8071 = ~1'b0 ;
  assign y8072 = ~1'b0 ;
  assign y8073 = ~1'b0 ;
  assign y8074 = ~1'b0 ;
  assign y8075 = n17849 ;
  assign y8076 = n17851 ;
  assign y8077 = n17852 ;
  assign y8078 = n17854 ;
  assign y8079 = ~n17856 ;
  assign y8080 = n17861 ;
  assign y8081 = ~n17862 ;
  assign y8082 = ~n17863 ;
  assign y8083 = n17865 ;
  assign y8084 = ~n17867 ;
  assign y8085 = n17870 ;
  assign y8086 = ~n17872 ;
  assign y8087 = ~n17875 ;
  assign y8088 = n17877 ;
  assign y8089 = ~1'b0 ;
  assign y8090 = n17882 ;
  assign y8091 = n17893 ;
  assign y8092 = ~n17894 ;
  assign y8093 = ~n17895 ;
  assign y8094 = ~n17896 ;
  assign y8095 = ~n17902 ;
  assign y8096 = ~n17904 ;
  assign y8097 = ~1'b0 ;
  assign y8098 = ~1'b0 ;
  assign y8099 = ~1'b0 ;
  assign y8100 = n17905 ;
  assign y8101 = ~1'b0 ;
  assign y8102 = n17906 ;
  assign y8103 = ~1'b0 ;
  assign y8104 = ~n17909 ;
  assign y8105 = n17915 ;
  assign y8106 = ~n17919 ;
  assign y8107 = ~1'b0 ;
  assign y8108 = n17921 ;
  assign y8109 = n17924 ;
  assign y8110 = 1'b0 ;
  assign y8111 = ~n17926 ;
  assign y8112 = ~1'b0 ;
  assign y8113 = n17930 ;
  assign y8114 = ~n17934 ;
  assign y8115 = ~1'b0 ;
  assign y8116 = n17938 ;
  assign y8117 = ~n17939 ;
  assign y8118 = ~1'b0 ;
  assign y8119 = ~n17945 ;
  assign y8120 = ~1'b0 ;
  assign y8121 = ~n17946 ;
  assign y8122 = n17947 ;
  assign y8123 = ~n7260 ;
  assign y8124 = n17949 ;
  assign y8125 = n17952 ;
  assign y8126 = ~1'b0 ;
  assign y8127 = n17953 ;
  assign y8128 = ~1'b0 ;
  assign y8129 = ~n17955 ;
  assign y8130 = n17958 ;
  assign y8131 = ~n17960 ;
  assign y8132 = n17962 ;
  assign y8133 = ~1'b0 ;
  assign y8134 = ~1'b0 ;
  assign y8135 = ~n17964 ;
  assign y8136 = ~n17966 ;
  assign y8137 = ~n17968 ;
  assign y8138 = n6829 ;
  assign y8139 = ~n17971 ;
  assign y8140 = n17979 ;
  assign y8141 = n17982 ;
  assign y8142 = ~n17988 ;
  assign y8143 = n17989 ;
  assign y8144 = ~1'b0 ;
  assign y8145 = ~n17978 ;
  assign y8146 = n17991 ;
  assign y8147 = ~1'b0 ;
  assign y8148 = n17994 ;
  assign y8149 = ~1'b0 ;
  assign y8150 = n17996 ;
  assign y8151 = ~1'b0 ;
  assign y8152 = ~n17997 ;
  assign y8153 = ~n17999 ;
  assign y8154 = ~1'b0 ;
  assign y8155 = ~n7444 ;
  assign y8156 = ~1'b0 ;
  assign y8157 = ~n18001 ;
  assign y8158 = ~n18002 ;
  assign y8159 = ~n269 ;
  assign y8160 = ~1'b0 ;
  assign y8161 = n18004 ;
  assign y8162 = ~1'b0 ;
  assign y8163 = n18005 ;
  assign y8164 = n12115 ;
  assign y8165 = ~1'b0 ;
  assign y8166 = ~n18007 ;
  assign y8167 = ~n18009 ;
  assign y8168 = ~n18011 ;
  assign y8169 = ~n18013 ;
  assign y8170 = n18016 ;
  assign y8171 = ~n18021 ;
  assign y8172 = ~n18022 ;
  assign y8173 = ~n18024 ;
  assign y8174 = n18025 ;
  assign y8175 = ~n18030 ;
  assign y8176 = ~n18038 ;
  assign y8177 = ~n18040 ;
  assign y8178 = ~1'b0 ;
  assign y8179 = ~n18047 ;
  assign y8180 = ~n18052 ;
  assign y8181 = ~1'b0 ;
  assign y8182 = ~n18054 ;
  assign y8183 = ~1'b0 ;
  assign y8184 = n18055 ;
  assign y8185 = ~1'b0 ;
  assign y8186 = n18056 ;
  assign y8187 = ~1'b0 ;
  assign y8188 = ~1'b0 ;
  assign y8189 = ~n18059 ;
  assign y8190 = n18063 ;
  assign y8191 = ~n18065 ;
  assign y8192 = n18067 ;
  assign y8193 = ~n18068 ;
  assign y8194 = ~n18069 ;
  assign y8195 = n18070 ;
  assign y8196 = ~1'b0 ;
  assign y8197 = ~1'b0 ;
  assign y8198 = ~1'b0 ;
  assign y8199 = ~1'b0 ;
  assign y8200 = ~n18072 ;
  assign y8201 = ~1'b0 ;
  assign y8202 = n18076 ;
  assign y8203 = n18078 ;
  assign y8204 = n18080 ;
  assign y8205 = ~n18086 ;
  assign y8206 = ~n18087 ;
  assign y8207 = ~n18088 ;
  assign y8208 = ~1'b0 ;
  assign y8209 = ~n18089 ;
  assign y8210 = ~n18092 ;
  assign y8211 = n18093 ;
  assign y8212 = ~1'b0 ;
  assign y8213 = ~1'b0 ;
  assign y8214 = n18094 ;
  assign y8215 = n18096 ;
  assign y8216 = n18099 ;
  assign y8217 = n18103 ;
  assign y8218 = ~1'b0 ;
  assign y8219 = ~n18107 ;
  assign y8220 = n18114 ;
  assign y8221 = n6346 ;
  assign y8222 = ~1'b0 ;
  assign y8223 = ~1'b0 ;
  assign y8224 = n18118 ;
  assign y8225 = n18120 ;
  assign y8226 = ~n18123 ;
  assign y8227 = n18124 ;
  assign y8228 = ~n18125 ;
  assign y8229 = n18126 ;
  assign y8230 = n18131 ;
  assign y8231 = ~1'b0 ;
  assign y8232 = ~n18141 ;
  assign y8233 = ~1'b0 ;
  assign y8234 = ~n18142 ;
  assign y8235 = n18147 ;
  assign y8236 = n18148 ;
  assign y8237 = ~n18149 ;
  assign y8238 = n18151 ;
  assign y8239 = ~1'b0 ;
  assign y8240 = ~n18153 ;
  assign y8241 = n18156 ;
  assign y8242 = ~1'b0 ;
  assign y8243 = n18160 ;
  assign y8244 = n18164 ;
  assign y8245 = ~n18165 ;
  assign y8246 = ~n6139 ;
  assign y8247 = ~1'b0 ;
  assign y8248 = n18170 ;
  assign y8249 = n18171 ;
  assign y8250 = ~n18175 ;
  assign y8251 = n18179 ;
  assign y8252 = n18180 ;
  assign y8253 = ~1'b0 ;
  assign y8254 = ~n18182 ;
  assign y8255 = ~1'b0 ;
  assign y8256 = ~n18185 ;
  assign y8257 = n13143 ;
  assign y8258 = ~n18190 ;
  assign y8259 = ~n18193 ;
  assign y8260 = ~1'b0 ;
  assign y8261 = n18194 ;
  assign y8262 = n18196 ;
  assign y8263 = n18198 ;
  assign y8264 = n18202 ;
  assign y8265 = ~n18206 ;
  assign y8266 = ~1'b0 ;
  assign y8267 = ~1'b0 ;
  assign y8268 = ~n18210 ;
  assign y8269 = n18211 ;
  assign y8270 = n18212 ;
  assign y8271 = 1'b0 ;
  assign y8272 = n18214 ;
  assign y8273 = ~1'b0 ;
  assign y8274 = ~1'b0 ;
  assign y8275 = n18215 ;
  assign y8276 = ~n18218 ;
  assign y8277 = n18219 ;
  assign y8278 = ~n18220 ;
  assign y8279 = n18222 ;
  assign y8280 = n18223 ;
  assign y8281 = n18224 ;
  assign y8282 = ~n18225 ;
  assign y8283 = ~1'b0 ;
  assign y8284 = ~n18227 ;
  assign y8285 = ~1'b0 ;
  assign y8286 = ~1'b0 ;
  assign y8287 = ~n18232 ;
  assign y8288 = n18234 ;
  assign y8289 = n18235 ;
  assign y8290 = ~n18241 ;
  assign y8291 = n18245 ;
  assign y8292 = 1'b0 ;
  assign y8293 = ~n18246 ;
  assign y8294 = n18247 ;
  assign y8295 = n18252 ;
  assign y8296 = ~n18255 ;
  assign y8297 = n18260 ;
  assign y8298 = n6218 ;
  assign y8299 = 1'b0 ;
  assign y8300 = ~1'b0 ;
  assign y8301 = ~n18262 ;
  assign y8302 = ~1'b0 ;
  assign y8303 = ~n18263 ;
  assign y8304 = n18264 ;
  assign y8305 = ~n18273 ;
  assign y8306 = ~n18275 ;
  assign y8307 = n18278 ;
  assign y8308 = ~n18279 ;
  assign y8309 = n18280 ;
  assign y8310 = ~1'b0 ;
  assign y8311 = ~1'b0 ;
  assign y8312 = ~n18284 ;
  assign y8313 = ~n18286 ;
  assign y8314 = n18290 ;
  assign y8315 = n18295 ;
  assign y8316 = ~1'b0 ;
  assign y8317 = n18300 ;
  assign y8318 = ~n18301 ;
  assign y8319 = n18305 ;
  assign y8320 = ~1'b0 ;
  assign y8321 = n18306 ;
  assign y8322 = ~1'b0 ;
  assign y8323 = ~1'b0 ;
  assign y8324 = ~n18308 ;
  assign y8325 = ~1'b0 ;
  assign y8326 = ~n18310 ;
  assign y8327 = n18313 ;
  assign y8328 = ~n18317 ;
  assign y8329 = ~1'b0 ;
  assign y8330 = ~n18319 ;
  assign y8331 = ~1'b0 ;
  assign y8332 = n18322 ;
  assign y8333 = n18323 ;
  assign y8334 = ~n18324 ;
  assign y8335 = n18327 ;
  assign y8336 = n18335 ;
  assign y8337 = ~1'b0 ;
  assign y8338 = ~1'b0 ;
  assign y8339 = ~1'b0 ;
  assign y8340 = ~1'b0 ;
  assign y8341 = ~n18336 ;
  assign y8342 = ~n18337 ;
  assign y8343 = ~1'b0 ;
  assign y8344 = ~n18338 ;
  assign y8345 = n18340 ;
  assign y8346 = ~n18341 ;
  assign y8347 = ~n18342 ;
  assign y8348 = ~1'b0 ;
  assign y8349 = ~n18345 ;
  assign y8350 = n18347 ;
  assign y8351 = ~1'b0 ;
  assign y8352 = ~n18348 ;
  assign y8353 = ~n18358 ;
  assign y8354 = ~n18359 ;
  assign y8355 = n18363 ;
  assign y8356 = n18364 ;
  assign y8357 = ~n13112 ;
  assign y8358 = ~1'b0 ;
  assign y8359 = ~n18365 ;
  assign y8360 = ~n18366 ;
  assign y8361 = n18370 ;
  assign y8362 = ~n18371 ;
  assign y8363 = n18372 ;
  assign y8364 = ~n8552 ;
  assign y8365 = ~n18375 ;
  assign y8366 = ~n18376 ;
  assign y8367 = n18377 ;
  assign y8368 = ~1'b0 ;
  assign y8369 = ~n18384 ;
  assign y8370 = n7546 ;
  assign y8371 = ~n18385 ;
  assign y8372 = n18387 ;
  assign y8373 = ~1'b0 ;
  assign y8374 = ~n18389 ;
  assign y8375 = n18390 ;
  assign y8376 = ~1'b0 ;
  assign y8377 = ~n18391 ;
  assign y8378 = ~1'b0 ;
  assign y8379 = ~n18396 ;
  assign y8380 = n18398 ;
  assign y8381 = ~1'b0 ;
  assign y8382 = ~1'b0 ;
  assign y8383 = ~n18402 ;
  assign y8384 = ~1'b0 ;
  assign y8385 = n18403 ;
  assign y8386 = ~n18404 ;
  assign y8387 = ~1'b0 ;
  assign y8388 = ~n18408 ;
  assign y8389 = ~n18409 ;
  assign y8390 = n18413 ;
  assign y8391 = ~n18418 ;
  assign y8392 = n18419 ;
  assign y8393 = ~n18422 ;
  assign y8394 = n18424 ;
  assign y8395 = n18426 ;
  assign y8396 = ~1'b0 ;
  assign y8397 = ~n18430 ;
  assign y8398 = ~n18431 ;
  assign y8399 = n18433 ;
  assign y8400 = ~1'b0 ;
  assign y8401 = ~1'b0 ;
  assign y8402 = ~1'b0 ;
  assign y8403 = n18435 ;
  assign y8404 = ~n18436 ;
  assign y8405 = ~n18437 ;
  assign y8406 = ~n18438 ;
  assign y8407 = ~n18444 ;
  assign y8408 = ~n18451 ;
  assign y8409 = n18457 ;
  assign y8410 = ~1'b0 ;
  assign y8411 = ~1'b0 ;
  assign y8412 = ~n18459 ;
  assign y8413 = ~n18460 ;
  assign y8414 = n18462 ;
  assign y8415 = ~1'b0 ;
  assign y8416 = ~n18467 ;
  assign y8417 = ~1'b0 ;
  assign y8418 = ~n18471 ;
  assign y8419 = n18473 ;
  assign y8420 = n18474 ;
  assign y8421 = n18479 ;
  assign y8422 = ~n18482 ;
  assign y8423 = ~1'b0 ;
  assign y8424 = ~1'b0 ;
  assign y8425 = ~1'b0 ;
  assign y8426 = ~n18484 ;
  assign y8427 = ~n18485 ;
  assign y8428 = ~n18486 ;
  assign y8429 = ~n18488 ;
  assign y8430 = n18489 ;
  assign y8431 = ~n18493 ;
  assign y8432 = ~n18494 ;
  assign y8433 = ~n18500 ;
  assign y8434 = ~n18505 ;
  assign y8435 = ~n18510 ;
  assign y8436 = ~n18514 ;
  assign y8437 = ~n1229 ;
  assign y8438 = ~n18515 ;
  assign y8439 = ~1'b0 ;
  assign y8440 = ~n18520 ;
  assign y8441 = ~n18523 ;
  assign y8442 = n18524 ;
  assign y8443 = n18526 ;
  assign y8444 = n18529 ;
  assign y8445 = n18531 ;
  assign y8446 = n18534 ;
  assign y8447 = n18536 ;
  assign y8448 = 1'b0 ;
  assign y8449 = ~1'b0 ;
  assign y8450 = ~1'b0 ;
  assign y8451 = ~n4374 ;
  assign y8452 = ~1'b0 ;
  assign y8453 = ~n18544 ;
  assign y8454 = n18549 ;
  assign y8455 = ~1'b0 ;
  assign y8456 = ~1'b0 ;
  assign y8457 = ~n17270 ;
  assign y8458 = n18550 ;
  assign y8459 = n18551 ;
  assign y8460 = ~n18552 ;
  assign y8461 = ~n18554 ;
  assign y8462 = ~n18558 ;
  assign y8463 = n18560 ;
  assign y8464 = n18561 ;
  assign y8465 = ~n18563 ;
  assign y8466 = ~n18568 ;
  assign y8467 = ~1'b0 ;
  assign y8468 = ~1'b0 ;
  assign y8469 = ~n18570 ;
  assign y8470 = n18573 ;
  assign y8471 = n18576 ;
  assign y8472 = ~n18578 ;
  assign y8473 = ~1'b0 ;
  assign y8474 = ~n11506 ;
  assign y8475 = n18580 ;
  assign y8476 = n18582 ;
  assign y8477 = ~1'b0 ;
  assign y8478 = ~n18583 ;
  assign y8479 = ~1'b0 ;
  assign y8480 = ~1'b0 ;
  assign y8481 = ~n18584 ;
  assign y8482 = ~1'b0 ;
  assign y8483 = ~n18587 ;
  assign y8484 = ~1'b0 ;
  assign y8485 = ~n18588 ;
  assign y8486 = n18591 ;
  assign y8487 = n13111 ;
  assign y8488 = ~n18592 ;
  assign y8489 = n18593 ;
  assign y8490 = ~n18595 ;
  assign y8491 = ~1'b0 ;
  assign y8492 = n1029 ;
  assign y8493 = ~n18599 ;
  assign y8494 = ~n18601 ;
  assign y8495 = ~n18606 ;
  assign y8496 = ~n18607 ;
  assign y8497 = ~1'b0 ;
  assign y8498 = ~n18612 ;
  assign y8499 = n18613 ;
  assign y8500 = ~n18614 ;
  assign y8501 = n18617 ;
  assign y8502 = n18619 ;
  assign y8503 = n18623 ;
  assign y8504 = n18624 ;
  assign y8505 = ~n484 ;
  assign y8506 = ~1'b0 ;
  assign y8507 = n18626 ;
  assign y8508 = ~n18633 ;
  assign y8509 = ~n18636 ;
  assign y8510 = n18641 ;
  assign y8511 = ~n18647 ;
  assign y8512 = ~1'b0 ;
  assign y8513 = n18652 ;
  assign y8514 = ~n18654 ;
  assign y8515 = ~1'b0 ;
  assign y8516 = n18655 ;
  assign y8517 = n18661 ;
  assign y8518 = ~n18662 ;
  assign y8519 = ~n18667 ;
  assign y8520 = n18675 ;
  assign y8521 = n18677 ;
  assign y8522 = ~n18681 ;
  assign y8523 = ~n18683 ;
  assign y8524 = ~n18686 ;
  assign y8525 = ~1'b0 ;
  assign y8526 = n18688 ;
  assign y8527 = n18691 ;
  assign y8528 = ~1'b0 ;
  assign y8529 = ~n18695 ;
  assign y8530 = 1'b0 ;
  assign y8531 = ~n9064 ;
  assign y8532 = ~n18700 ;
  assign y8533 = ~1'b0 ;
  assign y8534 = ~1'b0 ;
  assign y8535 = ~n18704 ;
  assign y8536 = n18708 ;
  assign y8537 = n18711 ;
  assign y8538 = ~n18716 ;
  assign y8539 = ~1'b0 ;
  assign y8540 = ~1'b0 ;
  assign y8541 = n2429 ;
  assign y8542 = ~n18717 ;
  assign y8543 = n18719 ;
  assign y8544 = n18720 ;
  assign y8545 = ~n18723 ;
  assign y8546 = ~1'b0 ;
  assign y8547 = n18725 ;
  assign y8548 = ~1'b0 ;
  assign y8549 = ~1'b0 ;
  assign y8550 = ~n18730 ;
  assign y8551 = ~1'b0 ;
  assign y8552 = n18733 ;
  assign y8553 = ~n18734 ;
  assign y8554 = ~1'b0 ;
  assign y8555 = n18737 ;
  assign y8556 = ~n7642 ;
  assign y8557 = n18738 ;
  assign y8558 = n18740 ;
  assign y8559 = n18742 ;
  assign y8560 = ~n18749 ;
  assign y8561 = ~1'b0 ;
  assign y8562 = ~n18750 ;
  assign y8563 = n8392 ;
  assign y8564 = n18751 ;
  assign y8565 = ~n18755 ;
  assign y8566 = ~1'b0 ;
  assign y8567 = n18756 ;
  assign y8568 = ~1'b0 ;
  assign y8569 = ~n18757 ;
  assign y8570 = ~n18764 ;
  assign y8571 = ~n18767 ;
  assign y8572 = ~n18769 ;
  assign y8573 = ~n18776 ;
  assign y8574 = n12489 ;
  assign y8575 = ~n18777 ;
  assign y8576 = ~1'b0 ;
  assign y8577 = ~n18778 ;
  assign y8578 = ~n18786 ;
  assign y8579 = ~1'b0 ;
  assign y8580 = ~1'b0 ;
  assign y8581 = ~1'b0 ;
  assign y8582 = ~n18787 ;
  assign y8583 = ~n18788 ;
  assign y8584 = n18790 ;
  assign y8585 = ~1'b0 ;
  assign y8586 = ~1'b0 ;
  assign y8587 = n18791 ;
  assign y8588 = ~n18793 ;
  assign y8589 = ~n18798 ;
  assign y8590 = n18800 ;
  assign y8591 = n18802 ;
  assign y8592 = ~n18803 ;
  assign y8593 = n18806 ;
  assign y8594 = ~1'b0 ;
  assign y8595 = ~n18807 ;
  assign y8596 = n18812 ;
  assign y8597 = n18816 ;
  assign y8598 = ~n18821 ;
  assign y8599 = ~n18824 ;
  assign y8600 = n18826 ;
  assign y8601 = n18827 ;
  assign y8602 = n18829 ;
  assign y8603 = n18832 ;
  assign y8604 = ~n8349 ;
  assign y8605 = n18839 ;
  assign y8606 = ~n18842 ;
  assign y8607 = n18849 ;
  assign y8608 = ~n18850 ;
  assign y8609 = ~1'b0 ;
  assign y8610 = ~1'b0 ;
  assign y8611 = ~n18852 ;
  assign y8612 = 1'b0 ;
  assign y8613 = ~n18855 ;
  assign y8614 = ~n18857 ;
  assign y8615 = ~n18859 ;
  assign y8616 = n18861 ;
  assign y8617 = ~n18865 ;
  assign y8618 = n18866 ;
  assign y8619 = n18867 ;
  assign y8620 = ~n18868 ;
  assign y8621 = ~n18873 ;
  assign y8622 = ~1'b0 ;
  assign y8623 = ~1'b0 ;
  assign y8624 = n15887 ;
  assign y8625 = n18875 ;
  assign y8626 = n18879 ;
  assign y8627 = ~n5567 ;
  assign y8628 = ~n18885 ;
  assign y8629 = ~1'b0 ;
  assign y8630 = n18893 ;
  assign y8631 = ~1'b0 ;
  assign y8632 = n18894 ;
  assign y8633 = n18895 ;
  assign y8634 = n18898 ;
  assign y8635 = ~1'b0 ;
  assign y8636 = ~n18903 ;
  assign y8637 = n18905 ;
  assign y8638 = ~1'b0 ;
  assign y8639 = ~n18906 ;
  assign y8640 = ~1'b0 ;
  assign y8641 = ~1'b0 ;
  assign y8642 = ~n18907 ;
  assign y8643 = ~1'b0 ;
  assign y8644 = ~n18913 ;
  assign y8645 = ~n18917 ;
  assign y8646 = ~n18920 ;
  assign y8647 = n18921 ;
  assign y8648 = ~1'b0 ;
  assign y8649 = ~n18922 ;
  assign y8650 = n18927 ;
  assign y8651 = ~1'b0 ;
  assign y8652 = ~n18932 ;
  assign y8653 = ~1'b0 ;
  assign y8654 = n18940 ;
  assign y8655 = n18941 ;
  assign y8656 = ~n18942 ;
  assign y8657 = n18943 ;
  assign y8658 = ~n18948 ;
  assign y8659 = n18954 ;
  assign y8660 = ~n18957 ;
  assign y8661 = ~n18965 ;
  assign y8662 = n18967 ;
  assign y8663 = n18974 ;
  assign y8664 = ~n18976 ;
  assign y8665 = n18977 ;
  assign y8666 = n2106 ;
  assign y8667 = n18980 ;
  assign y8668 = n18987 ;
  assign y8669 = ~n18988 ;
  assign y8670 = ~n18989 ;
  assign y8671 = ~n18990 ;
  assign y8672 = ~1'b0 ;
  assign y8673 = ~1'b0 ;
  assign y8674 = ~1'b0 ;
  assign y8675 = n2505 ;
  assign y8676 = ~1'b0 ;
  assign y8677 = n18993 ;
  assign y8678 = ~n18997 ;
  assign y8679 = ~1'b0 ;
  assign y8680 = ~1'b0 ;
  assign y8681 = ~n18998 ;
  assign y8682 = ~1'b0 ;
  assign y8683 = n18999 ;
  assign y8684 = ~n19001 ;
  assign y8685 = n19004 ;
  assign y8686 = n19006 ;
  assign y8687 = ~n19009 ;
  assign y8688 = ~n19010 ;
  assign y8689 = n19011 ;
  assign y8690 = n19013 ;
  assign y8691 = ~1'b0 ;
  assign y8692 = ~n19018 ;
  assign y8693 = n19022 ;
  assign y8694 = ~1'b0 ;
  assign y8695 = n9575 ;
  assign y8696 = n19025 ;
  assign y8697 = ~n19027 ;
  assign y8698 = n19034 ;
  assign y8699 = ~1'b0 ;
  assign y8700 = n19039 ;
  assign y8701 = n16357 ;
  assign y8702 = n19041 ;
  assign y8703 = ~1'b0 ;
  assign y8704 = ~n19043 ;
  assign y8705 = 1'b0 ;
  assign y8706 = ~n19044 ;
  assign y8707 = ~n19048 ;
  assign y8708 = ~n9005 ;
  assign y8709 = ~1'b0 ;
  assign y8710 = n19050 ;
  assign y8711 = n9865 ;
  assign y8712 = n19051 ;
  assign y8713 = ~n19052 ;
  assign y8714 = n19059 ;
  assign y8715 = ~n19062 ;
  assign y8716 = n19065 ;
  assign y8717 = n19066 ;
  assign y8718 = n19068 ;
  assign y8719 = ~n19071 ;
  assign y8720 = n19073 ;
  assign y8721 = n19074 ;
  assign y8722 = ~n19077 ;
  assign y8723 = ~1'b0 ;
  assign y8724 = n9982 ;
  assign y8725 = ~n19078 ;
  assign y8726 = n19080 ;
  assign y8727 = n5032 ;
  assign y8728 = 1'b0 ;
  assign y8729 = ~n19082 ;
  assign y8730 = n19083 ;
  assign y8731 = ~n19085 ;
  assign y8732 = ~n19091 ;
  assign y8733 = ~1'b0 ;
  assign y8734 = 1'b0 ;
  assign y8735 = ~1'b0 ;
  assign y8736 = ~n19096 ;
  assign y8737 = ~n19099 ;
  assign y8738 = ~n19101 ;
  assign y8739 = ~1'b0 ;
  assign y8740 = n19102 ;
  assign y8741 = ~n19115 ;
  assign y8742 = ~n19116 ;
  assign y8743 = n19122 ;
  assign y8744 = n19125 ;
  assign y8745 = ~n19127 ;
  assign y8746 = ~n19128 ;
  assign y8747 = ~n19129 ;
  assign y8748 = n15713 ;
  assign y8749 = ~n19132 ;
  assign y8750 = ~n19133 ;
  assign y8751 = n19134 ;
  assign y8752 = n19137 ;
  assign y8753 = ~1'b0 ;
  assign y8754 = n19139 ;
  assign y8755 = ~1'b0 ;
  assign y8756 = ~n19140 ;
  assign y8757 = ~n19141 ;
  assign y8758 = ~n19145 ;
  assign y8759 = ~1'b0 ;
  assign y8760 = ~n19146 ;
  assign y8761 = ~n19151 ;
  assign y8762 = ~1'b0 ;
  assign y8763 = ~1'b0 ;
  assign y8764 = ~n19156 ;
  assign y8765 = ~1'b0 ;
  assign y8766 = ~1'b0 ;
  assign y8767 = ~1'b0 ;
  assign y8768 = ~n9144 ;
  assign y8769 = 1'b0 ;
  assign y8770 = n19157 ;
  assign y8771 = ~n19158 ;
  assign y8772 = ~1'b0 ;
  assign y8773 = 1'b0 ;
  assign y8774 = n19160 ;
  assign y8775 = n19163 ;
  assign y8776 = n19166 ;
  assign y8777 = ~1'b0 ;
  assign y8778 = ~n7230 ;
  assign y8779 = ~n19167 ;
  assign y8780 = n19168 ;
  assign y8781 = n19169 ;
  assign y8782 = ~n19170 ;
  assign y8783 = ~1'b0 ;
  assign y8784 = ~n10701 ;
  assign y8785 = ~n15105 ;
  assign y8786 = ~1'b0 ;
  assign y8787 = ~n19172 ;
  assign y8788 = ~1'b0 ;
  assign y8789 = ~n19174 ;
  assign y8790 = n19182 ;
  assign y8791 = n19185 ;
  assign y8792 = ~n19186 ;
  assign y8793 = ~n19191 ;
  assign y8794 = ~n19194 ;
  assign y8795 = ~1'b0 ;
  assign y8796 = ~1'b0 ;
  assign y8797 = ~1'b0 ;
  assign y8798 = n19198 ;
  assign y8799 = n19200 ;
  assign y8800 = ~n19212 ;
  assign y8801 = n19213 ;
  assign y8802 = ~1'b0 ;
  assign y8803 = ~1'b0 ;
  assign y8804 = ~n19214 ;
  assign y8805 = n19234 ;
  assign y8806 = n19237 ;
  assign y8807 = n19239 ;
  assign y8808 = ~1'b0 ;
  assign y8809 = n19244 ;
  assign y8810 = ~n19248 ;
  assign y8811 = ~1'b0 ;
  assign y8812 = ~1'b0 ;
  assign y8813 = ~n19249 ;
  assign y8814 = ~n19250 ;
  assign y8815 = n19252 ;
  assign y8816 = ~n19253 ;
  assign y8817 = ~n19255 ;
  assign y8818 = n19257 ;
  assign y8819 = n19260 ;
  assign y8820 = ~1'b0 ;
  assign y8821 = ~n19262 ;
  assign y8822 = ~1'b0 ;
  assign y8823 = n19268 ;
  assign y8824 = ~1'b0 ;
  assign y8825 = n19270 ;
  assign y8826 = ~n1781 ;
  assign y8827 = n3448 ;
  assign y8828 = ~1'b0 ;
  assign y8829 = n19275 ;
  assign y8830 = n19276 ;
  assign y8831 = ~n19279 ;
  assign y8832 = n19280 ;
  assign y8833 = ~n19282 ;
  assign y8834 = ~1'b0 ;
  assign y8835 = n19285 ;
  assign y8836 = ~n19286 ;
  assign y8837 = ~n19289 ;
  assign y8838 = ~n19291 ;
  assign y8839 = ~n19294 ;
  assign y8840 = ~n19296 ;
  assign y8841 = ~n19297 ;
  assign y8842 = n19298 ;
  assign y8843 = ~n19300 ;
  assign y8844 = n19304 ;
  assign y8845 = ~n19308 ;
  assign y8846 = ~1'b0 ;
  assign y8847 = ~1'b0 ;
  assign y8848 = n19311 ;
  assign y8849 = n19312 ;
  assign y8850 = n19313 ;
  assign y8851 = ~n19314 ;
  assign y8852 = ~1'b0 ;
  assign y8853 = ~1'b0 ;
  assign y8854 = ~n19320 ;
  assign y8855 = n19322 ;
  assign y8856 = n19323 ;
  assign y8857 = n19326 ;
  assign y8858 = ~n19328 ;
  assign y8859 = n18794 ;
  assign y8860 = ~n19329 ;
  assign y8861 = n19330 ;
  assign y8862 = ~1'b0 ;
  assign y8863 = n19333 ;
  assign y8864 = ~1'b0 ;
  assign y8865 = ~n19337 ;
  assign y8866 = ~n19340 ;
  assign y8867 = n19341 ;
  assign y8868 = ~n19343 ;
  assign y8869 = ~1'b0 ;
  assign y8870 = n19344 ;
  assign y8871 = ~n19347 ;
  assign y8872 = ~n19348 ;
  assign y8873 = n19353 ;
  assign y8874 = ~n19356 ;
  assign y8875 = ~n19358 ;
  assign y8876 = n19359 ;
  assign y8877 = ~n19361 ;
  assign y8878 = ~1'b0 ;
  assign y8879 = n19366 ;
  assign y8880 = ~n19367 ;
  assign y8881 = n19370 ;
  assign y8882 = ~n19371 ;
  assign y8883 = ~n19375 ;
  assign y8884 = n19376 ;
  assign y8885 = ~1'b0 ;
  assign y8886 = n19377 ;
  assign y8887 = ~n19382 ;
  assign y8888 = ~n19383 ;
  assign y8889 = ~n19384 ;
  assign y8890 = ~1'b0 ;
  assign y8891 = ~n19386 ;
  assign y8892 = n19387 ;
  assign y8893 = n19390 ;
  assign y8894 = n19392 ;
  assign y8895 = ~n5275 ;
  assign y8896 = ~n19395 ;
  assign y8897 = n19396 ;
  assign y8898 = ~n19398 ;
  assign y8899 = ~n6148 ;
  assign y8900 = n19401 ;
  assign y8901 = ~n19403 ;
  assign y8902 = ~n19407 ;
  assign y8903 = ~1'b0 ;
  assign y8904 = ~n19412 ;
  assign y8905 = ~1'b0 ;
  assign y8906 = ~1'b0 ;
  assign y8907 = ~n19418 ;
  assign y8908 = ~n19420 ;
  assign y8909 = n8771 ;
  assign y8910 = n19424 ;
  assign y8911 = ~n19426 ;
  assign y8912 = n19428 ;
  assign y8913 = ~1'b0 ;
  assign y8914 = n19431 ;
  assign y8915 = n19432 ;
  assign y8916 = n19433 ;
  assign y8917 = n19437 ;
  assign y8918 = ~1'b0 ;
  assign y8919 = ~1'b0 ;
  assign y8920 = n19438 ;
  assign y8921 = ~1'b0 ;
  assign y8922 = ~1'b0 ;
  assign y8923 = n19264 ;
  assign y8924 = n19439 ;
  assign y8925 = ~n19441 ;
  assign y8926 = ~n4222 ;
  assign y8927 = ~n19446 ;
  assign y8928 = ~n19450 ;
  assign y8929 = 1'b0 ;
  assign y8930 = ~1'b0 ;
  assign y8931 = ~1'b0 ;
  assign y8932 = ~n19453 ;
  assign y8933 = ~n19456 ;
  assign y8934 = n19459 ;
  assign y8935 = n19461 ;
  assign y8936 = 1'b0 ;
  assign y8937 = ~1'b0 ;
  assign y8938 = n19462 ;
  assign y8939 = ~n19465 ;
  assign y8940 = n19466 ;
  assign y8941 = n19469 ;
  assign y8942 = ~n19471 ;
  assign y8943 = ~1'b0 ;
  assign y8944 = ~n19472 ;
  assign y8945 = ~1'b0 ;
  assign y8946 = ~n19474 ;
  assign y8947 = ~n19476 ;
  assign y8948 = ~1'b0 ;
  assign y8949 = ~1'b0 ;
  assign y8950 = n19477 ;
  assign y8951 = ~n19480 ;
  assign y8952 = ~n19484 ;
  assign y8953 = ~n19487 ;
  assign y8954 = ~n19490 ;
  assign y8955 = n19492 ;
  assign y8956 = ~n19493 ;
  assign y8957 = 1'b0 ;
  assign y8958 = ~1'b0 ;
  assign y8959 = ~n19494 ;
  assign y8960 = n19496 ;
  assign y8961 = n19504 ;
  assign y8962 = n19506 ;
  assign y8963 = ~n19511 ;
  assign y8964 = ~n19512 ;
  assign y8965 = ~1'b0 ;
  assign y8966 = ~1'b0 ;
  assign y8967 = ~n19515 ;
  assign y8968 = ~n19521 ;
  assign y8969 = n19522 ;
  assign y8970 = ~n19524 ;
  assign y8971 = n19528 ;
  assign y8972 = ~n18502 ;
  assign y8973 = n19529 ;
  assign y8974 = ~n19533 ;
  assign y8975 = ~1'b0 ;
  assign y8976 = n19537 ;
  assign y8977 = n19539 ;
  assign y8978 = n19540 ;
  assign y8979 = n19542 ;
  assign y8980 = n19545 ;
  assign y8981 = ~n19547 ;
  assign y8982 = ~1'b0 ;
  assign y8983 = ~1'b0 ;
  assign y8984 = 1'b0 ;
  assign y8985 = 1'b0 ;
  assign y8986 = ~n19551 ;
  assign y8987 = ~n19552 ;
  assign y8988 = ~1'b0 ;
  assign y8989 = n19554 ;
  assign y8990 = n19563 ;
  assign y8991 = ~1'b0 ;
  assign y8992 = n19565 ;
  assign y8993 = ~n19567 ;
  assign y8994 = n19573 ;
  assign y8995 = n9307 ;
  assign y8996 = n19576 ;
  assign y8997 = n19578 ;
  assign y8998 = ~n19586 ;
  assign y8999 = n19589 ;
  assign y9000 = n19595 ;
  assign y9001 = ~1'b0 ;
  assign y9002 = ~1'b0 ;
  assign y9003 = n19606 ;
  assign y9004 = ~1'b0 ;
  assign y9005 = ~n19607 ;
  assign y9006 = ~n6350 ;
  assign y9007 = ~n19608 ;
  assign y9008 = ~1'b0 ;
  assign y9009 = n19609 ;
  assign y9010 = ~1'b0 ;
  assign y9011 = ~n19611 ;
  assign y9012 = ~1'b0 ;
  assign y9013 = n19612 ;
  assign y9014 = ~n17790 ;
  assign y9015 = ~n19616 ;
  assign y9016 = ~n18632 ;
  assign y9017 = ~n19618 ;
  assign y9018 = ~1'b0 ;
  assign y9019 = n19620 ;
  assign y9020 = n19622 ;
  assign y9021 = n17052 ;
  assign y9022 = ~n19624 ;
  assign y9023 = ~n19625 ;
  assign y9024 = ~n19627 ;
  assign y9025 = n19628 ;
  assign y9026 = ~n19633 ;
  assign y9027 = ~n19638 ;
  assign y9028 = n19640 ;
  assign y9029 = ~1'b0 ;
  assign y9030 = ~n5721 ;
  assign y9031 = n19647 ;
  assign y9032 = n19648 ;
  assign y9033 = n19650 ;
  assign y9034 = n16835 ;
  assign y9035 = ~1'b0 ;
  assign y9036 = n19654 ;
  assign y9037 = ~1'b0 ;
  assign y9038 = ~1'b0 ;
  assign y9039 = ~n19656 ;
  assign y9040 = n19659 ;
  assign y9041 = n19664 ;
  assign y9042 = ~1'b0 ;
  assign y9043 = n19665 ;
  assign y9044 = ~n19670 ;
  assign y9045 = ~n19671 ;
  assign y9046 = ~n19673 ;
  assign y9047 = ~n19674 ;
  assign y9048 = n19676 ;
  assign y9049 = n19685 ;
  assign y9050 = ~1'b0 ;
  assign y9051 = ~n19686 ;
  assign y9052 = ~n2091 ;
  assign y9053 = n19687 ;
  assign y9054 = ~n19689 ;
  assign y9055 = ~n19690 ;
  assign y9056 = ~1'b0 ;
  assign y9057 = n19695 ;
  assign y9058 = ~n19696 ;
  assign y9059 = ~1'b0 ;
  assign y9060 = ~n16876 ;
  assign y9061 = ~1'b0 ;
  assign y9062 = ~1'b0 ;
  assign y9063 = ~n19698 ;
  assign y9064 = ~n14107 ;
  assign y9065 = ~n19701 ;
  assign y9066 = n19704 ;
  assign y9067 = n19712 ;
  assign y9068 = n19713 ;
  assign y9069 = ~1'b0 ;
  assign y9070 = n19715 ;
  assign y9071 = n19717 ;
  assign y9072 = ~n19720 ;
  assign y9073 = n19721 ;
  assign y9074 = n3037 ;
  assign y9075 = ~1'b0 ;
  assign y9076 = ~1'b0 ;
  assign y9077 = ~n19722 ;
  assign y9078 = n19723 ;
  assign y9079 = ~1'b0 ;
  assign y9080 = ~n19728 ;
  assign y9081 = n19731 ;
  assign y9082 = n19734 ;
  assign y9083 = n19735 ;
  assign y9084 = n11178 ;
  assign y9085 = n19736 ;
  assign y9086 = ~1'b0 ;
  assign y9087 = n19739 ;
  assign y9088 = ~n19741 ;
  assign y9089 = n19743 ;
  assign y9090 = ~n19744 ;
  assign y9091 = n19754 ;
  assign y9092 = n19756 ;
  assign y9093 = ~n19759 ;
  assign y9094 = n19763 ;
  assign y9095 = n19767 ;
  assign y9096 = n19774 ;
  assign y9097 = n285 ;
  assign y9098 = n19779 ;
  assign y9099 = n19780 ;
  assign y9100 = ~1'b0 ;
  assign y9101 = n19782 ;
  assign y9102 = ~n19784 ;
  assign y9103 = ~1'b0 ;
  assign y9104 = ~1'b0 ;
  assign y9105 = n19785 ;
  assign y9106 = ~n19786 ;
  assign y9107 = ~n19787 ;
  assign y9108 = ~n19792 ;
  assign y9109 = n19799 ;
  assign y9110 = ~1'b0 ;
  assign y9111 = ~n19800 ;
  assign y9112 = n19801 ;
  assign y9113 = n19802 ;
  assign y9114 = ~1'b0 ;
  assign y9115 = ~1'b0 ;
  assign y9116 = ~1'b0 ;
  assign y9117 = ~1'b0 ;
  assign y9118 = n19803 ;
  assign y9119 = n19805 ;
  assign y9120 = ~n19807 ;
  assign y9121 = ~1'b0 ;
  assign y9122 = n19808 ;
  assign y9123 = n19809 ;
  assign y9124 = ~n3113 ;
  assign y9125 = ~1'b0 ;
  assign y9126 = n19810 ;
  assign y9127 = n19811 ;
  assign y9128 = ~n19817 ;
  assign y9129 = ~n19818 ;
  assign y9130 = n19824 ;
  assign y9131 = ~n19825 ;
  assign y9132 = ~n19827 ;
  assign y9133 = ~n19829 ;
  assign y9134 = ~1'b0 ;
  assign y9135 = n19834 ;
  assign y9136 = ~n19837 ;
  assign y9137 = n19838 ;
  assign y9138 = ~n19839 ;
  assign y9139 = ~1'b0 ;
  assign y9140 = ~n19841 ;
  assign y9141 = n19843 ;
  assign y9142 = ~n19845 ;
  assign y9143 = n19848 ;
  assign y9144 = ~n19854 ;
  assign y9145 = n19856 ;
  assign y9146 = ~n19859 ;
  assign y9147 = ~n19861 ;
  assign y9148 = n4336 ;
  assign y9149 = ~n19863 ;
  assign y9150 = ~n19865 ;
  assign y9151 = n19867 ;
  assign y9152 = ~n19868 ;
  assign y9153 = ~n19870 ;
  assign y9154 = n19874 ;
  assign y9155 = ~1'b0 ;
  assign y9156 = ~n19875 ;
  assign y9157 = ~n19879 ;
  assign y9158 = ~n19880 ;
  assign y9159 = n19883 ;
  assign y9160 = ~n17815 ;
  assign y9161 = ~1'b0 ;
  assign y9162 = ~1'b0 ;
  assign y9163 = ~n19889 ;
  assign y9164 = ~1'b0 ;
  assign y9165 = ~1'b0 ;
  assign y9166 = n19891 ;
  assign y9167 = ~1'b0 ;
  assign y9168 = n19893 ;
  assign y9169 = ~1'b0 ;
  assign y9170 = ~n19897 ;
  assign y9171 = ~n19899 ;
  assign y9172 = ~n2253 ;
  assign y9173 = n19900 ;
  assign y9174 = ~n19903 ;
  assign y9175 = ~1'b0 ;
  assign y9176 = n19904 ;
  assign y9177 = n19905 ;
  assign y9178 = n19913 ;
  assign y9179 = ~n19915 ;
  assign y9180 = n19917 ;
  assign y9181 = ~n19918 ;
  assign y9182 = ~n19920 ;
  assign y9183 = ~n12843 ;
  assign y9184 = n19922 ;
  assign y9185 = ~n19923 ;
  assign y9186 = n19924 ;
  assign y9187 = ~1'b0 ;
  assign y9188 = n19925 ;
  assign y9189 = n19928 ;
  assign y9190 = n19930 ;
  assign y9191 = n19936 ;
  assign y9192 = n19940 ;
  assign y9193 = n19941 ;
  assign y9194 = ~1'b0 ;
  assign y9195 = ~n19942 ;
  assign y9196 = ~n19949 ;
  assign y9197 = ~n19952 ;
  assign y9198 = n19958 ;
  assign y9199 = ~n19963 ;
  assign y9200 = ~1'b0 ;
  assign y9201 = n19965 ;
  assign y9202 = ~1'b0 ;
  assign y9203 = ~1'b0 ;
  assign y9204 = ~n19966 ;
  assign y9205 = n19967 ;
  assign y9206 = ~n19968 ;
  assign y9207 = ~n19970 ;
  assign y9208 = ~n19972 ;
  assign y9209 = ~n19973 ;
  assign y9210 = ~1'b0 ;
  assign y9211 = n19974 ;
  assign y9212 = ~1'b0 ;
  assign y9213 = ~n19976 ;
  assign y9214 = n19983 ;
  assign y9215 = ~n19986 ;
  assign y9216 = ~n19988 ;
  assign y9217 = n19990 ;
  assign y9218 = ~n4085 ;
  assign y9219 = n19999 ;
  assign y9220 = ~1'b0 ;
  assign y9221 = ~n20000 ;
  assign y9222 = n20005 ;
  assign y9223 = ~1'b0 ;
  assign y9224 = n20009 ;
  assign y9225 = ~n20010 ;
  assign y9226 = ~1'b0 ;
  assign y9227 = ~n20012 ;
  assign y9228 = 1'b0 ;
  assign y9229 = ~1'b0 ;
  assign y9230 = ~1'b0 ;
  assign y9231 = ~n20014 ;
  assign y9232 = ~1'b0 ;
  assign y9233 = ~n20016 ;
  assign y9234 = ~1'b0 ;
  assign y9235 = ~1'b0 ;
  assign y9236 = ~n10626 ;
  assign y9237 = n20017 ;
  assign y9238 = n20018 ;
  assign y9239 = ~n20019 ;
  assign y9240 = ~n20023 ;
  assign y9241 = n20024 ;
  assign y9242 = ~n20027 ;
  assign y9243 = ~n20031 ;
  assign y9244 = ~1'b0 ;
  assign y9245 = ~1'b0 ;
  assign y9246 = ~n20033 ;
  assign y9247 = ~n20039 ;
  assign y9248 = n20041 ;
  assign y9249 = ~1'b0 ;
  assign y9250 = n20044 ;
  assign y9251 = n20045 ;
  assign y9252 = ~n20048 ;
  assign y9253 = ~1'b0 ;
  assign y9254 = n20052 ;
  assign y9255 = n20053 ;
  assign y9256 = ~n1683 ;
  assign y9257 = ~1'b0 ;
  assign y9258 = n20060 ;
  assign y9259 = ~n20069 ;
  assign y9260 = n20072 ;
  assign y9261 = ~n20074 ;
  assign y9262 = n20076 ;
  assign y9263 = n20079 ;
  assign y9264 = ~n20081 ;
  assign y9265 = ~n20082 ;
  assign y9266 = n20084 ;
  assign y9267 = ~n20086 ;
  assign y9268 = n20090 ;
  assign y9269 = ~n20092 ;
  assign y9270 = ~n3631 ;
  assign y9271 = n20095 ;
  assign y9272 = ~1'b0 ;
  assign y9273 = ~n20097 ;
  assign y9274 = ~n20100 ;
  assign y9275 = n20101 ;
  assign y9276 = ~1'b0 ;
  assign y9277 = ~n20109 ;
  assign y9278 = n20115 ;
  assign y9279 = ~n20117 ;
  assign y9280 = ~n20119 ;
  assign y9281 = n20123 ;
  assign y9282 = ~n20124 ;
  assign y9283 = n20125 ;
  assign y9284 = ~1'b0 ;
  assign y9285 = n20134 ;
  assign y9286 = n20138 ;
  assign y9287 = n20139 ;
  assign y9288 = n20143 ;
  assign y9289 = ~n20148 ;
  assign y9290 = ~n20149 ;
  assign y9291 = ~1'b0 ;
  assign y9292 = n20150 ;
  assign y9293 = ~n20154 ;
  assign y9294 = n20156 ;
  assign y9295 = n20157 ;
  assign y9296 = ~n20160 ;
  assign y9297 = ~1'b0 ;
  assign y9298 = ~n20163 ;
  assign y9299 = ~n20169 ;
  assign y9300 = ~1'b0 ;
  assign y9301 = ~n20170 ;
  assign y9302 = ~n20171 ;
  assign y9303 = ~1'b0 ;
  assign y9304 = n20176 ;
  assign y9305 = n20181 ;
  assign y9306 = n20193 ;
  assign y9307 = n20195 ;
  assign y9308 = ~1'b0 ;
  assign y9309 = ~n20196 ;
  assign y9310 = ~n20197 ;
  assign y9311 = ~n20204 ;
  assign y9312 = n20207 ;
  assign y9313 = ~n20208 ;
  assign y9314 = n20209 ;
  assign y9315 = ~1'b0 ;
  assign y9316 = ~n20211 ;
  assign y9317 = ~n20213 ;
  assign y9318 = n20217 ;
  assign y9319 = ~1'b0 ;
  assign y9320 = n20220 ;
  assign y9321 = n20221 ;
  assign y9322 = ~n15555 ;
  assign y9323 = ~1'b0 ;
  assign y9324 = ~n20223 ;
  assign y9325 = ~n20225 ;
  assign y9326 = ~n20227 ;
  assign y9327 = ~n20229 ;
  assign y9328 = ~1'b0 ;
  assign y9329 = ~1'b0 ;
  assign y9330 = ~n20230 ;
  assign y9331 = n20233 ;
  assign y9332 = n20235 ;
  assign y9333 = ~n20236 ;
  assign y9334 = n20237 ;
  assign y9335 = n20238 ;
  assign y9336 = n20241 ;
  assign y9337 = ~n20243 ;
  assign y9338 = ~1'b0 ;
  assign y9339 = ~n20245 ;
  assign y9340 = ~n20248 ;
  assign y9341 = n20250 ;
  assign y9342 = 1'b0 ;
  assign y9343 = ~1'b0 ;
  assign y9344 = n20254 ;
  assign y9345 = n20255 ;
  assign y9346 = n20258 ;
  assign y9347 = n20261 ;
  assign y9348 = ~n20265 ;
  assign y9349 = n9797 ;
  assign y9350 = n20268 ;
  assign y9351 = ~1'b0 ;
  assign y9352 = n20270 ;
  assign y9353 = ~1'b0 ;
  assign y9354 = ~1'b0 ;
  assign y9355 = ~n20271 ;
  assign y9356 = ~n20273 ;
  assign y9357 = ~n20275 ;
  assign y9358 = n20277 ;
  assign y9359 = n20281 ;
  assign y9360 = ~1'b0 ;
  assign y9361 = n5758 ;
  assign y9362 = n20286 ;
  assign y9363 = ~1'b0 ;
  assign y9364 = ~n20292 ;
  assign y9365 = ~n20294 ;
  assign y9366 = n20295 ;
  assign y9367 = n20296 ;
  assign y9368 = ~1'b0 ;
  assign y9369 = ~n20298 ;
  assign y9370 = ~1'b0 ;
  assign y9371 = ~n20305 ;
  assign y9372 = n20307 ;
  assign y9373 = 1'b0 ;
  assign y9374 = ~1'b0 ;
  assign y9375 = ~1'b0 ;
  assign y9376 = n20308 ;
  assign y9377 = n20310 ;
  assign y9378 = n20313 ;
  assign y9379 = n20314 ;
  assign y9380 = ~n20318 ;
  assign y9381 = ~n20321 ;
  assign y9382 = ~n20325 ;
  assign y9383 = n18796 ;
  assign y9384 = ~n20328 ;
  assign y9385 = ~n20329 ;
  assign y9386 = ~n20332 ;
  assign y9387 = n20335 ;
  assign y9388 = ~n20339 ;
  assign y9389 = ~n20341 ;
  assign y9390 = ~n20344 ;
  assign y9391 = n20345 ;
  assign y9392 = ~n20347 ;
  assign y9393 = ~1'b0 ;
  assign y9394 = ~n20352 ;
  assign y9395 = ~1'b0 ;
  assign y9396 = n20354 ;
  assign y9397 = ~1'b0 ;
  assign y9398 = ~1'b0 ;
  assign y9399 = ~1'b0 ;
  assign y9400 = ~1'b0 ;
  assign y9401 = ~n20355 ;
  assign y9402 = n20356 ;
  assign y9403 = n20359 ;
  assign y9404 = n20361 ;
  assign y9405 = ~1'b0 ;
  assign y9406 = n20363 ;
  assign y9407 = n20364 ;
  assign y9408 = ~n20365 ;
  assign y9409 = ~n20369 ;
  assign y9410 = n20371 ;
  assign y9411 = n20389 ;
  assign y9412 = ~n7139 ;
  assign y9413 = n20390 ;
  assign y9414 = ~n20394 ;
  assign y9415 = ~1'b0 ;
  assign y9416 = ~n20397 ;
  assign y9417 = ~n20398 ;
  assign y9418 = n14340 ;
  assign y9419 = n20399 ;
  assign y9420 = n20400 ;
  assign y9421 = ~n20403 ;
  assign y9422 = ~n20405 ;
  assign y9423 = n20410 ;
  assign y9424 = n17560 ;
  assign y9425 = n20411 ;
  assign y9426 = ~n20414 ;
  assign y9427 = ~1'b0 ;
  assign y9428 = n20418 ;
  assign y9429 = ~1'b0 ;
  assign y9430 = n20419 ;
  assign y9431 = n20420 ;
  assign y9432 = ~n20425 ;
  assign y9433 = ~n20426 ;
  assign y9434 = ~n20430 ;
  assign y9435 = n20435 ;
  assign y9436 = ~n20436 ;
  assign y9437 = ~1'b0 ;
  assign y9438 = ~n20439 ;
  assign y9439 = n20441 ;
  assign y9440 = ~n20442 ;
  assign y9441 = ~1'b0 ;
  assign y9442 = ~1'b0 ;
  assign y9443 = ~1'b0 ;
  assign y9444 = n20445 ;
  assign y9445 = n20448 ;
  assign y9446 = ~1'b0 ;
  assign y9447 = n20449 ;
  assign y9448 = n15432 ;
  assign y9449 = ~1'b0 ;
  assign y9450 = ~1'b0 ;
  assign y9451 = n20454 ;
  assign y9452 = ~1'b0 ;
  assign y9453 = n20457 ;
  assign y9454 = n20458 ;
  assign y9455 = ~n20459 ;
  assign y9456 = n20467 ;
  assign y9457 = n20468 ;
  assign y9458 = ~1'b0 ;
  assign y9459 = ~1'b0 ;
  assign y9460 = ~1'b0 ;
  assign y9461 = n20470 ;
  assign y9462 = ~n20474 ;
  assign y9463 = n20476 ;
  assign y9464 = n20479 ;
  assign y9465 = ~n20481 ;
  assign y9466 = ~1'b0 ;
  assign y9467 = ~1'b0 ;
  assign y9468 = ~n20494 ;
  assign y9469 = n20495 ;
  assign y9470 = ~n20499 ;
  assign y9471 = ~n20504 ;
  assign y9472 = n20511 ;
  assign y9473 = ~1'b0 ;
  assign y9474 = ~n20512 ;
  assign y9475 = n20515 ;
  assign y9476 = n20516 ;
  assign y9477 = n20517 ;
  assign y9478 = ~n1366 ;
  assign y9479 = ~n20519 ;
  assign y9480 = n20520 ;
  assign y9481 = ~1'b0 ;
  assign y9482 = n20521 ;
  assign y9483 = n20522 ;
  assign y9484 = n20523 ;
  assign y9485 = n5647 ;
  assign y9486 = ~n20524 ;
  assign y9487 = n20526 ;
  assign y9488 = n20530 ;
  assign y9489 = ~n20532 ;
  assign y9490 = ~1'b0 ;
  assign y9491 = n20534 ;
  assign y9492 = ~n20535 ;
  assign y9493 = ~n20537 ;
  assign y9494 = ~1'b0 ;
  assign y9495 = n20540 ;
  assign y9496 = n20542 ;
  assign y9497 = n20544 ;
  assign y9498 = n20546 ;
  assign y9499 = n20547 ;
  assign y9500 = n20552 ;
  assign y9501 = ~n20557 ;
  assign y9502 = ~n20561 ;
  assign y9503 = ~n7562 ;
  assign y9504 = 1'b0 ;
  assign y9505 = ~n20562 ;
  assign y9506 = ~1'b0 ;
  assign y9507 = ~1'b0 ;
  assign y9508 = ~n20568 ;
  assign y9509 = ~n20572 ;
  assign y9510 = ~1'b0 ;
  assign y9511 = ~1'b0 ;
  assign y9512 = ~n20573 ;
  assign y9513 = ~n20574 ;
  assign y9514 = ~n20581 ;
  assign y9515 = ~n20584 ;
  assign y9516 = ~n20587 ;
  assign y9517 = ~n20588 ;
  assign y9518 = n20589 ;
  assign y9519 = ~1'b0 ;
  assign y9520 = n20594 ;
  assign y9521 = ~n20596 ;
  assign y9522 = ~1'b0 ;
  assign y9523 = n20597 ;
  assign y9524 = ~n20598 ;
  assign y9525 = n20603 ;
  assign y9526 = n20608 ;
  assign y9527 = ~n20612 ;
  assign y9528 = ~n19169 ;
  assign y9529 = n20613 ;
  assign y9530 = ~n4342 ;
  assign y9531 = ~n20616 ;
  assign y9532 = ~n20619 ;
  assign y9533 = ~1'b0 ;
  assign y9534 = ~1'b0 ;
  assign y9535 = ~n20626 ;
  assign y9536 = ~1'b0 ;
  assign y9537 = ~1'b0 ;
  assign y9538 = ~n20630 ;
  assign y9539 = n9031 ;
  assign y9540 = ~1'b0 ;
  assign y9541 = n20633 ;
  assign y9542 = ~n20634 ;
  assign y9543 = ~1'b0 ;
  assign y9544 = n20635 ;
  assign y9545 = n20636 ;
  assign y9546 = ~n11043 ;
  assign y9547 = ~1'b0 ;
  assign y9548 = n20639 ;
  assign y9549 = n20641 ;
  assign y9550 = n20642 ;
  assign y9551 = ~1'b0 ;
  assign y9552 = ~n20646 ;
  assign y9553 = ~n20648 ;
  assign y9554 = n20652 ;
  assign y9555 = ~n20653 ;
  assign y9556 = ~n20654 ;
  assign y9557 = x16 ;
  assign y9558 = ~n20656 ;
  assign y9559 = ~1'b0 ;
  assign y9560 = ~n18920 ;
  assign y9561 = n20659 ;
  assign y9562 = n20663 ;
  assign y9563 = n20665 ;
  assign y9564 = ~1'b0 ;
  assign y9565 = ~n20670 ;
  assign y9566 = n20671 ;
  assign y9567 = ~n20672 ;
  assign y9568 = ~n20674 ;
  assign y9569 = n20675 ;
  assign y9570 = ~1'b0 ;
  assign y9571 = ~n14193 ;
  assign y9572 = ~1'b0 ;
  assign y9573 = ~n20679 ;
  assign y9574 = n20680 ;
  assign y9575 = n20681 ;
  assign y9576 = ~n20684 ;
  assign y9577 = ~1'b0 ;
  assign y9578 = ~n20687 ;
  assign y9579 = ~n20692 ;
  assign y9580 = ~n20694 ;
  assign y9581 = ~n20695 ;
  assign y9582 = ~n20701 ;
  assign y9583 = n20702 ;
  assign y9584 = ~n20703 ;
  assign y9585 = 1'b0 ;
  assign y9586 = ~1'b0 ;
  assign y9587 = n20704 ;
  assign y9588 = ~n20705 ;
  assign y9589 = n20707 ;
  assign y9590 = n20708 ;
  assign y9591 = ~1'b0 ;
  assign y9592 = ~n20709 ;
  assign y9593 = n20710 ;
  assign y9594 = n20716 ;
  assign y9595 = ~n20717 ;
  assign y9596 = ~n20718 ;
  assign y9597 = ~1'b0 ;
  assign y9598 = n20719 ;
  assign y9599 = n20721 ;
  assign y9600 = ~n20722 ;
  assign y9601 = ~n20724 ;
  assign y9602 = ~n20727 ;
  assign y9603 = ~n20730 ;
  assign y9604 = ~n20732 ;
  assign y9605 = ~n20733 ;
  assign y9606 = ~n20736 ;
  assign y9607 = ~1'b0 ;
  assign y9608 = n20737 ;
  assign y9609 = n20739 ;
  assign y9610 = n20741 ;
  assign y9611 = n20742 ;
  assign y9612 = n20745 ;
  assign y9613 = ~1'b0 ;
  assign y9614 = ~n20751 ;
  assign y9615 = ~1'b0 ;
  assign y9616 = n20754 ;
  assign y9617 = n20757 ;
  assign y9618 = n20758 ;
  assign y9619 = ~1'b0 ;
  assign y9620 = ~1'b0 ;
  assign y9621 = n13799 ;
  assign y9622 = n20760 ;
  assign y9623 = ~n20762 ;
  assign y9624 = ~1'b0 ;
  assign y9625 = ~n20767 ;
  assign y9626 = n20769 ;
  assign y9627 = ~n20777 ;
  assign y9628 = ~n20778 ;
  assign y9629 = n20779 ;
  assign y9630 = ~1'b0 ;
  assign y9631 = ~1'b0 ;
  assign y9632 = n20783 ;
  assign y9633 = n9067 ;
  assign y9634 = ~1'b0 ;
  assign y9635 = ~1'b0 ;
  assign y9636 = ~1'b0 ;
  assign y9637 = n20785 ;
  assign y9638 = ~1'b0 ;
  assign y9639 = n9653 ;
  assign y9640 = n20786 ;
  assign y9641 = n20787 ;
  assign y9642 = ~n20788 ;
  assign y9643 = n20791 ;
  assign y9644 = ~1'b0 ;
  assign y9645 = ~1'b0 ;
  assign y9646 = ~1'b0 ;
  assign y9647 = ~n20794 ;
  assign y9648 = n20795 ;
  assign y9649 = ~n20796 ;
  assign y9650 = n6516 ;
  assign y9651 = n20801 ;
  assign y9652 = ~1'b0 ;
  assign y9653 = ~n20802 ;
  assign y9654 = ~n20803 ;
  assign y9655 = ~n20809 ;
  assign y9656 = ~1'b0 ;
  assign y9657 = ~1'b0 ;
  assign y9658 = ~1'b0 ;
  assign y9659 = ~n12819 ;
  assign y9660 = ~1'b0 ;
  assign y9661 = ~n20813 ;
  assign y9662 = ~n20816 ;
  assign y9663 = ~n20819 ;
  assign y9664 = n20821 ;
  assign y9665 = ~1'b0 ;
  assign y9666 = ~1'b0 ;
  assign y9667 = ~n20822 ;
  assign y9668 = ~n20825 ;
  assign y9669 = n12969 ;
  assign y9670 = ~n20827 ;
  assign y9671 = ~n20831 ;
  assign y9672 = ~1'b0 ;
  assign y9673 = n20835 ;
  assign y9674 = ~n20838 ;
  assign y9675 = n20839 ;
  assign y9676 = n20843 ;
  assign y9677 = n20844 ;
  assign y9678 = ~n20845 ;
  assign y9679 = n20847 ;
  assign y9680 = n20851 ;
  assign y9681 = ~n20853 ;
  assign y9682 = ~1'b0 ;
  assign y9683 = ~1'b0 ;
  assign y9684 = ~1'b0 ;
  assign y9685 = n20854 ;
  assign y9686 = ~n20858 ;
  assign y9687 = n20860 ;
  assign y9688 = n20861 ;
  assign y9689 = n1300 ;
  assign y9690 = ~n20862 ;
  assign y9691 = n20866 ;
  assign y9692 = n20869 ;
  assign y9693 = 1'b0 ;
  assign y9694 = 1'b0 ;
  assign y9695 = ~n20875 ;
  assign y9696 = n20876 ;
  assign y9697 = n20877 ;
  assign y9698 = ~n20881 ;
  assign y9699 = ~1'b0 ;
  assign y9700 = ~1'b0 ;
  assign y9701 = n20882 ;
  assign y9702 = ~n20887 ;
  assign y9703 = ~1'b0 ;
  assign y9704 = n20889 ;
  assign y9705 = ~1'b0 ;
  assign y9706 = n5355 ;
  assign y9707 = ~n20896 ;
  assign y9708 = ~n20899 ;
  assign y9709 = ~n20903 ;
  assign y9710 = n6553 ;
  assign y9711 = ~1'b0 ;
  assign y9712 = n20906 ;
  assign y9713 = ~1'b0 ;
  assign y9714 = ~n20912 ;
  assign y9715 = ~1'b0 ;
  assign y9716 = n20915 ;
  assign y9717 = n20918 ;
  assign y9718 = n20920 ;
  assign y9719 = n20921 ;
  assign y9720 = n20923 ;
  assign y9721 = n20925 ;
  assign y9722 = ~1'b0 ;
  assign y9723 = ~n20927 ;
  assign y9724 = ~n20929 ;
  assign y9725 = ~n20934 ;
  assign y9726 = n20935 ;
  assign y9727 = ~n20938 ;
  assign y9728 = n20941 ;
  assign y9729 = ~n2256 ;
  assign y9730 = ~1'b0 ;
  assign y9731 = n20942 ;
  assign y9732 = ~n20947 ;
  assign y9733 = ~n20950 ;
  assign y9734 = ~1'b0 ;
  assign y9735 = ~n20953 ;
  assign y9736 = n20955 ;
  assign y9737 = ~n20957 ;
  assign y9738 = ~1'b0 ;
  assign y9739 = ~n20958 ;
  assign y9740 = ~n20960 ;
  assign y9741 = n20964 ;
  assign y9742 = ~n20967 ;
  assign y9743 = ~n20968 ;
  assign y9744 = ~n20970 ;
  assign y9745 = n20971 ;
  assign y9746 = ~1'b0 ;
  assign y9747 = ~n19913 ;
  assign y9748 = n20978 ;
  assign y9749 = n20981 ;
  assign y9750 = ~n20983 ;
  assign y9751 = n20986 ;
  assign y9752 = ~n20989 ;
  assign y9753 = ~1'b0 ;
  assign y9754 = ~n2736 ;
  assign y9755 = ~n3975 ;
  assign y9756 = ~1'b0 ;
  assign y9757 = ~1'b0 ;
  assign y9758 = n20991 ;
  assign y9759 = ~n20993 ;
  assign y9760 = ~n20996 ;
  assign y9761 = ~1'b0 ;
  assign y9762 = ~1'b0 ;
  assign y9763 = ~n21001 ;
  assign y9764 = ~1'b0 ;
  assign y9765 = n12293 ;
  assign y9766 = n21003 ;
  assign y9767 = n21008 ;
  assign y9768 = n21011 ;
  assign y9769 = ~n21012 ;
  assign y9770 = ~1'b0 ;
  assign y9771 = n21013 ;
  assign y9772 = n21014 ;
  assign y9773 = n21019 ;
  assign y9774 = 1'b0 ;
  assign y9775 = ~1'b0 ;
  assign y9776 = ~n21021 ;
  assign y9777 = n21023 ;
  assign y9778 = ~1'b0 ;
  assign y9779 = n21028 ;
  assign y9780 = ~n21031 ;
  assign y9781 = ~1'b0 ;
  assign y9782 = ~n21035 ;
  assign y9783 = ~n21046 ;
  assign y9784 = n21050 ;
  assign y9785 = ~n21053 ;
  assign y9786 = ~n21056 ;
  assign y9787 = ~1'b0 ;
  assign y9788 = n21060 ;
  assign y9789 = ~1'b0 ;
  assign y9790 = n15166 ;
  assign y9791 = ~n21063 ;
  assign y9792 = n21064 ;
  assign y9793 = ~n21065 ;
  assign y9794 = ~1'b0 ;
  assign y9795 = ~n21067 ;
  assign y9796 = ~1'b0 ;
  assign y9797 = ~1'b0 ;
  assign y9798 = ~1'b0 ;
  assign y9799 = n21069 ;
  assign y9800 = ~n18449 ;
  assign y9801 = ~n21073 ;
  assign y9802 = ~1'b0 ;
  assign y9803 = n21077 ;
  assign y9804 = ~n21086 ;
  assign y9805 = ~1'b0 ;
  assign y9806 = n1135 ;
  assign y9807 = ~n21087 ;
  assign y9808 = n21088 ;
  assign y9809 = n21089 ;
  assign y9810 = ~1'b0 ;
  assign y9811 = n21090 ;
  assign y9812 = ~n21092 ;
  assign y9813 = ~1'b0 ;
  assign y9814 = ~n21095 ;
  assign y9815 = ~1'b0 ;
  assign y9816 = ~n21096 ;
  assign y9817 = ~n21099 ;
  assign y9818 = ~1'b0 ;
  assign y9819 = ~1'b0 ;
  assign y9820 = ~n21101 ;
  assign y9821 = n21103 ;
  assign y9822 = n21106 ;
  assign y9823 = ~n8002 ;
  assign y9824 = ~1'b0 ;
  assign y9825 = n21108 ;
  assign y9826 = ~n21111 ;
  assign y9827 = ~n21112 ;
  assign y9828 = ~n21113 ;
  assign y9829 = n21115 ;
  assign y9830 = n21117 ;
  assign y9831 = n21119 ;
  assign y9832 = ~1'b0 ;
  assign y9833 = ~1'b0 ;
  assign y9834 = ~1'b0 ;
  assign y9835 = ~n21125 ;
  assign y9836 = ~n21127 ;
  assign y9837 = n21130 ;
  assign y9838 = ~1'b0 ;
  assign y9839 = ~n8120 ;
  assign y9840 = n21132 ;
  assign y9841 = n21133 ;
  assign y9842 = n21134 ;
  assign y9843 = ~n21138 ;
  assign y9844 = ~n21140 ;
  assign y9845 = n10778 ;
  assign y9846 = ~1'b0 ;
  assign y9847 = ~1'b0 ;
  assign y9848 = ~1'b0 ;
  assign y9849 = n21143 ;
  assign y9850 = ~n21146 ;
  assign y9851 = ~1'b0 ;
  assign y9852 = n21148 ;
  assign y9853 = n21152 ;
  assign y9854 = ~n21156 ;
  assign y9855 = ~n21160 ;
  assign y9856 = ~1'b0 ;
  assign y9857 = ~1'b0 ;
  assign y9858 = ~1'b0 ;
  assign y9859 = ~1'b0 ;
  assign y9860 = ~n21161 ;
  assign y9861 = ~n21162 ;
  assign y9862 = ~n21164 ;
  assign y9863 = n21165 ;
  assign y9864 = n21167 ;
  assign y9865 = n21169 ;
  assign y9866 = n21172 ;
  assign y9867 = ~n21174 ;
  assign y9868 = ~n21175 ;
  assign y9869 = ~n21176 ;
  assign y9870 = n21182 ;
  assign y9871 = n21185 ;
  assign y9872 = ~n21186 ;
  assign y9873 = n21188 ;
  assign y9874 = n21192 ;
  assign y9875 = n21193 ;
  assign y9876 = n21195 ;
  assign y9877 = ~n21197 ;
  assign y9878 = n6668 ;
  assign y9879 = n21198 ;
  assign y9880 = n20972 ;
  assign y9881 = n21205 ;
  assign y9882 = ~n21206 ;
  assign y9883 = ~n21211 ;
  assign y9884 = n21215 ;
  assign y9885 = ~n21217 ;
  assign y9886 = n21221 ;
  assign y9887 = ~n21222 ;
  assign y9888 = n21223 ;
  assign y9889 = n21230 ;
  assign y9890 = ~n21235 ;
  assign y9891 = ~1'b0 ;
  assign y9892 = ~1'b0 ;
  assign y9893 = n21240 ;
  assign y9894 = ~1'b0 ;
  assign y9895 = n21245 ;
  assign y9896 = n21246 ;
  assign y9897 = ~n21252 ;
  assign y9898 = ~n21253 ;
  assign y9899 = ~1'b0 ;
  assign y9900 = ~n21255 ;
  assign y9901 = n21259 ;
  assign y9902 = ~n21265 ;
  assign y9903 = 1'b0 ;
  assign y9904 = ~1'b0 ;
  assign y9905 = ~n21270 ;
  assign y9906 = ~n21272 ;
  assign y9907 = ~n21273 ;
  assign y9908 = n21277 ;
  assign y9909 = ~n21279 ;
  assign y9910 = ~1'b0 ;
  assign y9911 = ~1'b0 ;
  assign y9912 = ~1'b0 ;
  assign y9913 = ~n21283 ;
  assign y9914 = n21285 ;
  assign y9915 = ~x45 ;
  assign y9916 = n21286 ;
  assign y9917 = ~n21287 ;
  assign y9918 = n21290 ;
  assign y9919 = n21304 ;
  assign y9920 = ~1'b0 ;
  assign y9921 = ~n21306 ;
  assign y9922 = n21307 ;
  assign y9923 = ~1'b0 ;
  assign y9924 = n11995 ;
  assign y9925 = n21308 ;
  assign y9926 = ~n21311 ;
  assign y9927 = n21320 ;
  assign y9928 = n21321 ;
  assign y9929 = ~1'b0 ;
  assign y9930 = ~n21323 ;
  assign y9931 = n21325 ;
  assign y9932 = n21326 ;
  assign y9933 = n21328 ;
  assign y9934 = n21330 ;
  assign y9935 = n21336 ;
  assign y9936 = n21337 ;
  assign y9937 = ~1'b0 ;
  assign y9938 = ~n21338 ;
  assign y9939 = n9437 ;
  assign y9940 = ~n21339 ;
  assign y9941 = n21351 ;
  assign y9942 = ~n21353 ;
  assign y9943 = n14185 ;
  assign y9944 = ~n21355 ;
  assign y9945 = ~n21357 ;
  assign y9946 = n21362 ;
  assign y9947 = n20442 ;
  assign y9948 = ~n21363 ;
  assign y9949 = ~1'b0 ;
  assign y9950 = ~1'b0 ;
  assign y9951 = ~n21366 ;
  assign y9952 = n21367 ;
  assign y9953 = ~n21368 ;
  assign y9954 = ~1'b0 ;
  assign y9955 = ~n21370 ;
  assign y9956 = ~n21371 ;
  assign y9957 = n21375 ;
  assign y9958 = n21378 ;
  assign y9959 = ~1'b0 ;
  assign y9960 = ~n21382 ;
  assign y9961 = n21383 ;
  assign y9962 = n21384 ;
  assign y9963 = n21386 ;
  assign y9964 = n21388 ;
  assign y9965 = ~1'b0 ;
  assign y9966 = ~n21389 ;
  assign y9967 = n21391 ;
  assign y9968 = ~1'b0 ;
  assign y9969 = n21393 ;
  assign y9970 = ~n21404 ;
  assign y9971 = n21405 ;
  assign y9972 = n21410 ;
  assign y9973 = ~n21411 ;
  assign y9974 = ~n21412 ;
  assign y9975 = ~n21414 ;
  assign y9976 = ~n21416 ;
  assign y9977 = n21417 ;
  assign y9978 = ~n21420 ;
  assign y9979 = n21421 ;
  assign y9980 = ~n21427 ;
  assign y9981 = ~1'b0 ;
  assign y9982 = n21430 ;
  assign y9983 = ~1'b0 ;
  assign y9984 = n21432 ;
  assign y9985 = ~1'b0 ;
  assign y9986 = n21433 ;
  assign y9987 = n21434 ;
  assign y9988 = ~n21435 ;
  assign y9989 = ~n21439 ;
  assign y9990 = ~n21445 ;
  assign y9991 = ~1'b0 ;
  assign y9992 = ~n21446 ;
  assign y9993 = n21451 ;
  assign y9994 = ~n21453 ;
  assign y9995 = ~1'b0 ;
  assign y9996 = n8563 ;
  assign y9997 = 1'b0 ;
  assign y9998 = ~n21454 ;
  assign y9999 = ~n21457 ;
  assign y10000 = ~n13940 ;
  assign y10001 = n21458 ;
  assign y10002 = n21459 ;
  assign y10003 = ~1'b0 ;
  assign y10004 = ~n21461 ;
  assign y10005 = ~n12495 ;
  assign y10006 = n21463 ;
  assign y10007 = n21467 ;
  assign y10008 = n21468 ;
  assign y10009 = ~n21471 ;
  assign y10010 = ~n21472 ;
  assign y10011 = ~n21476 ;
  assign y10012 = ~n21478 ;
  assign y10013 = ~n21480 ;
  assign y10014 = n21482 ;
  assign y10015 = n21484 ;
  assign y10016 = ~1'b0 ;
  assign y10017 = ~1'b0 ;
  assign y10018 = ~n21487 ;
  assign y10019 = ~n21489 ;
  assign y10020 = ~n21492 ;
  assign y10021 = ~1'b0 ;
  assign y10022 = ~1'b0 ;
  assign y10023 = n21494 ;
  assign y10024 = n21497 ;
  assign y10025 = ~n21501 ;
  assign y10026 = ~1'b0 ;
  assign y10027 = n21503 ;
  assign y10028 = n21504 ;
  assign y10029 = ~n21507 ;
  assign y10030 = ~1'b0 ;
  assign y10031 = ~1'b0 ;
  assign y10032 = ~n1281 ;
  assign y10033 = ~n21510 ;
  assign y10034 = n21511 ;
  assign y10035 = n21513 ;
  assign y10036 = ~n21517 ;
  assign y10037 = ~n21518 ;
  assign y10038 = ~n21520 ;
  assign y10039 = ~n21521 ;
  assign y10040 = ~n21525 ;
  assign y10041 = n21526 ;
  assign y10042 = n21527 ;
  assign y10043 = ~1'b0 ;
  assign y10044 = n21532 ;
  assign y10045 = ~1'b0 ;
  assign y10046 = n21534 ;
  assign y10047 = ~n21535 ;
  assign y10048 = n21537 ;
  assign y10049 = ~1'b0 ;
  assign y10050 = ~n21539 ;
  assign y10051 = n21540 ;
  assign y10052 = n21542 ;
  assign y10053 = ~n21543 ;
  assign y10054 = n21544 ;
  assign y10055 = ~n21546 ;
  assign y10056 = ~1'b0 ;
  assign y10057 = ~n21548 ;
  assign y10058 = n21551 ;
  assign y10059 = ~n21553 ;
  assign y10060 = ~n21555 ;
  assign y10061 = ~n21556 ;
  assign y10062 = ~n21561 ;
  assign y10063 = ~1'b0 ;
  assign y10064 = n21562 ;
  assign y10065 = n21563 ;
  assign y10066 = ~1'b0 ;
  assign y10067 = ~n21564 ;
  assign y10068 = ~1'b0 ;
  assign y10069 = ~n21565 ;
  assign y10070 = n21566 ;
  assign y10071 = ~n21567 ;
  assign y10072 = ~1'b0 ;
  assign y10073 = n21569 ;
  assign y10074 = ~1'b0 ;
  assign y10075 = n21573 ;
  assign y10076 = ~n21575 ;
  assign y10077 = ~n21581 ;
  assign y10078 = ~n21583 ;
  assign y10079 = n21584 ;
  assign y10080 = ~n21586 ;
  assign y10081 = ~1'b0 ;
  assign y10082 = ~n21588 ;
  assign y10083 = n21589 ;
  assign y10084 = ~1'b0 ;
  assign y10085 = ~1'b0 ;
  assign y10086 = n8546 ;
  assign y10087 = n21592 ;
  assign y10088 = n21603 ;
  assign y10089 = ~n21605 ;
  assign y10090 = ~1'b0 ;
  assign y10091 = ~1'b0 ;
  assign y10092 = ~1'b0 ;
  assign y10093 = n3496 ;
  assign y10094 = 1'b0 ;
  assign y10095 = n21607 ;
  assign y10096 = ~n21610 ;
  assign y10097 = ~1'b0 ;
  assign y10098 = ~1'b0 ;
  assign y10099 = n21611 ;
  assign y10100 = ~n21612 ;
  assign y10101 = ~n21616 ;
  assign y10102 = 1'b0 ;
  assign y10103 = ~1'b0 ;
  assign y10104 = ~n21617 ;
  assign y10105 = n21618 ;
  assign y10106 = ~n21621 ;
  assign y10107 = n21622 ;
  assign y10108 = ~n21623 ;
  assign y10109 = n21625 ;
  assign y10110 = n21626 ;
  assign y10111 = ~n21627 ;
  assign y10112 = n21630 ;
  assign y10113 = n21632 ;
  assign y10114 = n21635 ;
  assign y10115 = ~1'b0 ;
  assign y10116 = ~1'b0 ;
  assign y10117 = ~n21637 ;
  assign y10118 = n21644 ;
  assign y10119 = ~1'b0 ;
  assign y10120 = ~n21646 ;
  assign y10121 = n21647 ;
  assign y10122 = ~1'b0 ;
  assign y10123 = ~n21648 ;
  assign y10124 = ~n21649 ;
  assign y10125 = n21652 ;
  assign y10126 = ~1'b0 ;
  assign y10127 = n21654 ;
  assign y10128 = ~1'b0 ;
  assign y10129 = n21658 ;
  assign y10130 = ~1'b0 ;
  assign y10131 = ~n21660 ;
  assign y10132 = n21663 ;
  assign y10133 = n21671 ;
  assign y10134 = n21672 ;
  assign y10135 = ~n21676 ;
  assign y10136 = n21678 ;
  assign y10137 = ~n21682 ;
  assign y10138 = ~1'b0 ;
  assign y10139 = n21684 ;
  assign y10140 = n19045 ;
  assign y10141 = n21685 ;
  assign y10142 = ~n21686 ;
  assign y10143 = ~n21687 ;
  assign y10144 = n21690 ;
  assign y10145 = ~1'b0 ;
  assign y10146 = n21695 ;
  assign y10147 = ~n21699 ;
  assign y10148 = ~1'b0 ;
  assign y10149 = 1'b0 ;
  assign y10150 = ~n21700 ;
  assign y10151 = ~1'b0 ;
  assign y10152 = ~n21708 ;
  assign y10153 = ~n21710 ;
  assign y10154 = ~n21712 ;
  assign y10155 = ~n21713 ;
  assign y10156 = ~n21715 ;
  assign y10157 = ~n21716 ;
  assign y10158 = ~1'b0 ;
  assign y10159 = n21718 ;
  assign y10160 = n21719 ;
  assign y10161 = ~n21720 ;
  assign y10162 = ~n21723 ;
  assign y10163 = n21724 ;
  assign y10164 = ~1'b0 ;
  assign y10165 = ~1'b0 ;
  assign y10166 = n21726 ;
  assign y10167 = n21728 ;
  assign y10168 = ~n21731 ;
  assign y10169 = n21732 ;
  assign y10170 = ~n21737 ;
  assign y10171 = n21744 ;
  assign y10172 = ~1'b0 ;
  assign y10173 = ~n21751 ;
  assign y10174 = ~1'b0 ;
  assign y10175 = ~n21753 ;
  assign y10176 = ~1'b0 ;
  assign y10177 = ~n21758 ;
  assign y10178 = n21760 ;
  assign y10179 = ~1'b0 ;
  assign y10180 = n21763 ;
  assign y10181 = n21766 ;
  assign y10182 = n21768 ;
  assign y10183 = ~n21770 ;
  assign y10184 = ~n21771 ;
  assign y10185 = n21772 ;
  assign y10186 = n21774 ;
  assign y10187 = 1'b0 ;
  assign y10188 = ~n21781 ;
  assign y10189 = ~n21782 ;
  assign y10190 = ~1'b0 ;
  assign y10191 = ~n21785 ;
  assign y10192 = n21786 ;
  assign y10193 = ~1'b0 ;
  assign y10194 = ~1'b0 ;
  assign y10195 = ~n21789 ;
  assign y10196 = ~n14171 ;
  assign y10197 = ~n21791 ;
  assign y10198 = n21792 ;
  assign y10199 = n21793 ;
  assign y10200 = ~n21796 ;
  assign y10201 = ~1'b0 ;
  assign y10202 = n21801 ;
  assign y10203 = ~1'b0 ;
  assign y10204 = n21802 ;
  assign y10205 = n21804 ;
  assign y10206 = ~n21805 ;
  assign y10207 = n19325 ;
  assign y10208 = n21809 ;
  assign y10209 = n21811 ;
  assign y10210 = ~1'b0 ;
  assign y10211 = ~1'b0 ;
  assign y10212 = n21814 ;
  assign y10213 = ~1'b0 ;
  assign y10214 = n21829 ;
  assign y10215 = ~n21833 ;
  assign y10216 = n21834 ;
  assign y10217 = ~1'b0 ;
  assign y10218 = ~1'b0 ;
  assign y10219 = n21836 ;
  assign y10220 = n21840 ;
  assign y10221 = ~n21845 ;
  assign y10222 = n21846 ;
  assign y10223 = n21847 ;
  assign y10224 = ~1'b0 ;
  assign y10225 = ~1'b0 ;
  assign y10226 = ~1'b0 ;
  assign y10227 = ~1'b0 ;
  assign y10228 = n21854 ;
  assign y10229 = ~n21855 ;
  assign y10230 = n21858 ;
  assign y10231 = ~n21860 ;
  assign y10232 = n12331 ;
  assign y10233 = n21861 ;
  assign y10234 = ~1'b0 ;
  assign y10235 = ~n21865 ;
  assign y10236 = ~1'b0 ;
  assign y10237 = ~1'b0 ;
  assign y10238 = n21868 ;
  assign y10239 = n21874 ;
  assign y10240 = ~n21877 ;
  assign y10241 = ~n21880 ;
  assign y10242 = ~n21881 ;
  assign y10243 = n21883 ;
  assign y10244 = ~n21888 ;
  assign y10245 = ~1'b0 ;
  assign y10246 = ~n21889 ;
  assign y10247 = n12482 ;
  assign y10248 = n21893 ;
  assign y10249 = ~1'b0 ;
  assign y10250 = ~n21894 ;
  assign y10251 = ~1'b0 ;
  assign y10252 = n17137 ;
  assign y10253 = ~n21897 ;
  assign y10254 = ~1'b0 ;
  assign y10255 = ~1'b0 ;
  assign y10256 = ~1'b0 ;
  assign y10257 = n21902 ;
  assign y10258 = ~n20795 ;
  assign y10259 = ~n21906 ;
  assign y10260 = n21913 ;
  assign y10261 = ~1'b0 ;
  assign y10262 = n21915 ;
  assign y10263 = n21918 ;
  assign y10264 = n21922 ;
  assign y10265 = n12419 ;
  assign y10266 = ~n21923 ;
  assign y10267 = n21929 ;
  assign y10268 = ~n21931 ;
  assign y10269 = ~n21936 ;
  assign y10270 = ~1'b0 ;
  assign y10271 = ~n21937 ;
  assign y10272 = ~n21940 ;
  assign y10273 = ~1'b0 ;
  assign y10274 = n21945 ;
  assign y10275 = ~n21949 ;
  assign y10276 = n21952 ;
  assign y10277 = n21953 ;
  assign y10278 = ~n21957 ;
  assign y10279 = n21961 ;
  assign y10280 = n21965 ;
  assign y10281 = ~1'b0 ;
  assign y10282 = ~n21966 ;
  assign y10283 = n21971 ;
  assign y10284 = ~n21972 ;
  assign y10285 = ~n21974 ;
  assign y10286 = n21980 ;
  assign y10287 = n21981 ;
  assign y10288 = ~1'b0 ;
  assign y10289 = n21986 ;
  assign y10290 = ~n4769 ;
  assign y10291 = ~n21988 ;
  assign y10292 = n21989 ;
  assign y10293 = n21995 ;
  assign y10294 = n21996 ;
  assign y10295 = 1'b0 ;
  assign y10296 = ~1'b0 ;
  assign y10297 = 1'b0 ;
  assign y10298 = n21997 ;
  assign y10299 = ~n21998 ;
  assign y10300 = ~n19836 ;
  assign y10301 = ~n22000 ;
  assign y10302 = n22001 ;
  assign y10303 = ~1'b0 ;
  assign y10304 = ~1'b0 ;
  assign y10305 = ~n22008 ;
  assign y10306 = n22009 ;
  assign y10307 = ~1'b0 ;
  assign y10308 = ~n22010 ;
  assign y10309 = ~n22013 ;
  assign y10310 = ~1'b0 ;
  assign y10311 = ~n22015 ;
  assign y10312 = ~1'b0 ;
  assign y10313 = ~1'b0 ;
  assign y10314 = n22017 ;
  assign y10315 = n22023 ;
  assign y10316 = ~n6257 ;
  assign y10317 = ~n22024 ;
  assign y10318 = ~1'b0 ;
  assign y10319 = ~n22026 ;
  assign y10320 = n22030 ;
  assign y10321 = ~n22031 ;
  assign y10322 = ~1'b0 ;
  assign y10323 = ~1'b0 ;
  assign y10324 = ~n22033 ;
  assign y10325 = 1'b0 ;
  assign y10326 = n1955 ;
  assign y10327 = ~n22034 ;
  assign y10328 = ~1'b0 ;
  assign y10329 = n22039 ;
  assign y10330 = 1'b0 ;
  assign y10331 = ~n22041 ;
  assign y10332 = ~1'b0 ;
  assign y10333 = ~n22046 ;
  assign y10334 = n22048 ;
  assign y10335 = n2901 ;
  assign y10336 = ~n22050 ;
  assign y10337 = ~n2603 ;
  assign y10338 = n22053 ;
  assign y10339 = n22056 ;
  assign y10340 = ~1'b0 ;
  assign y10341 = ~n22058 ;
  assign y10342 = ~1'b0 ;
  assign y10343 = ~n22060 ;
  assign y10344 = ~n22062 ;
  assign y10345 = n22064 ;
  assign y10346 = ~n22065 ;
  assign y10347 = ~n22069 ;
  assign y10348 = n22073 ;
  assign y10349 = ~n22075 ;
  assign y10350 = n22076 ;
  assign y10351 = n22077 ;
  assign y10352 = ~n22078 ;
  assign y10353 = ~1'b0 ;
  assign y10354 = ~n13912 ;
  assign y10355 = n22082 ;
  assign y10356 = n22085 ;
  assign y10357 = ~1'b0 ;
  assign y10358 = ~n22089 ;
  assign y10359 = ~1'b0 ;
  assign y10360 = n22090 ;
  assign y10361 = ~n22093 ;
  assign y10362 = n22094 ;
  assign y10363 = ~1'b0 ;
  assign y10364 = ~1'b0 ;
  assign y10365 = ~n22098 ;
  assign y10366 = ~n22102 ;
  assign y10367 = n22104 ;
  assign y10368 = ~1'b0 ;
  assign y10369 = n22105 ;
  assign y10370 = ~n22106 ;
  assign y10371 = ~1'b0 ;
  assign y10372 = n22107 ;
  assign y10373 = ~1'b0 ;
  assign y10374 = ~n22109 ;
  assign y10375 = ~n22110 ;
  assign y10376 = ~n22115 ;
  assign y10377 = n22118 ;
  assign y10378 = n22119 ;
  assign y10379 = ~n22120 ;
  assign y10380 = ~n22122 ;
  assign y10381 = n22123 ;
  assign y10382 = n22124 ;
  assign y10383 = ~1'b0 ;
  assign y10384 = ~n22126 ;
  assign y10385 = ~n22128 ;
  assign y10386 = 1'b0 ;
  assign y10387 = n22130 ;
  assign y10388 = ~1'b0 ;
  assign y10389 = n22136 ;
  assign y10390 = n22138 ;
  assign y10391 = ~n22141 ;
  assign y10392 = ~1'b0 ;
  assign y10393 = ~n22144 ;
  assign y10394 = ~n22145 ;
  assign y10395 = ~1'b0 ;
  assign y10396 = ~n22148 ;
  assign y10397 = ~n22150 ;
  assign y10398 = ~n22152 ;
  assign y10399 = ~1'b0 ;
  assign y10400 = ~n22153 ;
  assign y10401 = n22157 ;
  assign y10402 = n22158 ;
  assign y10403 = n22160 ;
  assign y10404 = n22163 ;
  assign y10405 = ~n22166 ;
  assign y10406 = ~1'b0 ;
  assign y10407 = n22169 ;
  assign y10408 = ~n22172 ;
  assign y10409 = n22173 ;
  assign y10410 = ~n22174 ;
  assign y10411 = ~n22176 ;
  assign y10412 = 1'b0 ;
  assign y10413 = n22177 ;
  assign y10414 = ~n22181 ;
  assign y10415 = n22184 ;
  assign y10416 = ~n22185 ;
  assign y10417 = ~n22188 ;
  assign y10418 = ~n22191 ;
  assign y10419 = n22193 ;
  assign y10420 = ~1'b0 ;
  assign y10421 = n22198 ;
  assign y10422 = ~n22202 ;
  assign y10423 = ~n22203 ;
  assign y10424 = ~1'b0 ;
  assign y10425 = n7588 ;
  assign y10426 = ~1'b0 ;
  assign y10427 = n22206 ;
  assign y10428 = ~1'b0 ;
  assign y10429 = n22207 ;
  assign y10430 = ~n22209 ;
  assign y10431 = ~n22212 ;
  assign y10432 = ~n14545 ;
  assign y10433 = n22213 ;
  assign y10434 = ~1'b0 ;
  assign y10435 = ~1'b0 ;
  assign y10436 = ~n22214 ;
  assign y10437 = ~1'b0 ;
  assign y10438 = n22222 ;
  assign y10439 = n22224 ;
  assign y10440 = n22229 ;
  assign y10441 = n22230 ;
  assign y10442 = ~n22235 ;
  assign y10443 = n22236 ;
  assign y10444 = n22238 ;
  assign y10445 = n22240 ;
  assign y10446 = ~1'b0 ;
  assign y10447 = n22243 ;
  assign y10448 = ~n22244 ;
  assign y10449 = ~n22246 ;
  assign y10450 = ~n22247 ;
  assign y10451 = ~n22249 ;
  assign y10452 = ~n12015 ;
  assign y10453 = ~1'b0 ;
  assign y10454 = n22250 ;
  assign y10455 = ~1'b0 ;
  assign y10456 = ~n22253 ;
  assign y10457 = ~n22254 ;
  assign y10458 = ~1'b0 ;
  assign y10459 = n22255 ;
  assign y10460 = n22256 ;
  assign y10461 = ~n22257 ;
  assign y10462 = ~1'b0 ;
  assign y10463 = ~n22265 ;
  assign y10464 = ~1'b0 ;
  assign y10465 = ~1'b0 ;
  assign y10466 = ~n22267 ;
  assign y10467 = ~1'b0 ;
  assign y10468 = n22269 ;
  assign y10469 = n10729 ;
  assign y10470 = n22275 ;
  assign y10471 = n22276 ;
  assign y10472 = ~n22278 ;
  assign y10473 = ~n22280 ;
  assign y10474 = ~1'b0 ;
  assign y10475 = ~1'b0 ;
  assign y10476 = ~n22281 ;
  assign y10477 = ~n22286 ;
  assign y10478 = n22290 ;
  assign y10479 = ~n22292 ;
  assign y10480 = ~n22296 ;
  assign y10481 = ~n22297 ;
  assign y10482 = n22298 ;
  assign y10483 = n22303 ;
  assign y10484 = n22306 ;
  assign y10485 = n22308 ;
  assign y10486 = ~1'b0 ;
  assign y10487 = n22309 ;
  assign y10488 = n22311 ;
  assign y10489 = n22313 ;
  assign y10490 = ~n22317 ;
  assign y10491 = ~1'b0 ;
  assign y10492 = ~n22320 ;
  assign y10493 = ~n22321 ;
  assign y10494 = ~n22323 ;
  assign y10495 = ~n22327 ;
  assign y10496 = ~1'b0 ;
  assign y10497 = ~1'b0 ;
  assign y10498 = n22328 ;
  assign y10499 = n22331 ;
  assign y10500 = n22332 ;
  assign y10501 = n22337 ;
  assign y10502 = ~n22339 ;
  assign y10503 = n22340 ;
  assign y10504 = ~1'b0 ;
  assign y10505 = ~n22343 ;
  assign y10506 = 1'b0 ;
  assign y10507 = ~1'b0 ;
  assign y10508 = ~n22345 ;
  assign y10509 = 1'b0 ;
  assign y10510 = ~n22349 ;
  assign y10511 = ~1'b0 ;
  assign y10512 = ~1'b0 ;
  assign y10513 = n22356 ;
  assign y10514 = ~1'b0 ;
  assign y10515 = n22357 ;
  assign y10516 = n22361 ;
  assign y10517 = n22366 ;
  assign y10518 = n22369 ;
  assign y10519 = ~1'b0 ;
  assign y10520 = ~1'b0 ;
  assign y10521 = ~n22371 ;
  assign y10522 = n22373 ;
  assign y10523 = ~n22377 ;
  assign y10524 = ~n22379 ;
  assign y10525 = ~n22381 ;
  assign y10526 = n22383 ;
  assign y10527 = ~n22384 ;
  assign y10528 = ~n22385 ;
  assign y10529 = ~n22387 ;
  assign y10530 = n1594 ;
  assign y10531 = ~1'b0 ;
  assign y10532 = 1'b0 ;
  assign y10533 = ~n22390 ;
  assign y10534 = ~n22391 ;
  assign y10535 = n22392 ;
  assign y10536 = n22395 ;
  assign y10537 = ~n22396 ;
  assign y10538 = ~n22397 ;
  assign y10539 = ~n22399 ;
  assign y10540 = n22402 ;
  assign y10541 = ~n22405 ;
  assign y10542 = ~1'b0 ;
  assign y10543 = n22407 ;
  assign y10544 = n22414 ;
  assign y10545 = ~n22417 ;
  assign y10546 = n22421 ;
  assign y10547 = ~1'b0 ;
  assign y10548 = ~1'b0 ;
  assign y10549 = ~1'b0 ;
  assign y10550 = ~1'b0 ;
  assign y10551 = ~1'b0 ;
  assign y10552 = n22424 ;
  assign y10553 = ~n22426 ;
  assign y10554 = ~n22427 ;
  assign y10555 = n2798 ;
  assign y10556 = n22428 ;
  assign y10557 = ~n22434 ;
  assign y10558 = ~1'b0 ;
  assign y10559 = n22436 ;
  assign y10560 = ~1'b0 ;
  assign y10561 = ~1'b0 ;
  assign y10562 = n22438 ;
  assign y10563 = ~n22442 ;
  assign y10564 = n22443 ;
  assign y10565 = ~n22447 ;
  assign y10566 = n8965 ;
  assign y10567 = 1'b0 ;
  assign y10568 = ~n22450 ;
  assign y10569 = ~n22451 ;
  assign y10570 = ~1'b0 ;
  assign y10571 = ~n22454 ;
  assign y10572 = ~1'b0 ;
  assign y10573 = n22455 ;
  assign y10574 = ~n22456 ;
  assign y10575 = ~n14354 ;
  assign y10576 = n22457 ;
  assign y10577 = ~n22460 ;
  assign y10578 = n22462 ;
  assign y10579 = ~n10268 ;
  assign y10580 = ~n22467 ;
  assign y10581 = ~n9466 ;
  assign y10582 = ~n22468 ;
  assign y10583 = n22469 ;
  assign y10584 = ~n22470 ;
  assign y10585 = n22471 ;
  assign y10586 = ~1'b0 ;
  assign y10587 = ~1'b0 ;
  assign y10588 = n22472 ;
  assign y10589 = ~n22477 ;
  assign y10590 = ~n22481 ;
  assign y10591 = ~n22485 ;
  assign y10592 = ~n22490 ;
  assign y10593 = ~n22492 ;
  assign y10594 = n22497 ;
  assign y10595 = ~n22499 ;
  assign y10596 = ~1'b0 ;
  assign y10597 = ~1'b0 ;
  assign y10598 = ~1'b0 ;
  assign y10599 = n22501 ;
  assign y10600 = ~n22503 ;
  assign y10601 = n22505 ;
  assign y10602 = ~n22506 ;
  assign y10603 = n22512 ;
  assign y10604 = ~n22514 ;
  assign y10605 = ~1'b0 ;
  assign y10606 = n22518 ;
  assign y10607 = ~1'b0 ;
  assign y10608 = n22522 ;
  assign y10609 = ~n22532 ;
  assign y10610 = ~1'b0 ;
  assign y10611 = ~n22535 ;
  assign y10612 = n22537 ;
  assign y10613 = n22544 ;
  assign y10614 = ~n22546 ;
  assign y10615 = ~n22548 ;
  assign y10616 = ~n22549 ;
  assign y10617 = ~n22553 ;
  assign y10618 = n22555 ;
  assign y10619 = n22556 ;
  assign y10620 = ~n22559 ;
  assign y10621 = ~n22560 ;
  assign y10622 = n22562 ;
  assign y10623 = ~n22565 ;
  assign y10624 = ~n22569 ;
  assign y10625 = ~1'b0 ;
  assign y10626 = ~n22571 ;
  assign y10627 = ~n22573 ;
  assign y10628 = ~1'b0 ;
  assign y10629 = n22586 ;
  assign y10630 = ~n22588 ;
  assign y10631 = ~n22590 ;
  assign y10632 = 1'b0 ;
  assign y10633 = n22593 ;
  assign y10634 = n22598 ;
  assign y10635 = n22600 ;
  assign y10636 = ~n22601 ;
  assign y10637 = ~n22605 ;
  assign y10638 = ~n22607 ;
  assign y10639 = ~n22608 ;
  assign y10640 = ~n22610 ;
  assign y10641 = ~1'b0 ;
  assign y10642 = ~1'b0 ;
  assign y10643 = ~1'b0 ;
  assign y10644 = n22614 ;
  assign y10645 = n22620 ;
  assign y10646 = ~1'b0 ;
  assign y10647 = ~1'b0 ;
  assign y10648 = ~n22621 ;
  assign y10649 = n22625 ;
  assign y10650 = ~n22631 ;
  assign y10651 = ~1'b0 ;
  assign y10652 = n22632 ;
  assign y10653 = n22634 ;
  assign y10654 = n22636 ;
  assign y10655 = n22638 ;
  assign y10656 = n22643 ;
  assign y10657 = n22645 ;
  assign y10658 = n22646 ;
  assign y10659 = ~1'b0 ;
  assign y10660 = ~n22648 ;
  assign y10661 = ~n22652 ;
  assign y10662 = ~1'b0 ;
  assign y10663 = ~n22654 ;
  assign y10664 = ~1'b0 ;
  assign y10665 = n22658 ;
  assign y10666 = n22663 ;
  assign y10667 = n22664 ;
  assign y10668 = n22666 ;
  assign y10669 = ~1'b0 ;
  assign y10670 = ~1'b0 ;
  assign y10671 = ~n22667 ;
  assign y10672 = ~n22673 ;
  assign y10673 = ~1'b0 ;
  assign y10674 = ~n22674 ;
  assign y10675 = ~n22675 ;
  assign y10676 = 1'b0 ;
  assign y10677 = n22677 ;
  assign y10678 = n22679 ;
  assign y10679 = ~1'b0 ;
  assign y10680 = ~n22683 ;
  assign y10681 = ~n22685 ;
  assign y10682 = ~1'b0 ;
  assign y10683 = n22689 ;
  assign y10684 = ~n22690 ;
  assign y10685 = n22691 ;
  assign y10686 = ~1'b0 ;
  assign y10687 = ~1'b0 ;
  assign y10688 = n22694 ;
  assign y10689 = ~n22696 ;
  assign y10690 = ~n22703 ;
  assign y10691 = ~n22706 ;
  assign y10692 = ~1'b0 ;
  assign y10693 = ~n22707 ;
  assign y10694 = ~n22708 ;
  assign y10695 = n22709 ;
  assign y10696 = n22713 ;
  assign y10697 = ~1'b0 ;
  assign y10698 = ~n5765 ;
  assign y10699 = ~n13912 ;
  assign y10700 = ~1'b0 ;
  assign y10701 = ~1'b0 ;
  assign y10702 = ~n3628 ;
  assign y10703 = ~1'b0 ;
  assign y10704 = ~n22718 ;
  assign y10705 = ~1'b0 ;
  assign y10706 = ~1'b0 ;
  assign y10707 = ~n22720 ;
  assign y10708 = n22725 ;
  assign y10709 = ~n22728 ;
  assign y10710 = ~1'b0 ;
  assign y10711 = ~n22731 ;
  assign y10712 = ~n22733 ;
  assign y10713 = n22734 ;
  assign y10714 = ~1'b0 ;
  assign y10715 = 1'b0 ;
  assign y10716 = ~1'b0 ;
  assign y10717 = ~1'b0 ;
  assign y10718 = ~n22736 ;
  assign y10719 = ~n22739 ;
  assign y10720 = n22740 ;
  assign y10721 = ~n22741 ;
  assign y10722 = ~n22747 ;
  assign y10723 = n22748 ;
  assign y10724 = ~1'b0 ;
  assign y10725 = n22751 ;
  assign y10726 = n22756 ;
  assign y10727 = ~n22759 ;
  assign y10728 = ~n22761 ;
  assign y10729 = ~n22762 ;
  assign y10730 = n22763 ;
  assign y10731 = ~1'b0 ;
  assign y10732 = n22769 ;
  assign y10733 = ~1'b0 ;
  assign y10734 = n22771 ;
  assign y10735 = ~1'b0 ;
  assign y10736 = n22774 ;
  assign y10737 = ~n22779 ;
  assign y10738 = ~n22780 ;
  assign y10739 = ~n22783 ;
  assign y10740 = n22785 ;
  assign y10741 = ~n22789 ;
  assign y10742 = n22790 ;
  assign y10743 = ~1'b0 ;
  assign y10744 = ~n22795 ;
  assign y10745 = n22797 ;
  assign y10746 = ~1'b0 ;
  assign y10747 = n22802 ;
  assign y10748 = n22803 ;
  assign y10749 = ~1'b0 ;
  assign y10750 = n22804 ;
  assign y10751 = ~n22808 ;
  assign y10752 = n22809 ;
  assign y10753 = n22811 ;
  assign y10754 = ~1'b0 ;
  assign y10755 = n22813 ;
  assign y10756 = ~n11813 ;
  assign y10757 = n22815 ;
  assign y10758 = ~1'b0 ;
  assign y10759 = ~n3802 ;
  assign y10760 = ~1'b0 ;
  assign y10761 = ~1'b0 ;
  assign y10762 = ~1'b0 ;
  assign y10763 = n16699 ;
  assign y10764 = ~1'b0 ;
  assign y10765 = ~n22818 ;
  assign y10766 = ~n22820 ;
  assign y10767 = n22821 ;
  assign y10768 = n22822 ;
  assign y10769 = ~n22826 ;
  assign y10770 = n22828 ;
  assign y10771 = n22831 ;
  assign y10772 = ~n22835 ;
  assign y10773 = n22841 ;
  assign y10774 = ~n22844 ;
  assign y10775 = ~n22846 ;
  assign y10776 = ~n22849 ;
  assign y10777 = n22851 ;
  assign y10778 = ~n22855 ;
  assign y10779 = ~n22856 ;
  assign y10780 = ~n22857 ;
  assign y10781 = ~n22860 ;
  assign y10782 = n22863 ;
  assign y10783 = ~n22866 ;
  assign y10784 = ~n22867 ;
  assign y10785 = ~1'b0 ;
  assign y10786 = ~n5046 ;
  assign y10787 = 1'b0 ;
  assign y10788 = n22873 ;
  assign y10789 = ~n22876 ;
  assign y10790 = ~n22878 ;
  assign y10791 = ~n9084 ;
  assign y10792 = n22881 ;
  assign y10793 = ~n22884 ;
  assign y10794 = ~n22889 ;
  assign y10795 = ~n22890 ;
  assign y10796 = ~n22892 ;
  assign y10797 = ~n22899 ;
  assign y10798 = ~1'b0 ;
  assign y10799 = n22905 ;
  assign y10800 = ~n22907 ;
  assign y10801 = ~1'b0 ;
  assign y10802 = ~1'b0 ;
  assign y10803 = ~n22913 ;
  assign y10804 = ~n22914 ;
  assign y10805 = ~1'b0 ;
  assign y10806 = ~1'b0 ;
  assign y10807 = ~n22916 ;
  assign y10808 = ~1'b0 ;
  assign y10809 = n22917 ;
  assign y10810 = ~n22826 ;
  assign y10811 = n22920 ;
  assign y10812 = n22922 ;
  assign y10813 = n22923 ;
  assign y10814 = ~n22925 ;
  assign y10815 = ~n22930 ;
  assign y10816 = n22934 ;
  assign y10817 = n22935 ;
  assign y10818 = ~n22937 ;
  assign y10819 = ~1'b0 ;
  assign y10820 = n22940 ;
  assign y10821 = ~n22941 ;
  assign y10822 = n22943 ;
  assign y10823 = ~n22944 ;
  assign y10824 = n22945 ;
  assign y10825 = ~1'b0 ;
  assign y10826 = n22949 ;
  assign y10827 = ~1'b0 ;
  assign y10828 = ~1'b0 ;
  assign y10829 = n22951 ;
  assign y10830 = ~1'b0 ;
  assign y10831 = n22953 ;
  assign y10832 = n22955 ;
  assign y10833 = n22958 ;
  assign y10834 = ~n22959 ;
  assign y10835 = n22960 ;
  assign y10836 = n22962 ;
  assign y10837 = ~n9717 ;
  assign y10838 = n22965 ;
  assign y10839 = ~1'b0 ;
  assign y10840 = ~n22967 ;
  assign y10841 = ~1'b0 ;
  assign y10842 = n22973 ;
  assign y10843 = ~1'b0 ;
  assign y10844 = ~n22974 ;
  assign y10845 = ~n22975 ;
  assign y10846 = ~1'b0 ;
  assign y10847 = ~1'b0 ;
  assign y10848 = ~1'b0 ;
  assign y10849 = ~n22980 ;
  assign y10850 = ~1'b0 ;
  assign y10851 = ~1'b0 ;
  assign y10852 = n22983 ;
  assign y10853 = ~n22984 ;
  assign y10854 = ~n22985 ;
  assign y10855 = ~1'b0 ;
  assign y10856 = ~1'b0 ;
  assign y10857 = ~1'b0 ;
  assign y10858 = ~n22987 ;
  assign y10859 = n2063 ;
  assign y10860 = ~1'b0 ;
  assign y10861 = n22990 ;
  assign y10862 = ~n22994 ;
  assign y10863 = ~n22997 ;
  assign y10864 = n22999 ;
  assign y10865 = ~n23001 ;
  assign y10866 = ~n23003 ;
  assign y10867 = ~1'b0 ;
  assign y10868 = ~n23007 ;
  assign y10869 = 1'b0 ;
  assign y10870 = n23011 ;
  assign y10871 = ~n23014 ;
  assign y10872 = ~n23015 ;
  assign y10873 = n23016 ;
  assign y10874 = ~n23020 ;
  assign y10875 = ~1'b0 ;
  assign y10876 = ~1'b0 ;
  assign y10877 = ~n23021 ;
  assign y10878 = n23025 ;
  assign y10879 = ~n23026 ;
  assign y10880 = ~n23027 ;
  assign y10881 = n23032 ;
  assign y10882 = ~n23033 ;
  assign y10883 = ~1'b0 ;
  assign y10884 = ~n23035 ;
  assign y10885 = ~1'b0 ;
  assign y10886 = ~1'b0 ;
  assign y10887 = n23036 ;
  assign y10888 = ~n23038 ;
  assign y10889 = ~1'b0 ;
  assign y10890 = n23041 ;
  assign y10891 = n23042 ;
  assign y10892 = n23043 ;
  assign y10893 = ~n23045 ;
  assign y10894 = n23047 ;
  assign y10895 = n23048 ;
  assign y10896 = n23053 ;
  assign y10897 = n23056 ;
  assign y10898 = ~n23058 ;
  assign y10899 = ~n23059 ;
  assign y10900 = ~n23061 ;
  assign y10901 = ~1'b0 ;
  assign y10902 = n23063 ;
  assign y10903 = ~n23067 ;
  assign y10904 = ~n23070 ;
  assign y10905 = ~n23071 ;
  assign y10906 = ~1'b0 ;
  assign y10907 = n14212 ;
  assign y10908 = ~n23072 ;
  assign y10909 = ~1'b0 ;
  assign y10910 = n23074 ;
  assign y10911 = ~n23076 ;
  assign y10912 = ~n23078 ;
  assign y10913 = n23079 ;
  assign y10914 = ~n23084 ;
  assign y10915 = n23086 ;
  assign y10916 = ~1'b0 ;
  assign y10917 = ~1'b0 ;
  assign y10918 = n23090 ;
  assign y10919 = ~n23091 ;
  assign y10920 = ~1'b0 ;
  assign y10921 = ~n23092 ;
  assign y10922 = n23097 ;
  assign y10923 = n23099 ;
  assign y10924 = ~n23100 ;
  assign y10925 = n23101 ;
  assign y10926 = ~n23102 ;
  assign y10927 = n23104 ;
  assign y10928 = n23105 ;
  assign y10929 = ~n23108 ;
  assign y10930 = ~1'b0 ;
  assign y10931 = ~n21538 ;
  assign y10932 = ~n23109 ;
  assign y10933 = ~n23112 ;
  assign y10934 = n23116 ;
  assign y10935 = n23118 ;
  assign y10936 = ~n23120 ;
  assign y10937 = n23122 ;
  assign y10938 = ~n23126 ;
  assign y10939 = ~1'b0 ;
  assign y10940 = ~n23129 ;
  assign y10941 = n18769 ;
  assign y10942 = ~n23130 ;
  assign y10943 = ~n23133 ;
  assign y10944 = n23134 ;
  assign y10945 = ~1'b0 ;
  assign y10946 = ~1'b0 ;
  assign y10947 = n23135 ;
  assign y10948 = n23137 ;
  assign y10949 = ~1'b0 ;
  assign y10950 = n23139 ;
  assign y10951 = n23142 ;
  assign y10952 = ~n23143 ;
  assign y10953 = ~n23146 ;
  assign y10954 = n23148 ;
  assign y10955 = n23152 ;
  assign y10956 = n23153 ;
  assign y10957 = ~n23157 ;
  assign y10958 = n23158 ;
  assign y10959 = n23160 ;
  assign y10960 = ~n23161 ;
  assign y10961 = n23163 ;
  assign y10962 = ~n23164 ;
  assign y10963 = n23165 ;
  assign y10964 = ~n23169 ;
  assign y10965 = ~n23171 ;
  assign y10966 = n23177 ;
  assign y10967 = ~1'b0 ;
  assign y10968 = ~n23179 ;
  assign y10969 = ~n23183 ;
  assign y10970 = ~n23187 ;
  assign y10971 = ~n23188 ;
  assign y10972 = n23190 ;
  assign y10973 = 1'b0 ;
  assign y10974 = ~1'b0 ;
  assign y10975 = ~1'b0 ;
  assign y10976 = ~1'b0 ;
  assign y10977 = ~n23193 ;
  assign y10978 = n23195 ;
  assign y10979 = ~n23196 ;
  assign y10980 = n23198 ;
  assign y10981 = ~n23204 ;
  assign y10982 = n23205 ;
  assign y10983 = n23206 ;
  assign y10984 = ~n23213 ;
  assign y10985 = ~1'b0 ;
  assign y10986 = n23215 ;
  assign y10987 = n10403 ;
  assign y10988 = ~n23217 ;
  assign y10989 = ~n23219 ;
  assign y10990 = ~n23220 ;
  assign y10991 = ~n23225 ;
  assign y10992 = ~n23226 ;
  assign y10993 = n23228 ;
  assign y10994 = n23229 ;
  assign y10995 = n23231 ;
  assign y10996 = ~n23232 ;
  assign y10997 = n23233 ;
  assign y10998 = n2362 ;
  assign y10999 = ~n23237 ;
  assign y11000 = n23238 ;
  assign y11001 = n23239 ;
  assign y11002 = ~1'b0 ;
  assign y11003 = ~n23242 ;
  assign y11004 = n23243 ;
  assign y11005 = n23244 ;
  assign y11006 = n23247 ;
  assign y11007 = ~1'b0 ;
  assign y11008 = n23251 ;
  assign y11009 = ~n23252 ;
  assign y11010 = ~1'b0 ;
  assign y11011 = ~n23253 ;
  assign y11012 = n23258 ;
  assign y11013 = ~n23260 ;
  assign y11014 = ~n23263 ;
  assign y11015 = ~1'b0 ;
  assign y11016 = ~1'b0 ;
  assign y11017 = ~n23266 ;
  assign y11018 = n23269 ;
  assign y11019 = n23272 ;
  assign y11020 = ~1'b0 ;
  assign y11021 = n175 ;
  assign y11022 = n23276 ;
  assign y11023 = ~n23277 ;
  assign y11024 = ~1'b0 ;
  assign y11025 = n23278 ;
  assign y11026 = ~n23279 ;
  assign y11027 = ~n23282 ;
  assign y11028 = n23286 ;
  assign y11029 = n23291 ;
  assign y11030 = ~1'b0 ;
  assign y11031 = ~n23294 ;
  assign y11032 = n23299 ;
  assign y11033 = n23301 ;
  assign y11034 = ~1'b0 ;
  assign y11035 = n10318 ;
  assign y11036 = ~n23307 ;
  assign y11037 = ~n23308 ;
  assign y11038 = ~n23309 ;
  assign y11039 = n23312 ;
  assign y11040 = ~1'b0 ;
  assign y11041 = ~n23315 ;
  assign y11042 = ~n23316 ;
  assign y11043 = ~n23318 ;
  assign y11044 = n23320 ;
  assign y11045 = n23321 ;
  assign y11046 = ~1'b0 ;
  assign y11047 = ~n23324 ;
  assign y11048 = ~n23332 ;
  assign y11049 = ~n23336 ;
  assign y11050 = ~n2404 ;
  assign y11051 = ~1'b0 ;
  assign y11052 = ~1'b0 ;
  assign y11053 = n23339 ;
  assign y11054 = ~1'b0 ;
  assign y11055 = n23341 ;
  assign y11056 = n10296 ;
  assign y11057 = n23354 ;
  assign y11058 = n23357 ;
  assign y11059 = ~n23359 ;
  assign y11060 = ~1'b0 ;
  assign y11061 = ~1'b0 ;
  assign y11062 = n6290 ;
  assign y11063 = ~n23360 ;
  assign y11064 = n23361 ;
  assign y11065 = ~n23363 ;
  assign y11066 = ~1'b0 ;
  assign y11067 = n23364 ;
  assign y11068 = n23365 ;
  assign y11069 = ~n23367 ;
  assign y11070 = ~1'b0 ;
  assign y11071 = ~n23368 ;
  assign y11072 = ~n23371 ;
  assign y11073 = ~n2194 ;
  assign y11074 = n23372 ;
  assign y11075 = n23373 ;
  assign y11076 = ~1'b0 ;
  assign y11077 = n1097 ;
  assign y11078 = n23375 ;
  assign y11079 = ~1'b0 ;
  assign y11080 = n23379 ;
  assign y11081 = ~1'b0 ;
  assign y11082 = ~n23381 ;
  assign y11083 = n23384 ;
  assign y11084 = ~n6068 ;
  assign y11085 = ~1'b0 ;
  assign y11086 = n23389 ;
  assign y11087 = ~1'b0 ;
  assign y11088 = n23390 ;
  assign y11089 = ~n23392 ;
  assign y11090 = ~n23394 ;
  assign y11091 = n21765 ;
  assign y11092 = ~n23397 ;
  assign y11093 = ~1'b0 ;
  assign y11094 = ~n13269 ;
  assign y11095 = ~n23398 ;
  assign y11096 = n23400 ;
  assign y11097 = ~n23403 ;
  assign y11098 = n23406 ;
  assign y11099 = n23411 ;
  assign y11100 = ~n23415 ;
  assign y11101 = ~n23416 ;
  assign y11102 = n23422 ;
  assign y11103 = ~1'b0 ;
  assign y11104 = ~1'b0 ;
  assign y11105 = n23423 ;
  assign y11106 = ~n23425 ;
  assign y11107 = ~1'b0 ;
  assign y11108 = ~n23426 ;
  assign y11109 = n23429 ;
  assign y11110 = n23435 ;
  assign y11111 = n23437 ;
  assign y11112 = ~1'b0 ;
  assign y11113 = n23438 ;
  assign y11114 = n23442 ;
  assign y11115 = ~1'b0 ;
  assign y11116 = ~1'b0 ;
  assign y11117 = ~1'b0 ;
  assign y11118 = ~n23444 ;
  assign y11119 = ~n23446 ;
  assign y11120 = ~n23451 ;
  assign y11121 = ~n23455 ;
  assign y11122 = n23458 ;
  assign y11123 = ~n23461 ;
  assign y11124 = n23462 ;
  assign y11125 = n23467 ;
  assign y11126 = ~1'b0 ;
  assign y11127 = ~n23473 ;
  assign y11128 = n23475 ;
  assign y11129 = ~n23476 ;
  assign y11130 = ~1'b0 ;
  assign y11131 = ~1'b0 ;
  assign y11132 = ~1'b0 ;
  assign y11133 = ~n23477 ;
  assign y11134 = ~n23480 ;
  assign y11135 = ~n23481 ;
  assign y11136 = ~n23482 ;
  assign y11137 = ~n23485 ;
  assign y11138 = n23486 ;
  assign y11139 = ~1'b0 ;
  assign y11140 = ~1'b0 ;
  assign y11141 = n23489 ;
  assign y11142 = ~1'b0 ;
  assign y11143 = ~n23492 ;
  assign y11144 = n23493 ;
  assign y11145 = ~n23495 ;
  assign y11146 = ~1'b0 ;
  assign y11147 = ~n23498 ;
  assign y11148 = ~n23500 ;
  assign y11149 = ~n23501 ;
  assign y11150 = n23506 ;
  assign y11151 = n12559 ;
  assign y11152 = n23507 ;
  assign y11153 = n23511 ;
  assign y11154 = ~n23514 ;
  assign y11155 = n23515 ;
  assign y11156 = ~n23521 ;
  assign y11157 = ~1'b0 ;
  assign y11158 = ~n23524 ;
  assign y11159 = ~n23525 ;
  assign y11160 = n23527 ;
  assign y11161 = ~n23529 ;
  assign y11162 = n23531 ;
  assign y11163 = ~n23537 ;
  assign y11164 = ~n23539 ;
  assign y11165 = n23541 ;
  assign y11166 = n23545 ;
  assign y11167 = n23547 ;
  assign y11168 = ~1'b0 ;
  assign y11169 = ~n23548 ;
  assign y11170 = ~1'b0 ;
  assign y11171 = n23549 ;
  assign y11172 = ~1'b0 ;
  assign y11173 = ~1'b0 ;
  assign y11174 = ~n23552 ;
  assign y11175 = ~n23555 ;
  assign y11176 = ~n23556 ;
  assign y11177 = ~n23561 ;
  assign y11178 = ~1'b0 ;
  assign y11179 = ~n23563 ;
  assign y11180 = ~1'b0 ;
  assign y11181 = ~1'b0 ;
  assign y11182 = ~1'b0 ;
  assign y11183 = ~n23564 ;
  assign y11184 = ~1'b0 ;
  assign y11185 = ~1'b0 ;
  assign y11186 = ~n23565 ;
  assign y11187 = ~1'b0 ;
  assign y11188 = ~1'b0 ;
  assign y11189 = ~n23568 ;
  assign y11190 = ~1'b0 ;
  assign y11191 = ~n23569 ;
  assign y11192 = ~1'b0 ;
  assign y11193 = n23571 ;
  assign y11194 = ~1'b0 ;
  assign y11195 = ~n23572 ;
  assign y11196 = ~n23575 ;
  assign y11197 = 1'b0 ;
  assign y11198 = ~1'b0 ;
  assign y11199 = n23579 ;
  assign y11200 = ~n23580 ;
  assign y11201 = ~1'b0 ;
  assign y11202 = ~n23581 ;
  assign y11203 = ~1'b0 ;
  assign y11204 = ~n23584 ;
  assign y11205 = ~n23585 ;
  assign y11206 = n23586 ;
  assign y11207 = ~n23588 ;
  assign y11208 = ~n23589 ;
  assign y11209 = n23591 ;
  assign y11210 = ~1'b0 ;
  assign y11211 = 1'b0 ;
  assign y11212 = ~1'b0 ;
  assign y11213 = ~n23592 ;
  assign y11214 = n23600 ;
  assign y11215 = ~1'b0 ;
  assign y11216 = 1'b0 ;
  assign y11217 = n23602 ;
  assign y11218 = n23605 ;
  assign y11219 = n23607 ;
  assign y11220 = ~n23608 ;
  assign y11221 = ~n23609 ;
  assign y11222 = n23614 ;
  assign y11223 = n23616 ;
  assign y11224 = ~n23618 ;
  assign y11225 = ~n23619 ;
  assign y11226 = ~n12338 ;
  assign y11227 = ~1'b0 ;
  assign y11228 = ~n23623 ;
  assign y11229 = ~n23624 ;
  assign y11230 = n23627 ;
  assign y11231 = ~n23628 ;
  assign y11232 = ~n23629 ;
  assign y11233 = n23631 ;
  assign y11234 = ~n16825 ;
  assign y11235 = n23633 ;
  assign y11236 = n23636 ;
  assign y11237 = n23641 ;
  assign y11238 = ~1'b0 ;
  assign y11239 = ~n23643 ;
  assign y11240 = n8721 ;
  assign y11241 = ~n23646 ;
  assign y11242 = ~n23648 ;
  assign y11243 = ~n23651 ;
  assign y11244 = ~1'b0 ;
  assign y11245 = ~n23652 ;
  assign y11246 = ~n23653 ;
  assign y11247 = ~1'b0 ;
  assign y11248 = n8162 ;
  assign y11249 = ~1'b0 ;
  assign y11250 = ~1'b0 ;
  assign y11251 = n23656 ;
  assign y11252 = n23659 ;
  assign y11253 = ~1'b0 ;
  assign y11254 = ~1'b0 ;
  assign y11255 = n23660 ;
  assign y11256 = n23662 ;
  assign y11257 = n23664 ;
  assign y11258 = n23665 ;
  assign y11259 = ~n23666 ;
  assign y11260 = n23668 ;
  assign y11261 = n23674 ;
  assign y11262 = n23676 ;
  assign y11263 = ~1'b0 ;
  assign y11264 = n23677 ;
  assign y11265 = ~n23678 ;
  assign y11266 = n23681 ;
  assign y11267 = ~n23684 ;
  assign y11268 = ~1'b0 ;
  assign y11269 = ~1'b0 ;
  assign y11270 = ~n23685 ;
  assign y11271 = ~1'b0 ;
  assign y11272 = ~n23686 ;
  assign y11273 = n23687 ;
  assign y11274 = n23689 ;
  assign y11275 = n23691 ;
  assign y11276 = n23692 ;
  assign y11277 = ~1'b0 ;
  assign y11278 = ~n23694 ;
  assign y11279 = ~n23696 ;
  assign y11280 = ~1'b0 ;
  assign y11281 = n2720 ;
  assign y11282 = n23699 ;
  assign y11283 = ~n23700 ;
  assign y11284 = n23701 ;
  assign y11285 = ~n23705 ;
  assign y11286 = n23707 ;
  assign y11287 = ~n23709 ;
  assign y11288 = n23715 ;
  assign y11289 = ~1'b0 ;
  assign y11290 = n23717 ;
  assign y11291 = n23718 ;
  assign y11292 = n23719 ;
  assign y11293 = n23723 ;
  assign y11294 = n23728 ;
  assign y11295 = ~n23729 ;
  assign y11296 = ~n23731 ;
  assign y11297 = ~n23734 ;
  assign y11298 = ~n23738 ;
  assign y11299 = n7514 ;
  assign y11300 = ~n23740 ;
  assign y11301 = ~1'b0 ;
  assign y11302 = ~1'b0 ;
  assign y11303 = ~n23744 ;
  assign y11304 = n11941 ;
  assign y11305 = ~1'b0 ;
  assign y11306 = ~1'b0 ;
  assign y11307 = n19371 ;
  assign y11308 = ~n23746 ;
  assign y11309 = ~n23748 ;
  assign y11310 = ~n23750 ;
  assign y11311 = ~n23752 ;
  assign y11312 = n23753 ;
  assign y11313 = ~n23754 ;
  assign y11314 = ~n23755 ;
  assign y11315 = n23757 ;
  assign y11316 = n23759 ;
  assign y11317 = ~1'b0 ;
  assign y11318 = ~1'b0 ;
  assign y11319 = n23761 ;
  assign y11320 = ~n5724 ;
  assign y11321 = ~n13768 ;
  assign y11322 = n23762 ;
  assign y11323 = ~n23764 ;
  assign y11324 = ~n12741 ;
  assign y11325 = ~n23772 ;
  assign y11326 = ~n23773 ;
  assign y11327 = ~n23774 ;
  assign y11328 = ~n23777 ;
  assign y11329 = ~n23778 ;
  assign y11330 = ~n23780 ;
  assign y11331 = ~1'b0 ;
  assign y11332 = ~n11327 ;
  assign y11333 = n23781 ;
  assign y11334 = n23782 ;
  assign y11335 = ~1'b0 ;
  assign y11336 = ~1'b0 ;
  assign y11337 = ~n23786 ;
  assign y11338 = n23790 ;
  assign y11339 = ~n23791 ;
  assign y11340 = n23793 ;
  assign y11341 = ~1'b0 ;
  assign y11342 = n23795 ;
  assign y11343 = ~n23800 ;
  assign y11344 = ~1'b0 ;
  assign y11345 = n23801 ;
  assign y11346 = ~n23804 ;
  assign y11347 = ~1'b0 ;
  assign y11348 = ~n23807 ;
  assign y11349 = ~n23808 ;
  assign y11350 = n23810 ;
  assign y11351 = ~1'b0 ;
  assign y11352 = n23811 ;
  assign y11353 = n23814 ;
  assign y11354 = ~n9564 ;
  assign y11355 = ~n141 ;
  assign y11356 = n23816 ;
  assign y11357 = n23819 ;
  assign y11358 = ~n23820 ;
  assign y11359 = n23823 ;
  assign y11360 = n13802 ;
  assign y11361 = n23824 ;
  assign y11362 = ~n23826 ;
  assign y11363 = ~n23827 ;
  assign y11364 = n23829 ;
  assign y11365 = ~n23830 ;
  assign y11366 = ~n23834 ;
  assign y11367 = ~n23840 ;
  assign y11368 = ~1'b0 ;
  assign y11369 = ~n23842 ;
  assign y11370 = n23843 ;
  assign y11371 = ~n23845 ;
  assign y11372 = ~n23847 ;
  assign y11373 = ~n23849 ;
  assign y11374 = ~1'b0 ;
  assign y11375 = ~1'b0 ;
  assign y11376 = ~n23851 ;
  assign y11377 = ~1'b0 ;
  assign y11378 = ~n23852 ;
  assign y11379 = n23855 ;
  assign y11380 = n23857 ;
  assign y11381 = ~1'b0 ;
  assign y11382 = n23859 ;
  assign y11383 = ~1'b0 ;
  assign y11384 = 1'b0 ;
  assign y11385 = ~1'b0 ;
  assign y11386 = ~1'b0 ;
  assign y11387 = ~1'b0 ;
  assign y11388 = ~1'b0 ;
  assign y11389 = n23861 ;
  assign y11390 = n23863 ;
  assign y11391 = ~n23876 ;
  assign y11392 = ~1'b0 ;
  assign y11393 = ~n23893 ;
  assign y11394 = n23895 ;
  assign y11395 = ~1'b0 ;
  assign y11396 = ~n23897 ;
  assign y11397 = ~1'b0 ;
  assign y11398 = ~n23903 ;
  assign y11399 = n23904 ;
  assign y11400 = ~n23905 ;
  assign y11401 = ~n23909 ;
  assign y11402 = n23910 ;
  assign y11403 = n23913 ;
  assign y11404 = ~1'b0 ;
  assign y11405 = 1'b0 ;
  assign y11406 = ~1'b0 ;
  assign y11407 = n23915 ;
  assign y11408 = n23918 ;
  assign y11409 = n3070 ;
  assign y11410 = ~n23926 ;
  assign y11411 = ~1'b0 ;
  assign y11412 = ~1'b0 ;
  assign y11413 = n23928 ;
  assign y11414 = ~n23929 ;
  assign y11415 = n23931 ;
  assign y11416 = ~1'b0 ;
  assign y11417 = ~n23935 ;
  assign y11418 = n23938 ;
  assign y11419 = ~n23942 ;
  assign y11420 = n23943 ;
  assign y11421 = n23944 ;
  assign y11422 = ~n23945 ;
  assign y11423 = n23947 ;
  assign y11424 = n23949 ;
  assign y11425 = ~n23953 ;
  assign y11426 = ~n23954 ;
  assign y11427 = ~n23957 ;
  assign y11428 = n23961 ;
  assign y11429 = ~1'b0 ;
  assign y11430 = n23963 ;
  assign y11431 = n23966 ;
  assign y11432 = ~1'b0 ;
  assign y11433 = ~n23970 ;
  assign y11434 = ~1'b0 ;
  assign y11435 = ~n23974 ;
  assign y11436 = ~n23977 ;
  assign y11437 = ~n23978 ;
  assign y11438 = ~n23981 ;
  assign y11439 = ~1'b0 ;
  assign y11440 = n23983 ;
  assign y11441 = ~n23985 ;
  assign y11442 = ~n23987 ;
  assign y11443 = ~1'b0 ;
  assign y11444 = ~n23989 ;
  assign y11445 = ~n23990 ;
  assign y11446 = ~n23993 ;
  assign y11447 = n23995 ;
  assign y11448 = n23996 ;
  assign y11449 = ~n23999 ;
  assign y11450 = 1'b0 ;
  assign y11451 = ~1'b0 ;
  assign y11452 = n24001 ;
  assign y11453 = n24003 ;
  assign y11454 = ~n24004 ;
  assign y11455 = n24007 ;
  assign y11456 = n24009 ;
  assign y11457 = ~1'b0 ;
  assign y11458 = n24010 ;
  assign y11459 = ~n24016 ;
  assign y11460 = n24019 ;
  assign y11461 = ~n24021 ;
  assign y11462 = ~n24022 ;
  assign y11463 = n24024 ;
  assign y11464 = ~n24025 ;
  assign y11465 = ~n24027 ;
  assign y11466 = n24030 ;
  assign y11467 = ~1'b0 ;
  assign y11468 = n24032 ;
  assign y11469 = ~n24033 ;
  assign y11470 = ~n24034 ;
  assign y11471 = n24037 ;
  assign y11472 = ~n24038 ;
  assign y11473 = ~n24040 ;
  assign y11474 = n24041 ;
  assign y11475 = ~n24042 ;
  assign y11476 = n24043 ;
  assign y11477 = ~n24044 ;
  assign y11478 = n24046 ;
  assign y11479 = ~1'b0 ;
  assign y11480 = ~1'b0 ;
  assign y11481 = ~n23008 ;
  assign y11482 = ~n24049 ;
  assign y11483 = ~n24055 ;
  assign y11484 = ~1'b0 ;
  assign y11485 = ~n24056 ;
  assign y11486 = n24058 ;
  assign y11487 = ~n24060 ;
  assign y11488 = ~1'b0 ;
  assign y11489 = ~n24061 ;
  assign y11490 = n24062 ;
  assign y11491 = ~n24063 ;
  assign y11492 = ~1'b0 ;
  assign y11493 = ~n24065 ;
  assign y11494 = ~1'b0 ;
  assign y11495 = ~1'b0 ;
  assign y11496 = ~1'b0 ;
  assign y11497 = n24067 ;
  assign y11498 = ~n24069 ;
  assign y11499 = ~n24070 ;
  assign y11500 = n24075 ;
  assign y11501 = n24077 ;
  assign y11502 = n24078 ;
  assign y11503 = ~n24079 ;
  assign y11504 = n24081 ;
  assign y11505 = ~n24088 ;
  assign y11506 = ~n24091 ;
  assign y11507 = ~n24092 ;
  assign y11508 = ~n24094 ;
  assign y11509 = n24096 ;
  assign y11510 = n24099 ;
  assign y11511 = n3874 ;
  assign y11512 = n24105 ;
  assign y11513 = ~n24106 ;
  assign y11514 = n24107 ;
  assign y11515 = n12915 ;
  assign y11516 = n6678 ;
  assign y11517 = ~n24111 ;
  assign y11518 = ~n24113 ;
  assign y11519 = n24117 ;
  assign y11520 = ~n24122 ;
  assign y11521 = ~n24123 ;
  assign y11522 = ~n24128 ;
  assign y11523 = ~1'b0 ;
  assign y11524 = ~1'b0 ;
  assign y11525 = ~n24133 ;
  assign y11526 = ~1'b0 ;
  assign y11527 = ~1'b0 ;
  assign y11528 = ~n8197 ;
  assign y11529 = ~n24134 ;
  assign y11530 = ~n24136 ;
  assign y11531 = n18952 ;
  assign y11532 = ~n24139 ;
  assign y11533 = n24143 ;
  assign y11534 = n24145 ;
  assign y11535 = ~n24147 ;
  assign y11536 = n24148 ;
  assign y11537 = n24151 ;
  assign y11538 = n24153 ;
  assign y11539 = n24156 ;
  assign y11540 = ~n24157 ;
  assign y11541 = n24158 ;
  assign y11542 = n24159 ;
  assign y11543 = ~n24161 ;
  assign y11544 = ~1'b0 ;
  assign y11545 = ~n24164 ;
  assign y11546 = n24166 ;
  assign y11547 = ~n24167 ;
  assign y11548 = ~1'b0 ;
  assign y11549 = ~n24175 ;
  assign y11550 = ~n24176 ;
  assign y11551 = n24178 ;
  assign y11552 = ~1'b0 ;
  assign y11553 = ~n24179 ;
  assign y11554 = n24185 ;
  assign y11555 = ~n24190 ;
  assign y11556 = ~1'b0 ;
  assign y11557 = ~n24195 ;
  assign y11558 = ~1'b0 ;
  assign y11559 = ~n24197 ;
  assign y11560 = n24200 ;
  assign y11561 = ~n24203 ;
  assign y11562 = ~n24204 ;
  assign y11563 = ~1'b0 ;
  assign y11564 = ~1'b0 ;
  assign y11565 = ~n24207 ;
  assign y11566 = ~1'b0 ;
  assign y11567 = ~1'b0 ;
  assign y11568 = n24214 ;
  assign y11569 = n1183 ;
  assign y11570 = n24215 ;
  assign y11571 = n24216 ;
  assign y11572 = ~n14196 ;
  assign y11573 = ~n24217 ;
  assign y11574 = n24218 ;
  assign y11575 = ~1'b0 ;
  assign y11576 = n24224 ;
  assign y11577 = n24226 ;
  assign y11578 = ~1'b0 ;
  assign y11579 = n24227 ;
  assign y11580 = n24228 ;
  assign y11581 = ~n24232 ;
  assign y11582 = ~n24237 ;
  assign y11583 = n24240 ;
  assign y11584 = n24243 ;
  assign y11585 = ~n24246 ;
  assign y11586 = ~n24251 ;
  assign y11587 = ~1'b0 ;
  assign y11588 = n24254 ;
  assign y11589 = ~n24259 ;
  assign y11590 = ~n24261 ;
  assign y11591 = ~n24264 ;
  assign y11592 = n24267 ;
  assign y11593 = n24269 ;
  assign y11594 = ~1'b0 ;
  assign y11595 = ~n24271 ;
  assign y11596 = 1'b0 ;
  assign y11597 = n24272 ;
  assign y11598 = ~1'b0 ;
  assign y11599 = ~n24275 ;
  assign y11600 = ~n24277 ;
  assign y11601 = n24278 ;
  assign y11602 = n24279 ;
  assign y11603 = ~1'b0 ;
  assign y11604 = n24281 ;
  assign y11605 = ~n24282 ;
  assign y11606 = ~n12135 ;
  assign y11607 = n24283 ;
  assign y11608 = n24286 ;
  assign y11609 = 1'b0 ;
  assign y11610 = n24288 ;
  assign y11611 = ~n24289 ;
  assign y11612 = n24291 ;
  assign y11613 = ~n24292 ;
  assign y11614 = ~n24296 ;
  assign y11615 = n24297 ;
  assign y11616 = ~1'b0 ;
  assign y11617 = ~1'b0 ;
  assign y11618 = ~n24301 ;
  assign y11619 = ~1'b0 ;
  assign y11620 = ~1'b0 ;
  assign y11621 = ~n24303 ;
  assign y11622 = n24304 ;
  assign y11623 = ~n24306 ;
  assign y11624 = ~1'b0 ;
  assign y11625 = ~n24310 ;
  assign y11626 = ~1'b0 ;
  assign y11627 = ~n24312 ;
  assign y11628 = n24315 ;
  assign y11629 = n24316 ;
  assign y11630 = ~n24318 ;
  assign y11631 = ~n1103 ;
  assign y11632 = n24319 ;
  assign y11633 = ~n24321 ;
  assign y11634 = ~n24324 ;
  assign y11635 = ~n24328 ;
  assign y11636 = n1217 ;
  assign y11637 = n8621 ;
  assign y11638 = n8733 ;
  assign y11639 = n24330 ;
  assign y11640 = n24332 ;
  assign y11641 = ~1'b0 ;
  assign y11642 = ~1'b0 ;
  assign y11643 = n24334 ;
  assign y11644 = ~n24338 ;
  assign y11645 = ~n24340 ;
  assign y11646 = ~n24342 ;
  assign y11647 = n24343 ;
  assign y11648 = ~1'b0 ;
  assign y11649 = ~1'b0 ;
  assign y11650 = ~n24346 ;
  assign y11651 = n24348 ;
  assign y11652 = n24352 ;
  assign y11653 = ~n24353 ;
  assign y11654 = ~n24356 ;
  assign y11655 = ~n24359 ;
  assign y11656 = ~n24365 ;
  assign y11657 = ~1'b0 ;
  assign y11658 = ~n24366 ;
  assign y11659 = ~1'b0 ;
  assign y11660 = n24370 ;
  assign y11661 = ~n20123 ;
  assign y11662 = n24371 ;
  assign y11663 = ~n24375 ;
  assign y11664 = ~n24378 ;
  assign y11665 = n24381 ;
  assign y11666 = ~1'b0 ;
  assign y11667 = n24383 ;
  assign y11668 = ~1'b0 ;
  assign y11669 = ~n24386 ;
  assign y11670 = n24387 ;
  assign y11671 = ~1'b0 ;
  assign y11672 = ~n3184 ;
  assign y11673 = ~n24388 ;
  assign y11674 = ~n24393 ;
  assign y11675 = n16679 ;
  assign y11676 = n6691 ;
  assign y11677 = ~n24394 ;
  assign y11678 = ~1'b0 ;
  assign y11679 = n24396 ;
  assign y11680 = ~n24398 ;
  assign y11681 = n24400 ;
  assign y11682 = ~n24401 ;
  assign y11683 = ~1'b0 ;
  assign y11684 = ~1'b0 ;
  assign y11685 = n4796 ;
  assign y11686 = n24405 ;
  assign y11687 = n24406 ;
  assign y11688 = ~n24410 ;
  assign y11689 = ~n24411 ;
  assign y11690 = n24413 ;
  assign y11691 = ~n24415 ;
  assign y11692 = ~n24421 ;
  assign y11693 = n24423 ;
  assign y11694 = n24424 ;
  assign y11695 = ~1'b0 ;
  assign y11696 = ~1'b0 ;
  assign y11697 = ~n24426 ;
  assign y11698 = ~n24427 ;
  assign y11699 = n24428 ;
  assign y11700 = n24429 ;
  assign y11701 = ~n24432 ;
  assign y11702 = n24435 ;
  assign y11703 = ~n24436 ;
  assign y11704 = ~n19978 ;
  assign y11705 = ~n24438 ;
  assign y11706 = ~n24440 ;
  assign y11707 = ~1'b0 ;
  assign y11708 = ~n24441 ;
  assign y11709 = n24442 ;
  assign y11710 = n24448 ;
  assign y11711 = n24456 ;
  assign y11712 = ~n24458 ;
  assign y11713 = ~n9952 ;
  assign y11714 = n24461 ;
  assign y11715 = ~1'b0 ;
  assign y11716 = n24464 ;
  assign y11717 = n24465 ;
  assign y11718 = ~1'b0 ;
  assign y11719 = ~n24468 ;
  assign y11720 = ~1'b0 ;
  assign y11721 = n24470 ;
  assign y11722 = ~n24471 ;
  assign y11723 = n24472 ;
  assign y11724 = n24477 ;
  assign y11725 = n24479 ;
  assign y11726 = n24483 ;
  assign y11727 = ~1'b0 ;
  assign y11728 = n24487 ;
  assign y11729 = ~n24488 ;
  assign y11730 = ~1'b0 ;
  assign y11731 = n895 ;
  assign y11732 = ~n24489 ;
  assign y11733 = n24494 ;
  assign y11734 = n24496 ;
  assign y11735 = n24498 ;
  assign y11736 = ~1'b0 ;
  assign y11737 = ~n24499 ;
  assign y11738 = ~n24500 ;
  assign y11739 = n24502 ;
  assign y11740 = ~n24503 ;
  assign y11741 = n24507 ;
  assign y11742 = ~n24510 ;
  assign y11743 = ~n24514 ;
  assign y11744 = ~n24518 ;
  assign y11745 = n24523 ;
  assign y11746 = n24039 ;
  assign y11747 = n24525 ;
  assign y11748 = n24527 ;
  assign y11749 = ~n24529 ;
  assign y11750 = n24531 ;
  assign y11751 = ~n5861 ;
  assign y11752 = ~n24534 ;
  assign y11753 = ~1'b0 ;
  assign y11754 = n24543 ;
  assign y11755 = ~1'b0 ;
  assign y11756 = ~1'b0 ;
  assign y11757 = n24545 ;
  assign y11758 = ~n24546 ;
  assign y11759 = ~n24548 ;
  assign y11760 = n24551 ;
  assign y11761 = ~n24556 ;
  assign y11762 = ~n24560 ;
  assign y11763 = ~1'b0 ;
  assign y11764 = ~1'b0 ;
  assign y11765 = n24561 ;
  assign y11766 = ~n24563 ;
  assign y11767 = ~1'b0 ;
  assign y11768 = ~n24567 ;
  assign y11769 = n24568 ;
  assign y11770 = ~n24569 ;
  assign y11771 = n24571 ;
  assign y11772 = ~n24572 ;
  assign y11773 = ~n24576 ;
  assign y11774 = ~n24577 ;
  assign y11775 = n24580 ;
  assign y11776 = n24583 ;
  assign y11777 = ~n24585 ;
  assign y11778 = ~n24586 ;
  assign y11779 = n24587 ;
  assign y11780 = n24588 ;
  assign y11781 = ~n24590 ;
  assign y11782 = ~n24593 ;
  assign y11783 = n24597 ;
  assign y11784 = ~n1568 ;
  assign y11785 = ~1'b0 ;
  assign y11786 = ~1'b0 ;
  assign y11787 = ~x7 ;
  assign y11788 = ~n24598 ;
  assign y11789 = n24599 ;
  assign y11790 = ~n24610 ;
  assign y11791 = ~1'b0 ;
  assign y11792 = n24612 ;
  assign y11793 = n24613 ;
  assign y11794 = ~n24615 ;
  assign y11795 = ~n24617 ;
  assign y11796 = ~1'b0 ;
  assign y11797 = 1'b0 ;
  assign y11798 = ~n24620 ;
  assign y11799 = n723 ;
  assign y11800 = ~n24621 ;
  assign y11801 = ~1'b0 ;
  assign y11802 = n10623 ;
  assign y11803 = ~n24624 ;
  assign y11804 = ~1'b0 ;
  assign y11805 = n24626 ;
  assign y11806 = ~n24628 ;
  assign y11807 = ~1'b0 ;
  assign y11808 = n24634 ;
  assign y11809 = ~n19566 ;
  assign y11810 = n24636 ;
  assign y11811 = ~n24638 ;
  assign y11812 = ~n24640 ;
  assign y11813 = ~n24643 ;
  assign y11814 = ~1'b0 ;
  assign y11815 = n24647 ;
  assign y11816 = ~n24649 ;
  assign y11817 = ~n24651 ;
  assign y11818 = ~n24652 ;
  assign y11819 = n24653 ;
  assign y11820 = n24656 ;
  assign y11821 = ~1'b0 ;
  assign y11822 = n24657 ;
  assign y11823 = ~n24659 ;
  assign y11824 = ~n24661 ;
  assign y11825 = n24663 ;
  assign y11826 = ~n24667 ;
  assign y11827 = ~1'b0 ;
  assign y11828 = n24669 ;
  assign y11829 = ~n24671 ;
  assign y11830 = ~n24672 ;
  assign y11831 = ~1'b0 ;
  assign y11832 = n24673 ;
  assign y11833 = n24674 ;
  assign y11834 = n977 ;
  assign y11835 = ~n24678 ;
  assign y11836 = ~n24680 ;
  assign y11837 = ~n24681 ;
  assign y11838 = n24682 ;
  assign y11839 = n20322 ;
  assign y11840 = ~1'b0 ;
  assign y11841 = ~n24686 ;
  assign y11842 = n24687 ;
  assign y11843 = n24688 ;
  assign y11844 = n24689 ;
  assign y11845 = n24690 ;
  assign y11846 = ~1'b0 ;
  assign y11847 = ~1'b0 ;
  assign y11848 = n24691 ;
  assign y11849 = n24696 ;
  assign y11850 = n24703 ;
  assign y11851 = ~n24707 ;
  assign y11852 = n24708 ;
  assign y11853 = n24710 ;
  assign y11854 = ~n24712 ;
  assign y11855 = n14078 ;
  assign y11856 = n24715 ;
  assign y11857 = ~n24720 ;
  assign y11858 = ~n24726 ;
  assign y11859 = n24727 ;
  assign y11860 = ~n24728 ;
  assign y11861 = ~1'b0 ;
  assign y11862 = n24729 ;
  assign y11863 = ~n24731 ;
  assign y11864 = ~1'b0 ;
  assign y11865 = ~n24733 ;
  assign y11866 = n24736 ;
  assign y11867 = ~1'b0 ;
  assign y11868 = ~n961 ;
  assign y11869 = n24737 ;
  assign y11870 = ~n24740 ;
  assign y11871 = ~n24744 ;
  assign y11872 = n24746 ;
  assign y11873 = n24752 ;
  assign y11874 = ~1'b0 ;
  assign y11875 = ~n24754 ;
  assign y11876 = ~n24755 ;
  assign y11877 = n24758 ;
  assign y11878 = n24759 ;
  assign y11879 = n24762 ;
  assign y11880 = ~1'b0 ;
  assign y11881 = ~n10662 ;
  assign y11882 = ~n24766 ;
  assign y11883 = n24768 ;
  assign y11884 = ~1'b0 ;
  assign y11885 = ~n24769 ;
  assign y11886 = ~1'b0 ;
  assign y11887 = n24775 ;
  assign y11888 = n24776 ;
  assign y11889 = n21852 ;
  assign y11890 = ~1'b0 ;
  assign y11891 = ~1'b0 ;
  assign y11892 = n24777 ;
  assign y11893 = n24781 ;
  assign y11894 = ~1'b0 ;
  assign y11895 = n24786 ;
  assign y11896 = n24787 ;
  assign y11897 = n24788 ;
  assign y11898 = n24790 ;
  assign y11899 = n24791 ;
  assign y11900 = ~1'b0 ;
  assign y11901 = ~n24793 ;
  assign y11902 = n24797 ;
  assign y11903 = ~n6638 ;
  assign y11904 = ~n24800 ;
  assign y11905 = n24802 ;
  assign y11906 = ~n24804 ;
  assign y11907 = ~n24807 ;
  assign y11908 = ~n24826 ;
  assign y11909 = n24830 ;
  assign y11910 = ~n24834 ;
  assign y11911 = n24836 ;
  assign y11912 = n24837 ;
  assign y11913 = n24839 ;
  assign y11914 = n24840 ;
  assign y11915 = n24842 ;
  assign y11916 = n24845 ;
  assign y11917 = ~n24848 ;
  assign y11918 = n24849 ;
  assign y11919 = ~n872 ;
  assign y11920 = ~1'b0 ;
  assign y11921 = ~1'b0 ;
  assign y11922 = n22857 ;
  assign y11923 = ~n24850 ;
  assign y11924 = n24853 ;
  assign y11925 = n24856 ;
  assign y11926 = ~n24858 ;
  assign y11927 = n24859 ;
  assign y11928 = n24861 ;
  assign y11929 = n24862 ;
  assign y11930 = 1'b0 ;
  assign y11931 = 1'b0 ;
  assign y11932 = ~1'b0 ;
  assign y11933 = ~1'b0 ;
  assign y11934 = ~n24865 ;
  assign y11935 = ~n24866 ;
  assign y11936 = n24873 ;
  assign y11937 = n24881 ;
  assign y11938 = ~1'b0 ;
  assign y11939 = ~n24885 ;
  assign y11940 = ~n24889 ;
  assign y11941 = ~1'b0 ;
  assign y11942 = n24890 ;
  assign y11943 = ~1'b0 ;
  assign y11944 = ~n24891 ;
  assign y11945 = ~n24894 ;
  assign y11946 = ~1'b0 ;
  assign y11947 = n24896 ;
  assign y11948 = n24897 ;
  assign y11949 = ~n24899 ;
  assign y11950 = ~n24902 ;
  assign y11951 = n24904 ;
  assign y11952 = ~n24906 ;
  assign y11953 = ~1'b0 ;
  assign y11954 = n24907 ;
  assign y11955 = ~n24910 ;
  assign y11956 = n24912 ;
  assign y11957 = ~n24913 ;
  assign y11958 = ~1'b0 ;
  assign y11959 = n24915 ;
  assign y11960 = n24918 ;
  assign y11961 = n24921 ;
  assign y11962 = ~n24922 ;
  assign y11963 = n24926 ;
  assign y11964 = n24930 ;
  assign y11965 = ~n24933 ;
  assign y11966 = ~n24936 ;
  assign y11967 = ~1'b0 ;
  assign y11968 = ~1'b0 ;
  assign y11969 = ~1'b0 ;
  assign y11970 = ~n24939 ;
  assign y11971 = ~n24941 ;
  assign y11972 = ~1'b0 ;
  assign y11973 = ~n24945 ;
  assign y11974 = n24950 ;
  assign y11975 = ~n24956 ;
  assign y11976 = ~n24959 ;
  assign y11977 = ~1'b0 ;
  assign y11978 = ~n24960 ;
  assign y11979 = ~1'b0 ;
  assign y11980 = ~n24962 ;
  assign y11981 = ~n24964 ;
  assign y11982 = ~n24969 ;
  assign y11983 = n24970 ;
  assign y11984 = ~1'b0 ;
  assign y11985 = n24977 ;
  assign y11986 = ~n24978 ;
  assign y11987 = n24982 ;
  assign y11988 = ~n24986 ;
  assign y11989 = ~1'b0 ;
  assign y11990 = n24987 ;
  assign y11991 = ~1'b0 ;
  assign y11992 = ~1'b0 ;
  assign y11993 = ~1'b0 ;
  assign y11994 = 1'b0 ;
  assign y11995 = n24988 ;
  assign y11996 = n24990 ;
  assign y11997 = ~n14371 ;
  assign y11998 = n24991 ;
  assign y11999 = n24997 ;
  assign y12000 = ~1'b0 ;
  assign y12001 = ~n25001 ;
  assign y12002 = n25004 ;
  assign y12003 = ~n25005 ;
  assign y12004 = ~x26 ;
  assign y12005 = n25006 ;
  assign y12006 = n25008 ;
  assign y12007 = n25009 ;
  assign y12008 = ~1'b0 ;
  assign y12009 = ~n25011 ;
  assign y12010 = n25015 ;
  assign y12011 = ~1'b0 ;
  assign y12012 = n25017 ;
  assign y12013 = ~n25018 ;
  assign y12014 = ~1'b0 ;
  assign y12015 = ~n25020 ;
  assign y12016 = n25021 ;
  assign y12017 = ~n25023 ;
  assign y12018 = ~n25024 ;
  assign y12019 = n25026 ;
  assign y12020 = n25031 ;
  assign y12021 = 1'b0 ;
  assign y12022 = ~1'b0 ;
  assign y12023 = n25032 ;
  assign y12024 = n25033 ;
  assign y12025 = ~1'b0 ;
  assign y12026 = n25035 ;
  assign y12027 = n25036 ;
  assign y12028 = n25038 ;
  assign y12029 = ~1'b0 ;
  assign y12030 = n25039 ;
  assign y12031 = n25042 ;
  assign y12032 = ~n25044 ;
  assign y12033 = ~n25045 ;
  assign y12034 = ~n25047 ;
  assign y12035 = ~n25051 ;
  assign y12036 = n25055 ;
  assign y12037 = n25056 ;
  assign y12038 = n25057 ;
  assign y12039 = n25059 ;
  assign y12040 = ~n25062 ;
  assign y12041 = n25067 ;
  assign y12042 = n25068 ;
  assign y12043 = ~n25072 ;
  assign y12044 = ~n25076 ;
  assign y12045 = ~1'b0 ;
  assign y12046 = ~1'b0 ;
  assign y12047 = n25079 ;
  assign y12048 = n25082 ;
  assign y12049 = ~n25087 ;
  assign y12050 = ~1'b0 ;
  assign y12051 = ~n25089 ;
  assign y12052 = ~1'b0 ;
  assign y12053 = ~n25091 ;
  assign y12054 = n17504 ;
  assign y12055 = ~n25102 ;
  assign y12056 = n25105 ;
  assign y12057 = n25113 ;
  assign y12058 = ~1'b0 ;
  assign y12059 = ~1'b0 ;
  assign y12060 = ~n25115 ;
  assign y12061 = n25116 ;
  assign y12062 = ~n25118 ;
  assign y12063 = n25120 ;
  assign y12064 = ~n25123 ;
  assign y12065 = ~n25125 ;
  assign y12066 = ~n25126 ;
  assign y12067 = n25127 ;
  assign y12068 = ~1'b0 ;
  assign y12069 = n25131 ;
  assign y12070 = ~n25134 ;
  assign y12071 = ~1'b0 ;
  assign y12072 = n25135 ;
  assign y12073 = n25137 ;
  assign y12074 = ~1'b0 ;
  assign y12075 = n25141 ;
  assign y12076 = ~1'b0 ;
  assign y12077 = ~n25144 ;
  assign y12078 = n25145 ;
  assign y12079 = ~1'b0 ;
  assign y12080 = ~n25147 ;
  assign y12081 = ~n25149 ;
  assign y12082 = ~n25151 ;
  assign y12083 = ~n25154 ;
  assign y12084 = ~n25156 ;
  assign y12085 = ~1'b0 ;
  assign y12086 = ~1'b0 ;
  assign y12087 = ~n25157 ;
  assign y12088 = n25158 ;
  assign y12089 = ~n25160 ;
  assign y12090 = n25161 ;
  assign y12091 = n25164 ;
  assign y12092 = ~1'b0 ;
  assign y12093 = n25166 ;
  assign y12094 = 1'b0 ;
  assign y12095 = ~1'b0 ;
  assign y12096 = ~1'b0 ;
  assign y12097 = ~1'b0 ;
  assign y12098 = ~n25167 ;
  assign y12099 = ~n25169 ;
  assign y12100 = n25170 ;
  assign y12101 = ~n25171 ;
  assign y12102 = n25179 ;
  assign y12103 = ~1'b0 ;
  assign y12104 = n25181 ;
  assign y12105 = ~1'b0 ;
  assign y12106 = ~n25182 ;
  assign y12107 = n25183 ;
  assign y12108 = n25184 ;
  assign y12109 = ~n25185 ;
  assign y12110 = n25186 ;
  assign y12111 = n25189 ;
  assign y12112 = ~1'b0 ;
  assign y12113 = ~1'b0 ;
  assign y12114 = ~1'b0 ;
  assign y12115 = ~n25191 ;
  assign y12116 = ~1'b0 ;
  assign y12117 = ~n25192 ;
  assign y12118 = n25199 ;
  assign y12119 = n25202 ;
  assign y12120 = n25205 ;
  assign y12121 = ~n25207 ;
  assign y12122 = ~1'b0 ;
  assign y12123 = ~n25208 ;
  assign y12124 = n25209 ;
  assign y12125 = ~1'b0 ;
  assign y12126 = n25211 ;
  assign y12127 = n25215 ;
  assign y12128 = n25216 ;
  assign y12129 = n25218 ;
  assign y12130 = ~n25219 ;
  assign y12131 = n25221 ;
  assign y12132 = n25222 ;
  assign y12133 = n25226 ;
  assign y12134 = ~1'b0 ;
  assign y12135 = ~n25228 ;
  assign y12136 = ~1'b0 ;
  assign y12137 = ~1'b0 ;
  assign y12138 = ~n25232 ;
  assign y12139 = ~n25233 ;
  assign y12140 = n25234 ;
  assign y12141 = n25235 ;
  assign y12142 = ~n25237 ;
  assign y12143 = ~n25238 ;
  assign y12144 = ~1'b0 ;
  assign y12145 = ~1'b0 ;
  assign y12146 = ~n25241 ;
  assign y12147 = ~1'b0 ;
  assign y12148 = ~1'b0 ;
  assign y12149 = n25245 ;
  assign y12150 = ~n25247 ;
  assign y12151 = ~n25249 ;
  assign y12152 = n25251 ;
  assign y12153 = ~n25255 ;
  assign y12154 = n25257 ;
  assign y12155 = n25259 ;
  assign y12156 = ~n25261 ;
  assign y12157 = n25262 ;
  assign y12158 = ~n25263 ;
  assign y12159 = ~n25265 ;
  assign y12160 = ~n25268 ;
  assign y12161 = n25272 ;
  assign y12162 = n25273 ;
  assign y12163 = ~1'b0 ;
  assign y12164 = ~n25275 ;
  assign y12165 = ~n25277 ;
  assign y12166 = n25279 ;
  assign y12167 = n25281 ;
  assign y12168 = n25286 ;
  assign y12169 = ~1'b0 ;
  assign y12170 = ~1'b0 ;
  assign y12171 = ~n25289 ;
  assign y12172 = n25295 ;
  assign y12173 = n25299 ;
  assign y12174 = ~1'b0 ;
  assign y12175 = ~n21481 ;
  assign y12176 = ~n25303 ;
  assign y12177 = n25307 ;
  assign y12178 = n25312 ;
  assign y12179 = ~1'b0 ;
  assign y12180 = n25319 ;
  assign y12181 = ~n22746 ;
  assign y12182 = n6007 ;
  assign y12183 = n25321 ;
  assign y12184 = n25322 ;
  assign y12185 = n25323 ;
  assign y12186 = ~1'b0 ;
  assign y12187 = ~n25327 ;
  assign y12188 = ~n25328 ;
  assign y12189 = ~n25332 ;
  assign y12190 = n25333 ;
  assign y12191 = n25334 ;
  assign y12192 = ~1'b0 ;
  assign y12193 = ~n25335 ;
  assign y12194 = ~1'b0 ;
  assign y12195 = ~n25336 ;
  assign y12196 = ~n25341 ;
  assign y12197 = ~n25347 ;
  assign y12198 = n25349 ;
  assign y12199 = ~n25351 ;
  assign y12200 = n25354 ;
  assign y12201 = n25356 ;
  assign y12202 = ~n25363 ;
  assign y12203 = n25364 ;
  assign y12204 = ~1'b0 ;
  assign y12205 = ~n25365 ;
  assign y12206 = ~1'b0 ;
  assign y12207 = ~n25366 ;
  assign y12208 = n25368 ;
  assign y12209 = n25370 ;
  assign y12210 = n25371 ;
  assign y12211 = ~n25374 ;
  assign y12212 = ~1'b0 ;
  assign y12213 = ~n25376 ;
  assign y12214 = ~n25377 ;
  assign y12215 = ~1'b0 ;
  assign y12216 = n12932 ;
  assign y12217 = ~1'b0 ;
  assign y12218 = n25380 ;
  assign y12219 = ~n25381 ;
  assign y12220 = ~n13003 ;
  assign y12221 = ~n25384 ;
  assign y12222 = ~1'b0 ;
  assign y12223 = ~1'b0 ;
  assign y12224 = ~1'b0 ;
  assign y12225 = n25386 ;
  assign y12226 = ~n25387 ;
  assign y12227 = n8509 ;
  assign y12228 = ~n25392 ;
  assign y12229 = ~1'b0 ;
  assign y12230 = n25396 ;
  assign y12231 = n25397 ;
  assign y12232 = n25401 ;
  assign y12233 = n25404 ;
  assign y12234 = n25406 ;
  assign y12235 = ~n25407 ;
  assign y12236 = n25408 ;
  assign y12237 = n25411 ;
  assign y12238 = n25416 ;
  assign y12239 = ~n25421 ;
  assign y12240 = ~1'b0 ;
  assign y12241 = ~1'b0 ;
  assign y12242 = n25423 ;
  assign y12243 = n25428 ;
  assign y12244 = ~n25431 ;
  assign y12245 = ~n25433 ;
  assign y12246 = ~n25435 ;
  assign y12247 = n3596 ;
  assign y12248 = ~n25437 ;
  assign y12249 = ~n25439 ;
  assign y12250 = ~n25442 ;
  assign y12251 = ~1'b0 ;
  assign y12252 = n25444 ;
  assign y12253 = ~n25449 ;
  assign y12254 = ~n25450 ;
  assign y12255 = ~n25451 ;
  assign y12256 = ~1'b0 ;
  assign y12257 = ~1'b0 ;
  assign y12258 = ~n25453 ;
  assign y12259 = ~n25457 ;
  assign y12260 = ~1'b0 ;
  assign y12261 = ~1'b0 ;
  assign y12262 = ~n25458 ;
  assign y12263 = n25461 ;
  assign y12264 = ~n19362 ;
  assign y12265 = ~1'b0 ;
  assign y12266 = n25463 ;
  assign y12267 = n25466 ;
  assign y12268 = ~1'b0 ;
  assign y12269 = ~1'b0 ;
  assign y12270 = ~1'b0 ;
  assign y12271 = ~n25469 ;
  assign y12272 = n25474 ;
  assign y12273 = n25475 ;
  assign y12274 = ~n25477 ;
  assign y12275 = n25479 ;
  assign y12276 = ~1'b0 ;
  assign y12277 = ~1'b0 ;
  assign y12278 = ~1'b0 ;
  assign y12279 = ~1'b0 ;
  assign y12280 = ~n25480 ;
  assign y12281 = n25481 ;
  assign y12282 = n25486 ;
  assign y12283 = n25489 ;
  assign y12284 = ~1'b0 ;
  assign y12285 = ~1'b0 ;
  assign y12286 = ~1'b0 ;
  assign y12287 = ~n25491 ;
  assign y12288 = ~n2706 ;
  assign y12289 = ~1'b0 ;
  assign y12290 = n25493 ;
  assign y12291 = n25496 ;
  assign y12292 = ~n25498 ;
  assign y12293 = n25499 ;
  assign y12294 = ~n25501 ;
  assign y12295 = ~n25503 ;
  assign y12296 = ~1'b0 ;
  assign y12297 = ~n25504 ;
  assign y12298 = ~1'b0 ;
  assign y12299 = ~1'b0 ;
  assign y12300 = ~1'b0 ;
  assign y12301 = ~1'b0 ;
  assign y12302 = ~1'b0 ;
  assign y12303 = 1'b0 ;
  assign y12304 = n25507 ;
  assign y12305 = ~n25508 ;
  assign y12306 = n25514 ;
  assign y12307 = n25517 ;
  assign y12308 = ~1'b0 ;
  assign y12309 = ~n25523 ;
  assign y12310 = ~1'b0 ;
  assign y12311 = ~1'b0 ;
  assign y12312 = ~1'b0 ;
  assign y12313 = ~n25524 ;
  assign y12314 = ~n25525 ;
  assign y12315 = ~n25528 ;
  assign y12316 = ~1'b0 ;
  assign y12317 = ~n25530 ;
  assign y12318 = n25531 ;
  assign y12319 = ~1'b0 ;
  assign y12320 = n6376 ;
  assign y12321 = n3402 ;
  assign y12322 = n12401 ;
  assign y12323 = n25533 ;
  assign y12324 = ~n25534 ;
  assign y12325 = ~1'b0 ;
  assign y12326 = n25536 ;
  assign y12327 = 1'b0 ;
  assign y12328 = ~n25539 ;
  assign y12329 = ~n25540 ;
  assign y12330 = ~n25543 ;
  assign y12331 = ~1'b0 ;
  assign y12332 = ~n25544 ;
  assign y12333 = n25546 ;
  assign y12334 = ~n25547 ;
  assign y12335 = n25550 ;
  assign y12336 = ~n25551 ;
  assign y12337 = ~n25553 ;
  assign y12338 = 1'b0 ;
  assign y12339 = ~n25555 ;
  assign y12340 = ~n25558 ;
  assign y12341 = n25562 ;
  assign y12342 = ~n25565 ;
  assign y12343 = n25566 ;
  assign y12344 = ~1'b0 ;
  assign y12345 = ~n25570 ;
  assign y12346 = ~n25573 ;
  assign y12347 = ~n25575 ;
  assign y12348 = ~1'b0 ;
  assign y12349 = ~1'b0 ;
  assign y12350 = ~n25577 ;
  assign y12351 = ~n4230 ;
  assign y12352 = ~n25579 ;
  assign y12353 = n25581 ;
  assign y12354 = ~n25585 ;
  assign y12355 = ~n25586 ;
  assign y12356 = n25589 ;
  assign y12357 = ~n25591 ;
  assign y12358 = ~n25592 ;
  assign y12359 = ~1'b0 ;
  assign y12360 = ~n25596 ;
  assign y12361 = ~1'b0 ;
  assign y12362 = ~1'b0 ;
  assign y12363 = ~1'b0 ;
  assign y12364 = ~1'b0 ;
  assign y12365 = ~n25597 ;
  assign y12366 = ~n25602 ;
  assign y12367 = n25604 ;
  assign y12368 = n25605 ;
  assign y12369 = n25607 ;
  assign y12370 = ~n25614 ;
  assign y12371 = ~1'b0 ;
  assign y12372 = ~n25616 ;
  assign y12373 = n25617 ;
  assign y12374 = ~n25618 ;
  assign y12375 = ~n25622 ;
  assign y12376 = n14889 ;
  assign y12377 = ~n25625 ;
  assign y12378 = n25626 ;
  assign y12379 = n25628 ;
  assign y12380 = ~n25629 ;
  assign y12381 = n25630 ;
  assign y12382 = ~1'b0 ;
  assign y12383 = ~1'b0 ;
  assign y12384 = ~n25633 ;
  assign y12385 = ~n7080 ;
  assign y12386 = n25634 ;
  assign y12387 = ~n25636 ;
  assign y12388 = ~n25641 ;
  assign y12389 = ~1'b0 ;
  assign y12390 = n25642 ;
  assign y12391 = ~1'b0 ;
  assign y12392 = ~1'b0 ;
  assign y12393 = n25646 ;
  assign y12394 = ~n25647 ;
  assign y12395 = n25649 ;
  assign y12396 = ~n25650 ;
  assign y12397 = n25651 ;
  assign y12398 = ~n25655 ;
  assign y12399 = n25659 ;
  assign y12400 = ~n25661 ;
  assign y12401 = n25662 ;
  assign y12402 = n25664 ;
  assign y12403 = ~1'b0 ;
  assign y12404 = ~n5640 ;
  assign y12405 = ~n25672 ;
  assign y12406 = n25674 ;
  assign y12407 = n25675 ;
  assign y12408 = ~n25676 ;
  assign y12409 = ~1'b0 ;
  assign y12410 = n25677 ;
  assign y12411 = n25678 ;
  assign y12412 = ~n25679 ;
  assign y12413 = n25681 ;
  assign y12414 = ~n25682 ;
  assign y12415 = ~n25683 ;
  assign y12416 = n25686 ;
  assign y12417 = ~1'b0 ;
  assign y12418 = ~n25687 ;
  assign y12419 = ~1'b0 ;
  assign y12420 = ~1'b0 ;
  assign y12421 = ~n25689 ;
  assign y12422 = n25691 ;
  assign y12423 = ~n25692 ;
  assign y12424 = ~1'b0 ;
  assign y12425 = ~1'b0 ;
  assign y12426 = ~n25695 ;
  assign y12427 = n25696 ;
  assign y12428 = ~n25697 ;
  assign y12429 = ~n25701 ;
  assign y12430 = n25702 ;
  assign y12431 = ~n25706 ;
  assign y12432 = ~n25707 ;
  assign y12433 = n25708 ;
  assign y12434 = n25712 ;
  assign y12435 = ~1'b0 ;
  assign y12436 = ~1'b0 ;
  assign y12437 = ~n25714 ;
  assign y12438 = ~1'b0 ;
  assign y12439 = ~1'b0 ;
  assign y12440 = n25715 ;
  assign y12441 = ~n25717 ;
  assign y12442 = ~1'b0 ;
  assign y12443 = ~1'b0 ;
  assign y12444 = ~n25720 ;
  assign y12445 = 1'b0 ;
  assign y12446 = ~n25723 ;
  assign y12447 = ~n25726 ;
  assign y12448 = n25730 ;
  assign y12449 = ~n25732 ;
  assign y12450 = ~1'b0 ;
  assign y12451 = n25733 ;
  assign y12452 = n25736 ;
  assign y12453 = ~1'b0 ;
  assign y12454 = n25738 ;
  assign y12455 = ~n25740 ;
  assign y12456 = ~n25746 ;
  assign y12457 = ~1'b0 ;
  assign y12458 = n25747 ;
  assign y12459 = ~n25748 ;
  assign y12460 = ~1'b0 ;
  assign y12461 = ~1'b0 ;
  assign y12462 = ~n25751 ;
  assign y12463 = n25754 ;
  assign y12464 = ~n25756 ;
  assign y12465 = ~n25757 ;
  assign y12466 = n25758 ;
  assign y12467 = ~n25763 ;
  assign y12468 = n25767 ;
  assign y12469 = ~n25768 ;
  assign y12470 = ~n25769 ;
  assign y12471 = ~1'b0 ;
  assign y12472 = ~n25770 ;
  assign y12473 = ~1'b0 ;
  assign y12474 = n21303 ;
  assign y12475 = ~n25772 ;
  assign y12476 = ~1'b0 ;
  assign y12477 = ~n25775 ;
  assign y12478 = ~n25777 ;
  assign y12479 = ~n25780 ;
  assign y12480 = ~n25782 ;
  assign y12481 = n25784 ;
  assign y12482 = n16274 ;
  assign y12483 = ~n25785 ;
  assign y12484 = n25791 ;
  assign y12485 = n25792 ;
  assign y12486 = ~n25796 ;
  assign y12487 = ~1'b0 ;
  assign y12488 = ~n25800 ;
  assign y12489 = n25803 ;
  assign y12490 = n25804 ;
  assign y12491 = ~1'b0 ;
  assign y12492 = n25805 ;
  assign y12493 = ~n22460 ;
  assign y12494 = n25807 ;
  assign y12495 = ~n25808 ;
  assign y12496 = n25809 ;
  assign y12497 = n25810 ;
  assign y12498 = n25812 ;
  assign y12499 = ~n25813 ;
  assign y12500 = ~n25819 ;
  assign y12501 = n4354 ;
  assign y12502 = n10281 ;
  assign y12503 = ~n25822 ;
  assign y12504 = ~n25824 ;
  assign y12505 = ~n25827 ;
  assign y12506 = ~1'b0 ;
  assign y12507 = ~1'b0 ;
  assign y12508 = n25829 ;
  assign y12509 = ~n25832 ;
  assign y12510 = n25833 ;
  assign y12511 = ~n25837 ;
  assign y12512 = ~n25839 ;
  assign y12513 = n25845 ;
  assign y12514 = n25848 ;
  assign y12515 = n25850 ;
  assign y12516 = ~1'b0 ;
  assign y12517 = n9925 ;
  assign y12518 = ~1'b0 ;
  assign y12519 = ~1'b0 ;
  assign y12520 = ~n25855 ;
  assign y12521 = n25860 ;
  assign y12522 = ~1'b0 ;
  assign y12523 = ~n25861 ;
  assign y12524 = ~n25862 ;
  assign y12525 = n25863 ;
  assign y12526 = ~1'b0 ;
  assign y12527 = n6010 ;
  assign y12528 = ~1'b0 ;
  assign y12529 = n20815 ;
  assign y12530 = n25866 ;
  assign y12531 = ~n25868 ;
  assign y12532 = ~1'b0 ;
  assign y12533 = n25870 ;
  assign y12534 = ~1'b0 ;
  assign y12535 = ~1'b0 ;
  assign y12536 = n25871 ;
  assign y12537 = n25875 ;
  assign y12538 = n25877 ;
  assign y12539 = n25878 ;
  assign y12540 = ~n22603 ;
  assign y12541 = n25881 ;
  assign y12542 = ~1'b0 ;
  assign y12543 = n17010 ;
  assign y12544 = n25886 ;
  assign y12545 = ~n25888 ;
  assign y12546 = ~1'b0 ;
  assign y12547 = ~1'b0 ;
  assign y12548 = ~1'b0 ;
  assign y12549 = ~n25891 ;
  assign y12550 = n25895 ;
  assign y12551 = n25899 ;
  assign y12552 = ~n25900 ;
  assign y12553 = ~n25904 ;
  assign y12554 = n25907 ;
  assign y12555 = n25909 ;
  assign y12556 = n25913 ;
  assign y12557 = ~1'b0 ;
  assign y12558 = n25916 ;
  assign y12559 = n25917 ;
  assign y12560 = n25921 ;
  assign y12561 = n25925 ;
  assign y12562 = ~n25928 ;
  assign y12563 = n16270 ;
  assign y12564 = ~n25932 ;
  assign y12565 = ~1'b0 ;
  assign y12566 = ~1'b0 ;
  assign y12567 = ~n25934 ;
  assign y12568 = n25936 ;
  assign y12569 = n25939 ;
  assign y12570 = n25943 ;
  assign y12571 = ~n25944 ;
  assign y12572 = n25947 ;
  assign y12573 = ~n25948 ;
  assign y12574 = ~1'b0 ;
  assign y12575 = n25949 ;
  assign y12576 = ~1'b0 ;
  assign y12577 = ~n25955 ;
  assign y12578 = ~1'b0 ;
  assign y12579 = n25957 ;
  assign y12580 = n10284 ;
  assign y12581 = ~n25963 ;
  assign y12582 = ~n25973 ;
  assign y12583 = n25974 ;
  assign y12584 = ~n25977 ;
  assign y12585 = ~1'b0 ;
  assign y12586 = ~1'b0 ;
  assign y12587 = ~1'b0 ;
  assign y12588 = n25978 ;
  assign y12589 = n25979 ;
  assign y12590 = ~1'b0 ;
  assign y12591 = ~1'b0 ;
  assign y12592 = ~n25981 ;
  assign y12593 = n8320 ;
  assign y12594 = n11396 ;
  assign y12595 = ~1'b0 ;
  assign y12596 = ~n25985 ;
  assign y12597 = 1'b0 ;
  assign y12598 = ~1'b0 ;
  assign y12599 = ~n25987 ;
  assign y12600 = ~1'b0 ;
  assign y12601 = ~n25989 ;
  assign y12602 = ~n25991 ;
  assign y12603 = n25992 ;
  assign y12604 = 1'b0 ;
  assign y12605 = ~n25993 ;
  assign y12606 = ~n25995 ;
  assign y12607 = ~n4024 ;
  assign y12608 = ~1'b0 ;
  assign y12609 = ~n25998 ;
  assign y12610 = ~1'b0 ;
  assign y12611 = n25999 ;
  assign y12612 = ~n1360 ;
  assign y12613 = n26001 ;
  assign y12614 = n23722 ;
  assign y12615 = ~n26002 ;
  assign y12616 = n26003 ;
  assign y12617 = ~1'b0 ;
  assign y12618 = ~1'b0 ;
  assign y12619 = ~1'b0 ;
  assign y12620 = ~n26007 ;
  assign y12621 = n26009 ;
  assign y12622 = ~1'b0 ;
  assign y12623 = n26010 ;
  assign y12624 = ~n26013 ;
  assign y12625 = ~n26016 ;
  assign y12626 = n26017 ;
  assign y12627 = ~n26019 ;
  assign y12628 = ~1'b0 ;
  assign y12629 = n26020 ;
  assign y12630 = ~1'b0 ;
  assign y12631 = ~n26021 ;
  assign y12632 = ~1'b0 ;
  assign y12633 = n26022 ;
  assign y12634 = ~n26024 ;
  assign y12635 = ~n26025 ;
  assign y12636 = n26028 ;
  assign y12637 = ~n26029 ;
  assign y12638 = ~n26031 ;
  assign y12639 = ~n20573 ;
  assign y12640 = ~1'b0 ;
  assign y12641 = n26033 ;
  assign y12642 = n26034 ;
  assign y12643 = ~1'b0 ;
  assign y12644 = ~n26035 ;
  assign y12645 = n2067 ;
  assign y12646 = ~n26038 ;
  assign y12647 = ~n17421 ;
  assign y12648 = n26040 ;
  assign y12649 = ~n26044 ;
  assign y12650 = n26049 ;
  assign y12651 = ~1'b0 ;
  assign y12652 = n26051 ;
  assign y12653 = n8261 ;
  assign y12654 = ~1'b0 ;
  assign y12655 = ~n26055 ;
  assign y12656 = ~n26057 ;
  assign y12657 = n26059 ;
  assign y12658 = ~1'b0 ;
  assign y12659 = n26061 ;
  assign y12660 = ~1'b0 ;
  assign y12661 = n26067 ;
  assign y12662 = 1'b0 ;
  assign y12663 = n26069 ;
  assign y12664 = ~1'b0 ;
  assign y12665 = ~1'b0 ;
  assign y12666 = n26070 ;
  assign y12667 = n24162 ;
  assign y12668 = n15260 ;
  assign y12669 = ~1'b0 ;
  assign y12670 = ~n26071 ;
  assign y12671 = n26072 ;
  assign y12672 = ~1'b0 ;
  assign y12673 = ~1'b0 ;
  assign y12674 = 1'b0 ;
  assign y12675 = n26078 ;
  assign y12676 = ~1'b0 ;
  assign y12677 = ~n26080 ;
  assign y12678 = ~n26083 ;
  assign y12679 = 1'b0 ;
  assign y12680 = ~n26087 ;
  assign y12681 = ~1'b0 ;
  assign y12682 = ~n26092 ;
  assign y12683 = n26093 ;
  assign y12684 = n26096 ;
  assign y12685 = n26102 ;
  assign y12686 = n26104 ;
  assign y12687 = ~1'b0 ;
  assign y12688 = ~n26106 ;
  assign y12689 = n26107 ;
  assign y12690 = n26109 ;
  assign y12691 = ~n26110 ;
  assign y12692 = n26112 ;
  assign y12693 = ~1'b0 ;
  assign y12694 = ~1'b0 ;
  assign y12695 = n26118 ;
  assign y12696 = ~1'b0 ;
  assign y12697 = ~1'b0 ;
  assign y12698 = n26119 ;
  assign y12699 = n21570 ;
  assign y12700 = ~n26122 ;
  assign y12701 = n26123 ;
  assign y12702 = 1'b0 ;
  assign y12703 = ~n5980 ;
  assign y12704 = n26125 ;
  assign y12705 = n26128 ;
  assign y12706 = ~n18628 ;
  assign y12707 = ~1'b0 ;
  assign y12708 = n26130 ;
  assign y12709 = ~n26131 ;
  assign y12710 = ~n26132 ;
  assign y12711 = ~1'b0 ;
  assign y12712 = ~1'b0 ;
  assign y12713 = ~1'b0 ;
  assign y12714 = ~1'b0 ;
  assign y12715 = n26134 ;
  assign y12716 = n26137 ;
  assign y12717 = n26140 ;
  assign y12718 = ~n26144 ;
  assign y12719 = ~n26145 ;
  assign y12720 = n26146 ;
  assign y12721 = ~n26147 ;
  assign y12722 = n20416 ;
  assign y12723 = n26149 ;
  assign y12724 = ~1'b0 ;
  assign y12725 = ~n26157 ;
  assign y12726 = ~1'b0 ;
  assign y12727 = ~n26158 ;
  assign y12728 = ~1'b0 ;
  assign y12729 = n26159 ;
  assign y12730 = n26160 ;
  assign y12731 = n26161 ;
  assign y12732 = n26163 ;
  assign y12733 = ~1'b0 ;
  assign y12734 = n26166 ;
  assign y12735 = ~1'b0 ;
  assign y12736 = ~n26167 ;
  assign y12737 = n18413 ;
  assign y12738 = n26168 ;
  assign y12739 = n26169 ;
  assign y12740 = n26173 ;
  assign y12741 = n26176 ;
  assign y12742 = n26179 ;
  assign y12743 = ~n26180 ;
  assign y12744 = ~1'b0 ;
  assign y12745 = ~n26181 ;
  assign y12746 = n26183 ;
  assign y12747 = ~1'b0 ;
  assign y12748 = n26185 ;
  assign y12749 = ~1'b0 ;
  assign y12750 = n26186 ;
  assign y12751 = n26191 ;
  assign y12752 = n26193 ;
  assign y12753 = ~1'b0 ;
  assign y12754 = ~1'b0 ;
  assign y12755 = ~n26194 ;
  assign y12756 = n26196 ;
  assign y12757 = n26199 ;
  assign y12758 = n26201 ;
  assign y12759 = n26203 ;
  assign y12760 = n26205 ;
  assign y12761 = ~n26206 ;
  assign y12762 = ~1'b0 ;
  assign y12763 = n26208 ;
  assign y12764 = n26209 ;
  assign y12765 = 1'b0 ;
  assign y12766 = n26212 ;
  assign y12767 = ~n26217 ;
  assign y12768 = ~1'b0 ;
  assign y12769 = ~1'b0 ;
  assign y12770 = ~n26218 ;
  assign y12771 = ~n26219 ;
  assign y12772 = n26221 ;
  assign y12773 = ~n26222 ;
  assign y12774 = ~1'b0 ;
  assign y12775 = ~n26224 ;
  assign y12776 = ~n26225 ;
  assign y12777 = ~1'b0 ;
  assign y12778 = n26227 ;
  assign y12779 = ~n26229 ;
  assign y12780 = n26234 ;
  assign y12781 = ~n26235 ;
  assign y12782 = n26239 ;
  assign y12783 = ~n16677 ;
  assign y12784 = n26241 ;
  assign y12785 = ~n26244 ;
  assign y12786 = ~n26250 ;
  assign y12787 = ~n26254 ;
  assign y12788 = ~1'b0 ;
  assign y12789 = ~n26257 ;
  assign y12790 = ~1'b0 ;
  assign y12791 = n26259 ;
  assign y12792 = ~n26261 ;
  assign y12793 = n26262 ;
  assign y12794 = n26265 ;
  assign y12795 = ~1'b0 ;
  assign y12796 = ~n9765 ;
  assign y12797 = ~n26269 ;
  assign y12798 = n26271 ;
  assign y12799 = ~n26273 ;
  assign y12800 = ~n26276 ;
  assign y12801 = ~1'b0 ;
  assign y12802 = ~n26279 ;
  assign y12803 = n7182 ;
  assign y12804 = ~n26280 ;
  assign y12805 = n26283 ;
  assign y12806 = ~1'b0 ;
  assign y12807 = n2506 ;
  assign y12808 = n26285 ;
  assign y12809 = ~1'b0 ;
  assign y12810 = ~1'b0 ;
  assign y12811 = ~1'b0 ;
  assign y12812 = ~1'b0 ;
  assign y12813 = ~n26286 ;
  assign y12814 = ~n26289 ;
  assign y12815 = n26290 ;
  assign y12816 = ~n26295 ;
  assign y12817 = ~1'b0 ;
  assign y12818 = ~n26298 ;
  assign y12819 = n26300 ;
  assign y12820 = n26302 ;
  assign y12821 = ~n26304 ;
  assign y12822 = ~1'b0 ;
  assign y12823 = ~n26305 ;
  assign y12824 = n26307 ;
  assign y12825 = ~n26308 ;
  assign y12826 = n26309 ;
  assign y12827 = n26311 ;
  assign y12828 = ~1'b0 ;
  assign y12829 = n26312 ;
  assign y12830 = n26313 ;
  assign y12831 = ~1'b0 ;
  assign y12832 = n26314 ;
  assign y12833 = ~n26315 ;
  assign y12834 = ~n26317 ;
  assign y12835 = ~n26321 ;
  assign y12836 = ~n26322 ;
  assign y12837 = ~n26323 ;
  assign y12838 = ~n26327 ;
  assign y12839 = ~1'b0 ;
  assign y12840 = ~1'b0 ;
  assign y12841 = ~n26329 ;
  assign y12842 = n26331 ;
  assign y12843 = n26333 ;
  assign y12844 = n26334 ;
  assign y12845 = ~n26336 ;
  assign y12846 = ~n26338 ;
  assign y12847 = ~n26339 ;
  assign y12848 = ~n26340 ;
  assign y12849 = ~1'b0 ;
  assign y12850 = ~1'b0 ;
  assign y12851 = ~1'b0 ;
  assign y12852 = ~n26347 ;
  assign y12853 = ~1'b0 ;
  assign y12854 = n26349 ;
  assign y12855 = n26351 ;
  assign y12856 = ~n26355 ;
  assign y12857 = n26356 ;
  assign y12858 = ~n26357 ;
  assign y12859 = ~n26361 ;
  assign y12860 = ~n26364 ;
  assign y12861 = n26367 ;
  assign y12862 = ~n26369 ;
  assign y12863 = ~1'b0 ;
  assign y12864 = ~n26373 ;
  assign y12865 = ~1'b0 ;
  assign y12866 = ~n26374 ;
  assign y12867 = ~n26377 ;
  assign y12868 = n12872 ;
  assign y12869 = ~n26381 ;
  assign y12870 = ~n26382 ;
  assign y12871 = ~1'b0 ;
  assign y12872 = ~1'b0 ;
  assign y12873 = ~1'b0 ;
  assign y12874 = ~n26384 ;
  assign y12875 = ~n26388 ;
  assign y12876 = n9094 ;
  assign y12877 = n26390 ;
  assign y12878 = ~1'b0 ;
  assign y12879 = n26391 ;
  assign y12880 = n26394 ;
  assign y12881 = n26396 ;
  assign y12882 = ~1'b0 ;
  assign y12883 = ~n26398 ;
  assign y12884 = n26402 ;
  assign y12885 = ~1'b0 ;
  assign y12886 = n26403 ;
  assign y12887 = ~n26406 ;
  assign y12888 = ~1'b0 ;
  assign y12889 = ~1'b0 ;
  assign y12890 = n26407 ;
  assign y12891 = ~n26408 ;
  assign y12892 = n8919 ;
  assign y12893 = n26410 ;
  assign y12894 = ~n26411 ;
  assign y12895 = ~n26413 ;
  assign y12896 = n26415 ;
  assign y12897 = n26420 ;
  assign y12898 = ~n26423 ;
  assign y12899 = ~n26426 ;
  assign y12900 = ~1'b0 ;
  assign y12901 = ~n26430 ;
  assign y12902 = ~n26433 ;
  assign y12903 = n2154 ;
  assign y12904 = ~n26434 ;
  assign y12905 = ~n26437 ;
  assign y12906 = ~1'b0 ;
  assign y12907 = ~n26438 ;
  assign y12908 = ~1'b0 ;
  assign y12909 = n26441 ;
  assign y12910 = n26449 ;
  assign y12911 = ~1'b0 ;
  assign y12912 = ~n21507 ;
  assign y12913 = ~n26453 ;
  assign y12914 = n26454 ;
  assign y12915 = n26455 ;
  assign y12916 = ~1'b0 ;
  assign y12917 = ~1'b0 ;
  assign y12918 = ~n26457 ;
  assign y12919 = ~1'b0 ;
  assign y12920 = ~n26472 ;
  assign y12921 = ~1'b0 ;
  assign y12922 = n26473 ;
  assign y12923 = n26484 ;
  assign y12924 = ~n26486 ;
  assign y12925 = n26492 ;
  assign y12926 = ~1'b0 ;
  assign y12927 = n26494 ;
  assign y12928 = 1'b0 ;
  assign y12929 = ~n26495 ;
  assign y12930 = ~n26496 ;
  assign y12931 = ~n26499 ;
  assign y12932 = ~n26500 ;
  assign y12933 = n26501 ;
  assign y12934 = n26502 ;
  assign y12935 = ~n26506 ;
  assign y12936 = n26509 ;
  assign y12937 = ~n26511 ;
  assign y12938 = ~1'b0 ;
  assign y12939 = ~n26516 ;
  assign y12940 = ~1'b0 ;
  assign y12941 = n4097 ;
  assign y12942 = ~1'b0 ;
  assign y12943 = n26521 ;
  assign y12944 = n26526 ;
  assign y12945 = ~n26527 ;
  assign y12946 = ~n26530 ;
  assign y12947 = 1'b0 ;
  assign y12948 = n26532 ;
  assign y12949 = n26533 ;
  assign y12950 = n26535 ;
  assign y12951 = n26537 ;
  assign y12952 = n26540 ;
  assign y12953 = 1'b0 ;
  assign y12954 = ~1'b0 ;
  assign y12955 = n26543 ;
  assign y12956 = n26544 ;
  assign y12957 = ~n26548 ;
  assign y12958 = n26550 ;
  assign y12959 = ~1'b0 ;
  assign y12960 = ~1'b0 ;
  assign y12961 = ~1'b0 ;
  assign y12962 = ~1'b0 ;
  assign y12963 = n26553 ;
  assign y12964 = ~1'b0 ;
  assign y12965 = n26557 ;
  assign y12966 = n26558 ;
  assign y12967 = n26559 ;
  assign y12968 = n26561 ;
  assign y12969 = ~1'b0 ;
  assign y12970 = n26562 ;
  assign y12971 = n26563 ;
  assign y12972 = ~1'b0 ;
  assign y12973 = n26566 ;
  assign y12974 = n26567 ;
  assign y12975 = ~n26568 ;
  assign y12976 = n26573 ;
  assign y12977 = n26579 ;
  assign y12978 = n26588 ;
  assign y12979 = ~n26590 ;
  assign y12980 = ~1'b0 ;
  assign y12981 = ~n26592 ;
  assign y12982 = n23677 ;
  assign y12983 = ~n8745 ;
  assign y12984 = n26593 ;
  assign y12985 = n956 ;
  assign y12986 = ~n9228 ;
  assign y12987 = ~n26598 ;
  assign y12988 = ~n3556 ;
  assign y12989 = ~n26600 ;
  assign y12990 = n26602 ;
  assign y12991 = ~n26604 ;
  assign y12992 = ~1'b0 ;
  assign y12993 = n26606 ;
  assign y12994 = 1'b0 ;
  assign y12995 = ~1'b0 ;
  assign y12996 = ~1'b0 ;
  assign y12997 = ~1'b0 ;
  assign y12998 = ~n26607 ;
  assign y12999 = ~n26612 ;
  assign y13000 = n26613 ;
  assign y13001 = n26614 ;
  assign y13002 = ~n26616 ;
  assign y13003 = n26619 ;
  assign y13004 = n26623 ;
  assign y13005 = n26624 ;
  assign y13006 = n26625 ;
  assign y13007 = 1'b0 ;
  assign y13008 = 1'b0 ;
  assign y13009 = ~n26630 ;
  assign y13010 = ~n26632 ;
  assign y13011 = ~n26636 ;
  assign y13012 = ~n14889 ;
  assign y13013 = n20375 ;
  assign y13014 = n26637 ;
  assign y13015 = ~n4264 ;
  assign y13016 = ~n26638 ;
  assign y13017 = ~n26639 ;
  assign y13018 = n26641 ;
  assign y13019 = n26642 ;
  assign y13020 = ~n17607 ;
  assign y13021 = ~n6076 ;
  assign y13022 = ~n26646 ;
  assign y13023 = n26652 ;
  assign y13024 = ~1'b0 ;
  assign y13025 = ~1'b0 ;
  assign y13026 = ~n26654 ;
  assign y13027 = ~1'b0 ;
  assign y13028 = ~n26655 ;
  assign y13029 = n26656 ;
  assign y13030 = ~1'b0 ;
  assign y13031 = ~n7934 ;
  assign y13032 = n11854 ;
  assign y13033 = n26657 ;
  assign y13034 = ~n26663 ;
  assign y13035 = ~1'b0 ;
  assign y13036 = ~1'b0 ;
  assign y13037 = n26666 ;
  assign y13038 = n26668 ;
  assign y13039 = ~n26670 ;
  assign y13040 = ~1'b0 ;
  assign y13041 = n26675 ;
  assign y13042 = n25936 ;
  assign y13043 = n26679 ;
  assign y13044 = ~n26682 ;
  assign y13045 = n26683 ;
  assign y13046 = ~1'b0 ;
  assign y13047 = ~1'b0 ;
  assign y13048 = ~1'b0 ;
  assign y13049 = ~1'b0 ;
  assign y13050 = n19720 ;
  assign y13051 = n26684 ;
  assign y13052 = ~n26687 ;
  assign y13053 = ~n26691 ;
  assign y13054 = ~n26694 ;
  assign y13055 = n26695 ;
  assign y13056 = n26696 ;
  assign y13057 = ~1'b0 ;
  assign y13058 = n26706 ;
  assign y13059 = n26707 ;
  assign y13060 = ~n26710 ;
  assign y13061 = n26715 ;
  assign y13062 = n26719 ;
  assign y13063 = ~1'b0 ;
  assign y13064 = n26720 ;
  assign y13065 = n26721 ;
  assign y13066 = n26722 ;
  assign y13067 = n26723 ;
  assign y13068 = n26725 ;
  assign y13069 = n6212 ;
  assign y13070 = n26727 ;
  assign y13071 = ~n26731 ;
  assign y13072 = ~1'b0 ;
  assign y13073 = 1'b0 ;
  assign y13074 = n26740 ;
  assign y13075 = ~n26742 ;
  assign y13076 = n26743 ;
  assign y13077 = ~1'b0 ;
  assign y13078 = ~1'b0 ;
  assign y13079 = ~1'b0 ;
  assign y13080 = ~1'b0 ;
  assign y13081 = ~n26744 ;
  assign y13082 = ~n26748 ;
  assign y13083 = ~1'b0 ;
  assign y13084 = ~n26749 ;
  assign y13085 = ~n26751 ;
  assign y13086 = ~n26752 ;
  assign y13087 = ~n26755 ;
  assign y13088 = ~1'b0 ;
  assign y13089 = ~n26757 ;
  assign y13090 = ~1'b0 ;
  assign y13091 = n26760 ;
  assign y13092 = n26763 ;
  assign y13093 = ~1'b0 ;
  assign y13094 = n26764 ;
  assign y13095 = ~1'b0 ;
  assign y13096 = n26771 ;
  assign y13097 = 1'b0 ;
  assign y13098 = n26772 ;
  assign y13099 = ~n26774 ;
  assign y13100 = ~n26776 ;
  assign y13101 = ~n26780 ;
  assign y13102 = n26781 ;
  assign y13103 = ~n25248 ;
  assign y13104 = n26783 ;
  assign y13105 = ~n26787 ;
  assign y13106 = ~1'b0 ;
  assign y13107 = ~n26788 ;
  assign y13108 = ~n26791 ;
  assign y13109 = ~n26792 ;
  assign y13110 = ~n26796 ;
  assign y13111 = ~1'b0 ;
  assign y13112 = ~n26801 ;
  assign y13113 = ~1'b0 ;
  assign y13114 = n26803 ;
  assign y13115 = ~n26805 ;
  assign y13116 = 1'b0 ;
  assign y13117 = ~1'b0 ;
  assign y13118 = n26809 ;
  assign y13119 = n26812 ;
  assign y13120 = ~n26813 ;
  assign y13121 = ~n26817 ;
  assign y13122 = n26819 ;
  assign y13123 = n26827 ;
  assign y13124 = n26829 ;
  assign y13125 = ~n26830 ;
  assign y13126 = n26832 ;
  assign y13127 = 1'b0 ;
  assign y13128 = ~n26834 ;
endmodule
