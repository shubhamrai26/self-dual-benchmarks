module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24448 , n24449 , n24450 ;
  assign n257 = x1 & ~x129 ;
  assign n258 = ~x2 & ~n257 ;
  assign n259 = ~x130 & ~x131 ;
  assign n260 = ~n258 & n259 ;
  assign n261 = x3 & ~x131 ;
  assign n262 = ~x4 & ~n261 ;
  assign n263 = ~x5 & n262 ;
  assign n264 = ~n260 & n263 ;
  assign n265 = ~x5 & x132 ;
  assign n266 = ~x133 & ~x134 ;
  assign n267 = ~n265 & n266 ;
  assign n268 = ~n264 & n267 ;
  assign n269 = x6 & ~x134 ;
  assign n270 = ~x7 & ~n269 ;
  assign n271 = ~x8 & n270 ;
  assign n272 = ~n268 & n271 ;
  assign n273 = ~x8 & x135 ;
  assign n274 = ~x136 & ~x137 ;
  assign n275 = ~n273 & n274 ;
  assign n276 = ~n272 & n275 ;
  assign n277 = x9 & ~x137 ;
  assign n278 = ~x10 & ~n277 ;
  assign n279 = ~x11 & n278 ;
  assign n280 = ~n276 & n279 ;
  assign n281 = ~x11 & x138 ;
  assign n282 = ~x139 & ~x140 ;
  assign n283 = ~n281 & n282 ;
  assign n284 = ~n280 & n283 ;
  assign n285 = x12 & ~x140 ;
  assign n286 = ~x13 & ~n285 ;
  assign n287 = ~x14 & n286 ;
  assign n288 = ~n284 & n287 ;
  assign n289 = ~x14 & x141 ;
  assign n290 = ~x142 & ~x143 ;
  assign n291 = ~n289 & n290 ;
  assign n292 = ~n288 & n291 ;
  assign n293 = x15 & ~x143 ;
  assign n294 = ~x16 & ~n293 ;
  assign n295 = ~x17 & n294 ;
  assign n296 = ~n292 & n295 ;
  assign n297 = ~x17 & x144 ;
  assign n298 = ~x145 & ~x146 ;
  assign n299 = ~n297 & n298 ;
  assign n300 = ~n296 & n299 ;
  assign n301 = x18 & ~x146 ;
  assign n302 = ~x19 & ~n301 ;
  assign n303 = ~x20 & n302 ;
  assign n304 = ~n300 & n303 ;
  assign n305 = ~x20 & x147 ;
  assign n306 = ~x148 & ~x149 ;
  assign n307 = ~n305 & n306 ;
  assign n308 = ~n304 & n307 ;
  assign n309 = x21 & ~x149 ;
  assign n310 = ~x22 & ~n309 ;
  assign n311 = ~x23 & n310 ;
  assign n312 = ~n308 & n311 ;
  assign n313 = ~x23 & x150 ;
  assign n314 = ~x151 & ~x152 ;
  assign n315 = ~n313 & n314 ;
  assign n316 = ~n312 & n315 ;
  assign n317 = x24 & ~x152 ;
  assign n318 = ~x25 & ~n317 ;
  assign n319 = ~x26 & n318 ;
  assign n320 = ~n316 & n319 ;
  assign n321 = ~x26 & x153 ;
  assign n322 = ~x154 & ~x155 ;
  assign n323 = ~n321 & n322 ;
  assign n324 = ~n320 & n323 ;
  assign n325 = x27 & ~x155 ;
  assign n326 = ~x28 & ~n325 ;
  assign n327 = ~x29 & n326 ;
  assign n328 = ~n324 & n327 ;
  assign n329 = ~x29 & x156 ;
  assign n330 = ~x157 & ~x158 ;
  assign n331 = ~n329 & n330 ;
  assign n332 = ~n328 & n331 ;
  assign n333 = x30 & ~x158 ;
  assign n334 = ~x31 & ~n333 ;
  assign n335 = ~x32 & n334 ;
  assign n336 = ~n332 & n335 ;
  assign n337 = ~x32 & x159 ;
  assign n338 = ~x160 & ~x161 ;
  assign n339 = ~n337 & n338 ;
  assign n340 = ~n336 & n339 ;
  assign n341 = x33 & ~x161 ;
  assign n342 = ~x34 & ~n341 ;
  assign n343 = ~x35 & n342 ;
  assign n344 = ~n340 & n343 ;
  assign n345 = ~x35 & x162 ;
  assign n346 = ~x163 & ~x164 ;
  assign n347 = ~n345 & n346 ;
  assign n348 = ~n344 & n347 ;
  assign n349 = x36 & ~x164 ;
  assign n350 = ~x37 & ~n349 ;
  assign n351 = ~x38 & n350 ;
  assign n352 = ~n348 & n351 ;
  assign n353 = ~x38 & x165 ;
  assign n354 = ~x166 & ~x167 ;
  assign n355 = ~n353 & n354 ;
  assign n356 = ~n352 & n355 ;
  assign n357 = x39 & ~x167 ;
  assign n358 = ~x40 & ~n357 ;
  assign n359 = ~x41 & n358 ;
  assign n360 = ~n356 & n359 ;
  assign n361 = ~x41 & x168 ;
  assign n362 = ~x169 & ~x170 ;
  assign n363 = ~n361 & n362 ;
  assign n364 = ~n360 & n363 ;
  assign n365 = x42 & ~x170 ;
  assign n366 = ~x43 & ~n365 ;
  assign n367 = ~x44 & n366 ;
  assign n368 = ~n364 & n367 ;
  assign n369 = ~x44 & x171 ;
  assign n370 = ~x172 & ~x173 ;
  assign n371 = ~n369 & n370 ;
  assign n372 = ~n368 & n371 ;
  assign n373 = x45 & ~x173 ;
  assign n374 = ~x46 & ~n373 ;
  assign n375 = ~x47 & n374 ;
  assign n376 = ~n372 & n375 ;
  assign n377 = ~x47 & x174 ;
  assign n378 = ~x175 & ~x176 ;
  assign n379 = ~n377 & n378 ;
  assign n380 = ~n376 & n379 ;
  assign n381 = x48 & ~x176 ;
  assign n382 = ~x49 & ~n381 ;
  assign n383 = ~x50 & n382 ;
  assign n384 = ~n380 & n383 ;
  assign n385 = ~x50 & x177 ;
  assign n386 = ~x178 & ~x179 ;
  assign n387 = ~n385 & n386 ;
  assign n388 = ~n384 & n387 ;
  assign n389 = x51 & ~x179 ;
  assign n390 = ~x52 & ~n389 ;
  assign n391 = ~x53 & n390 ;
  assign n392 = ~n388 & n391 ;
  assign n393 = ~x53 & x180 ;
  assign n394 = ~x181 & ~x182 ;
  assign n395 = ~n393 & n394 ;
  assign n396 = ~n392 & n395 ;
  assign n397 = x54 & ~x182 ;
  assign n398 = ~x55 & ~n397 ;
  assign n399 = ~x56 & n398 ;
  assign n400 = ~n396 & n399 ;
  assign n401 = ~x56 & x183 ;
  assign n402 = ~x184 & ~x185 ;
  assign n403 = ~n401 & n402 ;
  assign n404 = ~n400 & n403 ;
  assign n405 = x57 & ~x185 ;
  assign n406 = ~x58 & ~n405 ;
  assign n407 = ~x59 & n406 ;
  assign n408 = ~n404 & n407 ;
  assign n409 = ~x59 & x186 ;
  assign n410 = ~x187 & ~x188 ;
  assign n411 = ~n409 & n410 ;
  assign n412 = ~n408 & n411 ;
  assign n413 = x60 & ~x188 ;
  assign n414 = ~x61 & ~n413 ;
  assign n415 = ~x62 & n414 ;
  assign n416 = ~n412 & n415 ;
  assign n417 = ~x62 & x189 ;
  assign n418 = ~x190 & ~x191 ;
  assign n419 = ~n417 & n418 ;
  assign n420 = ~n416 & n419 ;
  assign n421 = x63 & ~x191 ;
  assign n422 = ~x64 & ~n421 ;
  assign n423 = ~x65 & n422 ;
  assign n424 = ~n420 & n423 ;
  assign n425 = ~x65 & x192 ;
  assign n426 = ~x193 & ~x194 ;
  assign n427 = ~n425 & n426 ;
  assign n428 = ~n424 & n427 ;
  assign n429 = x66 & ~x194 ;
  assign n430 = ~x67 & ~n429 ;
  assign n431 = ~x68 & n430 ;
  assign n432 = ~n428 & n431 ;
  assign n433 = ~x68 & x195 ;
  assign n434 = ~x196 & ~x197 ;
  assign n435 = ~n433 & n434 ;
  assign n436 = ~n432 & n435 ;
  assign n437 = x69 & ~x197 ;
  assign n438 = ~x70 & ~n437 ;
  assign n439 = ~x71 & n438 ;
  assign n440 = ~n436 & n439 ;
  assign n441 = ~x71 & x198 ;
  assign n442 = ~x199 & ~x200 ;
  assign n443 = ~n441 & n442 ;
  assign n444 = ~n440 & n443 ;
  assign n445 = x72 & ~x200 ;
  assign n446 = ~x73 & ~n445 ;
  assign n447 = ~x74 & n446 ;
  assign n448 = ~n444 & n447 ;
  assign n449 = ~x74 & x201 ;
  assign n450 = ~x202 & ~x203 ;
  assign n451 = ~n449 & n450 ;
  assign n452 = ~n448 & n451 ;
  assign n453 = x75 & ~x203 ;
  assign n454 = ~x76 & ~n453 ;
  assign n455 = ~x77 & n454 ;
  assign n456 = ~n452 & n455 ;
  assign n457 = ~x77 & x204 ;
  assign n458 = ~x205 & ~x206 ;
  assign n459 = ~n457 & n458 ;
  assign n460 = ~n456 & n459 ;
  assign n461 = x78 & ~x206 ;
  assign n462 = ~x79 & ~n461 ;
  assign n463 = ~x80 & n462 ;
  assign n464 = ~n460 & n463 ;
  assign n465 = ~x80 & x207 ;
  assign n466 = ~x208 & ~x209 ;
  assign n467 = ~n465 & n466 ;
  assign n468 = ~n464 & n467 ;
  assign n469 = x81 & ~x209 ;
  assign n470 = ~x82 & ~n469 ;
  assign n471 = ~x83 & n470 ;
  assign n472 = ~n468 & n471 ;
  assign n473 = ~x83 & x210 ;
  assign n474 = ~x211 & ~x212 ;
  assign n475 = ~n473 & n474 ;
  assign n476 = ~n472 & n475 ;
  assign n477 = x84 & ~x212 ;
  assign n478 = ~x85 & ~n477 ;
  assign n479 = ~x86 & n478 ;
  assign n480 = ~n476 & n479 ;
  assign n481 = ~x86 & x213 ;
  assign n482 = ~x214 & ~x215 ;
  assign n483 = ~n481 & n482 ;
  assign n484 = ~n480 & n483 ;
  assign n485 = x87 & ~x215 ;
  assign n486 = ~x88 & ~n485 ;
  assign n487 = ~x89 & n486 ;
  assign n488 = ~n484 & n487 ;
  assign n489 = ~x89 & x216 ;
  assign n490 = ~x217 & ~x218 ;
  assign n491 = ~n489 & n490 ;
  assign n492 = ~n488 & n491 ;
  assign n493 = x90 & ~x218 ;
  assign n494 = ~x91 & ~n493 ;
  assign n495 = ~x92 & n494 ;
  assign n496 = ~n492 & n495 ;
  assign n497 = ~x92 & x219 ;
  assign n498 = ~x220 & ~x221 ;
  assign n499 = ~n497 & n498 ;
  assign n500 = ~n496 & n499 ;
  assign n501 = x93 & ~x221 ;
  assign n502 = ~x94 & ~n501 ;
  assign n503 = ~x95 & n502 ;
  assign n504 = ~n500 & n503 ;
  assign n505 = ~x95 & x222 ;
  assign n506 = ~x223 & ~x224 ;
  assign n507 = ~n505 & n506 ;
  assign n508 = ~n504 & n507 ;
  assign n509 = x96 & ~x224 ;
  assign n510 = ~x97 & ~n509 ;
  assign n511 = ~x98 & n510 ;
  assign n512 = ~n508 & n511 ;
  assign n513 = ~x98 & x225 ;
  assign n514 = ~x226 & ~x227 ;
  assign n515 = ~n513 & n514 ;
  assign n516 = ~n512 & n515 ;
  assign n517 = x99 & ~x227 ;
  assign n518 = ~x100 & ~n517 ;
  assign n519 = ~x101 & n518 ;
  assign n520 = ~n516 & n519 ;
  assign n521 = ~x101 & x228 ;
  assign n522 = ~x229 & ~x230 ;
  assign n523 = ~n521 & n522 ;
  assign n524 = ~n520 & n523 ;
  assign n525 = x102 & ~x230 ;
  assign n526 = ~x103 & ~n525 ;
  assign n527 = ~x104 & n526 ;
  assign n528 = ~n524 & n527 ;
  assign n529 = ~x104 & x231 ;
  assign n530 = ~x232 & ~x233 ;
  assign n531 = ~n529 & n530 ;
  assign n532 = ~n528 & n531 ;
  assign n533 = x105 & ~x233 ;
  assign n534 = ~x106 & ~n533 ;
  assign n535 = ~x107 & n534 ;
  assign n536 = ~n532 & n535 ;
  assign n537 = ~x107 & x234 ;
  assign n538 = ~x235 & ~x236 ;
  assign n539 = ~n537 & n538 ;
  assign n540 = ~n536 & n539 ;
  assign n541 = x108 & ~x236 ;
  assign n542 = ~x109 & ~n541 ;
  assign n543 = ~x110 & n542 ;
  assign n544 = ~n540 & n543 ;
  assign n545 = ~x110 & x237 ;
  assign n546 = ~x238 & ~x239 ;
  assign n547 = ~n545 & n546 ;
  assign n548 = ~n544 & n547 ;
  assign n549 = x111 & ~x239 ;
  assign n550 = ~x112 & ~n549 ;
  assign n551 = ~x113 & n550 ;
  assign n552 = ~n548 & n551 ;
  assign n553 = ~x113 & x240 ;
  assign n554 = ~x241 & ~x242 ;
  assign n555 = ~n553 & n554 ;
  assign n556 = ~n552 & n555 ;
  assign n557 = x114 & ~x242 ;
  assign n558 = ~x115 & ~n557 ;
  assign n559 = ~x116 & n558 ;
  assign n560 = ~n556 & n559 ;
  assign n561 = ~x116 & x243 ;
  assign n562 = ~x244 & ~x245 ;
  assign n563 = ~n561 & n562 ;
  assign n564 = ~n560 & n563 ;
  assign n565 = x117 & ~x245 ;
  assign n566 = ~x118 & ~n565 ;
  assign n567 = ~x119 & n566 ;
  assign n568 = ~n564 & n567 ;
  assign n569 = ~x119 & x246 ;
  assign n570 = ~x247 & ~x248 ;
  assign n571 = ~n569 & n570 ;
  assign n572 = ~n568 & n571 ;
  assign n573 = x120 & ~x248 ;
  assign n574 = ~x121 & ~n573 ;
  assign n575 = ~x122 & n574 ;
  assign n576 = ~n572 & n575 ;
  assign n577 = ~x122 & x249 ;
  assign n578 = ~x250 & ~x251 ;
  assign n579 = ~n577 & n578 ;
  assign n580 = ~n576 & n579 ;
  assign n581 = x123 & ~x251 ;
  assign n582 = ~x124 & ~n581 ;
  assign n583 = ~x125 & n582 ;
  assign n584 = ~n580 & n583 ;
  assign n585 = ~x125 & x252 ;
  assign n586 = ~x253 & ~x254 ;
  assign n587 = ~n585 & n586 ;
  assign n588 = ~n584 & n587 ;
  assign n589 = x126 & ~x254 ;
  assign n590 = ~x127 & ~n589 ;
  assign n591 = ~x0 & n590 ;
  assign n592 = ~n588 & n591 ;
  assign n593 = ~x0 & x255 ;
  assign n594 = x128 & ~n593 ;
  assign n595 = ~n592 & n594 ;
  assign n936 = n595 & x256 ;
  assign n596 = ~x1 & x129 ;
  assign n597 = x2 & ~n596 ;
  assign n598 = x130 & x131 ;
  assign n599 = ~n597 & n598 ;
  assign n600 = ~x3 & x131 ;
  assign n601 = x4 & ~n600 ;
  assign n602 = x5 & n601 ;
  assign n603 = ~n599 & n602 ;
  assign n604 = x5 & ~x132 ;
  assign n605 = x133 & x134 ;
  assign n606 = ~n604 & n605 ;
  assign n607 = ~n603 & n606 ;
  assign n608 = ~x6 & x134 ;
  assign n609 = x7 & ~n608 ;
  assign n610 = x8 & n609 ;
  assign n611 = ~n607 & n610 ;
  assign n612 = x8 & ~x135 ;
  assign n613 = x136 & x137 ;
  assign n614 = ~n612 & n613 ;
  assign n615 = ~n611 & n614 ;
  assign n616 = ~x9 & x137 ;
  assign n617 = x10 & ~n616 ;
  assign n618 = x11 & n617 ;
  assign n619 = ~n615 & n618 ;
  assign n620 = x11 & ~x138 ;
  assign n621 = x139 & x140 ;
  assign n622 = ~n620 & n621 ;
  assign n623 = ~n619 & n622 ;
  assign n624 = ~x12 & x140 ;
  assign n625 = x13 & ~n624 ;
  assign n626 = x14 & n625 ;
  assign n627 = ~n623 & n626 ;
  assign n628 = x14 & ~x141 ;
  assign n629 = x142 & x143 ;
  assign n630 = ~n628 & n629 ;
  assign n631 = ~n627 & n630 ;
  assign n632 = ~x15 & x143 ;
  assign n633 = x16 & ~n632 ;
  assign n634 = x17 & n633 ;
  assign n635 = ~n631 & n634 ;
  assign n636 = x17 & ~x144 ;
  assign n637 = x145 & x146 ;
  assign n638 = ~n636 & n637 ;
  assign n639 = ~n635 & n638 ;
  assign n640 = ~x18 & x146 ;
  assign n641 = x19 & ~n640 ;
  assign n642 = x20 & n641 ;
  assign n643 = ~n639 & n642 ;
  assign n644 = x20 & ~x147 ;
  assign n645 = x148 & x149 ;
  assign n646 = ~n644 & n645 ;
  assign n647 = ~n643 & n646 ;
  assign n648 = ~x21 & x149 ;
  assign n649 = x22 & ~n648 ;
  assign n650 = x23 & n649 ;
  assign n651 = ~n647 & n650 ;
  assign n652 = x23 & ~x150 ;
  assign n653 = x151 & x152 ;
  assign n654 = ~n652 & n653 ;
  assign n655 = ~n651 & n654 ;
  assign n656 = ~x24 & x152 ;
  assign n657 = x25 & ~n656 ;
  assign n658 = x26 & n657 ;
  assign n659 = ~n655 & n658 ;
  assign n660 = x26 & ~x153 ;
  assign n661 = x154 & x155 ;
  assign n662 = ~n660 & n661 ;
  assign n663 = ~n659 & n662 ;
  assign n664 = ~x27 & x155 ;
  assign n665 = x28 & ~n664 ;
  assign n666 = x29 & n665 ;
  assign n667 = ~n663 & n666 ;
  assign n668 = x29 & ~x156 ;
  assign n669 = x157 & x158 ;
  assign n670 = ~n668 & n669 ;
  assign n671 = ~n667 & n670 ;
  assign n672 = ~x30 & x158 ;
  assign n673 = x31 & ~n672 ;
  assign n674 = x32 & n673 ;
  assign n675 = ~n671 & n674 ;
  assign n676 = x32 & ~x159 ;
  assign n677 = x160 & x161 ;
  assign n678 = ~n676 & n677 ;
  assign n679 = ~n675 & n678 ;
  assign n680 = ~x33 & x161 ;
  assign n681 = x34 & ~n680 ;
  assign n682 = x35 & n681 ;
  assign n683 = ~n679 & n682 ;
  assign n684 = x35 & ~x162 ;
  assign n685 = x163 & x164 ;
  assign n686 = ~n684 & n685 ;
  assign n687 = ~n683 & n686 ;
  assign n688 = ~x36 & x164 ;
  assign n689 = x37 & ~n688 ;
  assign n690 = x38 & n689 ;
  assign n691 = ~n687 & n690 ;
  assign n692 = x38 & ~x165 ;
  assign n693 = x166 & x167 ;
  assign n694 = ~n692 & n693 ;
  assign n695 = ~n691 & n694 ;
  assign n696 = ~x39 & x167 ;
  assign n697 = x40 & ~n696 ;
  assign n698 = x41 & n697 ;
  assign n699 = ~n695 & n698 ;
  assign n700 = x41 & ~x168 ;
  assign n701 = x169 & x170 ;
  assign n702 = ~n700 & n701 ;
  assign n703 = ~n699 & n702 ;
  assign n704 = ~x42 & x170 ;
  assign n705 = x43 & ~n704 ;
  assign n706 = x44 & n705 ;
  assign n707 = ~n703 & n706 ;
  assign n708 = x44 & ~x171 ;
  assign n709 = x172 & x173 ;
  assign n710 = ~n708 & n709 ;
  assign n711 = ~n707 & n710 ;
  assign n712 = ~x45 & x173 ;
  assign n713 = x46 & ~n712 ;
  assign n714 = x47 & n713 ;
  assign n715 = ~n711 & n714 ;
  assign n716 = x47 & ~x174 ;
  assign n717 = x175 & x176 ;
  assign n718 = ~n716 & n717 ;
  assign n719 = ~n715 & n718 ;
  assign n720 = ~x48 & x176 ;
  assign n721 = x49 & ~n720 ;
  assign n722 = x50 & n721 ;
  assign n723 = ~n719 & n722 ;
  assign n724 = x50 & ~x177 ;
  assign n725 = x178 & x179 ;
  assign n726 = ~n724 & n725 ;
  assign n727 = ~n723 & n726 ;
  assign n728 = ~x51 & x179 ;
  assign n729 = x52 & ~n728 ;
  assign n730 = x53 & n729 ;
  assign n731 = ~n727 & n730 ;
  assign n732 = x53 & ~x180 ;
  assign n733 = x181 & x182 ;
  assign n734 = ~n732 & n733 ;
  assign n735 = ~n731 & n734 ;
  assign n736 = ~x54 & x182 ;
  assign n737 = x55 & ~n736 ;
  assign n738 = x56 & n737 ;
  assign n739 = ~n735 & n738 ;
  assign n740 = x56 & ~x183 ;
  assign n741 = x184 & x185 ;
  assign n742 = ~n740 & n741 ;
  assign n743 = ~n739 & n742 ;
  assign n744 = ~x57 & x185 ;
  assign n745 = x58 & ~n744 ;
  assign n746 = x59 & n745 ;
  assign n747 = ~n743 & n746 ;
  assign n748 = x59 & ~x186 ;
  assign n749 = x187 & x188 ;
  assign n750 = ~n748 & n749 ;
  assign n751 = ~n747 & n750 ;
  assign n752 = ~x60 & x188 ;
  assign n753 = x61 & ~n752 ;
  assign n754 = x62 & n753 ;
  assign n755 = ~n751 & n754 ;
  assign n756 = x62 & ~x189 ;
  assign n757 = x190 & x191 ;
  assign n758 = ~n756 & n757 ;
  assign n759 = ~n755 & n758 ;
  assign n760 = ~x63 & x191 ;
  assign n761 = x64 & ~n760 ;
  assign n762 = x65 & n761 ;
  assign n763 = ~n759 & n762 ;
  assign n764 = x65 & ~x192 ;
  assign n765 = x193 & x194 ;
  assign n766 = ~n764 & n765 ;
  assign n767 = ~n763 & n766 ;
  assign n768 = ~x66 & x194 ;
  assign n769 = x67 & ~n768 ;
  assign n770 = x68 & n769 ;
  assign n771 = ~n767 & n770 ;
  assign n772 = x68 & ~x195 ;
  assign n773 = x196 & x197 ;
  assign n774 = ~n772 & n773 ;
  assign n775 = ~n771 & n774 ;
  assign n776 = ~x69 & x197 ;
  assign n777 = x70 & ~n776 ;
  assign n778 = x71 & n777 ;
  assign n779 = ~n775 & n778 ;
  assign n780 = x71 & ~x198 ;
  assign n781 = x199 & x200 ;
  assign n782 = ~n780 & n781 ;
  assign n783 = ~n779 & n782 ;
  assign n784 = ~x72 & x200 ;
  assign n785 = x73 & ~n784 ;
  assign n786 = x74 & n785 ;
  assign n787 = ~n783 & n786 ;
  assign n788 = x74 & ~x201 ;
  assign n789 = x202 & x203 ;
  assign n790 = ~n788 & n789 ;
  assign n791 = ~n787 & n790 ;
  assign n792 = ~x75 & x203 ;
  assign n793 = x76 & ~n792 ;
  assign n794 = x77 & n793 ;
  assign n795 = ~n791 & n794 ;
  assign n796 = x77 & ~x204 ;
  assign n797 = x205 & x206 ;
  assign n798 = ~n796 & n797 ;
  assign n799 = ~n795 & n798 ;
  assign n800 = ~x78 & x206 ;
  assign n801 = x79 & ~n800 ;
  assign n802 = x80 & n801 ;
  assign n803 = ~n799 & n802 ;
  assign n804 = x80 & ~x207 ;
  assign n805 = x208 & x209 ;
  assign n806 = ~n804 & n805 ;
  assign n807 = ~n803 & n806 ;
  assign n808 = ~x81 & x209 ;
  assign n809 = x82 & ~n808 ;
  assign n810 = x83 & n809 ;
  assign n811 = ~n807 & n810 ;
  assign n812 = x83 & ~x210 ;
  assign n813 = x211 & x212 ;
  assign n814 = ~n812 & n813 ;
  assign n815 = ~n811 & n814 ;
  assign n816 = ~x84 & x212 ;
  assign n817 = x85 & ~n816 ;
  assign n818 = x86 & n817 ;
  assign n819 = ~n815 & n818 ;
  assign n820 = x86 & ~x213 ;
  assign n821 = x214 & x215 ;
  assign n822 = ~n820 & n821 ;
  assign n823 = ~n819 & n822 ;
  assign n824 = ~x87 & x215 ;
  assign n825 = x88 & ~n824 ;
  assign n826 = x89 & n825 ;
  assign n827 = ~n823 & n826 ;
  assign n828 = x89 & ~x216 ;
  assign n829 = x217 & x218 ;
  assign n830 = ~n828 & n829 ;
  assign n831 = ~n827 & n830 ;
  assign n832 = ~x90 & x218 ;
  assign n833 = x91 & ~n832 ;
  assign n834 = x92 & n833 ;
  assign n835 = ~n831 & n834 ;
  assign n836 = x92 & ~x219 ;
  assign n837 = x220 & x221 ;
  assign n838 = ~n836 & n837 ;
  assign n839 = ~n835 & n838 ;
  assign n840 = ~x93 & x221 ;
  assign n841 = x94 & ~n840 ;
  assign n842 = x95 & n841 ;
  assign n843 = ~n839 & n842 ;
  assign n844 = x95 & ~x222 ;
  assign n845 = x223 & x224 ;
  assign n846 = ~n844 & n845 ;
  assign n847 = ~n843 & n846 ;
  assign n848 = ~x96 & x224 ;
  assign n849 = x97 & ~n848 ;
  assign n850 = x98 & n849 ;
  assign n851 = ~n847 & n850 ;
  assign n852 = x98 & ~x225 ;
  assign n853 = x226 & x227 ;
  assign n854 = ~n852 & n853 ;
  assign n855 = ~n851 & n854 ;
  assign n856 = ~x99 & x227 ;
  assign n857 = x100 & ~n856 ;
  assign n858 = x101 & n857 ;
  assign n859 = ~n855 & n858 ;
  assign n860 = x101 & ~x228 ;
  assign n861 = x229 & x230 ;
  assign n862 = ~n860 & n861 ;
  assign n863 = ~n859 & n862 ;
  assign n864 = ~x102 & x230 ;
  assign n865 = x103 & ~n864 ;
  assign n866 = x104 & n865 ;
  assign n867 = ~n863 & n866 ;
  assign n868 = x104 & ~x231 ;
  assign n869 = x232 & x233 ;
  assign n870 = ~n868 & n869 ;
  assign n871 = ~n867 & n870 ;
  assign n872 = ~x105 & x233 ;
  assign n873 = x106 & ~n872 ;
  assign n874 = x107 & n873 ;
  assign n875 = ~n871 & n874 ;
  assign n876 = x107 & ~x234 ;
  assign n877 = x235 & x236 ;
  assign n878 = ~n876 & n877 ;
  assign n879 = ~n875 & n878 ;
  assign n880 = ~x108 & x236 ;
  assign n881 = x109 & ~n880 ;
  assign n882 = x110 & n881 ;
  assign n883 = ~n879 & n882 ;
  assign n884 = x110 & ~x237 ;
  assign n885 = x238 & x239 ;
  assign n886 = ~n884 & n885 ;
  assign n887 = ~n883 & n886 ;
  assign n888 = ~x111 & x239 ;
  assign n889 = x112 & ~n888 ;
  assign n890 = x113 & n889 ;
  assign n891 = ~n887 & n890 ;
  assign n892 = x113 & ~x240 ;
  assign n893 = x241 & x242 ;
  assign n894 = ~n892 & n893 ;
  assign n895 = ~n891 & n894 ;
  assign n896 = ~x114 & x242 ;
  assign n897 = x115 & ~n896 ;
  assign n898 = x116 & n897 ;
  assign n899 = ~n895 & n898 ;
  assign n900 = x116 & ~x243 ;
  assign n901 = x244 & x245 ;
  assign n902 = ~n900 & n901 ;
  assign n903 = ~n899 & n902 ;
  assign n904 = ~x117 & x245 ;
  assign n905 = x118 & ~n904 ;
  assign n906 = x119 & n905 ;
  assign n907 = ~n903 & n906 ;
  assign n908 = x119 & ~x246 ;
  assign n909 = x247 & x248 ;
  assign n910 = ~n908 & n909 ;
  assign n911 = ~n907 & n910 ;
  assign n912 = ~x120 & x248 ;
  assign n913 = x121 & ~n912 ;
  assign n914 = x122 & n913 ;
  assign n915 = ~n911 & n914 ;
  assign n916 = x122 & ~x249 ;
  assign n917 = x250 & x251 ;
  assign n918 = ~n916 & n917 ;
  assign n919 = ~n915 & n918 ;
  assign n920 = ~x123 & x251 ;
  assign n921 = x124 & ~n920 ;
  assign n922 = x125 & n921 ;
  assign n923 = ~n919 & n922 ;
  assign n924 = x125 & ~x252 ;
  assign n925 = x253 & x254 ;
  assign n926 = ~n924 & n925 ;
  assign n927 = ~n923 & n926 ;
  assign n928 = ~x126 & x254 ;
  assign n929 = x127 & ~n928 ;
  assign n930 = x0 & n929 ;
  assign n931 = ~n927 & n930 ;
  assign n932 = x0 & ~x255 ;
  assign n933 = ~x128 & ~n932 ;
  assign n934 = ~n931 & n933 ;
  assign n937 = ~n934 & ~x256 ;
  assign n938 = ~n936 & ~n937 ;
  assign n939 = x2 & ~x130 ;
  assign n940 = ~x3 & ~n939 ;
  assign n941 = ~x131 & ~x132 ;
  assign n942 = ~n940 & n941 ;
  assign n943 = x4 & ~x132 ;
  assign n944 = ~x5 & ~n943 ;
  assign n945 = ~x6 & n944 ;
  assign n946 = ~n942 & n945 ;
  assign n947 = ~x6 & x133 ;
  assign n948 = ~x134 & ~x135 ;
  assign n949 = ~n947 & n948 ;
  assign n950 = ~n946 & n949 ;
  assign n951 = x7 & ~x135 ;
  assign n952 = ~x8 & ~n951 ;
  assign n953 = ~x9 & n952 ;
  assign n954 = ~n950 & n953 ;
  assign n955 = ~x9 & x136 ;
  assign n956 = ~x137 & ~x138 ;
  assign n957 = ~n955 & n956 ;
  assign n958 = ~n954 & n957 ;
  assign n959 = x10 & ~x138 ;
  assign n960 = ~x11 & ~n959 ;
  assign n961 = ~x12 & n960 ;
  assign n962 = ~n958 & n961 ;
  assign n963 = ~x12 & x139 ;
  assign n964 = ~x140 & ~x141 ;
  assign n965 = ~n963 & n964 ;
  assign n966 = ~n962 & n965 ;
  assign n967 = x13 & ~x141 ;
  assign n968 = ~x14 & ~n967 ;
  assign n969 = ~x15 & n968 ;
  assign n970 = ~n966 & n969 ;
  assign n971 = ~x15 & x142 ;
  assign n972 = ~x143 & ~x144 ;
  assign n973 = ~n971 & n972 ;
  assign n974 = ~n970 & n973 ;
  assign n975 = x16 & ~x144 ;
  assign n976 = ~x17 & ~n975 ;
  assign n977 = ~x18 & n976 ;
  assign n978 = ~n974 & n977 ;
  assign n979 = ~x18 & x145 ;
  assign n980 = ~x146 & ~x147 ;
  assign n981 = ~n979 & n980 ;
  assign n982 = ~n978 & n981 ;
  assign n983 = x19 & ~x147 ;
  assign n984 = ~x20 & ~n983 ;
  assign n985 = ~x21 & n984 ;
  assign n986 = ~n982 & n985 ;
  assign n987 = ~x21 & x148 ;
  assign n988 = ~x149 & ~x150 ;
  assign n989 = ~n987 & n988 ;
  assign n990 = ~n986 & n989 ;
  assign n991 = x22 & ~x150 ;
  assign n992 = ~x23 & ~n991 ;
  assign n993 = ~x24 & n992 ;
  assign n994 = ~n990 & n993 ;
  assign n995 = ~x24 & x151 ;
  assign n996 = ~x152 & ~x153 ;
  assign n997 = ~n995 & n996 ;
  assign n998 = ~n994 & n997 ;
  assign n999 = x25 & ~x153 ;
  assign n1000 = ~x26 & ~n999 ;
  assign n1001 = ~x27 & n1000 ;
  assign n1002 = ~n998 & n1001 ;
  assign n1003 = ~x27 & x154 ;
  assign n1004 = ~x155 & ~x156 ;
  assign n1005 = ~n1003 & n1004 ;
  assign n1006 = ~n1002 & n1005 ;
  assign n1007 = x28 & ~x156 ;
  assign n1008 = ~x29 & ~n1007 ;
  assign n1009 = ~x30 & n1008 ;
  assign n1010 = ~n1006 & n1009 ;
  assign n1011 = ~x30 & x157 ;
  assign n1012 = ~x158 & ~x159 ;
  assign n1013 = ~n1011 & n1012 ;
  assign n1014 = ~n1010 & n1013 ;
  assign n1015 = x31 & ~x159 ;
  assign n1016 = ~x32 & ~n1015 ;
  assign n1017 = ~x33 & n1016 ;
  assign n1018 = ~n1014 & n1017 ;
  assign n1019 = ~x33 & x160 ;
  assign n1020 = ~x161 & ~x162 ;
  assign n1021 = ~n1019 & n1020 ;
  assign n1022 = ~n1018 & n1021 ;
  assign n1023 = x34 & ~x162 ;
  assign n1024 = ~x35 & ~n1023 ;
  assign n1025 = ~x36 & n1024 ;
  assign n1026 = ~n1022 & n1025 ;
  assign n1027 = ~x36 & x163 ;
  assign n1028 = ~x164 & ~x165 ;
  assign n1029 = ~n1027 & n1028 ;
  assign n1030 = ~n1026 & n1029 ;
  assign n1031 = x37 & ~x165 ;
  assign n1032 = ~x38 & ~n1031 ;
  assign n1033 = ~x39 & n1032 ;
  assign n1034 = ~n1030 & n1033 ;
  assign n1035 = ~x39 & x166 ;
  assign n1036 = ~x167 & ~x168 ;
  assign n1037 = ~n1035 & n1036 ;
  assign n1038 = ~n1034 & n1037 ;
  assign n1039 = x40 & ~x168 ;
  assign n1040 = ~x41 & ~n1039 ;
  assign n1041 = ~x42 & n1040 ;
  assign n1042 = ~n1038 & n1041 ;
  assign n1043 = ~x42 & x169 ;
  assign n1044 = ~x170 & ~x171 ;
  assign n1045 = ~n1043 & n1044 ;
  assign n1046 = ~n1042 & n1045 ;
  assign n1047 = x43 & ~x171 ;
  assign n1048 = ~x44 & ~n1047 ;
  assign n1049 = ~x45 & n1048 ;
  assign n1050 = ~n1046 & n1049 ;
  assign n1051 = ~x45 & x172 ;
  assign n1052 = ~x173 & ~x174 ;
  assign n1053 = ~n1051 & n1052 ;
  assign n1054 = ~n1050 & n1053 ;
  assign n1055 = x46 & ~x174 ;
  assign n1056 = ~x47 & ~n1055 ;
  assign n1057 = ~x48 & n1056 ;
  assign n1058 = ~n1054 & n1057 ;
  assign n1059 = ~x48 & x175 ;
  assign n1060 = ~x176 & ~x177 ;
  assign n1061 = ~n1059 & n1060 ;
  assign n1062 = ~n1058 & n1061 ;
  assign n1063 = x49 & ~x177 ;
  assign n1064 = ~x50 & ~n1063 ;
  assign n1065 = ~x51 & n1064 ;
  assign n1066 = ~n1062 & n1065 ;
  assign n1067 = ~x51 & x178 ;
  assign n1068 = ~x179 & ~x180 ;
  assign n1069 = ~n1067 & n1068 ;
  assign n1070 = ~n1066 & n1069 ;
  assign n1071 = x52 & ~x180 ;
  assign n1072 = ~x53 & ~n1071 ;
  assign n1073 = ~x54 & n1072 ;
  assign n1074 = ~n1070 & n1073 ;
  assign n1075 = ~x54 & x181 ;
  assign n1076 = ~x182 & ~x183 ;
  assign n1077 = ~n1075 & n1076 ;
  assign n1078 = ~n1074 & n1077 ;
  assign n1079 = x55 & ~x183 ;
  assign n1080 = ~x56 & ~n1079 ;
  assign n1081 = ~x57 & n1080 ;
  assign n1082 = ~n1078 & n1081 ;
  assign n1083 = ~x57 & x184 ;
  assign n1084 = ~x185 & ~x186 ;
  assign n1085 = ~n1083 & n1084 ;
  assign n1086 = ~n1082 & n1085 ;
  assign n1087 = x58 & ~x186 ;
  assign n1088 = ~x59 & ~n1087 ;
  assign n1089 = ~x60 & n1088 ;
  assign n1090 = ~n1086 & n1089 ;
  assign n1091 = ~x60 & x187 ;
  assign n1092 = ~x188 & ~x189 ;
  assign n1093 = ~n1091 & n1092 ;
  assign n1094 = ~n1090 & n1093 ;
  assign n1095 = x61 & ~x189 ;
  assign n1096 = ~x62 & ~n1095 ;
  assign n1097 = ~x63 & n1096 ;
  assign n1098 = ~n1094 & n1097 ;
  assign n1099 = ~x63 & x190 ;
  assign n1100 = ~x191 & ~x192 ;
  assign n1101 = ~n1099 & n1100 ;
  assign n1102 = ~n1098 & n1101 ;
  assign n1103 = x64 & ~x192 ;
  assign n1104 = ~x65 & ~n1103 ;
  assign n1105 = ~x66 & n1104 ;
  assign n1106 = ~n1102 & n1105 ;
  assign n1107 = ~x66 & x193 ;
  assign n1108 = ~x194 & ~x195 ;
  assign n1109 = ~n1107 & n1108 ;
  assign n1110 = ~n1106 & n1109 ;
  assign n1111 = x67 & ~x195 ;
  assign n1112 = ~x68 & ~n1111 ;
  assign n1113 = ~x69 & n1112 ;
  assign n1114 = ~n1110 & n1113 ;
  assign n1115 = ~x69 & x196 ;
  assign n1116 = ~x197 & ~x198 ;
  assign n1117 = ~n1115 & n1116 ;
  assign n1118 = ~n1114 & n1117 ;
  assign n1119 = x70 & ~x198 ;
  assign n1120 = ~x71 & ~n1119 ;
  assign n1121 = ~x72 & n1120 ;
  assign n1122 = ~n1118 & n1121 ;
  assign n1123 = ~x72 & x199 ;
  assign n1124 = ~x200 & ~x201 ;
  assign n1125 = ~n1123 & n1124 ;
  assign n1126 = ~n1122 & n1125 ;
  assign n1127 = x73 & ~x201 ;
  assign n1128 = ~x74 & ~n1127 ;
  assign n1129 = ~x75 & n1128 ;
  assign n1130 = ~n1126 & n1129 ;
  assign n1131 = ~x75 & x202 ;
  assign n1132 = ~x203 & ~x204 ;
  assign n1133 = ~n1131 & n1132 ;
  assign n1134 = ~n1130 & n1133 ;
  assign n1135 = x76 & ~x204 ;
  assign n1136 = ~x77 & ~n1135 ;
  assign n1137 = ~x78 & n1136 ;
  assign n1138 = ~n1134 & n1137 ;
  assign n1139 = ~x78 & x205 ;
  assign n1140 = ~x206 & ~x207 ;
  assign n1141 = ~n1139 & n1140 ;
  assign n1142 = ~n1138 & n1141 ;
  assign n1143 = x79 & ~x207 ;
  assign n1144 = ~x80 & ~n1143 ;
  assign n1145 = ~x81 & n1144 ;
  assign n1146 = ~n1142 & n1145 ;
  assign n1147 = ~x81 & x208 ;
  assign n1148 = ~x209 & ~x210 ;
  assign n1149 = ~n1147 & n1148 ;
  assign n1150 = ~n1146 & n1149 ;
  assign n1151 = x82 & ~x210 ;
  assign n1152 = ~x83 & ~n1151 ;
  assign n1153 = ~x84 & n1152 ;
  assign n1154 = ~n1150 & n1153 ;
  assign n1155 = ~x84 & x211 ;
  assign n1156 = ~x212 & ~x213 ;
  assign n1157 = ~n1155 & n1156 ;
  assign n1158 = ~n1154 & n1157 ;
  assign n1159 = x85 & ~x213 ;
  assign n1160 = ~x86 & ~n1159 ;
  assign n1161 = ~x87 & n1160 ;
  assign n1162 = ~n1158 & n1161 ;
  assign n1163 = ~x87 & x214 ;
  assign n1164 = ~x215 & ~x216 ;
  assign n1165 = ~n1163 & n1164 ;
  assign n1166 = ~n1162 & n1165 ;
  assign n1167 = x88 & ~x216 ;
  assign n1168 = ~x89 & ~n1167 ;
  assign n1169 = ~x90 & n1168 ;
  assign n1170 = ~n1166 & n1169 ;
  assign n1171 = ~x90 & x217 ;
  assign n1172 = ~x218 & ~x219 ;
  assign n1173 = ~n1171 & n1172 ;
  assign n1174 = ~n1170 & n1173 ;
  assign n1175 = x91 & ~x219 ;
  assign n1176 = ~x92 & ~n1175 ;
  assign n1177 = ~x93 & n1176 ;
  assign n1178 = ~n1174 & n1177 ;
  assign n1179 = ~x93 & x220 ;
  assign n1180 = ~x221 & ~x222 ;
  assign n1181 = ~n1179 & n1180 ;
  assign n1182 = ~n1178 & n1181 ;
  assign n1183 = x94 & ~x222 ;
  assign n1184 = ~x95 & ~n1183 ;
  assign n1185 = ~x96 & n1184 ;
  assign n1186 = ~n1182 & n1185 ;
  assign n1187 = ~x96 & x223 ;
  assign n1188 = ~x224 & ~x225 ;
  assign n1189 = ~n1187 & n1188 ;
  assign n1190 = ~n1186 & n1189 ;
  assign n1191 = x97 & ~x225 ;
  assign n1192 = ~x98 & ~n1191 ;
  assign n1193 = ~x99 & n1192 ;
  assign n1194 = ~n1190 & n1193 ;
  assign n1195 = ~x99 & x226 ;
  assign n1196 = ~x227 & ~x228 ;
  assign n1197 = ~n1195 & n1196 ;
  assign n1198 = ~n1194 & n1197 ;
  assign n1199 = x100 & ~x228 ;
  assign n1200 = ~x101 & ~n1199 ;
  assign n1201 = ~x102 & n1200 ;
  assign n1202 = ~n1198 & n1201 ;
  assign n1203 = ~x102 & x229 ;
  assign n1204 = ~x230 & ~x231 ;
  assign n1205 = ~n1203 & n1204 ;
  assign n1206 = ~n1202 & n1205 ;
  assign n1207 = x103 & ~x231 ;
  assign n1208 = ~x104 & ~n1207 ;
  assign n1209 = ~x105 & n1208 ;
  assign n1210 = ~n1206 & n1209 ;
  assign n1211 = ~x105 & x232 ;
  assign n1212 = ~x233 & ~x234 ;
  assign n1213 = ~n1211 & n1212 ;
  assign n1214 = ~n1210 & n1213 ;
  assign n1215 = x106 & ~x234 ;
  assign n1216 = ~x107 & ~n1215 ;
  assign n1217 = ~x108 & n1216 ;
  assign n1218 = ~n1214 & n1217 ;
  assign n1219 = ~x108 & x235 ;
  assign n1220 = ~x236 & ~x237 ;
  assign n1221 = ~n1219 & n1220 ;
  assign n1222 = ~n1218 & n1221 ;
  assign n1223 = x109 & ~x237 ;
  assign n1224 = ~x110 & ~n1223 ;
  assign n1225 = ~x111 & n1224 ;
  assign n1226 = ~n1222 & n1225 ;
  assign n1227 = ~x111 & x238 ;
  assign n1228 = ~x239 & ~x240 ;
  assign n1229 = ~n1227 & n1228 ;
  assign n1230 = ~n1226 & n1229 ;
  assign n1231 = x112 & ~x240 ;
  assign n1232 = ~x113 & ~n1231 ;
  assign n1233 = ~x114 & n1232 ;
  assign n1234 = ~n1230 & n1233 ;
  assign n1235 = ~x114 & x241 ;
  assign n1236 = ~x242 & ~x243 ;
  assign n1237 = ~n1235 & n1236 ;
  assign n1238 = ~n1234 & n1237 ;
  assign n1239 = x115 & ~x243 ;
  assign n1240 = ~x116 & ~n1239 ;
  assign n1241 = ~x117 & n1240 ;
  assign n1242 = ~n1238 & n1241 ;
  assign n1243 = ~x117 & x244 ;
  assign n1244 = ~x245 & ~x246 ;
  assign n1245 = ~n1243 & n1244 ;
  assign n1246 = ~n1242 & n1245 ;
  assign n1247 = x118 & ~x246 ;
  assign n1248 = ~x119 & ~n1247 ;
  assign n1249 = ~x120 & n1248 ;
  assign n1250 = ~n1246 & n1249 ;
  assign n1251 = ~x120 & x247 ;
  assign n1252 = ~x248 & ~x249 ;
  assign n1253 = ~n1251 & n1252 ;
  assign n1254 = ~n1250 & n1253 ;
  assign n1255 = x121 & ~x249 ;
  assign n1256 = ~x122 & ~n1255 ;
  assign n1257 = ~x123 & n1256 ;
  assign n1258 = ~n1254 & n1257 ;
  assign n1259 = ~x123 & x250 ;
  assign n1260 = ~x251 & ~x252 ;
  assign n1261 = ~n1259 & n1260 ;
  assign n1262 = ~n1258 & n1261 ;
  assign n1263 = x124 & ~x252 ;
  assign n1264 = ~x125 & ~n1263 ;
  assign n1265 = ~x126 & n1264 ;
  assign n1266 = ~n1262 & n1265 ;
  assign n1267 = ~x126 & x253 ;
  assign n1268 = ~x254 & ~x255 ;
  assign n1269 = ~n1267 & n1268 ;
  assign n1270 = ~n1266 & n1269 ;
  assign n1271 = x127 & ~x255 ;
  assign n1272 = ~x0 & ~n1271 ;
  assign n1273 = ~x1 & n1272 ;
  assign n1274 = ~n1270 & n1273 ;
  assign n1275 = ~x1 & x128 ;
  assign n1276 = x129 & ~n1275 ;
  assign n1277 = ~n1274 & n1276 ;
  assign n1618 = n1277 & x257 ;
  assign n1278 = ~x2 & x130 ;
  assign n1279 = x3 & ~n1278 ;
  assign n1280 = x131 & x132 ;
  assign n1281 = ~n1279 & n1280 ;
  assign n1282 = ~x4 & x132 ;
  assign n1283 = x5 & ~n1282 ;
  assign n1284 = x6 & n1283 ;
  assign n1285 = ~n1281 & n1284 ;
  assign n1286 = x6 & ~x133 ;
  assign n1287 = x134 & x135 ;
  assign n1288 = ~n1286 & n1287 ;
  assign n1289 = ~n1285 & n1288 ;
  assign n1290 = ~x7 & x135 ;
  assign n1291 = x8 & ~n1290 ;
  assign n1292 = x9 & n1291 ;
  assign n1293 = ~n1289 & n1292 ;
  assign n1294 = x9 & ~x136 ;
  assign n1295 = x137 & x138 ;
  assign n1296 = ~n1294 & n1295 ;
  assign n1297 = ~n1293 & n1296 ;
  assign n1298 = ~x10 & x138 ;
  assign n1299 = x11 & ~n1298 ;
  assign n1300 = x12 & n1299 ;
  assign n1301 = ~n1297 & n1300 ;
  assign n1302 = x12 & ~x139 ;
  assign n1303 = x140 & x141 ;
  assign n1304 = ~n1302 & n1303 ;
  assign n1305 = ~n1301 & n1304 ;
  assign n1306 = ~x13 & x141 ;
  assign n1307 = x14 & ~n1306 ;
  assign n1308 = x15 & n1307 ;
  assign n1309 = ~n1305 & n1308 ;
  assign n1310 = x15 & ~x142 ;
  assign n1311 = x143 & x144 ;
  assign n1312 = ~n1310 & n1311 ;
  assign n1313 = ~n1309 & n1312 ;
  assign n1314 = ~x16 & x144 ;
  assign n1315 = x17 & ~n1314 ;
  assign n1316 = x18 & n1315 ;
  assign n1317 = ~n1313 & n1316 ;
  assign n1318 = x18 & ~x145 ;
  assign n1319 = x146 & x147 ;
  assign n1320 = ~n1318 & n1319 ;
  assign n1321 = ~n1317 & n1320 ;
  assign n1322 = ~x19 & x147 ;
  assign n1323 = x20 & ~n1322 ;
  assign n1324 = x21 & n1323 ;
  assign n1325 = ~n1321 & n1324 ;
  assign n1326 = x21 & ~x148 ;
  assign n1327 = x149 & x150 ;
  assign n1328 = ~n1326 & n1327 ;
  assign n1329 = ~n1325 & n1328 ;
  assign n1330 = ~x22 & x150 ;
  assign n1331 = x23 & ~n1330 ;
  assign n1332 = x24 & n1331 ;
  assign n1333 = ~n1329 & n1332 ;
  assign n1334 = x24 & ~x151 ;
  assign n1335 = x152 & x153 ;
  assign n1336 = ~n1334 & n1335 ;
  assign n1337 = ~n1333 & n1336 ;
  assign n1338 = ~x25 & x153 ;
  assign n1339 = x26 & ~n1338 ;
  assign n1340 = x27 & n1339 ;
  assign n1341 = ~n1337 & n1340 ;
  assign n1342 = x27 & ~x154 ;
  assign n1343 = x155 & x156 ;
  assign n1344 = ~n1342 & n1343 ;
  assign n1345 = ~n1341 & n1344 ;
  assign n1346 = ~x28 & x156 ;
  assign n1347 = x29 & ~n1346 ;
  assign n1348 = x30 & n1347 ;
  assign n1349 = ~n1345 & n1348 ;
  assign n1350 = x30 & ~x157 ;
  assign n1351 = x158 & x159 ;
  assign n1352 = ~n1350 & n1351 ;
  assign n1353 = ~n1349 & n1352 ;
  assign n1354 = ~x31 & x159 ;
  assign n1355 = x32 & ~n1354 ;
  assign n1356 = x33 & n1355 ;
  assign n1357 = ~n1353 & n1356 ;
  assign n1358 = x33 & ~x160 ;
  assign n1359 = x161 & x162 ;
  assign n1360 = ~n1358 & n1359 ;
  assign n1361 = ~n1357 & n1360 ;
  assign n1362 = ~x34 & x162 ;
  assign n1363 = x35 & ~n1362 ;
  assign n1364 = x36 & n1363 ;
  assign n1365 = ~n1361 & n1364 ;
  assign n1366 = x36 & ~x163 ;
  assign n1367 = x164 & x165 ;
  assign n1368 = ~n1366 & n1367 ;
  assign n1369 = ~n1365 & n1368 ;
  assign n1370 = ~x37 & x165 ;
  assign n1371 = x38 & ~n1370 ;
  assign n1372 = x39 & n1371 ;
  assign n1373 = ~n1369 & n1372 ;
  assign n1374 = x39 & ~x166 ;
  assign n1375 = x167 & x168 ;
  assign n1376 = ~n1374 & n1375 ;
  assign n1377 = ~n1373 & n1376 ;
  assign n1378 = ~x40 & x168 ;
  assign n1379 = x41 & ~n1378 ;
  assign n1380 = x42 & n1379 ;
  assign n1381 = ~n1377 & n1380 ;
  assign n1382 = x42 & ~x169 ;
  assign n1383 = x170 & x171 ;
  assign n1384 = ~n1382 & n1383 ;
  assign n1385 = ~n1381 & n1384 ;
  assign n1386 = ~x43 & x171 ;
  assign n1387 = x44 & ~n1386 ;
  assign n1388 = x45 & n1387 ;
  assign n1389 = ~n1385 & n1388 ;
  assign n1390 = x45 & ~x172 ;
  assign n1391 = x173 & x174 ;
  assign n1392 = ~n1390 & n1391 ;
  assign n1393 = ~n1389 & n1392 ;
  assign n1394 = ~x46 & x174 ;
  assign n1395 = x47 & ~n1394 ;
  assign n1396 = x48 & n1395 ;
  assign n1397 = ~n1393 & n1396 ;
  assign n1398 = x48 & ~x175 ;
  assign n1399 = x176 & x177 ;
  assign n1400 = ~n1398 & n1399 ;
  assign n1401 = ~n1397 & n1400 ;
  assign n1402 = ~x49 & x177 ;
  assign n1403 = x50 & ~n1402 ;
  assign n1404 = x51 & n1403 ;
  assign n1405 = ~n1401 & n1404 ;
  assign n1406 = x51 & ~x178 ;
  assign n1407 = x179 & x180 ;
  assign n1408 = ~n1406 & n1407 ;
  assign n1409 = ~n1405 & n1408 ;
  assign n1410 = ~x52 & x180 ;
  assign n1411 = x53 & ~n1410 ;
  assign n1412 = x54 & n1411 ;
  assign n1413 = ~n1409 & n1412 ;
  assign n1414 = x54 & ~x181 ;
  assign n1415 = x182 & x183 ;
  assign n1416 = ~n1414 & n1415 ;
  assign n1417 = ~n1413 & n1416 ;
  assign n1418 = ~x55 & x183 ;
  assign n1419 = x56 & ~n1418 ;
  assign n1420 = x57 & n1419 ;
  assign n1421 = ~n1417 & n1420 ;
  assign n1422 = x57 & ~x184 ;
  assign n1423 = x185 & x186 ;
  assign n1424 = ~n1422 & n1423 ;
  assign n1425 = ~n1421 & n1424 ;
  assign n1426 = ~x58 & x186 ;
  assign n1427 = x59 & ~n1426 ;
  assign n1428 = x60 & n1427 ;
  assign n1429 = ~n1425 & n1428 ;
  assign n1430 = x60 & ~x187 ;
  assign n1431 = x188 & x189 ;
  assign n1432 = ~n1430 & n1431 ;
  assign n1433 = ~n1429 & n1432 ;
  assign n1434 = ~x61 & x189 ;
  assign n1435 = x62 & ~n1434 ;
  assign n1436 = x63 & n1435 ;
  assign n1437 = ~n1433 & n1436 ;
  assign n1438 = x63 & ~x190 ;
  assign n1439 = x191 & x192 ;
  assign n1440 = ~n1438 & n1439 ;
  assign n1441 = ~n1437 & n1440 ;
  assign n1442 = ~x64 & x192 ;
  assign n1443 = x65 & ~n1442 ;
  assign n1444 = x66 & n1443 ;
  assign n1445 = ~n1441 & n1444 ;
  assign n1446 = x66 & ~x193 ;
  assign n1447 = x194 & x195 ;
  assign n1448 = ~n1446 & n1447 ;
  assign n1449 = ~n1445 & n1448 ;
  assign n1450 = ~x67 & x195 ;
  assign n1451 = x68 & ~n1450 ;
  assign n1452 = x69 & n1451 ;
  assign n1453 = ~n1449 & n1452 ;
  assign n1454 = x69 & ~x196 ;
  assign n1455 = x197 & x198 ;
  assign n1456 = ~n1454 & n1455 ;
  assign n1457 = ~n1453 & n1456 ;
  assign n1458 = ~x70 & x198 ;
  assign n1459 = x71 & ~n1458 ;
  assign n1460 = x72 & n1459 ;
  assign n1461 = ~n1457 & n1460 ;
  assign n1462 = x72 & ~x199 ;
  assign n1463 = x200 & x201 ;
  assign n1464 = ~n1462 & n1463 ;
  assign n1465 = ~n1461 & n1464 ;
  assign n1466 = ~x73 & x201 ;
  assign n1467 = x74 & ~n1466 ;
  assign n1468 = x75 & n1467 ;
  assign n1469 = ~n1465 & n1468 ;
  assign n1470 = x75 & ~x202 ;
  assign n1471 = x203 & x204 ;
  assign n1472 = ~n1470 & n1471 ;
  assign n1473 = ~n1469 & n1472 ;
  assign n1474 = ~x76 & x204 ;
  assign n1475 = x77 & ~n1474 ;
  assign n1476 = x78 & n1475 ;
  assign n1477 = ~n1473 & n1476 ;
  assign n1478 = x78 & ~x205 ;
  assign n1479 = x206 & x207 ;
  assign n1480 = ~n1478 & n1479 ;
  assign n1481 = ~n1477 & n1480 ;
  assign n1482 = ~x79 & x207 ;
  assign n1483 = x80 & ~n1482 ;
  assign n1484 = x81 & n1483 ;
  assign n1485 = ~n1481 & n1484 ;
  assign n1486 = x81 & ~x208 ;
  assign n1487 = x209 & x210 ;
  assign n1488 = ~n1486 & n1487 ;
  assign n1489 = ~n1485 & n1488 ;
  assign n1490 = ~x82 & x210 ;
  assign n1491 = x83 & ~n1490 ;
  assign n1492 = x84 & n1491 ;
  assign n1493 = ~n1489 & n1492 ;
  assign n1494 = x84 & ~x211 ;
  assign n1495 = x212 & x213 ;
  assign n1496 = ~n1494 & n1495 ;
  assign n1497 = ~n1493 & n1496 ;
  assign n1498 = ~x85 & x213 ;
  assign n1499 = x86 & ~n1498 ;
  assign n1500 = x87 & n1499 ;
  assign n1501 = ~n1497 & n1500 ;
  assign n1502 = x87 & ~x214 ;
  assign n1503 = x215 & x216 ;
  assign n1504 = ~n1502 & n1503 ;
  assign n1505 = ~n1501 & n1504 ;
  assign n1506 = ~x88 & x216 ;
  assign n1507 = x89 & ~n1506 ;
  assign n1508 = x90 & n1507 ;
  assign n1509 = ~n1505 & n1508 ;
  assign n1510 = x90 & ~x217 ;
  assign n1511 = x218 & x219 ;
  assign n1512 = ~n1510 & n1511 ;
  assign n1513 = ~n1509 & n1512 ;
  assign n1514 = ~x91 & x219 ;
  assign n1515 = x92 & ~n1514 ;
  assign n1516 = x93 & n1515 ;
  assign n1517 = ~n1513 & n1516 ;
  assign n1518 = x93 & ~x220 ;
  assign n1519 = x221 & x222 ;
  assign n1520 = ~n1518 & n1519 ;
  assign n1521 = ~n1517 & n1520 ;
  assign n1522 = ~x94 & x222 ;
  assign n1523 = x95 & ~n1522 ;
  assign n1524 = x96 & n1523 ;
  assign n1525 = ~n1521 & n1524 ;
  assign n1526 = x96 & ~x223 ;
  assign n1527 = x224 & x225 ;
  assign n1528 = ~n1526 & n1527 ;
  assign n1529 = ~n1525 & n1528 ;
  assign n1530 = ~x97 & x225 ;
  assign n1531 = x98 & ~n1530 ;
  assign n1532 = x99 & n1531 ;
  assign n1533 = ~n1529 & n1532 ;
  assign n1534 = x99 & ~x226 ;
  assign n1535 = x227 & x228 ;
  assign n1536 = ~n1534 & n1535 ;
  assign n1537 = ~n1533 & n1536 ;
  assign n1538 = ~x100 & x228 ;
  assign n1539 = x101 & ~n1538 ;
  assign n1540 = x102 & n1539 ;
  assign n1541 = ~n1537 & n1540 ;
  assign n1542 = x102 & ~x229 ;
  assign n1543 = x230 & x231 ;
  assign n1544 = ~n1542 & n1543 ;
  assign n1545 = ~n1541 & n1544 ;
  assign n1546 = ~x103 & x231 ;
  assign n1547 = x104 & ~n1546 ;
  assign n1548 = x105 & n1547 ;
  assign n1549 = ~n1545 & n1548 ;
  assign n1550 = x105 & ~x232 ;
  assign n1551 = x233 & x234 ;
  assign n1552 = ~n1550 & n1551 ;
  assign n1553 = ~n1549 & n1552 ;
  assign n1554 = ~x106 & x234 ;
  assign n1555 = x107 & ~n1554 ;
  assign n1556 = x108 & n1555 ;
  assign n1557 = ~n1553 & n1556 ;
  assign n1558 = x108 & ~x235 ;
  assign n1559 = x236 & x237 ;
  assign n1560 = ~n1558 & n1559 ;
  assign n1561 = ~n1557 & n1560 ;
  assign n1562 = ~x109 & x237 ;
  assign n1563 = x110 & ~n1562 ;
  assign n1564 = x111 & n1563 ;
  assign n1565 = ~n1561 & n1564 ;
  assign n1566 = x111 & ~x238 ;
  assign n1567 = x239 & x240 ;
  assign n1568 = ~n1566 & n1567 ;
  assign n1569 = ~n1565 & n1568 ;
  assign n1570 = ~x112 & x240 ;
  assign n1571 = x113 & ~n1570 ;
  assign n1572 = x114 & n1571 ;
  assign n1573 = ~n1569 & n1572 ;
  assign n1574 = x114 & ~x241 ;
  assign n1575 = x242 & x243 ;
  assign n1576 = ~n1574 & n1575 ;
  assign n1577 = ~n1573 & n1576 ;
  assign n1578 = ~x115 & x243 ;
  assign n1579 = x116 & ~n1578 ;
  assign n1580 = x117 & n1579 ;
  assign n1581 = ~n1577 & n1580 ;
  assign n1582 = x117 & ~x244 ;
  assign n1583 = x245 & x246 ;
  assign n1584 = ~n1582 & n1583 ;
  assign n1585 = ~n1581 & n1584 ;
  assign n1586 = ~x118 & x246 ;
  assign n1587 = x119 & ~n1586 ;
  assign n1588 = x120 & n1587 ;
  assign n1589 = ~n1585 & n1588 ;
  assign n1590 = x120 & ~x247 ;
  assign n1591 = x248 & x249 ;
  assign n1592 = ~n1590 & n1591 ;
  assign n1593 = ~n1589 & n1592 ;
  assign n1594 = ~x121 & x249 ;
  assign n1595 = x122 & ~n1594 ;
  assign n1596 = x123 & n1595 ;
  assign n1597 = ~n1593 & n1596 ;
  assign n1598 = x123 & ~x250 ;
  assign n1599 = x251 & x252 ;
  assign n1600 = ~n1598 & n1599 ;
  assign n1601 = ~n1597 & n1600 ;
  assign n1602 = ~x124 & x252 ;
  assign n1603 = x125 & ~n1602 ;
  assign n1604 = x126 & n1603 ;
  assign n1605 = ~n1601 & n1604 ;
  assign n1606 = x126 & ~x253 ;
  assign n1607 = x254 & x255 ;
  assign n1608 = ~n1606 & n1607 ;
  assign n1609 = ~n1605 & n1608 ;
  assign n1610 = ~x127 & x255 ;
  assign n1611 = x0 & ~n1610 ;
  assign n1612 = x1 & n1611 ;
  assign n1613 = ~n1609 & n1612 ;
  assign n1614 = x1 & ~x128 ;
  assign n1615 = ~x129 & ~n1614 ;
  assign n1616 = ~n1613 & n1615 ;
  assign n1619 = ~n1616 & ~x257 ;
  assign n1620 = ~n1618 & ~n1619 ;
  assign n1621 = ~x132 & ~x133 ;
  assign n1622 = ~n262 & n1621 ;
  assign n1623 = x5 & ~x133 ;
  assign n1624 = ~x6 & ~n1623 ;
  assign n1625 = ~x7 & n1624 ;
  assign n1626 = ~n1622 & n1625 ;
  assign n1627 = ~x7 & x134 ;
  assign n1628 = ~x135 & ~x136 ;
  assign n1629 = ~n1627 & n1628 ;
  assign n1630 = ~n1626 & n1629 ;
  assign n1631 = x8 & ~x136 ;
  assign n1632 = ~x9 & ~n1631 ;
  assign n1633 = ~x10 & n1632 ;
  assign n1634 = ~n1630 & n1633 ;
  assign n1635 = ~x10 & x137 ;
  assign n1636 = ~x138 & ~x139 ;
  assign n1637 = ~n1635 & n1636 ;
  assign n1638 = ~n1634 & n1637 ;
  assign n1639 = x11 & ~x139 ;
  assign n1640 = ~x12 & ~n1639 ;
  assign n1641 = ~x13 & n1640 ;
  assign n1642 = ~n1638 & n1641 ;
  assign n1643 = ~x13 & x140 ;
  assign n1644 = ~x141 & ~x142 ;
  assign n1645 = ~n1643 & n1644 ;
  assign n1646 = ~n1642 & n1645 ;
  assign n1647 = x14 & ~x142 ;
  assign n1648 = ~x15 & ~n1647 ;
  assign n1649 = ~x16 & n1648 ;
  assign n1650 = ~n1646 & n1649 ;
  assign n1651 = ~x16 & x143 ;
  assign n1652 = ~x144 & ~x145 ;
  assign n1653 = ~n1651 & n1652 ;
  assign n1654 = ~n1650 & n1653 ;
  assign n1655 = x17 & ~x145 ;
  assign n1656 = ~x18 & ~n1655 ;
  assign n1657 = ~x19 & n1656 ;
  assign n1658 = ~n1654 & n1657 ;
  assign n1659 = ~x19 & x146 ;
  assign n1660 = ~x147 & ~x148 ;
  assign n1661 = ~n1659 & n1660 ;
  assign n1662 = ~n1658 & n1661 ;
  assign n1663 = x20 & ~x148 ;
  assign n1664 = ~x21 & ~n1663 ;
  assign n1665 = ~x22 & n1664 ;
  assign n1666 = ~n1662 & n1665 ;
  assign n1667 = ~x22 & x149 ;
  assign n1668 = ~x150 & ~x151 ;
  assign n1669 = ~n1667 & n1668 ;
  assign n1670 = ~n1666 & n1669 ;
  assign n1671 = x23 & ~x151 ;
  assign n1672 = ~x24 & ~n1671 ;
  assign n1673 = ~x25 & n1672 ;
  assign n1674 = ~n1670 & n1673 ;
  assign n1675 = ~x25 & x152 ;
  assign n1676 = ~x153 & ~x154 ;
  assign n1677 = ~n1675 & n1676 ;
  assign n1678 = ~n1674 & n1677 ;
  assign n1679 = x26 & ~x154 ;
  assign n1680 = ~x27 & ~n1679 ;
  assign n1681 = ~x28 & n1680 ;
  assign n1682 = ~n1678 & n1681 ;
  assign n1683 = ~x28 & x155 ;
  assign n1684 = ~x156 & ~x157 ;
  assign n1685 = ~n1683 & n1684 ;
  assign n1686 = ~n1682 & n1685 ;
  assign n1687 = x29 & ~x157 ;
  assign n1688 = ~x30 & ~n1687 ;
  assign n1689 = ~x31 & n1688 ;
  assign n1690 = ~n1686 & n1689 ;
  assign n1691 = ~x31 & x158 ;
  assign n1692 = ~x159 & ~x160 ;
  assign n1693 = ~n1691 & n1692 ;
  assign n1694 = ~n1690 & n1693 ;
  assign n1695 = x32 & ~x160 ;
  assign n1696 = ~x33 & ~n1695 ;
  assign n1697 = ~x34 & n1696 ;
  assign n1698 = ~n1694 & n1697 ;
  assign n1699 = ~x34 & x161 ;
  assign n1700 = ~x162 & ~x163 ;
  assign n1701 = ~n1699 & n1700 ;
  assign n1702 = ~n1698 & n1701 ;
  assign n1703 = x35 & ~x163 ;
  assign n1704 = ~x36 & ~n1703 ;
  assign n1705 = ~x37 & n1704 ;
  assign n1706 = ~n1702 & n1705 ;
  assign n1707 = ~x37 & x164 ;
  assign n1708 = ~x165 & ~x166 ;
  assign n1709 = ~n1707 & n1708 ;
  assign n1710 = ~n1706 & n1709 ;
  assign n1711 = x38 & ~x166 ;
  assign n1712 = ~x39 & ~n1711 ;
  assign n1713 = ~x40 & n1712 ;
  assign n1714 = ~n1710 & n1713 ;
  assign n1715 = ~x40 & x167 ;
  assign n1716 = ~x168 & ~x169 ;
  assign n1717 = ~n1715 & n1716 ;
  assign n1718 = ~n1714 & n1717 ;
  assign n1719 = x41 & ~x169 ;
  assign n1720 = ~x42 & ~n1719 ;
  assign n1721 = ~x43 & n1720 ;
  assign n1722 = ~n1718 & n1721 ;
  assign n1723 = ~x43 & x170 ;
  assign n1724 = ~x171 & ~x172 ;
  assign n1725 = ~n1723 & n1724 ;
  assign n1726 = ~n1722 & n1725 ;
  assign n1727 = x44 & ~x172 ;
  assign n1728 = ~x45 & ~n1727 ;
  assign n1729 = ~x46 & n1728 ;
  assign n1730 = ~n1726 & n1729 ;
  assign n1731 = ~x46 & x173 ;
  assign n1732 = ~x174 & ~x175 ;
  assign n1733 = ~n1731 & n1732 ;
  assign n1734 = ~n1730 & n1733 ;
  assign n1735 = x47 & ~x175 ;
  assign n1736 = ~x48 & ~n1735 ;
  assign n1737 = ~x49 & n1736 ;
  assign n1738 = ~n1734 & n1737 ;
  assign n1739 = ~x49 & x176 ;
  assign n1740 = ~x177 & ~x178 ;
  assign n1741 = ~n1739 & n1740 ;
  assign n1742 = ~n1738 & n1741 ;
  assign n1743 = x50 & ~x178 ;
  assign n1744 = ~x51 & ~n1743 ;
  assign n1745 = ~x52 & n1744 ;
  assign n1746 = ~n1742 & n1745 ;
  assign n1747 = ~x52 & x179 ;
  assign n1748 = ~x180 & ~x181 ;
  assign n1749 = ~n1747 & n1748 ;
  assign n1750 = ~n1746 & n1749 ;
  assign n1751 = x53 & ~x181 ;
  assign n1752 = ~x54 & ~n1751 ;
  assign n1753 = ~x55 & n1752 ;
  assign n1754 = ~n1750 & n1753 ;
  assign n1755 = ~x55 & x182 ;
  assign n1756 = ~x183 & ~x184 ;
  assign n1757 = ~n1755 & n1756 ;
  assign n1758 = ~n1754 & n1757 ;
  assign n1759 = x56 & ~x184 ;
  assign n1760 = ~x57 & ~n1759 ;
  assign n1761 = ~x58 & n1760 ;
  assign n1762 = ~n1758 & n1761 ;
  assign n1763 = ~x58 & x185 ;
  assign n1764 = ~x186 & ~x187 ;
  assign n1765 = ~n1763 & n1764 ;
  assign n1766 = ~n1762 & n1765 ;
  assign n1767 = x59 & ~x187 ;
  assign n1768 = ~x60 & ~n1767 ;
  assign n1769 = ~x61 & n1768 ;
  assign n1770 = ~n1766 & n1769 ;
  assign n1771 = ~x61 & x188 ;
  assign n1772 = ~x189 & ~x190 ;
  assign n1773 = ~n1771 & n1772 ;
  assign n1774 = ~n1770 & n1773 ;
  assign n1775 = x62 & ~x190 ;
  assign n1776 = ~x63 & ~n1775 ;
  assign n1777 = ~x64 & n1776 ;
  assign n1778 = ~n1774 & n1777 ;
  assign n1779 = ~x64 & x191 ;
  assign n1780 = ~x192 & ~x193 ;
  assign n1781 = ~n1779 & n1780 ;
  assign n1782 = ~n1778 & n1781 ;
  assign n1783 = x65 & ~x193 ;
  assign n1784 = ~x66 & ~n1783 ;
  assign n1785 = ~x67 & n1784 ;
  assign n1786 = ~n1782 & n1785 ;
  assign n1787 = ~x67 & x194 ;
  assign n1788 = ~x195 & ~x196 ;
  assign n1789 = ~n1787 & n1788 ;
  assign n1790 = ~n1786 & n1789 ;
  assign n1791 = x68 & ~x196 ;
  assign n1792 = ~x69 & ~n1791 ;
  assign n1793 = ~x70 & n1792 ;
  assign n1794 = ~n1790 & n1793 ;
  assign n1795 = ~x70 & x197 ;
  assign n1796 = ~x198 & ~x199 ;
  assign n1797 = ~n1795 & n1796 ;
  assign n1798 = ~n1794 & n1797 ;
  assign n1799 = x71 & ~x199 ;
  assign n1800 = ~x72 & ~n1799 ;
  assign n1801 = ~x73 & n1800 ;
  assign n1802 = ~n1798 & n1801 ;
  assign n1803 = ~x73 & x200 ;
  assign n1804 = ~x201 & ~x202 ;
  assign n1805 = ~n1803 & n1804 ;
  assign n1806 = ~n1802 & n1805 ;
  assign n1807 = x74 & ~x202 ;
  assign n1808 = ~x75 & ~n1807 ;
  assign n1809 = ~x76 & n1808 ;
  assign n1810 = ~n1806 & n1809 ;
  assign n1811 = ~x76 & x203 ;
  assign n1812 = ~x204 & ~x205 ;
  assign n1813 = ~n1811 & n1812 ;
  assign n1814 = ~n1810 & n1813 ;
  assign n1815 = x77 & ~x205 ;
  assign n1816 = ~x78 & ~n1815 ;
  assign n1817 = ~x79 & n1816 ;
  assign n1818 = ~n1814 & n1817 ;
  assign n1819 = ~x79 & x206 ;
  assign n1820 = ~x207 & ~x208 ;
  assign n1821 = ~n1819 & n1820 ;
  assign n1822 = ~n1818 & n1821 ;
  assign n1823 = x80 & ~x208 ;
  assign n1824 = ~x81 & ~n1823 ;
  assign n1825 = ~x82 & n1824 ;
  assign n1826 = ~n1822 & n1825 ;
  assign n1827 = ~x82 & x209 ;
  assign n1828 = ~x210 & ~x211 ;
  assign n1829 = ~n1827 & n1828 ;
  assign n1830 = ~n1826 & n1829 ;
  assign n1831 = x83 & ~x211 ;
  assign n1832 = ~x84 & ~n1831 ;
  assign n1833 = ~x85 & n1832 ;
  assign n1834 = ~n1830 & n1833 ;
  assign n1835 = ~x85 & x212 ;
  assign n1836 = ~x213 & ~x214 ;
  assign n1837 = ~n1835 & n1836 ;
  assign n1838 = ~n1834 & n1837 ;
  assign n1839 = x86 & ~x214 ;
  assign n1840 = ~x87 & ~n1839 ;
  assign n1841 = ~x88 & n1840 ;
  assign n1842 = ~n1838 & n1841 ;
  assign n1843 = ~x88 & x215 ;
  assign n1844 = ~x216 & ~x217 ;
  assign n1845 = ~n1843 & n1844 ;
  assign n1846 = ~n1842 & n1845 ;
  assign n1847 = x89 & ~x217 ;
  assign n1848 = ~x90 & ~n1847 ;
  assign n1849 = ~x91 & n1848 ;
  assign n1850 = ~n1846 & n1849 ;
  assign n1851 = ~x91 & x218 ;
  assign n1852 = ~x219 & ~x220 ;
  assign n1853 = ~n1851 & n1852 ;
  assign n1854 = ~n1850 & n1853 ;
  assign n1855 = x92 & ~x220 ;
  assign n1856 = ~x93 & ~n1855 ;
  assign n1857 = ~x94 & n1856 ;
  assign n1858 = ~n1854 & n1857 ;
  assign n1859 = ~x94 & x221 ;
  assign n1860 = ~x222 & ~x223 ;
  assign n1861 = ~n1859 & n1860 ;
  assign n1862 = ~n1858 & n1861 ;
  assign n1863 = x95 & ~x223 ;
  assign n1864 = ~x96 & ~n1863 ;
  assign n1865 = ~x97 & n1864 ;
  assign n1866 = ~n1862 & n1865 ;
  assign n1867 = ~x97 & x224 ;
  assign n1868 = ~x225 & ~x226 ;
  assign n1869 = ~n1867 & n1868 ;
  assign n1870 = ~n1866 & n1869 ;
  assign n1871 = x98 & ~x226 ;
  assign n1872 = ~x99 & ~n1871 ;
  assign n1873 = ~x100 & n1872 ;
  assign n1874 = ~n1870 & n1873 ;
  assign n1875 = ~x100 & x227 ;
  assign n1876 = ~x228 & ~x229 ;
  assign n1877 = ~n1875 & n1876 ;
  assign n1878 = ~n1874 & n1877 ;
  assign n1879 = x101 & ~x229 ;
  assign n1880 = ~x102 & ~n1879 ;
  assign n1881 = ~x103 & n1880 ;
  assign n1882 = ~n1878 & n1881 ;
  assign n1883 = ~x103 & x230 ;
  assign n1884 = ~x231 & ~x232 ;
  assign n1885 = ~n1883 & n1884 ;
  assign n1886 = ~n1882 & n1885 ;
  assign n1887 = x104 & ~x232 ;
  assign n1888 = ~x105 & ~n1887 ;
  assign n1889 = ~x106 & n1888 ;
  assign n1890 = ~n1886 & n1889 ;
  assign n1891 = ~x106 & x233 ;
  assign n1892 = ~x234 & ~x235 ;
  assign n1893 = ~n1891 & n1892 ;
  assign n1894 = ~n1890 & n1893 ;
  assign n1895 = x107 & ~x235 ;
  assign n1896 = ~x108 & ~n1895 ;
  assign n1897 = ~x109 & n1896 ;
  assign n1898 = ~n1894 & n1897 ;
  assign n1899 = ~x109 & x236 ;
  assign n1900 = ~x237 & ~x238 ;
  assign n1901 = ~n1899 & n1900 ;
  assign n1902 = ~n1898 & n1901 ;
  assign n1903 = x110 & ~x238 ;
  assign n1904 = ~x111 & ~n1903 ;
  assign n1905 = ~x112 & n1904 ;
  assign n1906 = ~n1902 & n1905 ;
  assign n1907 = ~x112 & x239 ;
  assign n1908 = ~x240 & ~x241 ;
  assign n1909 = ~n1907 & n1908 ;
  assign n1910 = ~n1906 & n1909 ;
  assign n1911 = x113 & ~x241 ;
  assign n1912 = ~x114 & ~n1911 ;
  assign n1913 = ~x115 & n1912 ;
  assign n1914 = ~n1910 & n1913 ;
  assign n1915 = ~x115 & x242 ;
  assign n1916 = ~x243 & ~x244 ;
  assign n1917 = ~n1915 & n1916 ;
  assign n1918 = ~n1914 & n1917 ;
  assign n1919 = x116 & ~x244 ;
  assign n1920 = ~x117 & ~n1919 ;
  assign n1921 = ~x118 & n1920 ;
  assign n1922 = ~n1918 & n1921 ;
  assign n1923 = ~x118 & x245 ;
  assign n1924 = ~x246 & ~x247 ;
  assign n1925 = ~n1923 & n1924 ;
  assign n1926 = ~n1922 & n1925 ;
  assign n1927 = x119 & ~x247 ;
  assign n1928 = ~x120 & ~n1927 ;
  assign n1929 = ~x121 & n1928 ;
  assign n1930 = ~n1926 & n1929 ;
  assign n1931 = ~x121 & x248 ;
  assign n1932 = ~x249 & ~x250 ;
  assign n1933 = ~n1931 & n1932 ;
  assign n1934 = ~n1930 & n1933 ;
  assign n1935 = x122 & ~x250 ;
  assign n1936 = ~x123 & ~n1935 ;
  assign n1937 = ~x124 & n1936 ;
  assign n1938 = ~n1934 & n1937 ;
  assign n1939 = ~x124 & x251 ;
  assign n1940 = ~x252 & ~x253 ;
  assign n1941 = ~n1939 & n1940 ;
  assign n1942 = ~n1938 & n1941 ;
  assign n1943 = x125 & ~x253 ;
  assign n1944 = ~x126 & ~n1943 ;
  assign n1945 = ~x127 & n1944 ;
  assign n1946 = ~n1942 & n1945 ;
  assign n1947 = ~x127 & x254 ;
  assign n1948 = ~x128 & ~x255 ;
  assign n1949 = ~n1947 & n1948 ;
  assign n1950 = ~n1946 & n1949 ;
  assign n1951 = x0 & ~x128 ;
  assign n1952 = ~x1 & ~n1951 ;
  assign n1953 = ~x2 & n1952 ;
  assign n1954 = ~n1950 & n1953 ;
  assign n1955 = ~x2 & x129 ;
  assign n1956 = x130 & ~n1955 ;
  assign n1957 = ~n1954 & n1956 ;
  assign n2296 = n1957 & x258 ;
  assign n1958 = x132 & x133 ;
  assign n1959 = ~n601 & n1958 ;
  assign n1960 = ~x5 & x133 ;
  assign n1961 = x6 & ~n1960 ;
  assign n1962 = x7 & n1961 ;
  assign n1963 = ~n1959 & n1962 ;
  assign n1964 = x7 & ~x134 ;
  assign n1965 = x135 & x136 ;
  assign n1966 = ~n1964 & n1965 ;
  assign n1967 = ~n1963 & n1966 ;
  assign n1968 = ~x8 & x136 ;
  assign n1969 = x9 & ~n1968 ;
  assign n1970 = x10 & n1969 ;
  assign n1971 = ~n1967 & n1970 ;
  assign n1972 = x10 & ~x137 ;
  assign n1973 = x138 & x139 ;
  assign n1974 = ~n1972 & n1973 ;
  assign n1975 = ~n1971 & n1974 ;
  assign n1976 = ~x11 & x139 ;
  assign n1977 = x12 & ~n1976 ;
  assign n1978 = x13 & n1977 ;
  assign n1979 = ~n1975 & n1978 ;
  assign n1980 = x13 & ~x140 ;
  assign n1981 = x141 & x142 ;
  assign n1982 = ~n1980 & n1981 ;
  assign n1983 = ~n1979 & n1982 ;
  assign n1984 = ~x14 & x142 ;
  assign n1985 = x15 & ~n1984 ;
  assign n1986 = x16 & n1985 ;
  assign n1987 = ~n1983 & n1986 ;
  assign n1988 = x16 & ~x143 ;
  assign n1989 = x144 & x145 ;
  assign n1990 = ~n1988 & n1989 ;
  assign n1991 = ~n1987 & n1990 ;
  assign n1992 = ~x17 & x145 ;
  assign n1993 = x18 & ~n1992 ;
  assign n1994 = x19 & n1993 ;
  assign n1995 = ~n1991 & n1994 ;
  assign n1996 = x19 & ~x146 ;
  assign n1997 = x147 & x148 ;
  assign n1998 = ~n1996 & n1997 ;
  assign n1999 = ~n1995 & n1998 ;
  assign n2000 = ~x20 & x148 ;
  assign n2001 = x21 & ~n2000 ;
  assign n2002 = x22 & n2001 ;
  assign n2003 = ~n1999 & n2002 ;
  assign n2004 = x22 & ~x149 ;
  assign n2005 = x150 & x151 ;
  assign n2006 = ~n2004 & n2005 ;
  assign n2007 = ~n2003 & n2006 ;
  assign n2008 = ~x23 & x151 ;
  assign n2009 = x24 & ~n2008 ;
  assign n2010 = x25 & n2009 ;
  assign n2011 = ~n2007 & n2010 ;
  assign n2012 = x25 & ~x152 ;
  assign n2013 = x153 & x154 ;
  assign n2014 = ~n2012 & n2013 ;
  assign n2015 = ~n2011 & n2014 ;
  assign n2016 = ~x26 & x154 ;
  assign n2017 = x27 & ~n2016 ;
  assign n2018 = x28 & n2017 ;
  assign n2019 = ~n2015 & n2018 ;
  assign n2020 = x28 & ~x155 ;
  assign n2021 = x156 & x157 ;
  assign n2022 = ~n2020 & n2021 ;
  assign n2023 = ~n2019 & n2022 ;
  assign n2024 = ~x29 & x157 ;
  assign n2025 = x30 & ~n2024 ;
  assign n2026 = x31 & n2025 ;
  assign n2027 = ~n2023 & n2026 ;
  assign n2028 = x31 & ~x158 ;
  assign n2029 = x159 & x160 ;
  assign n2030 = ~n2028 & n2029 ;
  assign n2031 = ~n2027 & n2030 ;
  assign n2032 = ~x32 & x160 ;
  assign n2033 = x33 & ~n2032 ;
  assign n2034 = x34 & n2033 ;
  assign n2035 = ~n2031 & n2034 ;
  assign n2036 = x34 & ~x161 ;
  assign n2037 = x162 & x163 ;
  assign n2038 = ~n2036 & n2037 ;
  assign n2039 = ~n2035 & n2038 ;
  assign n2040 = ~x35 & x163 ;
  assign n2041 = x36 & ~n2040 ;
  assign n2042 = x37 & n2041 ;
  assign n2043 = ~n2039 & n2042 ;
  assign n2044 = x37 & ~x164 ;
  assign n2045 = x165 & x166 ;
  assign n2046 = ~n2044 & n2045 ;
  assign n2047 = ~n2043 & n2046 ;
  assign n2048 = ~x38 & x166 ;
  assign n2049 = x39 & ~n2048 ;
  assign n2050 = x40 & n2049 ;
  assign n2051 = ~n2047 & n2050 ;
  assign n2052 = x40 & ~x167 ;
  assign n2053 = x168 & x169 ;
  assign n2054 = ~n2052 & n2053 ;
  assign n2055 = ~n2051 & n2054 ;
  assign n2056 = ~x41 & x169 ;
  assign n2057 = x42 & ~n2056 ;
  assign n2058 = x43 & n2057 ;
  assign n2059 = ~n2055 & n2058 ;
  assign n2060 = x43 & ~x170 ;
  assign n2061 = x171 & x172 ;
  assign n2062 = ~n2060 & n2061 ;
  assign n2063 = ~n2059 & n2062 ;
  assign n2064 = ~x44 & x172 ;
  assign n2065 = x45 & ~n2064 ;
  assign n2066 = x46 & n2065 ;
  assign n2067 = ~n2063 & n2066 ;
  assign n2068 = x46 & ~x173 ;
  assign n2069 = x174 & x175 ;
  assign n2070 = ~n2068 & n2069 ;
  assign n2071 = ~n2067 & n2070 ;
  assign n2072 = ~x47 & x175 ;
  assign n2073 = x48 & ~n2072 ;
  assign n2074 = x49 & n2073 ;
  assign n2075 = ~n2071 & n2074 ;
  assign n2076 = x49 & ~x176 ;
  assign n2077 = x177 & x178 ;
  assign n2078 = ~n2076 & n2077 ;
  assign n2079 = ~n2075 & n2078 ;
  assign n2080 = ~x50 & x178 ;
  assign n2081 = x51 & ~n2080 ;
  assign n2082 = x52 & n2081 ;
  assign n2083 = ~n2079 & n2082 ;
  assign n2084 = x52 & ~x179 ;
  assign n2085 = x180 & x181 ;
  assign n2086 = ~n2084 & n2085 ;
  assign n2087 = ~n2083 & n2086 ;
  assign n2088 = ~x53 & x181 ;
  assign n2089 = x54 & ~n2088 ;
  assign n2090 = x55 & n2089 ;
  assign n2091 = ~n2087 & n2090 ;
  assign n2092 = x55 & ~x182 ;
  assign n2093 = x183 & x184 ;
  assign n2094 = ~n2092 & n2093 ;
  assign n2095 = ~n2091 & n2094 ;
  assign n2096 = ~x56 & x184 ;
  assign n2097 = x57 & ~n2096 ;
  assign n2098 = x58 & n2097 ;
  assign n2099 = ~n2095 & n2098 ;
  assign n2100 = x58 & ~x185 ;
  assign n2101 = x186 & x187 ;
  assign n2102 = ~n2100 & n2101 ;
  assign n2103 = ~n2099 & n2102 ;
  assign n2104 = ~x59 & x187 ;
  assign n2105 = x60 & ~n2104 ;
  assign n2106 = x61 & n2105 ;
  assign n2107 = ~n2103 & n2106 ;
  assign n2108 = x61 & ~x188 ;
  assign n2109 = x189 & x190 ;
  assign n2110 = ~n2108 & n2109 ;
  assign n2111 = ~n2107 & n2110 ;
  assign n2112 = ~x62 & x190 ;
  assign n2113 = x63 & ~n2112 ;
  assign n2114 = x64 & n2113 ;
  assign n2115 = ~n2111 & n2114 ;
  assign n2116 = x64 & ~x191 ;
  assign n2117 = x192 & x193 ;
  assign n2118 = ~n2116 & n2117 ;
  assign n2119 = ~n2115 & n2118 ;
  assign n2120 = ~x65 & x193 ;
  assign n2121 = x66 & ~n2120 ;
  assign n2122 = x67 & n2121 ;
  assign n2123 = ~n2119 & n2122 ;
  assign n2124 = x67 & ~x194 ;
  assign n2125 = x195 & x196 ;
  assign n2126 = ~n2124 & n2125 ;
  assign n2127 = ~n2123 & n2126 ;
  assign n2128 = ~x68 & x196 ;
  assign n2129 = x69 & ~n2128 ;
  assign n2130 = x70 & n2129 ;
  assign n2131 = ~n2127 & n2130 ;
  assign n2132 = x70 & ~x197 ;
  assign n2133 = x198 & x199 ;
  assign n2134 = ~n2132 & n2133 ;
  assign n2135 = ~n2131 & n2134 ;
  assign n2136 = ~x71 & x199 ;
  assign n2137 = x72 & ~n2136 ;
  assign n2138 = x73 & n2137 ;
  assign n2139 = ~n2135 & n2138 ;
  assign n2140 = x73 & ~x200 ;
  assign n2141 = x201 & x202 ;
  assign n2142 = ~n2140 & n2141 ;
  assign n2143 = ~n2139 & n2142 ;
  assign n2144 = ~x74 & x202 ;
  assign n2145 = x75 & ~n2144 ;
  assign n2146 = x76 & n2145 ;
  assign n2147 = ~n2143 & n2146 ;
  assign n2148 = x76 & ~x203 ;
  assign n2149 = x204 & x205 ;
  assign n2150 = ~n2148 & n2149 ;
  assign n2151 = ~n2147 & n2150 ;
  assign n2152 = ~x77 & x205 ;
  assign n2153 = x78 & ~n2152 ;
  assign n2154 = x79 & n2153 ;
  assign n2155 = ~n2151 & n2154 ;
  assign n2156 = x79 & ~x206 ;
  assign n2157 = x207 & x208 ;
  assign n2158 = ~n2156 & n2157 ;
  assign n2159 = ~n2155 & n2158 ;
  assign n2160 = ~x80 & x208 ;
  assign n2161 = x81 & ~n2160 ;
  assign n2162 = x82 & n2161 ;
  assign n2163 = ~n2159 & n2162 ;
  assign n2164 = x82 & ~x209 ;
  assign n2165 = x210 & x211 ;
  assign n2166 = ~n2164 & n2165 ;
  assign n2167 = ~n2163 & n2166 ;
  assign n2168 = ~x83 & x211 ;
  assign n2169 = x84 & ~n2168 ;
  assign n2170 = x85 & n2169 ;
  assign n2171 = ~n2167 & n2170 ;
  assign n2172 = x85 & ~x212 ;
  assign n2173 = x213 & x214 ;
  assign n2174 = ~n2172 & n2173 ;
  assign n2175 = ~n2171 & n2174 ;
  assign n2176 = ~x86 & x214 ;
  assign n2177 = x87 & ~n2176 ;
  assign n2178 = x88 & n2177 ;
  assign n2179 = ~n2175 & n2178 ;
  assign n2180 = x88 & ~x215 ;
  assign n2181 = x216 & x217 ;
  assign n2182 = ~n2180 & n2181 ;
  assign n2183 = ~n2179 & n2182 ;
  assign n2184 = ~x89 & x217 ;
  assign n2185 = x90 & ~n2184 ;
  assign n2186 = x91 & n2185 ;
  assign n2187 = ~n2183 & n2186 ;
  assign n2188 = x91 & ~x218 ;
  assign n2189 = x219 & x220 ;
  assign n2190 = ~n2188 & n2189 ;
  assign n2191 = ~n2187 & n2190 ;
  assign n2192 = ~x92 & x220 ;
  assign n2193 = x93 & ~n2192 ;
  assign n2194 = x94 & n2193 ;
  assign n2195 = ~n2191 & n2194 ;
  assign n2196 = x94 & ~x221 ;
  assign n2197 = x222 & x223 ;
  assign n2198 = ~n2196 & n2197 ;
  assign n2199 = ~n2195 & n2198 ;
  assign n2200 = ~x95 & x223 ;
  assign n2201 = x96 & ~n2200 ;
  assign n2202 = x97 & n2201 ;
  assign n2203 = ~n2199 & n2202 ;
  assign n2204 = x97 & ~x224 ;
  assign n2205 = x225 & x226 ;
  assign n2206 = ~n2204 & n2205 ;
  assign n2207 = ~n2203 & n2206 ;
  assign n2208 = ~x98 & x226 ;
  assign n2209 = x99 & ~n2208 ;
  assign n2210 = x100 & n2209 ;
  assign n2211 = ~n2207 & n2210 ;
  assign n2212 = x100 & ~x227 ;
  assign n2213 = x228 & x229 ;
  assign n2214 = ~n2212 & n2213 ;
  assign n2215 = ~n2211 & n2214 ;
  assign n2216 = ~x101 & x229 ;
  assign n2217 = x102 & ~n2216 ;
  assign n2218 = x103 & n2217 ;
  assign n2219 = ~n2215 & n2218 ;
  assign n2220 = x103 & ~x230 ;
  assign n2221 = x231 & x232 ;
  assign n2222 = ~n2220 & n2221 ;
  assign n2223 = ~n2219 & n2222 ;
  assign n2224 = ~x104 & x232 ;
  assign n2225 = x105 & ~n2224 ;
  assign n2226 = x106 & n2225 ;
  assign n2227 = ~n2223 & n2226 ;
  assign n2228 = x106 & ~x233 ;
  assign n2229 = x234 & x235 ;
  assign n2230 = ~n2228 & n2229 ;
  assign n2231 = ~n2227 & n2230 ;
  assign n2232 = ~x107 & x235 ;
  assign n2233 = x108 & ~n2232 ;
  assign n2234 = x109 & n2233 ;
  assign n2235 = ~n2231 & n2234 ;
  assign n2236 = x109 & ~x236 ;
  assign n2237 = x237 & x238 ;
  assign n2238 = ~n2236 & n2237 ;
  assign n2239 = ~n2235 & n2238 ;
  assign n2240 = ~x110 & x238 ;
  assign n2241 = x111 & ~n2240 ;
  assign n2242 = x112 & n2241 ;
  assign n2243 = ~n2239 & n2242 ;
  assign n2244 = x112 & ~x239 ;
  assign n2245 = x240 & x241 ;
  assign n2246 = ~n2244 & n2245 ;
  assign n2247 = ~n2243 & n2246 ;
  assign n2248 = ~x113 & x241 ;
  assign n2249 = x114 & ~n2248 ;
  assign n2250 = x115 & n2249 ;
  assign n2251 = ~n2247 & n2250 ;
  assign n2252 = x115 & ~x242 ;
  assign n2253 = x243 & x244 ;
  assign n2254 = ~n2252 & n2253 ;
  assign n2255 = ~n2251 & n2254 ;
  assign n2256 = ~x116 & x244 ;
  assign n2257 = x117 & ~n2256 ;
  assign n2258 = x118 & n2257 ;
  assign n2259 = ~n2255 & n2258 ;
  assign n2260 = x118 & ~x245 ;
  assign n2261 = x246 & x247 ;
  assign n2262 = ~n2260 & n2261 ;
  assign n2263 = ~n2259 & n2262 ;
  assign n2264 = ~x119 & x247 ;
  assign n2265 = x120 & ~n2264 ;
  assign n2266 = x121 & n2265 ;
  assign n2267 = ~n2263 & n2266 ;
  assign n2268 = x121 & ~x248 ;
  assign n2269 = x249 & x250 ;
  assign n2270 = ~n2268 & n2269 ;
  assign n2271 = ~n2267 & n2270 ;
  assign n2272 = ~x122 & x250 ;
  assign n2273 = x123 & ~n2272 ;
  assign n2274 = x124 & n2273 ;
  assign n2275 = ~n2271 & n2274 ;
  assign n2276 = x124 & ~x251 ;
  assign n2277 = x252 & x253 ;
  assign n2278 = ~n2276 & n2277 ;
  assign n2279 = ~n2275 & n2278 ;
  assign n2280 = ~x125 & x253 ;
  assign n2281 = x126 & ~n2280 ;
  assign n2282 = x127 & n2281 ;
  assign n2283 = ~n2279 & n2282 ;
  assign n2284 = x127 & ~x254 ;
  assign n2285 = x128 & x255 ;
  assign n2286 = ~n2284 & n2285 ;
  assign n2287 = ~n2283 & n2286 ;
  assign n2288 = ~x0 & x128 ;
  assign n2289 = x1 & ~n2288 ;
  assign n2290 = x2 & n2289 ;
  assign n2291 = ~n2287 & n2290 ;
  assign n2292 = x2 & ~x129 ;
  assign n2293 = ~x130 & ~n2292 ;
  assign n2294 = ~n2291 & n2293 ;
  assign n2297 = ~n2294 & ~x258 ;
  assign n2298 = ~n2296 & ~n2297 ;
  assign n2299 = n266 & ~n944 ;
  assign n2300 = n271 & ~n2299 ;
  assign n2301 = n275 & ~n2300 ;
  assign n2302 = n279 & ~n2301 ;
  assign n2303 = n283 & ~n2302 ;
  assign n2304 = n287 & ~n2303 ;
  assign n2305 = n291 & ~n2304 ;
  assign n2306 = n295 & ~n2305 ;
  assign n2307 = n299 & ~n2306 ;
  assign n2308 = n303 & ~n2307 ;
  assign n2309 = n307 & ~n2308 ;
  assign n2310 = n311 & ~n2309 ;
  assign n2311 = n315 & ~n2310 ;
  assign n2312 = n319 & ~n2311 ;
  assign n2313 = n323 & ~n2312 ;
  assign n2314 = n327 & ~n2313 ;
  assign n2315 = n331 & ~n2314 ;
  assign n2316 = n335 & ~n2315 ;
  assign n2317 = n339 & ~n2316 ;
  assign n2318 = n343 & ~n2317 ;
  assign n2319 = n347 & ~n2318 ;
  assign n2320 = n351 & ~n2319 ;
  assign n2321 = n355 & ~n2320 ;
  assign n2322 = n359 & ~n2321 ;
  assign n2323 = n363 & ~n2322 ;
  assign n2324 = n367 & ~n2323 ;
  assign n2325 = n371 & ~n2324 ;
  assign n2326 = n375 & ~n2325 ;
  assign n2327 = n379 & ~n2326 ;
  assign n2328 = n383 & ~n2327 ;
  assign n2329 = n387 & ~n2328 ;
  assign n2330 = n391 & ~n2329 ;
  assign n2331 = n395 & ~n2330 ;
  assign n2332 = n399 & ~n2331 ;
  assign n2333 = n403 & ~n2332 ;
  assign n2334 = n407 & ~n2333 ;
  assign n2335 = n411 & ~n2334 ;
  assign n2336 = n415 & ~n2335 ;
  assign n2337 = n419 & ~n2336 ;
  assign n2338 = n423 & ~n2337 ;
  assign n2339 = n427 & ~n2338 ;
  assign n2340 = n431 & ~n2339 ;
  assign n2341 = n435 & ~n2340 ;
  assign n2342 = n439 & ~n2341 ;
  assign n2343 = n443 & ~n2342 ;
  assign n2344 = n447 & ~n2343 ;
  assign n2345 = n451 & ~n2344 ;
  assign n2346 = n455 & ~n2345 ;
  assign n2347 = n459 & ~n2346 ;
  assign n2348 = n463 & ~n2347 ;
  assign n2349 = n467 & ~n2348 ;
  assign n2350 = n471 & ~n2349 ;
  assign n2351 = n475 & ~n2350 ;
  assign n2352 = n479 & ~n2351 ;
  assign n2353 = n483 & ~n2352 ;
  assign n2354 = n487 & ~n2353 ;
  assign n2355 = n491 & ~n2354 ;
  assign n2356 = n495 & ~n2355 ;
  assign n2357 = n499 & ~n2356 ;
  assign n2358 = n503 & ~n2357 ;
  assign n2359 = n507 & ~n2358 ;
  assign n2360 = n511 & ~n2359 ;
  assign n2361 = n515 & ~n2360 ;
  assign n2362 = n519 & ~n2361 ;
  assign n2363 = n523 & ~n2362 ;
  assign n2364 = n527 & ~n2363 ;
  assign n2365 = n531 & ~n2364 ;
  assign n2366 = n535 & ~n2365 ;
  assign n2367 = n539 & ~n2366 ;
  assign n2368 = n543 & ~n2367 ;
  assign n2369 = n547 & ~n2368 ;
  assign n2370 = n551 & ~n2369 ;
  assign n2371 = n555 & ~n2370 ;
  assign n2372 = n559 & ~n2371 ;
  assign n2373 = n563 & ~n2372 ;
  assign n2374 = n567 & ~n2373 ;
  assign n2375 = n571 & ~n2374 ;
  assign n2376 = n575 & ~n2375 ;
  assign n2377 = n579 & ~n2376 ;
  assign n2378 = n583 & ~n2377 ;
  assign n2379 = n587 & ~n2378 ;
  assign n2380 = n591 & ~n2379 ;
  assign n2381 = ~x128 & ~x129 ;
  assign n2382 = ~n593 & n2381 ;
  assign n2383 = ~n2380 & n2382 ;
  assign n2384 = ~x3 & n258 ;
  assign n2385 = ~n2383 & n2384 ;
  assign n2386 = ~x3 & x130 ;
  assign n2387 = x131 & ~n2386 ;
  assign n2388 = ~n2385 & n2387 ;
  assign n2480 = n2388 & x259 ;
  assign n2389 = n605 & ~n1283 ;
  assign n2390 = n610 & ~n2389 ;
  assign n2391 = n614 & ~n2390 ;
  assign n2392 = n618 & ~n2391 ;
  assign n2393 = n622 & ~n2392 ;
  assign n2394 = n626 & ~n2393 ;
  assign n2395 = n630 & ~n2394 ;
  assign n2396 = n634 & ~n2395 ;
  assign n2397 = n638 & ~n2396 ;
  assign n2398 = n642 & ~n2397 ;
  assign n2399 = n646 & ~n2398 ;
  assign n2400 = n650 & ~n2399 ;
  assign n2401 = n654 & ~n2400 ;
  assign n2402 = n658 & ~n2401 ;
  assign n2403 = n662 & ~n2402 ;
  assign n2404 = n666 & ~n2403 ;
  assign n2405 = n670 & ~n2404 ;
  assign n2406 = n674 & ~n2405 ;
  assign n2407 = n678 & ~n2406 ;
  assign n2408 = n682 & ~n2407 ;
  assign n2409 = n686 & ~n2408 ;
  assign n2410 = n690 & ~n2409 ;
  assign n2411 = n694 & ~n2410 ;
  assign n2412 = n698 & ~n2411 ;
  assign n2413 = n702 & ~n2412 ;
  assign n2414 = n706 & ~n2413 ;
  assign n2415 = n710 & ~n2414 ;
  assign n2416 = n714 & ~n2415 ;
  assign n2417 = n718 & ~n2416 ;
  assign n2418 = n722 & ~n2417 ;
  assign n2419 = n726 & ~n2418 ;
  assign n2420 = n730 & ~n2419 ;
  assign n2421 = n734 & ~n2420 ;
  assign n2422 = n738 & ~n2421 ;
  assign n2423 = n742 & ~n2422 ;
  assign n2424 = n746 & ~n2423 ;
  assign n2425 = n750 & ~n2424 ;
  assign n2426 = n754 & ~n2425 ;
  assign n2427 = n758 & ~n2426 ;
  assign n2428 = n762 & ~n2427 ;
  assign n2429 = n766 & ~n2428 ;
  assign n2430 = n770 & ~n2429 ;
  assign n2431 = n774 & ~n2430 ;
  assign n2432 = n778 & ~n2431 ;
  assign n2433 = n782 & ~n2432 ;
  assign n2434 = n786 & ~n2433 ;
  assign n2435 = n790 & ~n2434 ;
  assign n2436 = n794 & ~n2435 ;
  assign n2437 = n798 & ~n2436 ;
  assign n2438 = n802 & ~n2437 ;
  assign n2439 = n806 & ~n2438 ;
  assign n2440 = n810 & ~n2439 ;
  assign n2441 = n814 & ~n2440 ;
  assign n2442 = n818 & ~n2441 ;
  assign n2443 = n822 & ~n2442 ;
  assign n2444 = n826 & ~n2443 ;
  assign n2445 = n830 & ~n2444 ;
  assign n2446 = n834 & ~n2445 ;
  assign n2447 = n838 & ~n2446 ;
  assign n2448 = n842 & ~n2447 ;
  assign n2449 = n846 & ~n2448 ;
  assign n2450 = n850 & ~n2449 ;
  assign n2451 = n854 & ~n2450 ;
  assign n2452 = n858 & ~n2451 ;
  assign n2453 = n862 & ~n2452 ;
  assign n2454 = n866 & ~n2453 ;
  assign n2455 = n870 & ~n2454 ;
  assign n2456 = n874 & ~n2455 ;
  assign n2457 = n878 & ~n2456 ;
  assign n2458 = n882 & ~n2457 ;
  assign n2459 = n886 & ~n2458 ;
  assign n2460 = n890 & ~n2459 ;
  assign n2461 = n894 & ~n2460 ;
  assign n2462 = n898 & ~n2461 ;
  assign n2463 = n902 & ~n2462 ;
  assign n2464 = n906 & ~n2463 ;
  assign n2465 = n910 & ~n2464 ;
  assign n2466 = n914 & ~n2465 ;
  assign n2467 = n918 & ~n2466 ;
  assign n2468 = n922 & ~n2467 ;
  assign n2469 = n926 & ~n2468 ;
  assign n2470 = n930 & ~n2469 ;
  assign n2471 = x128 & x129 ;
  assign n2472 = ~n932 & n2471 ;
  assign n2473 = ~n2470 & n2472 ;
  assign n2474 = x3 & n597 ;
  assign n2475 = ~n2473 & n2474 ;
  assign n2476 = x3 & ~x130 ;
  assign n2477 = ~x131 & ~n2476 ;
  assign n2478 = ~n2475 & n2477 ;
  assign n2481 = ~n2478 & ~x259 ;
  assign n2482 = ~n2480 & ~n2481 ;
  assign n2483 = n948 & ~n1624 ;
  assign n2484 = n953 & ~n2483 ;
  assign n2485 = n957 & ~n2484 ;
  assign n2486 = n961 & ~n2485 ;
  assign n2487 = n965 & ~n2486 ;
  assign n2488 = n969 & ~n2487 ;
  assign n2489 = n973 & ~n2488 ;
  assign n2490 = n977 & ~n2489 ;
  assign n2491 = n981 & ~n2490 ;
  assign n2492 = n985 & ~n2491 ;
  assign n2493 = n989 & ~n2492 ;
  assign n2494 = n993 & ~n2493 ;
  assign n2495 = n997 & ~n2494 ;
  assign n2496 = n1001 & ~n2495 ;
  assign n2497 = n1005 & ~n2496 ;
  assign n2498 = n1009 & ~n2497 ;
  assign n2499 = n1013 & ~n2498 ;
  assign n2500 = n1017 & ~n2499 ;
  assign n2501 = n1021 & ~n2500 ;
  assign n2502 = n1025 & ~n2501 ;
  assign n2503 = n1029 & ~n2502 ;
  assign n2504 = n1033 & ~n2503 ;
  assign n2505 = n1037 & ~n2504 ;
  assign n2506 = n1041 & ~n2505 ;
  assign n2507 = n1045 & ~n2506 ;
  assign n2508 = n1049 & ~n2507 ;
  assign n2509 = n1053 & ~n2508 ;
  assign n2510 = n1057 & ~n2509 ;
  assign n2511 = n1061 & ~n2510 ;
  assign n2512 = n1065 & ~n2511 ;
  assign n2513 = n1069 & ~n2512 ;
  assign n2514 = n1073 & ~n2513 ;
  assign n2515 = n1077 & ~n2514 ;
  assign n2516 = n1081 & ~n2515 ;
  assign n2517 = n1085 & ~n2516 ;
  assign n2518 = n1089 & ~n2517 ;
  assign n2519 = n1093 & ~n2518 ;
  assign n2520 = n1097 & ~n2519 ;
  assign n2521 = n1101 & ~n2520 ;
  assign n2522 = n1105 & ~n2521 ;
  assign n2523 = n1109 & ~n2522 ;
  assign n2524 = n1113 & ~n2523 ;
  assign n2525 = n1117 & ~n2524 ;
  assign n2526 = n1121 & ~n2525 ;
  assign n2527 = n1125 & ~n2526 ;
  assign n2528 = n1129 & ~n2527 ;
  assign n2529 = n1133 & ~n2528 ;
  assign n2530 = n1137 & ~n2529 ;
  assign n2531 = n1141 & ~n2530 ;
  assign n2532 = n1145 & ~n2531 ;
  assign n2533 = n1149 & ~n2532 ;
  assign n2534 = n1153 & ~n2533 ;
  assign n2535 = n1157 & ~n2534 ;
  assign n2536 = n1161 & ~n2535 ;
  assign n2537 = n1165 & ~n2536 ;
  assign n2538 = n1169 & ~n2537 ;
  assign n2539 = n1173 & ~n2538 ;
  assign n2540 = n1177 & ~n2539 ;
  assign n2541 = n1181 & ~n2540 ;
  assign n2542 = n1185 & ~n2541 ;
  assign n2543 = n1189 & ~n2542 ;
  assign n2544 = n1193 & ~n2543 ;
  assign n2545 = n1197 & ~n2544 ;
  assign n2546 = n1201 & ~n2545 ;
  assign n2547 = n1205 & ~n2546 ;
  assign n2548 = n1209 & ~n2547 ;
  assign n2549 = n1213 & ~n2548 ;
  assign n2550 = n1217 & ~n2549 ;
  assign n2551 = n1221 & ~n2550 ;
  assign n2552 = n1225 & ~n2551 ;
  assign n2553 = n1229 & ~n2552 ;
  assign n2554 = n1233 & ~n2553 ;
  assign n2555 = n1237 & ~n2554 ;
  assign n2556 = n1241 & ~n2555 ;
  assign n2557 = n1245 & ~n2556 ;
  assign n2558 = n1249 & ~n2557 ;
  assign n2559 = n1253 & ~n2558 ;
  assign n2560 = n1257 & ~n2559 ;
  assign n2561 = n1261 & ~n2560 ;
  assign n2562 = n1265 & ~n2561 ;
  assign n2563 = n1269 & ~n2562 ;
  assign n2564 = n1273 & ~n2563 ;
  assign n2565 = ~x129 & ~x130 ;
  assign n2566 = ~n1275 & n2565 ;
  assign n2567 = ~n2564 & n2566 ;
  assign n2568 = ~x4 & n940 ;
  assign n2569 = ~n2567 & n2568 ;
  assign n2570 = ~x4 & x131 ;
  assign n2571 = x132 & ~n2570 ;
  assign n2572 = ~n2569 & n2571 ;
  assign n2664 = n2572 & x260 ;
  assign n2573 = n1287 & ~n1961 ;
  assign n2574 = n1292 & ~n2573 ;
  assign n2575 = n1296 & ~n2574 ;
  assign n2576 = n1300 & ~n2575 ;
  assign n2577 = n1304 & ~n2576 ;
  assign n2578 = n1308 & ~n2577 ;
  assign n2579 = n1312 & ~n2578 ;
  assign n2580 = n1316 & ~n2579 ;
  assign n2581 = n1320 & ~n2580 ;
  assign n2582 = n1324 & ~n2581 ;
  assign n2583 = n1328 & ~n2582 ;
  assign n2584 = n1332 & ~n2583 ;
  assign n2585 = n1336 & ~n2584 ;
  assign n2586 = n1340 & ~n2585 ;
  assign n2587 = n1344 & ~n2586 ;
  assign n2588 = n1348 & ~n2587 ;
  assign n2589 = n1352 & ~n2588 ;
  assign n2590 = n1356 & ~n2589 ;
  assign n2591 = n1360 & ~n2590 ;
  assign n2592 = n1364 & ~n2591 ;
  assign n2593 = n1368 & ~n2592 ;
  assign n2594 = n1372 & ~n2593 ;
  assign n2595 = n1376 & ~n2594 ;
  assign n2596 = n1380 & ~n2595 ;
  assign n2597 = n1384 & ~n2596 ;
  assign n2598 = n1388 & ~n2597 ;
  assign n2599 = n1392 & ~n2598 ;
  assign n2600 = n1396 & ~n2599 ;
  assign n2601 = n1400 & ~n2600 ;
  assign n2602 = n1404 & ~n2601 ;
  assign n2603 = n1408 & ~n2602 ;
  assign n2604 = n1412 & ~n2603 ;
  assign n2605 = n1416 & ~n2604 ;
  assign n2606 = n1420 & ~n2605 ;
  assign n2607 = n1424 & ~n2606 ;
  assign n2608 = n1428 & ~n2607 ;
  assign n2609 = n1432 & ~n2608 ;
  assign n2610 = n1436 & ~n2609 ;
  assign n2611 = n1440 & ~n2610 ;
  assign n2612 = n1444 & ~n2611 ;
  assign n2613 = n1448 & ~n2612 ;
  assign n2614 = n1452 & ~n2613 ;
  assign n2615 = n1456 & ~n2614 ;
  assign n2616 = n1460 & ~n2615 ;
  assign n2617 = n1464 & ~n2616 ;
  assign n2618 = n1468 & ~n2617 ;
  assign n2619 = n1472 & ~n2618 ;
  assign n2620 = n1476 & ~n2619 ;
  assign n2621 = n1480 & ~n2620 ;
  assign n2622 = n1484 & ~n2621 ;
  assign n2623 = n1488 & ~n2622 ;
  assign n2624 = n1492 & ~n2623 ;
  assign n2625 = n1496 & ~n2624 ;
  assign n2626 = n1500 & ~n2625 ;
  assign n2627 = n1504 & ~n2626 ;
  assign n2628 = n1508 & ~n2627 ;
  assign n2629 = n1512 & ~n2628 ;
  assign n2630 = n1516 & ~n2629 ;
  assign n2631 = n1520 & ~n2630 ;
  assign n2632 = n1524 & ~n2631 ;
  assign n2633 = n1528 & ~n2632 ;
  assign n2634 = n1532 & ~n2633 ;
  assign n2635 = n1536 & ~n2634 ;
  assign n2636 = n1540 & ~n2635 ;
  assign n2637 = n1544 & ~n2636 ;
  assign n2638 = n1548 & ~n2637 ;
  assign n2639 = n1552 & ~n2638 ;
  assign n2640 = n1556 & ~n2639 ;
  assign n2641 = n1560 & ~n2640 ;
  assign n2642 = n1564 & ~n2641 ;
  assign n2643 = n1568 & ~n2642 ;
  assign n2644 = n1572 & ~n2643 ;
  assign n2645 = n1576 & ~n2644 ;
  assign n2646 = n1580 & ~n2645 ;
  assign n2647 = n1584 & ~n2646 ;
  assign n2648 = n1588 & ~n2647 ;
  assign n2649 = n1592 & ~n2648 ;
  assign n2650 = n1596 & ~n2649 ;
  assign n2651 = n1600 & ~n2650 ;
  assign n2652 = n1604 & ~n2651 ;
  assign n2653 = n1608 & ~n2652 ;
  assign n2654 = n1612 & ~n2653 ;
  assign n2655 = x129 & x130 ;
  assign n2656 = ~n1614 & n2655 ;
  assign n2657 = ~n2654 & n2656 ;
  assign n2658 = x4 & n1279 ;
  assign n2659 = ~n2657 & n2658 ;
  assign n2660 = x4 & ~x131 ;
  assign n2661 = ~x132 & ~n2660 ;
  assign n2662 = ~n2659 & n2661 ;
  assign n2665 = ~n2662 & ~x260 ;
  assign n2666 = ~n2664 & ~n2665 ;
  assign n2667 = ~n270 & n1628 ;
  assign n2668 = n1633 & ~n2667 ;
  assign n2669 = n1637 & ~n2668 ;
  assign n2670 = n1641 & ~n2669 ;
  assign n2671 = n1645 & ~n2670 ;
  assign n2672 = n1649 & ~n2671 ;
  assign n2673 = n1653 & ~n2672 ;
  assign n2674 = n1657 & ~n2673 ;
  assign n2675 = n1661 & ~n2674 ;
  assign n2676 = n1665 & ~n2675 ;
  assign n2677 = n1669 & ~n2676 ;
  assign n2678 = n1673 & ~n2677 ;
  assign n2679 = n1677 & ~n2678 ;
  assign n2680 = n1681 & ~n2679 ;
  assign n2681 = n1685 & ~n2680 ;
  assign n2682 = n1689 & ~n2681 ;
  assign n2683 = n1693 & ~n2682 ;
  assign n2684 = n1697 & ~n2683 ;
  assign n2685 = n1701 & ~n2684 ;
  assign n2686 = n1705 & ~n2685 ;
  assign n2687 = n1709 & ~n2686 ;
  assign n2688 = n1713 & ~n2687 ;
  assign n2689 = n1717 & ~n2688 ;
  assign n2690 = n1721 & ~n2689 ;
  assign n2691 = n1725 & ~n2690 ;
  assign n2692 = n1729 & ~n2691 ;
  assign n2693 = n1733 & ~n2692 ;
  assign n2694 = n1737 & ~n2693 ;
  assign n2695 = n1741 & ~n2694 ;
  assign n2696 = n1745 & ~n2695 ;
  assign n2697 = n1749 & ~n2696 ;
  assign n2698 = n1753 & ~n2697 ;
  assign n2699 = n1757 & ~n2698 ;
  assign n2700 = n1761 & ~n2699 ;
  assign n2701 = n1765 & ~n2700 ;
  assign n2702 = n1769 & ~n2701 ;
  assign n2703 = n1773 & ~n2702 ;
  assign n2704 = n1777 & ~n2703 ;
  assign n2705 = n1781 & ~n2704 ;
  assign n2706 = n1785 & ~n2705 ;
  assign n2707 = n1789 & ~n2706 ;
  assign n2708 = n1793 & ~n2707 ;
  assign n2709 = n1797 & ~n2708 ;
  assign n2710 = n1801 & ~n2709 ;
  assign n2711 = n1805 & ~n2710 ;
  assign n2712 = n1809 & ~n2711 ;
  assign n2713 = n1813 & ~n2712 ;
  assign n2714 = n1817 & ~n2713 ;
  assign n2715 = n1821 & ~n2714 ;
  assign n2716 = n1825 & ~n2715 ;
  assign n2717 = n1829 & ~n2716 ;
  assign n2718 = n1833 & ~n2717 ;
  assign n2719 = n1837 & ~n2718 ;
  assign n2720 = n1841 & ~n2719 ;
  assign n2721 = n1845 & ~n2720 ;
  assign n2722 = n1849 & ~n2721 ;
  assign n2723 = n1853 & ~n2722 ;
  assign n2724 = n1857 & ~n2723 ;
  assign n2725 = n1861 & ~n2724 ;
  assign n2726 = n1865 & ~n2725 ;
  assign n2727 = n1869 & ~n2726 ;
  assign n2728 = n1873 & ~n2727 ;
  assign n2729 = n1877 & ~n2728 ;
  assign n2730 = n1881 & ~n2729 ;
  assign n2731 = n1885 & ~n2730 ;
  assign n2732 = n1889 & ~n2731 ;
  assign n2733 = n1893 & ~n2732 ;
  assign n2734 = n1897 & ~n2733 ;
  assign n2735 = n1901 & ~n2734 ;
  assign n2736 = n1905 & ~n2735 ;
  assign n2737 = n1909 & ~n2736 ;
  assign n2738 = n1913 & ~n2737 ;
  assign n2739 = n1917 & ~n2738 ;
  assign n2740 = n1921 & ~n2739 ;
  assign n2741 = n1925 & ~n2740 ;
  assign n2742 = n1929 & ~n2741 ;
  assign n2743 = n1933 & ~n2742 ;
  assign n2744 = n1937 & ~n2743 ;
  assign n2745 = n1941 & ~n2744 ;
  assign n2746 = n1945 & ~n2745 ;
  assign n2747 = n1949 & ~n2746 ;
  assign n2748 = n1953 & ~n2747 ;
  assign n2749 = n259 & ~n1955 ;
  assign n2750 = ~n2748 & n2749 ;
  assign n2751 = n263 & ~n2750 ;
  assign n2752 = x133 & ~n265 ;
  assign n2753 = ~n2751 & n2752 ;
  assign n2842 = n2753 & x261 ;
  assign n2754 = ~n609 & n1965 ;
  assign n2755 = n1970 & ~n2754 ;
  assign n2756 = n1974 & ~n2755 ;
  assign n2757 = n1978 & ~n2756 ;
  assign n2758 = n1982 & ~n2757 ;
  assign n2759 = n1986 & ~n2758 ;
  assign n2760 = n1990 & ~n2759 ;
  assign n2761 = n1994 & ~n2760 ;
  assign n2762 = n1998 & ~n2761 ;
  assign n2763 = n2002 & ~n2762 ;
  assign n2764 = n2006 & ~n2763 ;
  assign n2765 = n2010 & ~n2764 ;
  assign n2766 = n2014 & ~n2765 ;
  assign n2767 = n2018 & ~n2766 ;
  assign n2768 = n2022 & ~n2767 ;
  assign n2769 = n2026 & ~n2768 ;
  assign n2770 = n2030 & ~n2769 ;
  assign n2771 = n2034 & ~n2770 ;
  assign n2772 = n2038 & ~n2771 ;
  assign n2773 = n2042 & ~n2772 ;
  assign n2774 = n2046 & ~n2773 ;
  assign n2775 = n2050 & ~n2774 ;
  assign n2776 = n2054 & ~n2775 ;
  assign n2777 = n2058 & ~n2776 ;
  assign n2778 = n2062 & ~n2777 ;
  assign n2779 = n2066 & ~n2778 ;
  assign n2780 = n2070 & ~n2779 ;
  assign n2781 = n2074 & ~n2780 ;
  assign n2782 = n2078 & ~n2781 ;
  assign n2783 = n2082 & ~n2782 ;
  assign n2784 = n2086 & ~n2783 ;
  assign n2785 = n2090 & ~n2784 ;
  assign n2786 = n2094 & ~n2785 ;
  assign n2787 = n2098 & ~n2786 ;
  assign n2788 = n2102 & ~n2787 ;
  assign n2789 = n2106 & ~n2788 ;
  assign n2790 = n2110 & ~n2789 ;
  assign n2791 = n2114 & ~n2790 ;
  assign n2792 = n2118 & ~n2791 ;
  assign n2793 = n2122 & ~n2792 ;
  assign n2794 = n2126 & ~n2793 ;
  assign n2795 = n2130 & ~n2794 ;
  assign n2796 = n2134 & ~n2795 ;
  assign n2797 = n2138 & ~n2796 ;
  assign n2798 = n2142 & ~n2797 ;
  assign n2799 = n2146 & ~n2798 ;
  assign n2800 = n2150 & ~n2799 ;
  assign n2801 = n2154 & ~n2800 ;
  assign n2802 = n2158 & ~n2801 ;
  assign n2803 = n2162 & ~n2802 ;
  assign n2804 = n2166 & ~n2803 ;
  assign n2805 = n2170 & ~n2804 ;
  assign n2806 = n2174 & ~n2805 ;
  assign n2807 = n2178 & ~n2806 ;
  assign n2808 = n2182 & ~n2807 ;
  assign n2809 = n2186 & ~n2808 ;
  assign n2810 = n2190 & ~n2809 ;
  assign n2811 = n2194 & ~n2810 ;
  assign n2812 = n2198 & ~n2811 ;
  assign n2813 = n2202 & ~n2812 ;
  assign n2814 = n2206 & ~n2813 ;
  assign n2815 = n2210 & ~n2814 ;
  assign n2816 = n2214 & ~n2815 ;
  assign n2817 = n2218 & ~n2816 ;
  assign n2818 = n2222 & ~n2817 ;
  assign n2819 = n2226 & ~n2818 ;
  assign n2820 = n2230 & ~n2819 ;
  assign n2821 = n2234 & ~n2820 ;
  assign n2822 = n2238 & ~n2821 ;
  assign n2823 = n2242 & ~n2822 ;
  assign n2824 = n2246 & ~n2823 ;
  assign n2825 = n2250 & ~n2824 ;
  assign n2826 = n2254 & ~n2825 ;
  assign n2827 = n2258 & ~n2826 ;
  assign n2828 = n2262 & ~n2827 ;
  assign n2829 = n2266 & ~n2828 ;
  assign n2830 = n2270 & ~n2829 ;
  assign n2831 = n2274 & ~n2830 ;
  assign n2832 = n2278 & ~n2831 ;
  assign n2833 = n2282 & ~n2832 ;
  assign n2834 = n2286 & ~n2833 ;
  assign n2835 = n2290 & ~n2834 ;
  assign n2836 = n598 & ~n2292 ;
  assign n2837 = ~n2835 & n2836 ;
  assign n2838 = n602 & ~n2837 ;
  assign n2839 = ~x133 & ~n604 ;
  assign n2840 = ~n2838 & n2839 ;
  assign n2843 = ~n2840 & ~x261 ;
  assign n2844 = ~n2842 & ~n2843 ;
  assign n2845 = n274 & ~n952 ;
  assign n2846 = n279 & ~n2845 ;
  assign n2847 = n283 & ~n2846 ;
  assign n2848 = n287 & ~n2847 ;
  assign n2849 = n291 & ~n2848 ;
  assign n2850 = n295 & ~n2849 ;
  assign n2851 = n299 & ~n2850 ;
  assign n2852 = n303 & ~n2851 ;
  assign n2853 = n307 & ~n2852 ;
  assign n2854 = n311 & ~n2853 ;
  assign n2855 = n315 & ~n2854 ;
  assign n2856 = n319 & ~n2855 ;
  assign n2857 = n323 & ~n2856 ;
  assign n2858 = n327 & ~n2857 ;
  assign n2859 = n331 & ~n2858 ;
  assign n2860 = n335 & ~n2859 ;
  assign n2861 = n339 & ~n2860 ;
  assign n2862 = n343 & ~n2861 ;
  assign n2863 = n347 & ~n2862 ;
  assign n2864 = n351 & ~n2863 ;
  assign n2865 = n355 & ~n2864 ;
  assign n2866 = n359 & ~n2865 ;
  assign n2867 = n363 & ~n2866 ;
  assign n2868 = n367 & ~n2867 ;
  assign n2869 = n371 & ~n2868 ;
  assign n2870 = n375 & ~n2869 ;
  assign n2871 = n379 & ~n2870 ;
  assign n2872 = n383 & ~n2871 ;
  assign n2873 = n387 & ~n2872 ;
  assign n2874 = n391 & ~n2873 ;
  assign n2875 = n395 & ~n2874 ;
  assign n2876 = n399 & ~n2875 ;
  assign n2877 = n403 & ~n2876 ;
  assign n2878 = n407 & ~n2877 ;
  assign n2879 = n411 & ~n2878 ;
  assign n2880 = n415 & ~n2879 ;
  assign n2881 = n419 & ~n2880 ;
  assign n2882 = n423 & ~n2881 ;
  assign n2883 = n427 & ~n2882 ;
  assign n2884 = n431 & ~n2883 ;
  assign n2885 = n435 & ~n2884 ;
  assign n2886 = n439 & ~n2885 ;
  assign n2887 = n443 & ~n2886 ;
  assign n2888 = n447 & ~n2887 ;
  assign n2889 = n451 & ~n2888 ;
  assign n2890 = n455 & ~n2889 ;
  assign n2891 = n459 & ~n2890 ;
  assign n2892 = n463 & ~n2891 ;
  assign n2893 = n467 & ~n2892 ;
  assign n2894 = n471 & ~n2893 ;
  assign n2895 = n475 & ~n2894 ;
  assign n2896 = n479 & ~n2895 ;
  assign n2897 = n483 & ~n2896 ;
  assign n2898 = n487 & ~n2897 ;
  assign n2899 = n491 & ~n2898 ;
  assign n2900 = n495 & ~n2899 ;
  assign n2901 = n499 & ~n2900 ;
  assign n2902 = n503 & ~n2901 ;
  assign n2903 = n507 & ~n2902 ;
  assign n2904 = n511 & ~n2903 ;
  assign n2905 = n515 & ~n2904 ;
  assign n2906 = n519 & ~n2905 ;
  assign n2907 = n523 & ~n2906 ;
  assign n2908 = n527 & ~n2907 ;
  assign n2909 = n531 & ~n2908 ;
  assign n2910 = n535 & ~n2909 ;
  assign n2911 = n539 & ~n2910 ;
  assign n2912 = n543 & ~n2911 ;
  assign n2913 = n547 & ~n2912 ;
  assign n2914 = n551 & ~n2913 ;
  assign n2915 = n555 & ~n2914 ;
  assign n2916 = n559 & ~n2915 ;
  assign n2917 = n563 & ~n2916 ;
  assign n2918 = n567 & ~n2917 ;
  assign n2919 = n571 & ~n2918 ;
  assign n2920 = n575 & ~n2919 ;
  assign n2921 = n579 & ~n2920 ;
  assign n2922 = n583 & ~n2921 ;
  assign n2923 = n587 & ~n2922 ;
  assign n2924 = n591 & ~n2923 ;
  assign n2925 = n2382 & ~n2924 ;
  assign n2926 = n2384 & ~n2925 ;
  assign n2927 = n941 & ~n2386 ;
  assign n2928 = ~n2926 & n2927 ;
  assign n2929 = n945 & ~n2928 ;
  assign n2930 = x134 & ~n947 ;
  assign n2931 = ~n2929 & n2930 ;
  assign n3020 = n2931 & x262 ;
  assign n2932 = n613 & ~n1291 ;
  assign n2933 = n618 & ~n2932 ;
  assign n2934 = n622 & ~n2933 ;
  assign n2935 = n626 & ~n2934 ;
  assign n2936 = n630 & ~n2935 ;
  assign n2937 = n634 & ~n2936 ;
  assign n2938 = n638 & ~n2937 ;
  assign n2939 = n642 & ~n2938 ;
  assign n2940 = n646 & ~n2939 ;
  assign n2941 = n650 & ~n2940 ;
  assign n2942 = n654 & ~n2941 ;
  assign n2943 = n658 & ~n2942 ;
  assign n2944 = n662 & ~n2943 ;
  assign n2945 = n666 & ~n2944 ;
  assign n2946 = n670 & ~n2945 ;
  assign n2947 = n674 & ~n2946 ;
  assign n2948 = n678 & ~n2947 ;
  assign n2949 = n682 & ~n2948 ;
  assign n2950 = n686 & ~n2949 ;
  assign n2951 = n690 & ~n2950 ;
  assign n2952 = n694 & ~n2951 ;
  assign n2953 = n698 & ~n2952 ;
  assign n2954 = n702 & ~n2953 ;
  assign n2955 = n706 & ~n2954 ;
  assign n2956 = n710 & ~n2955 ;
  assign n2957 = n714 & ~n2956 ;
  assign n2958 = n718 & ~n2957 ;
  assign n2959 = n722 & ~n2958 ;
  assign n2960 = n726 & ~n2959 ;
  assign n2961 = n730 & ~n2960 ;
  assign n2962 = n734 & ~n2961 ;
  assign n2963 = n738 & ~n2962 ;
  assign n2964 = n742 & ~n2963 ;
  assign n2965 = n746 & ~n2964 ;
  assign n2966 = n750 & ~n2965 ;
  assign n2967 = n754 & ~n2966 ;
  assign n2968 = n758 & ~n2967 ;
  assign n2969 = n762 & ~n2968 ;
  assign n2970 = n766 & ~n2969 ;
  assign n2971 = n770 & ~n2970 ;
  assign n2972 = n774 & ~n2971 ;
  assign n2973 = n778 & ~n2972 ;
  assign n2974 = n782 & ~n2973 ;
  assign n2975 = n786 & ~n2974 ;
  assign n2976 = n790 & ~n2975 ;
  assign n2977 = n794 & ~n2976 ;
  assign n2978 = n798 & ~n2977 ;
  assign n2979 = n802 & ~n2978 ;
  assign n2980 = n806 & ~n2979 ;
  assign n2981 = n810 & ~n2980 ;
  assign n2982 = n814 & ~n2981 ;
  assign n2983 = n818 & ~n2982 ;
  assign n2984 = n822 & ~n2983 ;
  assign n2985 = n826 & ~n2984 ;
  assign n2986 = n830 & ~n2985 ;
  assign n2987 = n834 & ~n2986 ;
  assign n2988 = n838 & ~n2987 ;
  assign n2989 = n842 & ~n2988 ;
  assign n2990 = n846 & ~n2989 ;
  assign n2991 = n850 & ~n2990 ;
  assign n2992 = n854 & ~n2991 ;
  assign n2993 = n858 & ~n2992 ;
  assign n2994 = n862 & ~n2993 ;
  assign n2995 = n866 & ~n2994 ;
  assign n2996 = n870 & ~n2995 ;
  assign n2997 = n874 & ~n2996 ;
  assign n2998 = n878 & ~n2997 ;
  assign n2999 = n882 & ~n2998 ;
  assign n3000 = n886 & ~n2999 ;
  assign n3001 = n890 & ~n3000 ;
  assign n3002 = n894 & ~n3001 ;
  assign n3003 = n898 & ~n3002 ;
  assign n3004 = n902 & ~n3003 ;
  assign n3005 = n906 & ~n3004 ;
  assign n3006 = n910 & ~n3005 ;
  assign n3007 = n914 & ~n3006 ;
  assign n3008 = n918 & ~n3007 ;
  assign n3009 = n922 & ~n3008 ;
  assign n3010 = n926 & ~n3009 ;
  assign n3011 = n930 & ~n3010 ;
  assign n3012 = n2472 & ~n3011 ;
  assign n3013 = n2474 & ~n3012 ;
  assign n3014 = n1280 & ~n2476 ;
  assign n3015 = ~n3013 & n3014 ;
  assign n3016 = n1284 & ~n3015 ;
  assign n3017 = ~x134 & ~n1286 ;
  assign n3018 = ~n3016 & n3017 ;
  assign n3021 = ~n3018 & ~x262 ;
  assign n3022 = ~n3020 & ~n3021 ;
  assign n3023 = n956 & ~n1632 ;
  assign n3024 = n961 & ~n3023 ;
  assign n3025 = n965 & ~n3024 ;
  assign n3026 = n969 & ~n3025 ;
  assign n3027 = n973 & ~n3026 ;
  assign n3028 = n977 & ~n3027 ;
  assign n3029 = n981 & ~n3028 ;
  assign n3030 = n985 & ~n3029 ;
  assign n3031 = n989 & ~n3030 ;
  assign n3032 = n993 & ~n3031 ;
  assign n3033 = n997 & ~n3032 ;
  assign n3034 = n1001 & ~n3033 ;
  assign n3035 = n1005 & ~n3034 ;
  assign n3036 = n1009 & ~n3035 ;
  assign n3037 = n1013 & ~n3036 ;
  assign n3038 = n1017 & ~n3037 ;
  assign n3039 = n1021 & ~n3038 ;
  assign n3040 = n1025 & ~n3039 ;
  assign n3041 = n1029 & ~n3040 ;
  assign n3042 = n1033 & ~n3041 ;
  assign n3043 = n1037 & ~n3042 ;
  assign n3044 = n1041 & ~n3043 ;
  assign n3045 = n1045 & ~n3044 ;
  assign n3046 = n1049 & ~n3045 ;
  assign n3047 = n1053 & ~n3046 ;
  assign n3048 = n1057 & ~n3047 ;
  assign n3049 = n1061 & ~n3048 ;
  assign n3050 = n1065 & ~n3049 ;
  assign n3051 = n1069 & ~n3050 ;
  assign n3052 = n1073 & ~n3051 ;
  assign n3053 = n1077 & ~n3052 ;
  assign n3054 = n1081 & ~n3053 ;
  assign n3055 = n1085 & ~n3054 ;
  assign n3056 = n1089 & ~n3055 ;
  assign n3057 = n1093 & ~n3056 ;
  assign n3058 = n1097 & ~n3057 ;
  assign n3059 = n1101 & ~n3058 ;
  assign n3060 = n1105 & ~n3059 ;
  assign n3061 = n1109 & ~n3060 ;
  assign n3062 = n1113 & ~n3061 ;
  assign n3063 = n1117 & ~n3062 ;
  assign n3064 = n1121 & ~n3063 ;
  assign n3065 = n1125 & ~n3064 ;
  assign n3066 = n1129 & ~n3065 ;
  assign n3067 = n1133 & ~n3066 ;
  assign n3068 = n1137 & ~n3067 ;
  assign n3069 = n1141 & ~n3068 ;
  assign n3070 = n1145 & ~n3069 ;
  assign n3071 = n1149 & ~n3070 ;
  assign n3072 = n1153 & ~n3071 ;
  assign n3073 = n1157 & ~n3072 ;
  assign n3074 = n1161 & ~n3073 ;
  assign n3075 = n1165 & ~n3074 ;
  assign n3076 = n1169 & ~n3075 ;
  assign n3077 = n1173 & ~n3076 ;
  assign n3078 = n1177 & ~n3077 ;
  assign n3079 = n1181 & ~n3078 ;
  assign n3080 = n1185 & ~n3079 ;
  assign n3081 = n1189 & ~n3080 ;
  assign n3082 = n1193 & ~n3081 ;
  assign n3083 = n1197 & ~n3082 ;
  assign n3084 = n1201 & ~n3083 ;
  assign n3085 = n1205 & ~n3084 ;
  assign n3086 = n1209 & ~n3085 ;
  assign n3087 = n1213 & ~n3086 ;
  assign n3088 = n1217 & ~n3087 ;
  assign n3089 = n1221 & ~n3088 ;
  assign n3090 = n1225 & ~n3089 ;
  assign n3091 = n1229 & ~n3090 ;
  assign n3092 = n1233 & ~n3091 ;
  assign n3093 = n1237 & ~n3092 ;
  assign n3094 = n1241 & ~n3093 ;
  assign n3095 = n1245 & ~n3094 ;
  assign n3096 = n1249 & ~n3095 ;
  assign n3097 = n1253 & ~n3096 ;
  assign n3098 = n1257 & ~n3097 ;
  assign n3099 = n1261 & ~n3098 ;
  assign n3100 = n1265 & ~n3099 ;
  assign n3101 = n1269 & ~n3100 ;
  assign n3102 = n1273 & ~n3101 ;
  assign n3103 = n2566 & ~n3102 ;
  assign n3104 = n2568 & ~n3103 ;
  assign n3105 = n1621 & ~n2570 ;
  assign n3106 = ~n3104 & n3105 ;
  assign n3107 = n1625 & ~n3106 ;
  assign n3108 = x135 & ~n1627 ;
  assign n3109 = ~n3107 & n3108 ;
  assign n3198 = n3109 & x263 ;
  assign n3110 = n1295 & ~n1969 ;
  assign n3111 = n1300 & ~n3110 ;
  assign n3112 = n1304 & ~n3111 ;
  assign n3113 = n1308 & ~n3112 ;
  assign n3114 = n1312 & ~n3113 ;
  assign n3115 = n1316 & ~n3114 ;
  assign n3116 = n1320 & ~n3115 ;
  assign n3117 = n1324 & ~n3116 ;
  assign n3118 = n1328 & ~n3117 ;
  assign n3119 = n1332 & ~n3118 ;
  assign n3120 = n1336 & ~n3119 ;
  assign n3121 = n1340 & ~n3120 ;
  assign n3122 = n1344 & ~n3121 ;
  assign n3123 = n1348 & ~n3122 ;
  assign n3124 = n1352 & ~n3123 ;
  assign n3125 = n1356 & ~n3124 ;
  assign n3126 = n1360 & ~n3125 ;
  assign n3127 = n1364 & ~n3126 ;
  assign n3128 = n1368 & ~n3127 ;
  assign n3129 = n1372 & ~n3128 ;
  assign n3130 = n1376 & ~n3129 ;
  assign n3131 = n1380 & ~n3130 ;
  assign n3132 = n1384 & ~n3131 ;
  assign n3133 = n1388 & ~n3132 ;
  assign n3134 = n1392 & ~n3133 ;
  assign n3135 = n1396 & ~n3134 ;
  assign n3136 = n1400 & ~n3135 ;
  assign n3137 = n1404 & ~n3136 ;
  assign n3138 = n1408 & ~n3137 ;
  assign n3139 = n1412 & ~n3138 ;
  assign n3140 = n1416 & ~n3139 ;
  assign n3141 = n1420 & ~n3140 ;
  assign n3142 = n1424 & ~n3141 ;
  assign n3143 = n1428 & ~n3142 ;
  assign n3144 = n1432 & ~n3143 ;
  assign n3145 = n1436 & ~n3144 ;
  assign n3146 = n1440 & ~n3145 ;
  assign n3147 = n1444 & ~n3146 ;
  assign n3148 = n1448 & ~n3147 ;
  assign n3149 = n1452 & ~n3148 ;
  assign n3150 = n1456 & ~n3149 ;
  assign n3151 = n1460 & ~n3150 ;
  assign n3152 = n1464 & ~n3151 ;
  assign n3153 = n1468 & ~n3152 ;
  assign n3154 = n1472 & ~n3153 ;
  assign n3155 = n1476 & ~n3154 ;
  assign n3156 = n1480 & ~n3155 ;
  assign n3157 = n1484 & ~n3156 ;
  assign n3158 = n1488 & ~n3157 ;
  assign n3159 = n1492 & ~n3158 ;
  assign n3160 = n1496 & ~n3159 ;
  assign n3161 = n1500 & ~n3160 ;
  assign n3162 = n1504 & ~n3161 ;
  assign n3163 = n1508 & ~n3162 ;
  assign n3164 = n1512 & ~n3163 ;
  assign n3165 = n1516 & ~n3164 ;
  assign n3166 = n1520 & ~n3165 ;
  assign n3167 = n1524 & ~n3166 ;
  assign n3168 = n1528 & ~n3167 ;
  assign n3169 = n1532 & ~n3168 ;
  assign n3170 = n1536 & ~n3169 ;
  assign n3171 = n1540 & ~n3170 ;
  assign n3172 = n1544 & ~n3171 ;
  assign n3173 = n1548 & ~n3172 ;
  assign n3174 = n1552 & ~n3173 ;
  assign n3175 = n1556 & ~n3174 ;
  assign n3176 = n1560 & ~n3175 ;
  assign n3177 = n1564 & ~n3176 ;
  assign n3178 = n1568 & ~n3177 ;
  assign n3179 = n1572 & ~n3178 ;
  assign n3180 = n1576 & ~n3179 ;
  assign n3181 = n1580 & ~n3180 ;
  assign n3182 = n1584 & ~n3181 ;
  assign n3183 = n1588 & ~n3182 ;
  assign n3184 = n1592 & ~n3183 ;
  assign n3185 = n1596 & ~n3184 ;
  assign n3186 = n1600 & ~n3185 ;
  assign n3187 = n1604 & ~n3186 ;
  assign n3188 = n1608 & ~n3187 ;
  assign n3189 = n1612 & ~n3188 ;
  assign n3190 = n2656 & ~n3189 ;
  assign n3191 = n2658 & ~n3190 ;
  assign n3192 = n1958 & ~n2660 ;
  assign n3193 = ~n3191 & n3192 ;
  assign n3194 = n1962 & ~n3193 ;
  assign n3195 = ~x135 & ~n1964 ;
  assign n3196 = ~n3194 & n3195 ;
  assign n3199 = ~n3196 & ~x263 ;
  assign n3200 = ~n3198 & ~n3199 ;
  assign n3201 = ~n278 & n1636 ;
  assign n3202 = n1641 & ~n3201 ;
  assign n3203 = n1645 & ~n3202 ;
  assign n3204 = n1649 & ~n3203 ;
  assign n3205 = n1653 & ~n3204 ;
  assign n3206 = n1657 & ~n3205 ;
  assign n3207 = n1661 & ~n3206 ;
  assign n3208 = n1665 & ~n3207 ;
  assign n3209 = n1669 & ~n3208 ;
  assign n3210 = n1673 & ~n3209 ;
  assign n3211 = n1677 & ~n3210 ;
  assign n3212 = n1681 & ~n3211 ;
  assign n3213 = n1685 & ~n3212 ;
  assign n3214 = n1689 & ~n3213 ;
  assign n3215 = n1693 & ~n3214 ;
  assign n3216 = n1697 & ~n3215 ;
  assign n3217 = n1701 & ~n3216 ;
  assign n3218 = n1705 & ~n3217 ;
  assign n3219 = n1709 & ~n3218 ;
  assign n3220 = n1713 & ~n3219 ;
  assign n3221 = n1717 & ~n3220 ;
  assign n3222 = n1721 & ~n3221 ;
  assign n3223 = n1725 & ~n3222 ;
  assign n3224 = n1729 & ~n3223 ;
  assign n3225 = n1733 & ~n3224 ;
  assign n3226 = n1737 & ~n3225 ;
  assign n3227 = n1741 & ~n3226 ;
  assign n3228 = n1745 & ~n3227 ;
  assign n3229 = n1749 & ~n3228 ;
  assign n3230 = n1753 & ~n3229 ;
  assign n3231 = n1757 & ~n3230 ;
  assign n3232 = n1761 & ~n3231 ;
  assign n3233 = n1765 & ~n3232 ;
  assign n3234 = n1769 & ~n3233 ;
  assign n3235 = n1773 & ~n3234 ;
  assign n3236 = n1777 & ~n3235 ;
  assign n3237 = n1781 & ~n3236 ;
  assign n3238 = n1785 & ~n3237 ;
  assign n3239 = n1789 & ~n3238 ;
  assign n3240 = n1793 & ~n3239 ;
  assign n3241 = n1797 & ~n3240 ;
  assign n3242 = n1801 & ~n3241 ;
  assign n3243 = n1805 & ~n3242 ;
  assign n3244 = n1809 & ~n3243 ;
  assign n3245 = n1813 & ~n3244 ;
  assign n3246 = n1817 & ~n3245 ;
  assign n3247 = n1821 & ~n3246 ;
  assign n3248 = n1825 & ~n3247 ;
  assign n3249 = n1829 & ~n3248 ;
  assign n3250 = n1833 & ~n3249 ;
  assign n3251 = n1837 & ~n3250 ;
  assign n3252 = n1841 & ~n3251 ;
  assign n3253 = n1845 & ~n3252 ;
  assign n3254 = n1849 & ~n3253 ;
  assign n3255 = n1853 & ~n3254 ;
  assign n3256 = n1857 & ~n3255 ;
  assign n3257 = n1861 & ~n3256 ;
  assign n3258 = n1865 & ~n3257 ;
  assign n3259 = n1869 & ~n3258 ;
  assign n3260 = n1873 & ~n3259 ;
  assign n3261 = n1877 & ~n3260 ;
  assign n3262 = n1881 & ~n3261 ;
  assign n3263 = n1885 & ~n3262 ;
  assign n3264 = n1889 & ~n3263 ;
  assign n3265 = n1893 & ~n3264 ;
  assign n3266 = n1897 & ~n3265 ;
  assign n3267 = n1901 & ~n3266 ;
  assign n3268 = n1905 & ~n3267 ;
  assign n3269 = n1909 & ~n3268 ;
  assign n3270 = n1913 & ~n3269 ;
  assign n3271 = n1917 & ~n3270 ;
  assign n3272 = n1921 & ~n3271 ;
  assign n3273 = n1925 & ~n3272 ;
  assign n3274 = n1929 & ~n3273 ;
  assign n3275 = n1933 & ~n3274 ;
  assign n3276 = n1937 & ~n3275 ;
  assign n3277 = n1941 & ~n3276 ;
  assign n3278 = n1945 & ~n3277 ;
  assign n3279 = n1949 & ~n3278 ;
  assign n3280 = n1953 & ~n3279 ;
  assign n3281 = n2749 & ~n3280 ;
  assign n3282 = n263 & ~n3281 ;
  assign n3283 = n267 & ~n3282 ;
  assign n3284 = n271 & ~n3283 ;
  assign n3285 = x136 & ~n273 ;
  assign n3286 = ~n3284 & n3285 ;
  assign n3374 = n3286 & x264 ;
  assign n3287 = ~n617 & n1973 ;
  assign n3288 = n1978 & ~n3287 ;
  assign n3289 = n1982 & ~n3288 ;
  assign n3290 = n1986 & ~n3289 ;
  assign n3291 = n1990 & ~n3290 ;
  assign n3292 = n1994 & ~n3291 ;
  assign n3293 = n1998 & ~n3292 ;
  assign n3294 = n2002 & ~n3293 ;
  assign n3295 = n2006 & ~n3294 ;
  assign n3296 = n2010 & ~n3295 ;
  assign n3297 = n2014 & ~n3296 ;
  assign n3298 = n2018 & ~n3297 ;
  assign n3299 = n2022 & ~n3298 ;
  assign n3300 = n2026 & ~n3299 ;
  assign n3301 = n2030 & ~n3300 ;
  assign n3302 = n2034 & ~n3301 ;
  assign n3303 = n2038 & ~n3302 ;
  assign n3304 = n2042 & ~n3303 ;
  assign n3305 = n2046 & ~n3304 ;
  assign n3306 = n2050 & ~n3305 ;
  assign n3307 = n2054 & ~n3306 ;
  assign n3308 = n2058 & ~n3307 ;
  assign n3309 = n2062 & ~n3308 ;
  assign n3310 = n2066 & ~n3309 ;
  assign n3311 = n2070 & ~n3310 ;
  assign n3312 = n2074 & ~n3311 ;
  assign n3313 = n2078 & ~n3312 ;
  assign n3314 = n2082 & ~n3313 ;
  assign n3315 = n2086 & ~n3314 ;
  assign n3316 = n2090 & ~n3315 ;
  assign n3317 = n2094 & ~n3316 ;
  assign n3318 = n2098 & ~n3317 ;
  assign n3319 = n2102 & ~n3318 ;
  assign n3320 = n2106 & ~n3319 ;
  assign n3321 = n2110 & ~n3320 ;
  assign n3322 = n2114 & ~n3321 ;
  assign n3323 = n2118 & ~n3322 ;
  assign n3324 = n2122 & ~n3323 ;
  assign n3325 = n2126 & ~n3324 ;
  assign n3326 = n2130 & ~n3325 ;
  assign n3327 = n2134 & ~n3326 ;
  assign n3328 = n2138 & ~n3327 ;
  assign n3329 = n2142 & ~n3328 ;
  assign n3330 = n2146 & ~n3329 ;
  assign n3331 = n2150 & ~n3330 ;
  assign n3332 = n2154 & ~n3331 ;
  assign n3333 = n2158 & ~n3332 ;
  assign n3334 = n2162 & ~n3333 ;
  assign n3335 = n2166 & ~n3334 ;
  assign n3336 = n2170 & ~n3335 ;
  assign n3337 = n2174 & ~n3336 ;
  assign n3338 = n2178 & ~n3337 ;
  assign n3339 = n2182 & ~n3338 ;
  assign n3340 = n2186 & ~n3339 ;
  assign n3341 = n2190 & ~n3340 ;
  assign n3342 = n2194 & ~n3341 ;
  assign n3343 = n2198 & ~n3342 ;
  assign n3344 = n2202 & ~n3343 ;
  assign n3345 = n2206 & ~n3344 ;
  assign n3346 = n2210 & ~n3345 ;
  assign n3347 = n2214 & ~n3346 ;
  assign n3348 = n2218 & ~n3347 ;
  assign n3349 = n2222 & ~n3348 ;
  assign n3350 = n2226 & ~n3349 ;
  assign n3351 = n2230 & ~n3350 ;
  assign n3352 = n2234 & ~n3351 ;
  assign n3353 = n2238 & ~n3352 ;
  assign n3354 = n2242 & ~n3353 ;
  assign n3355 = n2246 & ~n3354 ;
  assign n3356 = n2250 & ~n3355 ;
  assign n3357 = n2254 & ~n3356 ;
  assign n3358 = n2258 & ~n3357 ;
  assign n3359 = n2262 & ~n3358 ;
  assign n3360 = n2266 & ~n3359 ;
  assign n3361 = n2270 & ~n3360 ;
  assign n3362 = n2274 & ~n3361 ;
  assign n3363 = n2278 & ~n3362 ;
  assign n3364 = n2282 & ~n3363 ;
  assign n3365 = n2286 & ~n3364 ;
  assign n3366 = n2290 & ~n3365 ;
  assign n3367 = n2836 & ~n3366 ;
  assign n3368 = n602 & ~n3367 ;
  assign n3369 = n606 & ~n3368 ;
  assign n3370 = n610 & ~n3369 ;
  assign n3371 = ~x136 & ~n612 ;
  assign n3372 = ~n3370 & n3371 ;
  assign n3375 = ~n3372 & ~x264 ;
  assign n3376 = ~n3374 & ~n3375 ;
  assign n3377 = n282 & ~n960 ;
  assign n3378 = n287 & ~n3377 ;
  assign n3379 = n291 & ~n3378 ;
  assign n3380 = n295 & ~n3379 ;
  assign n3381 = n299 & ~n3380 ;
  assign n3382 = n303 & ~n3381 ;
  assign n3383 = n307 & ~n3382 ;
  assign n3384 = n311 & ~n3383 ;
  assign n3385 = n315 & ~n3384 ;
  assign n3386 = n319 & ~n3385 ;
  assign n3387 = n323 & ~n3386 ;
  assign n3388 = n327 & ~n3387 ;
  assign n3389 = n331 & ~n3388 ;
  assign n3390 = n335 & ~n3389 ;
  assign n3391 = n339 & ~n3390 ;
  assign n3392 = n343 & ~n3391 ;
  assign n3393 = n347 & ~n3392 ;
  assign n3394 = n351 & ~n3393 ;
  assign n3395 = n355 & ~n3394 ;
  assign n3396 = n359 & ~n3395 ;
  assign n3397 = n363 & ~n3396 ;
  assign n3398 = n367 & ~n3397 ;
  assign n3399 = n371 & ~n3398 ;
  assign n3400 = n375 & ~n3399 ;
  assign n3401 = n379 & ~n3400 ;
  assign n3402 = n383 & ~n3401 ;
  assign n3403 = n387 & ~n3402 ;
  assign n3404 = n391 & ~n3403 ;
  assign n3405 = n395 & ~n3404 ;
  assign n3406 = n399 & ~n3405 ;
  assign n3407 = n403 & ~n3406 ;
  assign n3408 = n407 & ~n3407 ;
  assign n3409 = n411 & ~n3408 ;
  assign n3410 = n415 & ~n3409 ;
  assign n3411 = n419 & ~n3410 ;
  assign n3412 = n423 & ~n3411 ;
  assign n3413 = n427 & ~n3412 ;
  assign n3414 = n431 & ~n3413 ;
  assign n3415 = n435 & ~n3414 ;
  assign n3416 = n439 & ~n3415 ;
  assign n3417 = n443 & ~n3416 ;
  assign n3418 = n447 & ~n3417 ;
  assign n3419 = n451 & ~n3418 ;
  assign n3420 = n455 & ~n3419 ;
  assign n3421 = n459 & ~n3420 ;
  assign n3422 = n463 & ~n3421 ;
  assign n3423 = n467 & ~n3422 ;
  assign n3424 = n471 & ~n3423 ;
  assign n3425 = n475 & ~n3424 ;
  assign n3426 = n479 & ~n3425 ;
  assign n3427 = n483 & ~n3426 ;
  assign n3428 = n487 & ~n3427 ;
  assign n3429 = n491 & ~n3428 ;
  assign n3430 = n495 & ~n3429 ;
  assign n3431 = n499 & ~n3430 ;
  assign n3432 = n503 & ~n3431 ;
  assign n3433 = n507 & ~n3432 ;
  assign n3434 = n511 & ~n3433 ;
  assign n3435 = n515 & ~n3434 ;
  assign n3436 = n519 & ~n3435 ;
  assign n3437 = n523 & ~n3436 ;
  assign n3438 = n527 & ~n3437 ;
  assign n3439 = n531 & ~n3438 ;
  assign n3440 = n535 & ~n3439 ;
  assign n3441 = n539 & ~n3440 ;
  assign n3442 = n543 & ~n3441 ;
  assign n3443 = n547 & ~n3442 ;
  assign n3444 = n551 & ~n3443 ;
  assign n3445 = n555 & ~n3444 ;
  assign n3446 = n559 & ~n3445 ;
  assign n3447 = n563 & ~n3446 ;
  assign n3448 = n567 & ~n3447 ;
  assign n3449 = n571 & ~n3448 ;
  assign n3450 = n575 & ~n3449 ;
  assign n3451 = n579 & ~n3450 ;
  assign n3452 = n583 & ~n3451 ;
  assign n3453 = n587 & ~n3452 ;
  assign n3454 = n591 & ~n3453 ;
  assign n3455 = n2382 & ~n3454 ;
  assign n3456 = n2384 & ~n3455 ;
  assign n3457 = n2927 & ~n3456 ;
  assign n3458 = n945 & ~n3457 ;
  assign n3459 = n949 & ~n3458 ;
  assign n3460 = n953 & ~n3459 ;
  assign n3461 = x137 & ~n955 ;
  assign n3462 = ~n3460 & n3461 ;
  assign n3550 = n3462 & x265 ;
  assign n3463 = n621 & ~n1299 ;
  assign n3464 = n626 & ~n3463 ;
  assign n3465 = n630 & ~n3464 ;
  assign n3466 = n634 & ~n3465 ;
  assign n3467 = n638 & ~n3466 ;
  assign n3468 = n642 & ~n3467 ;
  assign n3469 = n646 & ~n3468 ;
  assign n3470 = n650 & ~n3469 ;
  assign n3471 = n654 & ~n3470 ;
  assign n3472 = n658 & ~n3471 ;
  assign n3473 = n662 & ~n3472 ;
  assign n3474 = n666 & ~n3473 ;
  assign n3475 = n670 & ~n3474 ;
  assign n3476 = n674 & ~n3475 ;
  assign n3477 = n678 & ~n3476 ;
  assign n3478 = n682 & ~n3477 ;
  assign n3479 = n686 & ~n3478 ;
  assign n3480 = n690 & ~n3479 ;
  assign n3481 = n694 & ~n3480 ;
  assign n3482 = n698 & ~n3481 ;
  assign n3483 = n702 & ~n3482 ;
  assign n3484 = n706 & ~n3483 ;
  assign n3485 = n710 & ~n3484 ;
  assign n3486 = n714 & ~n3485 ;
  assign n3487 = n718 & ~n3486 ;
  assign n3488 = n722 & ~n3487 ;
  assign n3489 = n726 & ~n3488 ;
  assign n3490 = n730 & ~n3489 ;
  assign n3491 = n734 & ~n3490 ;
  assign n3492 = n738 & ~n3491 ;
  assign n3493 = n742 & ~n3492 ;
  assign n3494 = n746 & ~n3493 ;
  assign n3495 = n750 & ~n3494 ;
  assign n3496 = n754 & ~n3495 ;
  assign n3497 = n758 & ~n3496 ;
  assign n3498 = n762 & ~n3497 ;
  assign n3499 = n766 & ~n3498 ;
  assign n3500 = n770 & ~n3499 ;
  assign n3501 = n774 & ~n3500 ;
  assign n3502 = n778 & ~n3501 ;
  assign n3503 = n782 & ~n3502 ;
  assign n3504 = n786 & ~n3503 ;
  assign n3505 = n790 & ~n3504 ;
  assign n3506 = n794 & ~n3505 ;
  assign n3507 = n798 & ~n3506 ;
  assign n3508 = n802 & ~n3507 ;
  assign n3509 = n806 & ~n3508 ;
  assign n3510 = n810 & ~n3509 ;
  assign n3511 = n814 & ~n3510 ;
  assign n3512 = n818 & ~n3511 ;
  assign n3513 = n822 & ~n3512 ;
  assign n3514 = n826 & ~n3513 ;
  assign n3515 = n830 & ~n3514 ;
  assign n3516 = n834 & ~n3515 ;
  assign n3517 = n838 & ~n3516 ;
  assign n3518 = n842 & ~n3517 ;
  assign n3519 = n846 & ~n3518 ;
  assign n3520 = n850 & ~n3519 ;
  assign n3521 = n854 & ~n3520 ;
  assign n3522 = n858 & ~n3521 ;
  assign n3523 = n862 & ~n3522 ;
  assign n3524 = n866 & ~n3523 ;
  assign n3525 = n870 & ~n3524 ;
  assign n3526 = n874 & ~n3525 ;
  assign n3527 = n878 & ~n3526 ;
  assign n3528 = n882 & ~n3527 ;
  assign n3529 = n886 & ~n3528 ;
  assign n3530 = n890 & ~n3529 ;
  assign n3531 = n894 & ~n3530 ;
  assign n3532 = n898 & ~n3531 ;
  assign n3533 = n902 & ~n3532 ;
  assign n3534 = n906 & ~n3533 ;
  assign n3535 = n910 & ~n3534 ;
  assign n3536 = n914 & ~n3535 ;
  assign n3537 = n918 & ~n3536 ;
  assign n3538 = n922 & ~n3537 ;
  assign n3539 = n926 & ~n3538 ;
  assign n3540 = n930 & ~n3539 ;
  assign n3541 = n2472 & ~n3540 ;
  assign n3542 = n2474 & ~n3541 ;
  assign n3543 = n3014 & ~n3542 ;
  assign n3544 = n1284 & ~n3543 ;
  assign n3545 = n1288 & ~n3544 ;
  assign n3546 = n1292 & ~n3545 ;
  assign n3547 = ~x137 & ~n1294 ;
  assign n3548 = ~n3546 & n3547 ;
  assign n3551 = ~n3548 & ~x265 ;
  assign n3552 = ~n3550 & ~n3551 ;
  assign n3553 = n964 & ~n1640 ;
  assign n3554 = n969 & ~n3553 ;
  assign n3555 = n973 & ~n3554 ;
  assign n3556 = n977 & ~n3555 ;
  assign n3557 = n981 & ~n3556 ;
  assign n3558 = n985 & ~n3557 ;
  assign n3559 = n989 & ~n3558 ;
  assign n3560 = n993 & ~n3559 ;
  assign n3561 = n997 & ~n3560 ;
  assign n3562 = n1001 & ~n3561 ;
  assign n3563 = n1005 & ~n3562 ;
  assign n3564 = n1009 & ~n3563 ;
  assign n3565 = n1013 & ~n3564 ;
  assign n3566 = n1017 & ~n3565 ;
  assign n3567 = n1021 & ~n3566 ;
  assign n3568 = n1025 & ~n3567 ;
  assign n3569 = n1029 & ~n3568 ;
  assign n3570 = n1033 & ~n3569 ;
  assign n3571 = n1037 & ~n3570 ;
  assign n3572 = n1041 & ~n3571 ;
  assign n3573 = n1045 & ~n3572 ;
  assign n3574 = n1049 & ~n3573 ;
  assign n3575 = n1053 & ~n3574 ;
  assign n3576 = n1057 & ~n3575 ;
  assign n3577 = n1061 & ~n3576 ;
  assign n3578 = n1065 & ~n3577 ;
  assign n3579 = n1069 & ~n3578 ;
  assign n3580 = n1073 & ~n3579 ;
  assign n3581 = n1077 & ~n3580 ;
  assign n3582 = n1081 & ~n3581 ;
  assign n3583 = n1085 & ~n3582 ;
  assign n3584 = n1089 & ~n3583 ;
  assign n3585 = n1093 & ~n3584 ;
  assign n3586 = n1097 & ~n3585 ;
  assign n3587 = n1101 & ~n3586 ;
  assign n3588 = n1105 & ~n3587 ;
  assign n3589 = n1109 & ~n3588 ;
  assign n3590 = n1113 & ~n3589 ;
  assign n3591 = n1117 & ~n3590 ;
  assign n3592 = n1121 & ~n3591 ;
  assign n3593 = n1125 & ~n3592 ;
  assign n3594 = n1129 & ~n3593 ;
  assign n3595 = n1133 & ~n3594 ;
  assign n3596 = n1137 & ~n3595 ;
  assign n3597 = n1141 & ~n3596 ;
  assign n3598 = n1145 & ~n3597 ;
  assign n3599 = n1149 & ~n3598 ;
  assign n3600 = n1153 & ~n3599 ;
  assign n3601 = n1157 & ~n3600 ;
  assign n3602 = n1161 & ~n3601 ;
  assign n3603 = n1165 & ~n3602 ;
  assign n3604 = n1169 & ~n3603 ;
  assign n3605 = n1173 & ~n3604 ;
  assign n3606 = n1177 & ~n3605 ;
  assign n3607 = n1181 & ~n3606 ;
  assign n3608 = n1185 & ~n3607 ;
  assign n3609 = n1189 & ~n3608 ;
  assign n3610 = n1193 & ~n3609 ;
  assign n3611 = n1197 & ~n3610 ;
  assign n3612 = n1201 & ~n3611 ;
  assign n3613 = n1205 & ~n3612 ;
  assign n3614 = n1209 & ~n3613 ;
  assign n3615 = n1213 & ~n3614 ;
  assign n3616 = n1217 & ~n3615 ;
  assign n3617 = n1221 & ~n3616 ;
  assign n3618 = n1225 & ~n3617 ;
  assign n3619 = n1229 & ~n3618 ;
  assign n3620 = n1233 & ~n3619 ;
  assign n3621 = n1237 & ~n3620 ;
  assign n3622 = n1241 & ~n3621 ;
  assign n3623 = n1245 & ~n3622 ;
  assign n3624 = n1249 & ~n3623 ;
  assign n3625 = n1253 & ~n3624 ;
  assign n3626 = n1257 & ~n3625 ;
  assign n3627 = n1261 & ~n3626 ;
  assign n3628 = n1265 & ~n3627 ;
  assign n3629 = n1269 & ~n3628 ;
  assign n3630 = n1273 & ~n3629 ;
  assign n3631 = n2566 & ~n3630 ;
  assign n3632 = n2568 & ~n3631 ;
  assign n3633 = n3105 & ~n3632 ;
  assign n3634 = n1625 & ~n3633 ;
  assign n3635 = n1629 & ~n3634 ;
  assign n3636 = n1633 & ~n3635 ;
  assign n3637 = x138 & ~n1635 ;
  assign n3638 = ~n3636 & n3637 ;
  assign n3726 = n3638 & x266 ;
  assign n3639 = n1303 & ~n1977 ;
  assign n3640 = n1308 & ~n3639 ;
  assign n3641 = n1312 & ~n3640 ;
  assign n3642 = n1316 & ~n3641 ;
  assign n3643 = n1320 & ~n3642 ;
  assign n3644 = n1324 & ~n3643 ;
  assign n3645 = n1328 & ~n3644 ;
  assign n3646 = n1332 & ~n3645 ;
  assign n3647 = n1336 & ~n3646 ;
  assign n3648 = n1340 & ~n3647 ;
  assign n3649 = n1344 & ~n3648 ;
  assign n3650 = n1348 & ~n3649 ;
  assign n3651 = n1352 & ~n3650 ;
  assign n3652 = n1356 & ~n3651 ;
  assign n3653 = n1360 & ~n3652 ;
  assign n3654 = n1364 & ~n3653 ;
  assign n3655 = n1368 & ~n3654 ;
  assign n3656 = n1372 & ~n3655 ;
  assign n3657 = n1376 & ~n3656 ;
  assign n3658 = n1380 & ~n3657 ;
  assign n3659 = n1384 & ~n3658 ;
  assign n3660 = n1388 & ~n3659 ;
  assign n3661 = n1392 & ~n3660 ;
  assign n3662 = n1396 & ~n3661 ;
  assign n3663 = n1400 & ~n3662 ;
  assign n3664 = n1404 & ~n3663 ;
  assign n3665 = n1408 & ~n3664 ;
  assign n3666 = n1412 & ~n3665 ;
  assign n3667 = n1416 & ~n3666 ;
  assign n3668 = n1420 & ~n3667 ;
  assign n3669 = n1424 & ~n3668 ;
  assign n3670 = n1428 & ~n3669 ;
  assign n3671 = n1432 & ~n3670 ;
  assign n3672 = n1436 & ~n3671 ;
  assign n3673 = n1440 & ~n3672 ;
  assign n3674 = n1444 & ~n3673 ;
  assign n3675 = n1448 & ~n3674 ;
  assign n3676 = n1452 & ~n3675 ;
  assign n3677 = n1456 & ~n3676 ;
  assign n3678 = n1460 & ~n3677 ;
  assign n3679 = n1464 & ~n3678 ;
  assign n3680 = n1468 & ~n3679 ;
  assign n3681 = n1472 & ~n3680 ;
  assign n3682 = n1476 & ~n3681 ;
  assign n3683 = n1480 & ~n3682 ;
  assign n3684 = n1484 & ~n3683 ;
  assign n3685 = n1488 & ~n3684 ;
  assign n3686 = n1492 & ~n3685 ;
  assign n3687 = n1496 & ~n3686 ;
  assign n3688 = n1500 & ~n3687 ;
  assign n3689 = n1504 & ~n3688 ;
  assign n3690 = n1508 & ~n3689 ;
  assign n3691 = n1512 & ~n3690 ;
  assign n3692 = n1516 & ~n3691 ;
  assign n3693 = n1520 & ~n3692 ;
  assign n3694 = n1524 & ~n3693 ;
  assign n3695 = n1528 & ~n3694 ;
  assign n3696 = n1532 & ~n3695 ;
  assign n3697 = n1536 & ~n3696 ;
  assign n3698 = n1540 & ~n3697 ;
  assign n3699 = n1544 & ~n3698 ;
  assign n3700 = n1548 & ~n3699 ;
  assign n3701 = n1552 & ~n3700 ;
  assign n3702 = n1556 & ~n3701 ;
  assign n3703 = n1560 & ~n3702 ;
  assign n3704 = n1564 & ~n3703 ;
  assign n3705 = n1568 & ~n3704 ;
  assign n3706 = n1572 & ~n3705 ;
  assign n3707 = n1576 & ~n3706 ;
  assign n3708 = n1580 & ~n3707 ;
  assign n3709 = n1584 & ~n3708 ;
  assign n3710 = n1588 & ~n3709 ;
  assign n3711 = n1592 & ~n3710 ;
  assign n3712 = n1596 & ~n3711 ;
  assign n3713 = n1600 & ~n3712 ;
  assign n3714 = n1604 & ~n3713 ;
  assign n3715 = n1608 & ~n3714 ;
  assign n3716 = n1612 & ~n3715 ;
  assign n3717 = n2656 & ~n3716 ;
  assign n3718 = n2658 & ~n3717 ;
  assign n3719 = n3192 & ~n3718 ;
  assign n3720 = n1962 & ~n3719 ;
  assign n3721 = n1966 & ~n3720 ;
  assign n3722 = n1970 & ~n3721 ;
  assign n3723 = ~x138 & ~n1972 ;
  assign n3724 = ~n3722 & n3723 ;
  assign n3727 = ~n3724 & ~x266 ;
  assign n3728 = ~n3726 & ~n3727 ;
  assign n3729 = ~n286 & n1644 ;
  assign n3730 = n1649 & ~n3729 ;
  assign n3731 = n1653 & ~n3730 ;
  assign n3732 = n1657 & ~n3731 ;
  assign n3733 = n1661 & ~n3732 ;
  assign n3734 = n1665 & ~n3733 ;
  assign n3735 = n1669 & ~n3734 ;
  assign n3736 = n1673 & ~n3735 ;
  assign n3737 = n1677 & ~n3736 ;
  assign n3738 = n1681 & ~n3737 ;
  assign n3739 = n1685 & ~n3738 ;
  assign n3740 = n1689 & ~n3739 ;
  assign n3741 = n1693 & ~n3740 ;
  assign n3742 = n1697 & ~n3741 ;
  assign n3743 = n1701 & ~n3742 ;
  assign n3744 = n1705 & ~n3743 ;
  assign n3745 = n1709 & ~n3744 ;
  assign n3746 = n1713 & ~n3745 ;
  assign n3747 = n1717 & ~n3746 ;
  assign n3748 = n1721 & ~n3747 ;
  assign n3749 = n1725 & ~n3748 ;
  assign n3750 = n1729 & ~n3749 ;
  assign n3751 = n1733 & ~n3750 ;
  assign n3752 = n1737 & ~n3751 ;
  assign n3753 = n1741 & ~n3752 ;
  assign n3754 = n1745 & ~n3753 ;
  assign n3755 = n1749 & ~n3754 ;
  assign n3756 = n1753 & ~n3755 ;
  assign n3757 = n1757 & ~n3756 ;
  assign n3758 = n1761 & ~n3757 ;
  assign n3759 = n1765 & ~n3758 ;
  assign n3760 = n1769 & ~n3759 ;
  assign n3761 = n1773 & ~n3760 ;
  assign n3762 = n1777 & ~n3761 ;
  assign n3763 = n1781 & ~n3762 ;
  assign n3764 = n1785 & ~n3763 ;
  assign n3765 = n1789 & ~n3764 ;
  assign n3766 = n1793 & ~n3765 ;
  assign n3767 = n1797 & ~n3766 ;
  assign n3768 = n1801 & ~n3767 ;
  assign n3769 = n1805 & ~n3768 ;
  assign n3770 = n1809 & ~n3769 ;
  assign n3771 = n1813 & ~n3770 ;
  assign n3772 = n1817 & ~n3771 ;
  assign n3773 = n1821 & ~n3772 ;
  assign n3774 = n1825 & ~n3773 ;
  assign n3775 = n1829 & ~n3774 ;
  assign n3776 = n1833 & ~n3775 ;
  assign n3777 = n1837 & ~n3776 ;
  assign n3778 = n1841 & ~n3777 ;
  assign n3779 = n1845 & ~n3778 ;
  assign n3780 = n1849 & ~n3779 ;
  assign n3781 = n1853 & ~n3780 ;
  assign n3782 = n1857 & ~n3781 ;
  assign n3783 = n1861 & ~n3782 ;
  assign n3784 = n1865 & ~n3783 ;
  assign n3785 = n1869 & ~n3784 ;
  assign n3786 = n1873 & ~n3785 ;
  assign n3787 = n1877 & ~n3786 ;
  assign n3788 = n1881 & ~n3787 ;
  assign n3789 = n1885 & ~n3788 ;
  assign n3790 = n1889 & ~n3789 ;
  assign n3791 = n1893 & ~n3790 ;
  assign n3792 = n1897 & ~n3791 ;
  assign n3793 = n1901 & ~n3792 ;
  assign n3794 = n1905 & ~n3793 ;
  assign n3795 = n1909 & ~n3794 ;
  assign n3796 = n1913 & ~n3795 ;
  assign n3797 = n1917 & ~n3796 ;
  assign n3798 = n1921 & ~n3797 ;
  assign n3799 = n1925 & ~n3798 ;
  assign n3800 = n1929 & ~n3799 ;
  assign n3801 = n1933 & ~n3800 ;
  assign n3802 = n1937 & ~n3801 ;
  assign n3803 = n1941 & ~n3802 ;
  assign n3804 = n1945 & ~n3803 ;
  assign n3805 = n1949 & ~n3804 ;
  assign n3806 = n1953 & ~n3805 ;
  assign n3807 = n2749 & ~n3806 ;
  assign n3808 = n263 & ~n3807 ;
  assign n3809 = n267 & ~n3808 ;
  assign n3810 = n271 & ~n3809 ;
  assign n3811 = n275 & ~n3810 ;
  assign n3812 = n279 & ~n3811 ;
  assign n3813 = x139 & ~n281 ;
  assign n3814 = ~n3812 & n3813 ;
  assign n3902 = n3814 & x267 ;
  assign n3815 = ~n625 & n1981 ;
  assign n3816 = n1986 & ~n3815 ;
  assign n3817 = n1990 & ~n3816 ;
  assign n3818 = n1994 & ~n3817 ;
  assign n3819 = n1998 & ~n3818 ;
  assign n3820 = n2002 & ~n3819 ;
  assign n3821 = n2006 & ~n3820 ;
  assign n3822 = n2010 & ~n3821 ;
  assign n3823 = n2014 & ~n3822 ;
  assign n3824 = n2018 & ~n3823 ;
  assign n3825 = n2022 & ~n3824 ;
  assign n3826 = n2026 & ~n3825 ;
  assign n3827 = n2030 & ~n3826 ;
  assign n3828 = n2034 & ~n3827 ;
  assign n3829 = n2038 & ~n3828 ;
  assign n3830 = n2042 & ~n3829 ;
  assign n3831 = n2046 & ~n3830 ;
  assign n3832 = n2050 & ~n3831 ;
  assign n3833 = n2054 & ~n3832 ;
  assign n3834 = n2058 & ~n3833 ;
  assign n3835 = n2062 & ~n3834 ;
  assign n3836 = n2066 & ~n3835 ;
  assign n3837 = n2070 & ~n3836 ;
  assign n3838 = n2074 & ~n3837 ;
  assign n3839 = n2078 & ~n3838 ;
  assign n3840 = n2082 & ~n3839 ;
  assign n3841 = n2086 & ~n3840 ;
  assign n3842 = n2090 & ~n3841 ;
  assign n3843 = n2094 & ~n3842 ;
  assign n3844 = n2098 & ~n3843 ;
  assign n3845 = n2102 & ~n3844 ;
  assign n3846 = n2106 & ~n3845 ;
  assign n3847 = n2110 & ~n3846 ;
  assign n3848 = n2114 & ~n3847 ;
  assign n3849 = n2118 & ~n3848 ;
  assign n3850 = n2122 & ~n3849 ;
  assign n3851 = n2126 & ~n3850 ;
  assign n3852 = n2130 & ~n3851 ;
  assign n3853 = n2134 & ~n3852 ;
  assign n3854 = n2138 & ~n3853 ;
  assign n3855 = n2142 & ~n3854 ;
  assign n3856 = n2146 & ~n3855 ;
  assign n3857 = n2150 & ~n3856 ;
  assign n3858 = n2154 & ~n3857 ;
  assign n3859 = n2158 & ~n3858 ;
  assign n3860 = n2162 & ~n3859 ;
  assign n3861 = n2166 & ~n3860 ;
  assign n3862 = n2170 & ~n3861 ;
  assign n3863 = n2174 & ~n3862 ;
  assign n3864 = n2178 & ~n3863 ;
  assign n3865 = n2182 & ~n3864 ;
  assign n3866 = n2186 & ~n3865 ;
  assign n3867 = n2190 & ~n3866 ;
  assign n3868 = n2194 & ~n3867 ;
  assign n3869 = n2198 & ~n3868 ;
  assign n3870 = n2202 & ~n3869 ;
  assign n3871 = n2206 & ~n3870 ;
  assign n3872 = n2210 & ~n3871 ;
  assign n3873 = n2214 & ~n3872 ;
  assign n3874 = n2218 & ~n3873 ;
  assign n3875 = n2222 & ~n3874 ;
  assign n3876 = n2226 & ~n3875 ;
  assign n3877 = n2230 & ~n3876 ;
  assign n3878 = n2234 & ~n3877 ;
  assign n3879 = n2238 & ~n3878 ;
  assign n3880 = n2242 & ~n3879 ;
  assign n3881 = n2246 & ~n3880 ;
  assign n3882 = n2250 & ~n3881 ;
  assign n3883 = n2254 & ~n3882 ;
  assign n3884 = n2258 & ~n3883 ;
  assign n3885 = n2262 & ~n3884 ;
  assign n3886 = n2266 & ~n3885 ;
  assign n3887 = n2270 & ~n3886 ;
  assign n3888 = n2274 & ~n3887 ;
  assign n3889 = n2278 & ~n3888 ;
  assign n3890 = n2282 & ~n3889 ;
  assign n3891 = n2286 & ~n3890 ;
  assign n3892 = n2290 & ~n3891 ;
  assign n3893 = n2836 & ~n3892 ;
  assign n3894 = n602 & ~n3893 ;
  assign n3895 = n606 & ~n3894 ;
  assign n3896 = n610 & ~n3895 ;
  assign n3897 = n614 & ~n3896 ;
  assign n3898 = n618 & ~n3897 ;
  assign n3899 = ~x139 & ~n620 ;
  assign n3900 = ~n3898 & n3899 ;
  assign n3903 = ~n3900 & ~x267 ;
  assign n3904 = ~n3902 & ~n3903 ;
  assign n3905 = n290 & ~n968 ;
  assign n3906 = n295 & ~n3905 ;
  assign n3907 = n299 & ~n3906 ;
  assign n3908 = n303 & ~n3907 ;
  assign n3909 = n307 & ~n3908 ;
  assign n3910 = n311 & ~n3909 ;
  assign n3911 = n315 & ~n3910 ;
  assign n3912 = n319 & ~n3911 ;
  assign n3913 = n323 & ~n3912 ;
  assign n3914 = n327 & ~n3913 ;
  assign n3915 = n331 & ~n3914 ;
  assign n3916 = n335 & ~n3915 ;
  assign n3917 = n339 & ~n3916 ;
  assign n3918 = n343 & ~n3917 ;
  assign n3919 = n347 & ~n3918 ;
  assign n3920 = n351 & ~n3919 ;
  assign n3921 = n355 & ~n3920 ;
  assign n3922 = n359 & ~n3921 ;
  assign n3923 = n363 & ~n3922 ;
  assign n3924 = n367 & ~n3923 ;
  assign n3925 = n371 & ~n3924 ;
  assign n3926 = n375 & ~n3925 ;
  assign n3927 = n379 & ~n3926 ;
  assign n3928 = n383 & ~n3927 ;
  assign n3929 = n387 & ~n3928 ;
  assign n3930 = n391 & ~n3929 ;
  assign n3931 = n395 & ~n3930 ;
  assign n3932 = n399 & ~n3931 ;
  assign n3933 = n403 & ~n3932 ;
  assign n3934 = n407 & ~n3933 ;
  assign n3935 = n411 & ~n3934 ;
  assign n3936 = n415 & ~n3935 ;
  assign n3937 = n419 & ~n3936 ;
  assign n3938 = n423 & ~n3937 ;
  assign n3939 = n427 & ~n3938 ;
  assign n3940 = n431 & ~n3939 ;
  assign n3941 = n435 & ~n3940 ;
  assign n3942 = n439 & ~n3941 ;
  assign n3943 = n443 & ~n3942 ;
  assign n3944 = n447 & ~n3943 ;
  assign n3945 = n451 & ~n3944 ;
  assign n3946 = n455 & ~n3945 ;
  assign n3947 = n459 & ~n3946 ;
  assign n3948 = n463 & ~n3947 ;
  assign n3949 = n467 & ~n3948 ;
  assign n3950 = n471 & ~n3949 ;
  assign n3951 = n475 & ~n3950 ;
  assign n3952 = n479 & ~n3951 ;
  assign n3953 = n483 & ~n3952 ;
  assign n3954 = n487 & ~n3953 ;
  assign n3955 = n491 & ~n3954 ;
  assign n3956 = n495 & ~n3955 ;
  assign n3957 = n499 & ~n3956 ;
  assign n3958 = n503 & ~n3957 ;
  assign n3959 = n507 & ~n3958 ;
  assign n3960 = n511 & ~n3959 ;
  assign n3961 = n515 & ~n3960 ;
  assign n3962 = n519 & ~n3961 ;
  assign n3963 = n523 & ~n3962 ;
  assign n3964 = n527 & ~n3963 ;
  assign n3965 = n531 & ~n3964 ;
  assign n3966 = n535 & ~n3965 ;
  assign n3967 = n539 & ~n3966 ;
  assign n3968 = n543 & ~n3967 ;
  assign n3969 = n547 & ~n3968 ;
  assign n3970 = n551 & ~n3969 ;
  assign n3971 = n555 & ~n3970 ;
  assign n3972 = n559 & ~n3971 ;
  assign n3973 = n563 & ~n3972 ;
  assign n3974 = n567 & ~n3973 ;
  assign n3975 = n571 & ~n3974 ;
  assign n3976 = n575 & ~n3975 ;
  assign n3977 = n579 & ~n3976 ;
  assign n3978 = n583 & ~n3977 ;
  assign n3979 = n587 & ~n3978 ;
  assign n3980 = n591 & ~n3979 ;
  assign n3981 = n2382 & ~n3980 ;
  assign n3982 = n2384 & ~n3981 ;
  assign n3983 = n2927 & ~n3982 ;
  assign n3984 = n945 & ~n3983 ;
  assign n3985 = n949 & ~n3984 ;
  assign n3986 = n953 & ~n3985 ;
  assign n3987 = n957 & ~n3986 ;
  assign n3988 = n961 & ~n3987 ;
  assign n3989 = x140 & ~n963 ;
  assign n3990 = ~n3988 & n3989 ;
  assign n4078 = n3990 & x268 ;
  assign n3991 = n629 & ~n1307 ;
  assign n3992 = n634 & ~n3991 ;
  assign n3993 = n638 & ~n3992 ;
  assign n3994 = n642 & ~n3993 ;
  assign n3995 = n646 & ~n3994 ;
  assign n3996 = n650 & ~n3995 ;
  assign n3997 = n654 & ~n3996 ;
  assign n3998 = n658 & ~n3997 ;
  assign n3999 = n662 & ~n3998 ;
  assign n4000 = n666 & ~n3999 ;
  assign n4001 = n670 & ~n4000 ;
  assign n4002 = n674 & ~n4001 ;
  assign n4003 = n678 & ~n4002 ;
  assign n4004 = n682 & ~n4003 ;
  assign n4005 = n686 & ~n4004 ;
  assign n4006 = n690 & ~n4005 ;
  assign n4007 = n694 & ~n4006 ;
  assign n4008 = n698 & ~n4007 ;
  assign n4009 = n702 & ~n4008 ;
  assign n4010 = n706 & ~n4009 ;
  assign n4011 = n710 & ~n4010 ;
  assign n4012 = n714 & ~n4011 ;
  assign n4013 = n718 & ~n4012 ;
  assign n4014 = n722 & ~n4013 ;
  assign n4015 = n726 & ~n4014 ;
  assign n4016 = n730 & ~n4015 ;
  assign n4017 = n734 & ~n4016 ;
  assign n4018 = n738 & ~n4017 ;
  assign n4019 = n742 & ~n4018 ;
  assign n4020 = n746 & ~n4019 ;
  assign n4021 = n750 & ~n4020 ;
  assign n4022 = n754 & ~n4021 ;
  assign n4023 = n758 & ~n4022 ;
  assign n4024 = n762 & ~n4023 ;
  assign n4025 = n766 & ~n4024 ;
  assign n4026 = n770 & ~n4025 ;
  assign n4027 = n774 & ~n4026 ;
  assign n4028 = n778 & ~n4027 ;
  assign n4029 = n782 & ~n4028 ;
  assign n4030 = n786 & ~n4029 ;
  assign n4031 = n790 & ~n4030 ;
  assign n4032 = n794 & ~n4031 ;
  assign n4033 = n798 & ~n4032 ;
  assign n4034 = n802 & ~n4033 ;
  assign n4035 = n806 & ~n4034 ;
  assign n4036 = n810 & ~n4035 ;
  assign n4037 = n814 & ~n4036 ;
  assign n4038 = n818 & ~n4037 ;
  assign n4039 = n822 & ~n4038 ;
  assign n4040 = n826 & ~n4039 ;
  assign n4041 = n830 & ~n4040 ;
  assign n4042 = n834 & ~n4041 ;
  assign n4043 = n838 & ~n4042 ;
  assign n4044 = n842 & ~n4043 ;
  assign n4045 = n846 & ~n4044 ;
  assign n4046 = n850 & ~n4045 ;
  assign n4047 = n854 & ~n4046 ;
  assign n4048 = n858 & ~n4047 ;
  assign n4049 = n862 & ~n4048 ;
  assign n4050 = n866 & ~n4049 ;
  assign n4051 = n870 & ~n4050 ;
  assign n4052 = n874 & ~n4051 ;
  assign n4053 = n878 & ~n4052 ;
  assign n4054 = n882 & ~n4053 ;
  assign n4055 = n886 & ~n4054 ;
  assign n4056 = n890 & ~n4055 ;
  assign n4057 = n894 & ~n4056 ;
  assign n4058 = n898 & ~n4057 ;
  assign n4059 = n902 & ~n4058 ;
  assign n4060 = n906 & ~n4059 ;
  assign n4061 = n910 & ~n4060 ;
  assign n4062 = n914 & ~n4061 ;
  assign n4063 = n918 & ~n4062 ;
  assign n4064 = n922 & ~n4063 ;
  assign n4065 = n926 & ~n4064 ;
  assign n4066 = n930 & ~n4065 ;
  assign n4067 = n2472 & ~n4066 ;
  assign n4068 = n2474 & ~n4067 ;
  assign n4069 = n3014 & ~n4068 ;
  assign n4070 = n1284 & ~n4069 ;
  assign n4071 = n1288 & ~n4070 ;
  assign n4072 = n1292 & ~n4071 ;
  assign n4073 = n1296 & ~n4072 ;
  assign n4074 = n1300 & ~n4073 ;
  assign n4075 = ~x140 & ~n1302 ;
  assign n4076 = ~n4074 & n4075 ;
  assign n4079 = ~n4076 & ~x268 ;
  assign n4080 = ~n4078 & ~n4079 ;
  assign n4081 = n972 & ~n1648 ;
  assign n4082 = n977 & ~n4081 ;
  assign n4083 = n981 & ~n4082 ;
  assign n4084 = n985 & ~n4083 ;
  assign n4085 = n989 & ~n4084 ;
  assign n4086 = n993 & ~n4085 ;
  assign n4087 = n997 & ~n4086 ;
  assign n4088 = n1001 & ~n4087 ;
  assign n4089 = n1005 & ~n4088 ;
  assign n4090 = n1009 & ~n4089 ;
  assign n4091 = n1013 & ~n4090 ;
  assign n4092 = n1017 & ~n4091 ;
  assign n4093 = n1021 & ~n4092 ;
  assign n4094 = n1025 & ~n4093 ;
  assign n4095 = n1029 & ~n4094 ;
  assign n4096 = n1033 & ~n4095 ;
  assign n4097 = n1037 & ~n4096 ;
  assign n4098 = n1041 & ~n4097 ;
  assign n4099 = n1045 & ~n4098 ;
  assign n4100 = n1049 & ~n4099 ;
  assign n4101 = n1053 & ~n4100 ;
  assign n4102 = n1057 & ~n4101 ;
  assign n4103 = n1061 & ~n4102 ;
  assign n4104 = n1065 & ~n4103 ;
  assign n4105 = n1069 & ~n4104 ;
  assign n4106 = n1073 & ~n4105 ;
  assign n4107 = n1077 & ~n4106 ;
  assign n4108 = n1081 & ~n4107 ;
  assign n4109 = n1085 & ~n4108 ;
  assign n4110 = n1089 & ~n4109 ;
  assign n4111 = n1093 & ~n4110 ;
  assign n4112 = n1097 & ~n4111 ;
  assign n4113 = n1101 & ~n4112 ;
  assign n4114 = n1105 & ~n4113 ;
  assign n4115 = n1109 & ~n4114 ;
  assign n4116 = n1113 & ~n4115 ;
  assign n4117 = n1117 & ~n4116 ;
  assign n4118 = n1121 & ~n4117 ;
  assign n4119 = n1125 & ~n4118 ;
  assign n4120 = n1129 & ~n4119 ;
  assign n4121 = n1133 & ~n4120 ;
  assign n4122 = n1137 & ~n4121 ;
  assign n4123 = n1141 & ~n4122 ;
  assign n4124 = n1145 & ~n4123 ;
  assign n4125 = n1149 & ~n4124 ;
  assign n4126 = n1153 & ~n4125 ;
  assign n4127 = n1157 & ~n4126 ;
  assign n4128 = n1161 & ~n4127 ;
  assign n4129 = n1165 & ~n4128 ;
  assign n4130 = n1169 & ~n4129 ;
  assign n4131 = n1173 & ~n4130 ;
  assign n4132 = n1177 & ~n4131 ;
  assign n4133 = n1181 & ~n4132 ;
  assign n4134 = n1185 & ~n4133 ;
  assign n4135 = n1189 & ~n4134 ;
  assign n4136 = n1193 & ~n4135 ;
  assign n4137 = n1197 & ~n4136 ;
  assign n4138 = n1201 & ~n4137 ;
  assign n4139 = n1205 & ~n4138 ;
  assign n4140 = n1209 & ~n4139 ;
  assign n4141 = n1213 & ~n4140 ;
  assign n4142 = n1217 & ~n4141 ;
  assign n4143 = n1221 & ~n4142 ;
  assign n4144 = n1225 & ~n4143 ;
  assign n4145 = n1229 & ~n4144 ;
  assign n4146 = n1233 & ~n4145 ;
  assign n4147 = n1237 & ~n4146 ;
  assign n4148 = n1241 & ~n4147 ;
  assign n4149 = n1245 & ~n4148 ;
  assign n4150 = n1249 & ~n4149 ;
  assign n4151 = n1253 & ~n4150 ;
  assign n4152 = n1257 & ~n4151 ;
  assign n4153 = n1261 & ~n4152 ;
  assign n4154 = n1265 & ~n4153 ;
  assign n4155 = n1269 & ~n4154 ;
  assign n4156 = n1273 & ~n4155 ;
  assign n4157 = n2566 & ~n4156 ;
  assign n4158 = n2568 & ~n4157 ;
  assign n4159 = n3105 & ~n4158 ;
  assign n4160 = n1625 & ~n4159 ;
  assign n4161 = n1629 & ~n4160 ;
  assign n4162 = n1633 & ~n4161 ;
  assign n4163 = n1637 & ~n4162 ;
  assign n4164 = n1641 & ~n4163 ;
  assign n4165 = x141 & ~n1643 ;
  assign n4166 = ~n4164 & n4165 ;
  assign n4254 = n4166 & x269 ;
  assign n4167 = n1311 & ~n1985 ;
  assign n4168 = n1316 & ~n4167 ;
  assign n4169 = n1320 & ~n4168 ;
  assign n4170 = n1324 & ~n4169 ;
  assign n4171 = n1328 & ~n4170 ;
  assign n4172 = n1332 & ~n4171 ;
  assign n4173 = n1336 & ~n4172 ;
  assign n4174 = n1340 & ~n4173 ;
  assign n4175 = n1344 & ~n4174 ;
  assign n4176 = n1348 & ~n4175 ;
  assign n4177 = n1352 & ~n4176 ;
  assign n4178 = n1356 & ~n4177 ;
  assign n4179 = n1360 & ~n4178 ;
  assign n4180 = n1364 & ~n4179 ;
  assign n4181 = n1368 & ~n4180 ;
  assign n4182 = n1372 & ~n4181 ;
  assign n4183 = n1376 & ~n4182 ;
  assign n4184 = n1380 & ~n4183 ;
  assign n4185 = n1384 & ~n4184 ;
  assign n4186 = n1388 & ~n4185 ;
  assign n4187 = n1392 & ~n4186 ;
  assign n4188 = n1396 & ~n4187 ;
  assign n4189 = n1400 & ~n4188 ;
  assign n4190 = n1404 & ~n4189 ;
  assign n4191 = n1408 & ~n4190 ;
  assign n4192 = n1412 & ~n4191 ;
  assign n4193 = n1416 & ~n4192 ;
  assign n4194 = n1420 & ~n4193 ;
  assign n4195 = n1424 & ~n4194 ;
  assign n4196 = n1428 & ~n4195 ;
  assign n4197 = n1432 & ~n4196 ;
  assign n4198 = n1436 & ~n4197 ;
  assign n4199 = n1440 & ~n4198 ;
  assign n4200 = n1444 & ~n4199 ;
  assign n4201 = n1448 & ~n4200 ;
  assign n4202 = n1452 & ~n4201 ;
  assign n4203 = n1456 & ~n4202 ;
  assign n4204 = n1460 & ~n4203 ;
  assign n4205 = n1464 & ~n4204 ;
  assign n4206 = n1468 & ~n4205 ;
  assign n4207 = n1472 & ~n4206 ;
  assign n4208 = n1476 & ~n4207 ;
  assign n4209 = n1480 & ~n4208 ;
  assign n4210 = n1484 & ~n4209 ;
  assign n4211 = n1488 & ~n4210 ;
  assign n4212 = n1492 & ~n4211 ;
  assign n4213 = n1496 & ~n4212 ;
  assign n4214 = n1500 & ~n4213 ;
  assign n4215 = n1504 & ~n4214 ;
  assign n4216 = n1508 & ~n4215 ;
  assign n4217 = n1512 & ~n4216 ;
  assign n4218 = n1516 & ~n4217 ;
  assign n4219 = n1520 & ~n4218 ;
  assign n4220 = n1524 & ~n4219 ;
  assign n4221 = n1528 & ~n4220 ;
  assign n4222 = n1532 & ~n4221 ;
  assign n4223 = n1536 & ~n4222 ;
  assign n4224 = n1540 & ~n4223 ;
  assign n4225 = n1544 & ~n4224 ;
  assign n4226 = n1548 & ~n4225 ;
  assign n4227 = n1552 & ~n4226 ;
  assign n4228 = n1556 & ~n4227 ;
  assign n4229 = n1560 & ~n4228 ;
  assign n4230 = n1564 & ~n4229 ;
  assign n4231 = n1568 & ~n4230 ;
  assign n4232 = n1572 & ~n4231 ;
  assign n4233 = n1576 & ~n4232 ;
  assign n4234 = n1580 & ~n4233 ;
  assign n4235 = n1584 & ~n4234 ;
  assign n4236 = n1588 & ~n4235 ;
  assign n4237 = n1592 & ~n4236 ;
  assign n4238 = n1596 & ~n4237 ;
  assign n4239 = n1600 & ~n4238 ;
  assign n4240 = n1604 & ~n4239 ;
  assign n4241 = n1608 & ~n4240 ;
  assign n4242 = n1612 & ~n4241 ;
  assign n4243 = n2656 & ~n4242 ;
  assign n4244 = n2658 & ~n4243 ;
  assign n4245 = n3192 & ~n4244 ;
  assign n4246 = n1962 & ~n4245 ;
  assign n4247 = n1966 & ~n4246 ;
  assign n4248 = n1970 & ~n4247 ;
  assign n4249 = n1974 & ~n4248 ;
  assign n4250 = n1978 & ~n4249 ;
  assign n4251 = ~x141 & ~n1980 ;
  assign n4252 = ~n4250 & n4251 ;
  assign n4255 = ~n4252 & ~x269 ;
  assign n4256 = ~n4254 & ~n4255 ;
  assign n4257 = ~n294 & n1652 ;
  assign n4258 = n1657 & ~n4257 ;
  assign n4259 = n1661 & ~n4258 ;
  assign n4260 = n1665 & ~n4259 ;
  assign n4261 = n1669 & ~n4260 ;
  assign n4262 = n1673 & ~n4261 ;
  assign n4263 = n1677 & ~n4262 ;
  assign n4264 = n1681 & ~n4263 ;
  assign n4265 = n1685 & ~n4264 ;
  assign n4266 = n1689 & ~n4265 ;
  assign n4267 = n1693 & ~n4266 ;
  assign n4268 = n1697 & ~n4267 ;
  assign n4269 = n1701 & ~n4268 ;
  assign n4270 = n1705 & ~n4269 ;
  assign n4271 = n1709 & ~n4270 ;
  assign n4272 = n1713 & ~n4271 ;
  assign n4273 = n1717 & ~n4272 ;
  assign n4274 = n1721 & ~n4273 ;
  assign n4275 = n1725 & ~n4274 ;
  assign n4276 = n1729 & ~n4275 ;
  assign n4277 = n1733 & ~n4276 ;
  assign n4278 = n1737 & ~n4277 ;
  assign n4279 = n1741 & ~n4278 ;
  assign n4280 = n1745 & ~n4279 ;
  assign n4281 = n1749 & ~n4280 ;
  assign n4282 = n1753 & ~n4281 ;
  assign n4283 = n1757 & ~n4282 ;
  assign n4284 = n1761 & ~n4283 ;
  assign n4285 = n1765 & ~n4284 ;
  assign n4286 = n1769 & ~n4285 ;
  assign n4287 = n1773 & ~n4286 ;
  assign n4288 = n1777 & ~n4287 ;
  assign n4289 = n1781 & ~n4288 ;
  assign n4290 = n1785 & ~n4289 ;
  assign n4291 = n1789 & ~n4290 ;
  assign n4292 = n1793 & ~n4291 ;
  assign n4293 = n1797 & ~n4292 ;
  assign n4294 = n1801 & ~n4293 ;
  assign n4295 = n1805 & ~n4294 ;
  assign n4296 = n1809 & ~n4295 ;
  assign n4297 = n1813 & ~n4296 ;
  assign n4298 = n1817 & ~n4297 ;
  assign n4299 = n1821 & ~n4298 ;
  assign n4300 = n1825 & ~n4299 ;
  assign n4301 = n1829 & ~n4300 ;
  assign n4302 = n1833 & ~n4301 ;
  assign n4303 = n1837 & ~n4302 ;
  assign n4304 = n1841 & ~n4303 ;
  assign n4305 = n1845 & ~n4304 ;
  assign n4306 = n1849 & ~n4305 ;
  assign n4307 = n1853 & ~n4306 ;
  assign n4308 = n1857 & ~n4307 ;
  assign n4309 = n1861 & ~n4308 ;
  assign n4310 = n1865 & ~n4309 ;
  assign n4311 = n1869 & ~n4310 ;
  assign n4312 = n1873 & ~n4311 ;
  assign n4313 = n1877 & ~n4312 ;
  assign n4314 = n1881 & ~n4313 ;
  assign n4315 = n1885 & ~n4314 ;
  assign n4316 = n1889 & ~n4315 ;
  assign n4317 = n1893 & ~n4316 ;
  assign n4318 = n1897 & ~n4317 ;
  assign n4319 = n1901 & ~n4318 ;
  assign n4320 = n1905 & ~n4319 ;
  assign n4321 = n1909 & ~n4320 ;
  assign n4322 = n1913 & ~n4321 ;
  assign n4323 = n1917 & ~n4322 ;
  assign n4324 = n1921 & ~n4323 ;
  assign n4325 = n1925 & ~n4324 ;
  assign n4326 = n1929 & ~n4325 ;
  assign n4327 = n1933 & ~n4326 ;
  assign n4328 = n1937 & ~n4327 ;
  assign n4329 = n1941 & ~n4328 ;
  assign n4330 = n1945 & ~n4329 ;
  assign n4331 = n1949 & ~n4330 ;
  assign n4332 = n1953 & ~n4331 ;
  assign n4333 = n2749 & ~n4332 ;
  assign n4334 = n263 & ~n4333 ;
  assign n4335 = n267 & ~n4334 ;
  assign n4336 = n271 & ~n4335 ;
  assign n4337 = n275 & ~n4336 ;
  assign n4338 = n279 & ~n4337 ;
  assign n4339 = n283 & ~n4338 ;
  assign n4340 = n287 & ~n4339 ;
  assign n4341 = x142 & ~n289 ;
  assign n4342 = ~n4340 & n4341 ;
  assign n4430 = n4342 & x270 ;
  assign n4343 = ~n633 & n1989 ;
  assign n4344 = n1994 & ~n4343 ;
  assign n4345 = n1998 & ~n4344 ;
  assign n4346 = n2002 & ~n4345 ;
  assign n4347 = n2006 & ~n4346 ;
  assign n4348 = n2010 & ~n4347 ;
  assign n4349 = n2014 & ~n4348 ;
  assign n4350 = n2018 & ~n4349 ;
  assign n4351 = n2022 & ~n4350 ;
  assign n4352 = n2026 & ~n4351 ;
  assign n4353 = n2030 & ~n4352 ;
  assign n4354 = n2034 & ~n4353 ;
  assign n4355 = n2038 & ~n4354 ;
  assign n4356 = n2042 & ~n4355 ;
  assign n4357 = n2046 & ~n4356 ;
  assign n4358 = n2050 & ~n4357 ;
  assign n4359 = n2054 & ~n4358 ;
  assign n4360 = n2058 & ~n4359 ;
  assign n4361 = n2062 & ~n4360 ;
  assign n4362 = n2066 & ~n4361 ;
  assign n4363 = n2070 & ~n4362 ;
  assign n4364 = n2074 & ~n4363 ;
  assign n4365 = n2078 & ~n4364 ;
  assign n4366 = n2082 & ~n4365 ;
  assign n4367 = n2086 & ~n4366 ;
  assign n4368 = n2090 & ~n4367 ;
  assign n4369 = n2094 & ~n4368 ;
  assign n4370 = n2098 & ~n4369 ;
  assign n4371 = n2102 & ~n4370 ;
  assign n4372 = n2106 & ~n4371 ;
  assign n4373 = n2110 & ~n4372 ;
  assign n4374 = n2114 & ~n4373 ;
  assign n4375 = n2118 & ~n4374 ;
  assign n4376 = n2122 & ~n4375 ;
  assign n4377 = n2126 & ~n4376 ;
  assign n4378 = n2130 & ~n4377 ;
  assign n4379 = n2134 & ~n4378 ;
  assign n4380 = n2138 & ~n4379 ;
  assign n4381 = n2142 & ~n4380 ;
  assign n4382 = n2146 & ~n4381 ;
  assign n4383 = n2150 & ~n4382 ;
  assign n4384 = n2154 & ~n4383 ;
  assign n4385 = n2158 & ~n4384 ;
  assign n4386 = n2162 & ~n4385 ;
  assign n4387 = n2166 & ~n4386 ;
  assign n4388 = n2170 & ~n4387 ;
  assign n4389 = n2174 & ~n4388 ;
  assign n4390 = n2178 & ~n4389 ;
  assign n4391 = n2182 & ~n4390 ;
  assign n4392 = n2186 & ~n4391 ;
  assign n4393 = n2190 & ~n4392 ;
  assign n4394 = n2194 & ~n4393 ;
  assign n4395 = n2198 & ~n4394 ;
  assign n4396 = n2202 & ~n4395 ;
  assign n4397 = n2206 & ~n4396 ;
  assign n4398 = n2210 & ~n4397 ;
  assign n4399 = n2214 & ~n4398 ;
  assign n4400 = n2218 & ~n4399 ;
  assign n4401 = n2222 & ~n4400 ;
  assign n4402 = n2226 & ~n4401 ;
  assign n4403 = n2230 & ~n4402 ;
  assign n4404 = n2234 & ~n4403 ;
  assign n4405 = n2238 & ~n4404 ;
  assign n4406 = n2242 & ~n4405 ;
  assign n4407 = n2246 & ~n4406 ;
  assign n4408 = n2250 & ~n4407 ;
  assign n4409 = n2254 & ~n4408 ;
  assign n4410 = n2258 & ~n4409 ;
  assign n4411 = n2262 & ~n4410 ;
  assign n4412 = n2266 & ~n4411 ;
  assign n4413 = n2270 & ~n4412 ;
  assign n4414 = n2274 & ~n4413 ;
  assign n4415 = n2278 & ~n4414 ;
  assign n4416 = n2282 & ~n4415 ;
  assign n4417 = n2286 & ~n4416 ;
  assign n4418 = n2290 & ~n4417 ;
  assign n4419 = n2836 & ~n4418 ;
  assign n4420 = n602 & ~n4419 ;
  assign n4421 = n606 & ~n4420 ;
  assign n4422 = n610 & ~n4421 ;
  assign n4423 = n614 & ~n4422 ;
  assign n4424 = n618 & ~n4423 ;
  assign n4425 = n622 & ~n4424 ;
  assign n4426 = n626 & ~n4425 ;
  assign n4427 = ~x142 & ~n628 ;
  assign n4428 = ~n4426 & n4427 ;
  assign n4431 = ~n4428 & ~x270 ;
  assign n4432 = ~n4430 & ~n4431 ;
  assign n4433 = n298 & ~n976 ;
  assign n4434 = n303 & ~n4433 ;
  assign n4435 = n307 & ~n4434 ;
  assign n4436 = n311 & ~n4435 ;
  assign n4437 = n315 & ~n4436 ;
  assign n4438 = n319 & ~n4437 ;
  assign n4439 = n323 & ~n4438 ;
  assign n4440 = n327 & ~n4439 ;
  assign n4441 = n331 & ~n4440 ;
  assign n4442 = n335 & ~n4441 ;
  assign n4443 = n339 & ~n4442 ;
  assign n4444 = n343 & ~n4443 ;
  assign n4445 = n347 & ~n4444 ;
  assign n4446 = n351 & ~n4445 ;
  assign n4447 = n355 & ~n4446 ;
  assign n4448 = n359 & ~n4447 ;
  assign n4449 = n363 & ~n4448 ;
  assign n4450 = n367 & ~n4449 ;
  assign n4451 = n371 & ~n4450 ;
  assign n4452 = n375 & ~n4451 ;
  assign n4453 = n379 & ~n4452 ;
  assign n4454 = n383 & ~n4453 ;
  assign n4455 = n387 & ~n4454 ;
  assign n4456 = n391 & ~n4455 ;
  assign n4457 = n395 & ~n4456 ;
  assign n4458 = n399 & ~n4457 ;
  assign n4459 = n403 & ~n4458 ;
  assign n4460 = n407 & ~n4459 ;
  assign n4461 = n411 & ~n4460 ;
  assign n4462 = n415 & ~n4461 ;
  assign n4463 = n419 & ~n4462 ;
  assign n4464 = n423 & ~n4463 ;
  assign n4465 = n427 & ~n4464 ;
  assign n4466 = n431 & ~n4465 ;
  assign n4467 = n435 & ~n4466 ;
  assign n4468 = n439 & ~n4467 ;
  assign n4469 = n443 & ~n4468 ;
  assign n4470 = n447 & ~n4469 ;
  assign n4471 = n451 & ~n4470 ;
  assign n4472 = n455 & ~n4471 ;
  assign n4473 = n459 & ~n4472 ;
  assign n4474 = n463 & ~n4473 ;
  assign n4475 = n467 & ~n4474 ;
  assign n4476 = n471 & ~n4475 ;
  assign n4477 = n475 & ~n4476 ;
  assign n4478 = n479 & ~n4477 ;
  assign n4479 = n483 & ~n4478 ;
  assign n4480 = n487 & ~n4479 ;
  assign n4481 = n491 & ~n4480 ;
  assign n4482 = n495 & ~n4481 ;
  assign n4483 = n499 & ~n4482 ;
  assign n4484 = n503 & ~n4483 ;
  assign n4485 = n507 & ~n4484 ;
  assign n4486 = n511 & ~n4485 ;
  assign n4487 = n515 & ~n4486 ;
  assign n4488 = n519 & ~n4487 ;
  assign n4489 = n523 & ~n4488 ;
  assign n4490 = n527 & ~n4489 ;
  assign n4491 = n531 & ~n4490 ;
  assign n4492 = n535 & ~n4491 ;
  assign n4493 = n539 & ~n4492 ;
  assign n4494 = n543 & ~n4493 ;
  assign n4495 = n547 & ~n4494 ;
  assign n4496 = n551 & ~n4495 ;
  assign n4497 = n555 & ~n4496 ;
  assign n4498 = n559 & ~n4497 ;
  assign n4499 = n563 & ~n4498 ;
  assign n4500 = n567 & ~n4499 ;
  assign n4501 = n571 & ~n4500 ;
  assign n4502 = n575 & ~n4501 ;
  assign n4503 = n579 & ~n4502 ;
  assign n4504 = n583 & ~n4503 ;
  assign n4505 = n587 & ~n4504 ;
  assign n4506 = n591 & ~n4505 ;
  assign n4507 = n2382 & ~n4506 ;
  assign n4508 = n2384 & ~n4507 ;
  assign n4509 = n2927 & ~n4508 ;
  assign n4510 = n945 & ~n4509 ;
  assign n4511 = n949 & ~n4510 ;
  assign n4512 = n953 & ~n4511 ;
  assign n4513 = n957 & ~n4512 ;
  assign n4514 = n961 & ~n4513 ;
  assign n4515 = n965 & ~n4514 ;
  assign n4516 = n969 & ~n4515 ;
  assign n4517 = x143 & ~n971 ;
  assign n4518 = ~n4516 & n4517 ;
  assign n4606 = n4518 & x271 ;
  assign n4519 = n637 & ~n1315 ;
  assign n4520 = n642 & ~n4519 ;
  assign n4521 = n646 & ~n4520 ;
  assign n4522 = n650 & ~n4521 ;
  assign n4523 = n654 & ~n4522 ;
  assign n4524 = n658 & ~n4523 ;
  assign n4525 = n662 & ~n4524 ;
  assign n4526 = n666 & ~n4525 ;
  assign n4527 = n670 & ~n4526 ;
  assign n4528 = n674 & ~n4527 ;
  assign n4529 = n678 & ~n4528 ;
  assign n4530 = n682 & ~n4529 ;
  assign n4531 = n686 & ~n4530 ;
  assign n4532 = n690 & ~n4531 ;
  assign n4533 = n694 & ~n4532 ;
  assign n4534 = n698 & ~n4533 ;
  assign n4535 = n702 & ~n4534 ;
  assign n4536 = n706 & ~n4535 ;
  assign n4537 = n710 & ~n4536 ;
  assign n4538 = n714 & ~n4537 ;
  assign n4539 = n718 & ~n4538 ;
  assign n4540 = n722 & ~n4539 ;
  assign n4541 = n726 & ~n4540 ;
  assign n4542 = n730 & ~n4541 ;
  assign n4543 = n734 & ~n4542 ;
  assign n4544 = n738 & ~n4543 ;
  assign n4545 = n742 & ~n4544 ;
  assign n4546 = n746 & ~n4545 ;
  assign n4547 = n750 & ~n4546 ;
  assign n4548 = n754 & ~n4547 ;
  assign n4549 = n758 & ~n4548 ;
  assign n4550 = n762 & ~n4549 ;
  assign n4551 = n766 & ~n4550 ;
  assign n4552 = n770 & ~n4551 ;
  assign n4553 = n774 & ~n4552 ;
  assign n4554 = n778 & ~n4553 ;
  assign n4555 = n782 & ~n4554 ;
  assign n4556 = n786 & ~n4555 ;
  assign n4557 = n790 & ~n4556 ;
  assign n4558 = n794 & ~n4557 ;
  assign n4559 = n798 & ~n4558 ;
  assign n4560 = n802 & ~n4559 ;
  assign n4561 = n806 & ~n4560 ;
  assign n4562 = n810 & ~n4561 ;
  assign n4563 = n814 & ~n4562 ;
  assign n4564 = n818 & ~n4563 ;
  assign n4565 = n822 & ~n4564 ;
  assign n4566 = n826 & ~n4565 ;
  assign n4567 = n830 & ~n4566 ;
  assign n4568 = n834 & ~n4567 ;
  assign n4569 = n838 & ~n4568 ;
  assign n4570 = n842 & ~n4569 ;
  assign n4571 = n846 & ~n4570 ;
  assign n4572 = n850 & ~n4571 ;
  assign n4573 = n854 & ~n4572 ;
  assign n4574 = n858 & ~n4573 ;
  assign n4575 = n862 & ~n4574 ;
  assign n4576 = n866 & ~n4575 ;
  assign n4577 = n870 & ~n4576 ;
  assign n4578 = n874 & ~n4577 ;
  assign n4579 = n878 & ~n4578 ;
  assign n4580 = n882 & ~n4579 ;
  assign n4581 = n886 & ~n4580 ;
  assign n4582 = n890 & ~n4581 ;
  assign n4583 = n894 & ~n4582 ;
  assign n4584 = n898 & ~n4583 ;
  assign n4585 = n902 & ~n4584 ;
  assign n4586 = n906 & ~n4585 ;
  assign n4587 = n910 & ~n4586 ;
  assign n4588 = n914 & ~n4587 ;
  assign n4589 = n918 & ~n4588 ;
  assign n4590 = n922 & ~n4589 ;
  assign n4591 = n926 & ~n4590 ;
  assign n4592 = n930 & ~n4591 ;
  assign n4593 = n2472 & ~n4592 ;
  assign n4594 = n2474 & ~n4593 ;
  assign n4595 = n3014 & ~n4594 ;
  assign n4596 = n1284 & ~n4595 ;
  assign n4597 = n1288 & ~n4596 ;
  assign n4598 = n1292 & ~n4597 ;
  assign n4599 = n1296 & ~n4598 ;
  assign n4600 = n1300 & ~n4599 ;
  assign n4601 = n1304 & ~n4600 ;
  assign n4602 = n1308 & ~n4601 ;
  assign n4603 = ~x143 & ~n1310 ;
  assign n4604 = ~n4602 & n4603 ;
  assign n4607 = ~n4604 & ~x271 ;
  assign n4608 = ~n4606 & ~n4607 ;
  assign n4609 = n980 & ~n1656 ;
  assign n4610 = n985 & ~n4609 ;
  assign n4611 = n989 & ~n4610 ;
  assign n4612 = n993 & ~n4611 ;
  assign n4613 = n997 & ~n4612 ;
  assign n4614 = n1001 & ~n4613 ;
  assign n4615 = n1005 & ~n4614 ;
  assign n4616 = n1009 & ~n4615 ;
  assign n4617 = n1013 & ~n4616 ;
  assign n4618 = n1017 & ~n4617 ;
  assign n4619 = n1021 & ~n4618 ;
  assign n4620 = n1025 & ~n4619 ;
  assign n4621 = n1029 & ~n4620 ;
  assign n4622 = n1033 & ~n4621 ;
  assign n4623 = n1037 & ~n4622 ;
  assign n4624 = n1041 & ~n4623 ;
  assign n4625 = n1045 & ~n4624 ;
  assign n4626 = n1049 & ~n4625 ;
  assign n4627 = n1053 & ~n4626 ;
  assign n4628 = n1057 & ~n4627 ;
  assign n4629 = n1061 & ~n4628 ;
  assign n4630 = n1065 & ~n4629 ;
  assign n4631 = n1069 & ~n4630 ;
  assign n4632 = n1073 & ~n4631 ;
  assign n4633 = n1077 & ~n4632 ;
  assign n4634 = n1081 & ~n4633 ;
  assign n4635 = n1085 & ~n4634 ;
  assign n4636 = n1089 & ~n4635 ;
  assign n4637 = n1093 & ~n4636 ;
  assign n4638 = n1097 & ~n4637 ;
  assign n4639 = n1101 & ~n4638 ;
  assign n4640 = n1105 & ~n4639 ;
  assign n4641 = n1109 & ~n4640 ;
  assign n4642 = n1113 & ~n4641 ;
  assign n4643 = n1117 & ~n4642 ;
  assign n4644 = n1121 & ~n4643 ;
  assign n4645 = n1125 & ~n4644 ;
  assign n4646 = n1129 & ~n4645 ;
  assign n4647 = n1133 & ~n4646 ;
  assign n4648 = n1137 & ~n4647 ;
  assign n4649 = n1141 & ~n4648 ;
  assign n4650 = n1145 & ~n4649 ;
  assign n4651 = n1149 & ~n4650 ;
  assign n4652 = n1153 & ~n4651 ;
  assign n4653 = n1157 & ~n4652 ;
  assign n4654 = n1161 & ~n4653 ;
  assign n4655 = n1165 & ~n4654 ;
  assign n4656 = n1169 & ~n4655 ;
  assign n4657 = n1173 & ~n4656 ;
  assign n4658 = n1177 & ~n4657 ;
  assign n4659 = n1181 & ~n4658 ;
  assign n4660 = n1185 & ~n4659 ;
  assign n4661 = n1189 & ~n4660 ;
  assign n4662 = n1193 & ~n4661 ;
  assign n4663 = n1197 & ~n4662 ;
  assign n4664 = n1201 & ~n4663 ;
  assign n4665 = n1205 & ~n4664 ;
  assign n4666 = n1209 & ~n4665 ;
  assign n4667 = n1213 & ~n4666 ;
  assign n4668 = n1217 & ~n4667 ;
  assign n4669 = n1221 & ~n4668 ;
  assign n4670 = n1225 & ~n4669 ;
  assign n4671 = n1229 & ~n4670 ;
  assign n4672 = n1233 & ~n4671 ;
  assign n4673 = n1237 & ~n4672 ;
  assign n4674 = n1241 & ~n4673 ;
  assign n4675 = n1245 & ~n4674 ;
  assign n4676 = n1249 & ~n4675 ;
  assign n4677 = n1253 & ~n4676 ;
  assign n4678 = n1257 & ~n4677 ;
  assign n4679 = n1261 & ~n4678 ;
  assign n4680 = n1265 & ~n4679 ;
  assign n4681 = n1269 & ~n4680 ;
  assign n4682 = n1273 & ~n4681 ;
  assign n4683 = n2566 & ~n4682 ;
  assign n4684 = n2568 & ~n4683 ;
  assign n4685 = n3105 & ~n4684 ;
  assign n4686 = n1625 & ~n4685 ;
  assign n4687 = n1629 & ~n4686 ;
  assign n4688 = n1633 & ~n4687 ;
  assign n4689 = n1637 & ~n4688 ;
  assign n4690 = n1641 & ~n4689 ;
  assign n4691 = n1645 & ~n4690 ;
  assign n4692 = n1649 & ~n4691 ;
  assign n4693 = x144 & ~n1651 ;
  assign n4694 = ~n4692 & n4693 ;
  assign n4782 = n4694 & x272 ;
  assign n4695 = n1319 & ~n1993 ;
  assign n4696 = n1324 & ~n4695 ;
  assign n4697 = n1328 & ~n4696 ;
  assign n4698 = n1332 & ~n4697 ;
  assign n4699 = n1336 & ~n4698 ;
  assign n4700 = n1340 & ~n4699 ;
  assign n4701 = n1344 & ~n4700 ;
  assign n4702 = n1348 & ~n4701 ;
  assign n4703 = n1352 & ~n4702 ;
  assign n4704 = n1356 & ~n4703 ;
  assign n4705 = n1360 & ~n4704 ;
  assign n4706 = n1364 & ~n4705 ;
  assign n4707 = n1368 & ~n4706 ;
  assign n4708 = n1372 & ~n4707 ;
  assign n4709 = n1376 & ~n4708 ;
  assign n4710 = n1380 & ~n4709 ;
  assign n4711 = n1384 & ~n4710 ;
  assign n4712 = n1388 & ~n4711 ;
  assign n4713 = n1392 & ~n4712 ;
  assign n4714 = n1396 & ~n4713 ;
  assign n4715 = n1400 & ~n4714 ;
  assign n4716 = n1404 & ~n4715 ;
  assign n4717 = n1408 & ~n4716 ;
  assign n4718 = n1412 & ~n4717 ;
  assign n4719 = n1416 & ~n4718 ;
  assign n4720 = n1420 & ~n4719 ;
  assign n4721 = n1424 & ~n4720 ;
  assign n4722 = n1428 & ~n4721 ;
  assign n4723 = n1432 & ~n4722 ;
  assign n4724 = n1436 & ~n4723 ;
  assign n4725 = n1440 & ~n4724 ;
  assign n4726 = n1444 & ~n4725 ;
  assign n4727 = n1448 & ~n4726 ;
  assign n4728 = n1452 & ~n4727 ;
  assign n4729 = n1456 & ~n4728 ;
  assign n4730 = n1460 & ~n4729 ;
  assign n4731 = n1464 & ~n4730 ;
  assign n4732 = n1468 & ~n4731 ;
  assign n4733 = n1472 & ~n4732 ;
  assign n4734 = n1476 & ~n4733 ;
  assign n4735 = n1480 & ~n4734 ;
  assign n4736 = n1484 & ~n4735 ;
  assign n4737 = n1488 & ~n4736 ;
  assign n4738 = n1492 & ~n4737 ;
  assign n4739 = n1496 & ~n4738 ;
  assign n4740 = n1500 & ~n4739 ;
  assign n4741 = n1504 & ~n4740 ;
  assign n4742 = n1508 & ~n4741 ;
  assign n4743 = n1512 & ~n4742 ;
  assign n4744 = n1516 & ~n4743 ;
  assign n4745 = n1520 & ~n4744 ;
  assign n4746 = n1524 & ~n4745 ;
  assign n4747 = n1528 & ~n4746 ;
  assign n4748 = n1532 & ~n4747 ;
  assign n4749 = n1536 & ~n4748 ;
  assign n4750 = n1540 & ~n4749 ;
  assign n4751 = n1544 & ~n4750 ;
  assign n4752 = n1548 & ~n4751 ;
  assign n4753 = n1552 & ~n4752 ;
  assign n4754 = n1556 & ~n4753 ;
  assign n4755 = n1560 & ~n4754 ;
  assign n4756 = n1564 & ~n4755 ;
  assign n4757 = n1568 & ~n4756 ;
  assign n4758 = n1572 & ~n4757 ;
  assign n4759 = n1576 & ~n4758 ;
  assign n4760 = n1580 & ~n4759 ;
  assign n4761 = n1584 & ~n4760 ;
  assign n4762 = n1588 & ~n4761 ;
  assign n4763 = n1592 & ~n4762 ;
  assign n4764 = n1596 & ~n4763 ;
  assign n4765 = n1600 & ~n4764 ;
  assign n4766 = n1604 & ~n4765 ;
  assign n4767 = n1608 & ~n4766 ;
  assign n4768 = n1612 & ~n4767 ;
  assign n4769 = n2656 & ~n4768 ;
  assign n4770 = n2658 & ~n4769 ;
  assign n4771 = n3192 & ~n4770 ;
  assign n4772 = n1962 & ~n4771 ;
  assign n4773 = n1966 & ~n4772 ;
  assign n4774 = n1970 & ~n4773 ;
  assign n4775 = n1974 & ~n4774 ;
  assign n4776 = n1978 & ~n4775 ;
  assign n4777 = n1982 & ~n4776 ;
  assign n4778 = n1986 & ~n4777 ;
  assign n4779 = ~x144 & ~n1988 ;
  assign n4780 = ~n4778 & n4779 ;
  assign n4783 = ~n4780 & ~x272 ;
  assign n4784 = ~n4782 & ~n4783 ;
  assign n4785 = ~n302 & n1660 ;
  assign n4786 = n1665 & ~n4785 ;
  assign n4787 = n1669 & ~n4786 ;
  assign n4788 = n1673 & ~n4787 ;
  assign n4789 = n1677 & ~n4788 ;
  assign n4790 = n1681 & ~n4789 ;
  assign n4791 = n1685 & ~n4790 ;
  assign n4792 = n1689 & ~n4791 ;
  assign n4793 = n1693 & ~n4792 ;
  assign n4794 = n1697 & ~n4793 ;
  assign n4795 = n1701 & ~n4794 ;
  assign n4796 = n1705 & ~n4795 ;
  assign n4797 = n1709 & ~n4796 ;
  assign n4798 = n1713 & ~n4797 ;
  assign n4799 = n1717 & ~n4798 ;
  assign n4800 = n1721 & ~n4799 ;
  assign n4801 = n1725 & ~n4800 ;
  assign n4802 = n1729 & ~n4801 ;
  assign n4803 = n1733 & ~n4802 ;
  assign n4804 = n1737 & ~n4803 ;
  assign n4805 = n1741 & ~n4804 ;
  assign n4806 = n1745 & ~n4805 ;
  assign n4807 = n1749 & ~n4806 ;
  assign n4808 = n1753 & ~n4807 ;
  assign n4809 = n1757 & ~n4808 ;
  assign n4810 = n1761 & ~n4809 ;
  assign n4811 = n1765 & ~n4810 ;
  assign n4812 = n1769 & ~n4811 ;
  assign n4813 = n1773 & ~n4812 ;
  assign n4814 = n1777 & ~n4813 ;
  assign n4815 = n1781 & ~n4814 ;
  assign n4816 = n1785 & ~n4815 ;
  assign n4817 = n1789 & ~n4816 ;
  assign n4818 = n1793 & ~n4817 ;
  assign n4819 = n1797 & ~n4818 ;
  assign n4820 = n1801 & ~n4819 ;
  assign n4821 = n1805 & ~n4820 ;
  assign n4822 = n1809 & ~n4821 ;
  assign n4823 = n1813 & ~n4822 ;
  assign n4824 = n1817 & ~n4823 ;
  assign n4825 = n1821 & ~n4824 ;
  assign n4826 = n1825 & ~n4825 ;
  assign n4827 = n1829 & ~n4826 ;
  assign n4828 = n1833 & ~n4827 ;
  assign n4829 = n1837 & ~n4828 ;
  assign n4830 = n1841 & ~n4829 ;
  assign n4831 = n1845 & ~n4830 ;
  assign n4832 = n1849 & ~n4831 ;
  assign n4833 = n1853 & ~n4832 ;
  assign n4834 = n1857 & ~n4833 ;
  assign n4835 = n1861 & ~n4834 ;
  assign n4836 = n1865 & ~n4835 ;
  assign n4837 = n1869 & ~n4836 ;
  assign n4838 = n1873 & ~n4837 ;
  assign n4839 = n1877 & ~n4838 ;
  assign n4840 = n1881 & ~n4839 ;
  assign n4841 = n1885 & ~n4840 ;
  assign n4842 = n1889 & ~n4841 ;
  assign n4843 = n1893 & ~n4842 ;
  assign n4844 = n1897 & ~n4843 ;
  assign n4845 = n1901 & ~n4844 ;
  assign n4846 = n1905 & ~n4845 ;
  assign n4847 = n1909 & ~n4846 ;
  assign n4848 = n1913 & ~n4847 ;
  assign n4849 = n1917 & ~n4848 ;
  assign n4850 = n1921 & ~n4849 ;
  assign n4851 = n1925 & ~n4850 ;
  assign n4852 = n1929 & ~n4851 ;
  assign n4853 = n1933 & ~n4852 ;
  assign n4854 = n1937 & ~n4853 ;
  assign n4855 = n1941 & ~n4854 ;
  assign n4856 = n1945 & ~n4855 ;
  assign n4857 = n1949 & ~n4856 ;
  assign n4858 = n1953 & ~n4857 ;
  assign n4859 = n2749 & ~n4858 ;
  assign n4860 = n263 & ~n4859 ;
  assign n4861 = n267 & ~n4860 ;
  assign n4862 = n271 & ~n4861 ;
  assign n4863 = n275 & ~n4862 ;
  assign n4864 = n279 & ~n4863 ;
  assign n4865 = n283 & ~n4864 ;
  assign n4866 = n287 & ~n4865 ;
  assign n4867 = n291 & ~n4866 ;
  assign n4868 = n295 & ~n4867 ;
  assign n4869 = x145 & ~n297 ;
  assign n4870 = ~n4868 & n4869 ;
  assign n4958 = n4870 & x273 ;
  assign n4871 = ~n641 & n1997 ;
  assign n4872 = n2002 & ~n4871 ;
  assign n4873 = n2006 & ~n4872 ;
  assign n4874 = n2010 & ~n4873 ;
  assign n4875 = n2014 & ~n4874 ;
  assign n4876 = n2018 & ~n4875 ;
  assign n4877 = n2022 & ~n4876 ;
  assign n4878 = n2026 & ~n4877 ;
  assign n4879 = n2030 & ~n4878 ;
  assign n4880 = n2034 & ~n4879 ;
  assign n4881 = n2038 & ~n4880 ;
  assign n4882 = n2042 & ~n4881 ;
  assign n4883 = n2046 & ~n4882 ;
  assign n4884 = n2050 & ~n4883 ;
  assign n4885 = n2054 & ~n4884 ;
  assign n4886 = n2058 & ~n4885 ;
  assign n4887 = n2062 & ~n4886 ;
  assign n4888 = n2066 & ~n4887 ;
  assign n4889 = n2070 & ~n4888 ;
  assign n4890 = n2074 & ~n4889 ;
  assign n4891 = n2078 & ~n4890 ;
  assign n4892 = n2082 & ~n4891 ;
  assign n4893 = n2086 & ~n4892 ;
  assign n4894 = n2090 & ~n4893 ;
  assign n4895 = n2094 & ~n4894 ;
  assign n4896 = n2098 & ~n4895 ;
  assign n4897 = n2102 & ~n4896 ;
  assign n4898 = n2106 & ~n4897 ;
  assign n4899 = n2110 & ~n4898 ;
  assign n4900 = n2114 & ~n4899 ;
  assign n4901 = n2118 & ~n4900 ;
  assign n4902 = n2122 & ~n4901 ;
  assign n4903 = n2126 & ~n4902 ;
  assign n4904 = n2130 & ~n4903 ;
  assign n4905 = n2134 & ~n4904 ;
  assign n4906 = n2138 & ~n4905 ;
  assign n4907 = n2142 & ~n4906 ;
  assign n4908 = n2146 & ~n4907 ;
  assign n4909 = n2150 & ~n4908 ;
  assign n4910 = n2154 & ~n4909 ;
  assign n4911 = n2158 & ~n4910 ;
  assign n4912 = n2162 & ~n4911 ;
  assign n4913 = n2166 & ~n4912 ;
  assign n4914 = n2170 & ~n4913 ;
  assign n4915 = n2174 & ~n4914 ;
  assign n4916 = n2178 & ~n4915 ;
  assign n4917 = n2182 & ~n4916 ;
  assign n4918 = n2186 & ~n4917 ;
  assign n4919 = n2190 & ~n4918 ;
  assign n4920 = n2194 & ~n4919 ;
  assign n4921 = n2198 & ~n4920 ;
  assign n4922 = n2202 & ~n4921 ;
  assign n4923 = n2206 & ~n4922 ;
  assign n4924 = n2210 & ~n4923 ;
  assign n4925 = n2214 & ~n4924 ;
  assign n4926 = n2218 & ~n4925 ;
  assign n4927 = n2222 & ~n4926 ;
  assign n4928 = n2226 & ~n4927 ;
  assign n4929 = n2230 & ~n4928 ;
  assign n4930 = n2234 & ~n4929 ;
  assign n4931 = n2238 & ~n4930 ;
  assign n4932 = n2242 & ~n4931 ;
  assign n4933 = n2246 & ~n4932 ;
  assign n4934 = n2250 & ~n4933 ;
  assign n4935 = n2254 & ~n4934 ;
  assign n4936 = n2258 & ~n4935 ;
  assign n4937 = n2262 & ~n4936 ;
  assign n4938 = n2266 & ~n4937 ;
  assign n4939 = n2270 & ~n4938 ;
  assign n4940 = n2274 & ~n4939 ;
  assign n4941 = n2278 & ~n4940 ;
  assign n4942 = n2282 & ~n4941 ;
  assign n4943 = n2286 & ~n4942 ;
  assign n4944 = n2290 & ~n4943 ;
  assign n4945 = n2836 & ~n4944 ;
  assign n4946 = n602 & ~n4945 ;
  assign n4947 = n606 & ~n4946 ;
  assign n4948 = n610 & ~n4947 ;
  assign n4949 = n614 & ~n4948 ;
  assign n4950 = n618 & ~n4949 ;
  assign n4951 = n622 & ~n4950 ;
  assign n4952 = n626 & ~n4951 ;
  assign n4953 = n630 & ~n4952 ;
  assign n4954 = n634 & ~n4953 ;
  assign n4955 = ~x145 & ~n636 ;
  assign n4956 = ~n4954 & n4955 ;
  assign n4959 = ~n4956 & ~x273 ;
  assign n4960 = ~n4958 & ~n4959 ;
  assign n4961 = n306 & ~n984 ;
  assign n4962 = n311 & ~n4961 ;
  assign n4963 = n315 & ~n4962 ;
  assign n4964 = n319 & ~n4963 ;
  assign n4965 = n323 & ~n4964 ;
  assign n4966 = n327 & ~n4965 ;
  assign n4967 = n331 & ~n4966 ;
  assign n4968 = n335 & ~n4967 ;
  assign n4969 = n339 & ~n4968 ;
  assign n4970 = n343 & ~n4969 ;
  assign n4971 = n347 & ~n4970 ;
  assign n4972 = n351 & ~n4971 ;
  assign n4973 = n355 & ~n4972 ;
  assign n4974 = n359 & ~n4973 ;
  assign n4975 = n363 & ~n4974 ;
  assign n4976 = n367 & ~n4975 ;
  assign n4977 = n371 & ~n4976 ;
  assign n4978 = n375 & ~n4977 ;
  assign n4979 = n379 & ~n4978 ;
  assign n4980 = n383 & ~n4979 ;
  assign n4981 = n387 & ~n4980 ;
  assign n4982 = n391 & ~n4981 ;
  assign n4983 = n395 & ~n4982 ;
  assign n4984 = n399 & ~n4983 ;
  assign n4985 = n403 & ~n4984 ;
  assign n4986 = n407 & ~n4985 ;
  assign n4987 = n411 & ~n4986 ;
  assign n4988 = n415 & ~n4987 ;
  assign n4989 = n419 & ~n4988 ;
  assign n4990 = n423 & ~n4989 ;
  assign n4991 = n427 & ~n4990 ;
  assign n4992 = n431 & ~n4991 ;
  assign n4993 = n435 & ~n4992 ;
  assign n4994 = n439 & ~n4993 ;
  assign n4995 = n443 & ~n4994 ;
  assign n4996 = n447 & ~n4995 ;
  assign n4997 = n451 & ~n4996 ;
  assign n4998 = n455 & ~n4997 ;
  assign n4999 = n459 & ~n4998 ;
  assign n5000 = n463 & ~n4999 ;
  assign n5001 = n467 & ~n5000 ;
  assign n5002 = n471 & ~n5001 ;
  assign n5003 = n475 & ~n5002 ;
  assign n5004 = n479 & ~n5003 ;
  assign n5005 = n483 & ~n5004 ;
  assign n5006 = n487 & ~n5005 ;
  assign n5007 = n491 & ~n5006 ;
  assign n5008 = n495 & ~n5007 ;
  assign n5009 = n499 & ~n5008 ;
  assign n5010 = n503 & ~n5009 ;
  assign n5011 = n507 & ~n5010 ;
  assign n5012 = n511 & ~n5011 ;
  assign n5013 = n515 & ~n5012 ;
  assign n5014 = n519 & ~n5013 ;
  assign n5015 = n523 & ~n5014 ;
  assign n5016 = n527 & ~n5015 ;
  assign n5017 = n531 & ~n5016 ;
  assign n5018 = n535 & ~n5017 ;
  assign n5019 = n539 & ~n5018 ;
  assign n5020 = n543 & ~n5019 ;
  assign n5021 = n547 & ~n5020 ;
  assign n5022 = n551 & ~n5021 ;
  assign n5023 = n555 & ~n5022 ;
  assign n5024 = n559 & ~n5023 ;
  assign n5025 = n563 & ~n5024 ;
  assign n5026 = n567 & ~n5025 ;
  assign n5027 = n571 & ~n5026 ;
  assign n5028 = n575 & ~n5027 ;
  assign n5029 = n579 & ~n5028 ;
  assign n5030 = n583 & ~n5029 ;
  assign n5031 = n587 & ~n5030 ;
  assign n5032 = n591 & ~n5031 ;
  assign n5033 = n2382 & ~n5032 ;
  assign n5034 = n2384 & ~n5033 ;
  assign n5035 = n2927 & ~n5034 ;
  assign n5036 = n945 & ~n5035 ;
  assign n5037 = n949 & ~n5036 ;
  assign n5038 = n953 & ~n5037 ;
  assign n5039 = n957 & ~n5038 ;
  assign n5040 = n961 & ~n5039 ;
  assign n5041 = n965 & ~n5040 ;
  assign n5042 = n969 & ~n5041 ;
  assign n5043 = n973 & ~n5042 ;
  assign n5044 = n977 & ~n5043 ;
  assign n5045 = x146 & ~n979 ;
  assign n5046 = ~n5044 & n5045 ;
  assign n5134 = n5046 & x274 ;
  assign n5047 = n645 & ~n1323 ;
  assign n5048 = n650 & ~n5047 ;
  assign n5049 = n654 & ~n5048 ;
  assign n5050 = n658 & ~n5049 ;
  assign n5051 = n662 & ~n5050 ;
  assign n5052 = n666 & ~n5051 ;
  assign n5053 = n670 & ~n5052 ;
  assign n5054 = n674 & ~n5053 ;
  assign n5055 = n678 & ~n5054 ;
  assign n5056 = n682 & ~n5055 ;
  assign n5057 = n686 & ~n5056 ;
  assign n5058 = n690 & ~n5057 ;
  assign n5059 = n694 & ~n5058 ;
  assign n5060 = n698 & ~n5059 ;
  assign n5061 = n702 & ~n5060 ;
  assign n5062 = n706 & ~n5061 ;
  assign n5063 = n710 & ~n5062 ;
  assign n5064 = n714 & ~n5063 ;
  assign n5065 = n718 & ~n5064 ;
  assign n5066 = n722 & ~n5065 ;
  assign n5067 = n726 & ~n5066 ;
  assign n5068 = n730 & ~n5067 ;
  assign n5069 = n734 & ~n5068 ;
  assign n5070 = n738 & ~n5069 ;
  assign n5071 = n742 & ~n5070 ;
  assign n5072 = n746 & ~n5071 ;
  assign n5073 = n750 & ~n5072 ;
  assign n5074 = n754 & ~n5073 ;
  assign n5075 = n758 & ~n5074 ;
  assign n5076 = n762 & ~n5075 ;
  assign n5077 = n766 & ~n5076 ;
  assign n5078 = n770 & ~n5077 ;
  assign n5079 = n774 & ~n5078 ;
  assign n5080 = n778 & ~n5079 ;
  assign n5081 = n782 & ~n5080 ;
  assign n5082 = n786 & ~n5081 ;
  assign n5083 = n790 & ~n5082 ;
  assign n5084 = n794 & ~n5083 ;
  assign n5085 = n798 & ~n5084 ;
  assign n5086 = n802 & ~n5085 ;
  assign n5087 = n806 & ~n5086 ;
  assign n5088 = n810 & ~n5087 ;
  assign n5089 = n814 & ~n5088 ;
  assign n5090 = n818 & ~n5089 ;
  assign n5091 = n822 & ~n5090 ;
  assign n5092 = n826 & ~n5091 ;
  assign n5093 = n830 & ~n5092 ;
  assign n5094 = n834 & ~n5093 ;
  assign n5095 = n838 & ~n5094 ;
  assign n5096 = n842 & ~n5095 ;
  assign n5097 = n846 & ~n5096 ;
  assign n5098 = n850 & ~n5097 ;
  assign n5099 = n854 & ~n5098 ;
  assign n5100 = n858 & ~n5099 ;
  assign n5101 = n862 & ~n5100 ;
  assign n5102 = n866 & ~n5101 ;
  assign n5103 = n870 & ~n5102 ;
  assign n5104 = n874 & ~n5103 ;
  assign n5105 = n878 & ~n5104 ;
  assign n5106 = n882 & ~n5105 ;
  assign n5107 = n886 & ~n5106 ;
  assign n5108 = n890 & ~n5107 ;
  assign n5109 = n894 & ~n5108 ;
  assign n5110 = n898 & ~n5109 ;
  assign n5111 = n902 & ~n5110 ;
  assign n5112 = n906 & ~n5111 ;
  assign n5113 = n910 & ~n5112 ;
  assign n5114 = n914 & ~n5113 ;
  assign n5115 = n918 & ~n5114 ;
  assign n5116 = n922 & ~n5115 ;
  assign n5117 = n926 & ~n5116 ;
  assign n5118 = n930 & ~n5117 ;
  assign n5119 = n2472 & ~n5118 ;
  assign n5120 = n2474 & ~n5119 ;
  assign n5121 = n3014 & ~n5120 ;
  assign n5122 = n1284 & ~n5121 ;
  assign n5123 = n1288 & ~n5122 ;
  assign n5124 = n1292 & ~n5123 ;
  assign n5125 = n1296 & ~n5124 ;
  assign n5126 = n1300 & ~n5125 ;
  assign n5127 = n1304 & ~n5126 ;
  assign n5128 = n1308 & ~n5127 ;
  assign n5129 = n1312 & ~n5128 ;
  assign n5130 = n1316 & ~n5129 ;
  assign n5131 = ~x146 & ~n1318 ;
  assign n5132 = ~n5130 & n5131 ;
  assign n5135 = ~n5132 & ~x274 ;
  assign n5136 = ~n5134 & ~n5135 ;
  assign n5137 = n988 & ~n1664 ;
  assign n5138 = n993 & ~n5137 ;
  assign n5139 = n997 & ~n5138 ;
  assign n5140 = n1001 & ~n5139 ;
  assign n5141 = n1005 & ~n5140 ;
  assign n5142 = n1009 & ~n5141 ;
  assign n5143 = n1013 & ~n5142 ;
  assign n5144 = n1017 & ~n5143 ;
  assign n5145 = n1021 & ~n5144 ;
  assign n5146 = n1025 & ~n5145 ;
  assign n5147 = n1029 & ~n5146 ;
  assign n5148 = n1033 & ~n5147 ;
  assign n5149 = n1037 & ~n5148 ;
  assign n5150 = n1041 & ~n5149 ;
  assign n5151 = n1045 & ~n5150 ;
  assign n5152 = n1049 & ~n5151 ;
  assign n5153 = n1053 & ~n5152 ;
  assign n5154 = n1057 & ~n5153 ;
  assign n5155 = n1061 & ~n5154 ;
  assign n5156 = n1065 & ~n5155 ;
  assign n5157 = n1069 & ~n5156 ;
  assign n5158 = n1073 & ~n5157 ;
  assign n5159 = n1077 & ~n5158 ;
  assign n5160 = n1081 & ~n5159 ;
  assign n5161 = n1085 & ~n5160 ;
  assign n5162 = n1089 & ~n5161 ;
  assign n5163 = n1093 & ~n5162 ;
  assign n5164 = n1097 & ~n5163 ;
  assign n5165 = n1101 & ~n5164 ;
  assign n5166 = n1105 & ~n5165 ;
  assign n5167 = n1109 & ~n5166 ;
  assign n5168 = n1113 & ~n5167 ;
  assign n5169 = n1117 & ~n5168 ;
  assign n5170 = n1121 & ~n5169 ;
  assign n5171 = n1125 & ~n5170 ;
  assign n5172 = n1129 & ~n5171 ;
  assign n5173 = n1133 & ~n5172 ;
  assign n5174 = n1137 & ~n5173 ;
  assign n5175 = n1141 & ~n5174 ;
  assign n5176 = n1145 & ~n5175 ;
  assign n5177 = n1149 & ~n5176 ;
  assign n5178 = n1153 & ~n5177 ;
  assign n5179 = n1157 & ~n5178 ;
  assign n5180 = n1161 & ~n5179 ;
  assign n5181 = n1165 & ~n5180 ;
  assign n5182 = n1169 & ~n5181 ;
  assign n5183 = n1173 & ~n5182 ;
  assign n5184 = n1177 & ~n5183 ;
  assign n5185 = n1181 & ~n5184 ;
  assign n5186 = n1185 & ~n5185 ;
  assign n5187 = n1189 & ~n5186 ;
  assign n5188 = n1193 & ~n5187 ;
  assign n5189 = n1197 & ~n5188 ;
  assign n5190 = n1201 & ~n5189 ;
  assign n5191 = n1205 & ~n5190 ;
  assign n5192 = n1209 & ~n5191 ;
  assign n5193 = n1213 & ~n5192 ;
  assign n5194 = n1217 & ~n5193 ;
  assign n5195 = n1221 & ~n5194 ;
  assign n5196 = n1225 & ~n5195 ;
  assign n5197 = n1229 & ~n5196 ;
  assign n5198 = n1233 & ~n5197 ;
  assign n5199 = n1237 & ~n5198 ;
  assign n5200 = n1241 & ~n5199 ;
  assign n5201 = n1245 & ~n5200 ;
  assign n5202 = n1249 & ~n5201 ;
  assign n5203 = n1253 & ~n5202 ;
  assign n5204 = n1257 & ~n5203 ;
  assign n5205 = n1261 & ~n5204 ;
  assign n5206 = n1265 & ~n5205 ;
  assign n5207 = n1269 & ~n5206 ;
  assign n5208 = n1273 & ~n5207 ;
  assign n5209 = n2566 & ~n5208 ;
  assign n5210 = n2568 & ~n5209 ;
  assign n5211 = n3105 & ~n5210 ;
  assign n5212 = n1625 & ~n5211 ;
  assign n5213 = n1629 & ~n5212 ;
  assign n5214 = n1633 & ~n5213 ;
  assign n5215 = n1637 & ~n5214 ;
  assign n5216 = n1641 & ~n5215 ;
  assign n5217 = n1645 & ~n5216 ;
  assign n5218 = n1649 & ~n5217 ;
  assign n5219 = n1653 & ~n5218 ;
  assign n5220 = n1657 & ~n5219 ;
  assign n5221 = x147 & ~n1659 ;
  assign n5222 = ~n5220 & n5221 ;
  assign n5310 = n5222 & x275 ;
  assign n5223 = n1327 & ~n2001 ;
  assign n5224 = n1332 & ~n5223 ;
  assign n5225 = n1336 & ~n5224 ;
  assign n5226 = n1340 & ~n5225 ;
  assign n5227 = n1344 & ~n5226 ;
  assign n5228 = n1348 & ~n5227 ;
  assign n5229 = n1352 & ~n5228 ;
  assign n5230 = n1356 & ~n5229 ;
  assign n5231 = n1360 & ~n5230 ;
  assign n5232 = n1364 & ~n5231 ;
  assign n5233 = n1368 & ~n5232 ;
  assign n5234 = n1372 & ~n5233 ;
  assign n5235 = n1376 & ~n5234 ;
  assign n5236 = n1380 & ~n5235 ;
  assign n5237 = n1384 & ~n5236 ;
  assign n5238 = n1388 & ~n5237 ;
  assign n5239 = n1392 & ~n5238 ;
  assign n5240 = n1396 & ~n5239 ;
  assign n5241 = n1400 & ~n5240 ;
  assign n5242 = n1404 & ~n5241 ;
  assign n5243 = n1408 & ~n5242 ;
  assign n5244 = n1412 & ~n5243 ;
  assign n5245 = n1416 & ~n5244 ;
  assign n5246 = n1420 & ~n5245 ;
  assign n5247 = n1424 & ~n5246 ;
  assign n5248 = n1428 & ~n5247 ;
  assign n5249 = n1432 & ~n5248 ;
  assign n5250 = n1436 & ~n5249 ;
  assign n5251 = n1440 & ~n5250 ;
  assign n5252 = n1444 & ~n5251 ;
  assign n5253 = n1448 & ~n5252 ;
  assign n5254 = n1452 & ~n5253 ;
  assign n5255 = n1456 & ~n5254 ;
  assign n5256 = n1460 & ~n5255 ;
  assign n5257 = n1464 & ~n5256 ;
  assign n5258 = n1468 & ~n5257 ;
  assign n5259 = n1472 & ~n5258 ;
  assign n5260 = n1476 & ~n5259 ;
  assign n5261 = n1480 & ~n5260 ;
  assign n5262 = n1484 & ~n5261 ;
  assign n5263 = n1488 & ~n5262 ;
  assign n5264 = n1492 & ~n5263 ;
  assign n5265 = n1496 & ~n5264 ;
  assign n5266 = n1500 & ~n5265 ;
  assign n5267 = n1504 & ~n5266 ;
  assign n5268 = n1508 & ~n5267 ;
  assign n5269 = n1512 & ~n5268 ;
  assign n5270 = n1516 & ~n5269 ;
  assign n5271 = n1520 & ~n5270 ;
  assign n5272 = n1524 & ~n5271 ;
  assign n5273 = n1528 & ~n5272 ;
  assign n5274 = n1532 & ~n5273 ;
  assign n5275 = n1536 & ~n5274 ;
  assign n5276 = n1540 & ~n5275 ;
  assign n5277 = n1544 & ~n5276 ;
  assign n5278 = n1548 & ~n5277 ;
  assign n5279 = n1552 & ~n5278 ;
  assign n5280 = n1556 & ~n5279 ;
  assign n5281 = n1560 & ~n5280 ;
  assign n5282 = n1564 & ~n5281 ;
  assign n5283 = n1568 & ~n5282 ;
  assign n5284 = n1572 & ~n5283 ;
  assign n5285 = n1576 & ~n5284 ;
  assign n5286 = n1580 & ~n5285 ;
  assign n5287 = n1584 & ~n5286 ;
  assign n5288 = n1588 & ~n5287 ;
  assign n5289 = n1592 & ~n5288 ;
  assign n5290 = n1596 & ~n5289 ;
  assign n5291 = n1600 & ~n5290 ;
  assign n5292 = n1604 & ~n5291 ;
  assign n5293 = n1608 & ~n5292 ;
  assign n5294 = n1612 & ~n5293 ;
  assign n5295 = n2656 & ~n5294 ;
  assign n5296 = n2658 & ~n5295 ;
  assign n5297 = n3192 & ~n5296 ;
  assign n5298 = n1962 & ~n5297 ;
  assign n5299 = n1966 & ~n5298 ;
  assign n5300 = n1970 & ~n5299 ;
  assign n5301 = n1974 & ~n5300 ;
  assign n5302 = n1978 & ~n5301 ;
  assign n5303 = n1982 & ~n5302 ;
  assign n5304 = n1986 & ~n5303 ;
  assign n5305 = n1990 & ~n5304 ;
  assign n5306 = n1994 & ~n5305 ;
  assign n5307 = ~x147 & ~n1996 ;
  assign n5308 = ~n5306 & n5307 ;
  assign n5311 = ~n5308 & ~x275 ;
  assign n5312 = ~n5310 & ~n5311 ;
  assign n5313 = ~n310 & n1668 ;
  assign n5314 = n1673 & ~n5313 ;
  assign n5315 = n1677 & ~n5314 ;
  assign n5316 = n1681 & ~n5315 ;
  assign n5317 = n1685 & ~n5316 ;
  assign n5318 = n1689 & ~n5317 ;
  assign n5319 = n1693 & ~n5318 ;
  assign n5320 = n1697 & ~n5319 ;
  assign n5321 = n1701 & ~n5320 ;
  assign n5322 = n1705 & ~n5321 ;
  assign n5323 = n1709 & ~n5322 ;
  assign n5324 = n1713 & ~n5323 ;
  assign n5325 = n1717 & ~n5324 ;
  assign n5326 = n1721 & ~n5325 ;
  assign n5327 = n1725 & ~n5326 ;
  assign n5328 = n1729 & ~n5327 ;
  assign n5329 = n1733 & ~n5328 ;
  assign n5330 = n1737 & ~n5329 ;
  assign n5331 = n1741 & ~n5330 ;
  assign n5332 = n1745 & ~n5331 ;
  assign n5333 = n1749 & ~n5332 ;
  assign n5334 = n1753 & ~n5333 ;
  assign n5335 = n1757 & ~n5334 ;
  assign n5336 = n1761 & ~n5335 ;
  assign n5337 = n1765 & ~n5336 ;
  assign n5338 = n1769 & ~n5337 ;
  assign n5339 = n1773 & ~n5338 ;
  assign n5340 = n1777 & ~n5339 ;
  assign n5341 = n1781 & ~n5340 ;
  assign n5342 = n1785 & ~n5341 ;
  assign n5343 = n1789 & ~n5342 ;
  assign n5344 = n1793 & ~n5343 ;
  assign n5345 = n1797 & ~n5344 ;
  assign n5346 = n1801 & ~n5345 ;
  assign n5347 = n1805 & ~n5346 ;
  assign n5348 = n1809 & ~n5347 ;
  assign n5349 = n1813 & ~n5348 ;
  assign n5350 = n1817 & ~n5349 ;
  assign n5351 = n1821 & ~n5350 ;
  assign n5352 = n1825 & ~n5351 ;
  assign n5353 = n1829 & ~n5352 ;
  assign n5354 = n1833 & ~n5353 ;
  assign n5355 = n1837 & ~n5354 ;
  assign n5356 = n1841 & ~n5355 ;
  assign n5357 = n1845 & ~n5356 ;
  assign n5358 = n1849 & ~n5357 ;
  assign n5359 = n1853 & ~n5358 ;
  assign n5360 = n1857 & ~n5359 ;
  assign n5361 = n1861 & ~n5360 ;
  assign n5362 = n1865 & ~n5361 ;
  assign n5363 = n1869 & ~n5362 ;
  assign n5364 = n1873 & ~n5363 ;
  assign n5365 = n1877 & ~n5364 ;
  assign n5366 = n1881 & ~n5365 ;
  assign n5367 = n1885 & ~n5366 ;
  assign n5368 = n1889 & ~n5367 ;
  assign n5369 = n1893 & ~n5368 ;
  assign n5370 = n1897 & ~n5369 ;
  assign n5371 = n1901 & ~n5370 ;
  assign n5372 = n1905 & ~n5371 ;
  assign n5373 = n1909 & ~n5372 ;
  assign n5374 = n1913 & ~n5373 ;
  assign n5375 = n1917 & ~n5374 ;
  assign n5376 = n1921 & ~n5375 ;
  assign n5377 = n1925 & ~n5376 ;
  assign n5378 = n1929 & ~n5377 ;
  assign n5379 = n1933 & ~n5378 ;
  assign n5380 = n1937 & ~n5379 ;
  assign n5381 = n1941 & ~n5380 ;
  assign n5382 = n1945 & ~n5381 ;
  assign n5383 = n1949 & ~n5382 ;
  assign n5384 = n1953 & ~n5383 ;
  assign n5385 = n2749 & ~n5384 ;
  assign n5386 = n263 & ~n5385 ;
  assign n5387 = n267 & ~n5386 ;
  assign n5388 = n271 & ~n5387 ;
  assign n5389 = n275 & ~n5388 ;
  assign n5390 = n279 & ~n5389 ;
  assign n5391 = n283 & ~n5390 ;
  assign n5392 = n287 & ~n5391 ;
  assign n5393 = n291 & ~n5392 ;
  assign n5394 = n295 & ~n5393 ;
  assign n5395 = n299 & ~n5394 ;
  assign n5396 = n303 & ~n5395 ;
  assign n5397 = x148 & ~n305 ;
  assign n5398 = ~n5396 & n5397 ;
  assign n5486 = n5398 & x276 ;
  assign n5399 = ~n649 & n2005 ;
  assign n5400 = n2010 & ~n5399 ;
  assign n5401 = n2014 & ~n5400 ;
  assign n5402 = n2018 & ~n5401 ;
  assign n5403 = n2022 & ~n5402 ;
  assign n5404 = n2026 & ~n5403 ;
  assign n5405 = n2030 & ~n5404 ;
  assign n5406 = n2034 & ~n5405 ;
  assign n5407 = n2038 & ~n5406 ;
  assign n5408 = n2042 & ~n5407 ;
  assign n5409 = n2046 & ~n5408 ;
  assign n5410 = n2050 & ~n5409 ;
  assign n5411 = n2054 & ~n5410 ;
  assign n5412 = n2058 & ~n5411 ;
  assign n5413 = n2062 & ~n5412 ;
  assign n5414 = n2066 & ~n5413 ;
  assign n5415 = n2070 & ~n5414 ;
  assign n5416 = n2074 & ~n5415 ;
  assign n5417 = n2078 & ~n5416 ;
  assign n5418 = n2082 & ~n5417 ;
  assign n5419 = n2086 & ~n5418 ;
  assign n5420 = n2090 & ~n5419 ;
  assign n5421 = n2094 & ~n5420 ;
  assign n5422 = n2098 & ~n5421 ;
  assign n5423 = n2102 & ~n5422 ;
  assign n5424 = n2106 & ~n5423 ;
  assign n5425 = n2110 & ~n5424 ;
  assign n5426 = n2114 & ~n5425 ;
  assign n5427 = n2118 & ~n5426 ;
  assign n5428 = n2122 & ~n5427 ;
  assign n5429 = n2126 & ~n5428 ;
  assign n5430 = n2130 & ~n5429 ;
  assign n5431 = n2134 & ~n5430 ;
  assign n5432 = n2138 & ~n5431 ;
  assign n5433 = n2142 & ~n5432 ;
  assign n5434 = n2146 & ~n5433 ;
  assign n5435 = n2150 & ~n5434 ;
  assign n5436 = n2154 & ~n5435 ;
  assign n5437 = n2158 & ~n5436 ;
  assign n5438 = n2162 & ~n5437 ;
  assign n5439 = n2166 & ~n5438 ;
  assign n5440 = n2170 & ~n5439 ;
  assign n5441 = n2174 & ~n5440 ;
  assign n5442 = n2178 & ~n5441 ;
  assign n5443 = n2182 & ~n5442 ;
  assign n5444 = n2186 & ~n5443 ;
  assign n5445 = n2190 & ~n5444 ;
  assign n5446 = n2194 & ~n5445 ;
  assign n5447 = n2198 & ~n5446 ;
  assign n5448 = n2202 & ~n5447 ;
  assign n5449 = n2206 & ~n5448 ;
  assign n5450 = n2210 & ~n5449 ;
  assign n5451 = n2214 & ~n5450 ;
  assign n5452 = n2218 & ~n5451 ;
  assign n5453 = n2222 & ~n5452 ;
  assign n5454 = n2226 & ~n5453 ;
  assign n5455 = n2230 & ~n5454 ;
  assign n5456 = n2234 & ~n5455 ;
  assign n5457 = n2238 & ~n5456 ;
  assign n5458 = n2242 & ~n5457 ;
  assign n5459 = n2246 & ~n5458 ;
  assign n5460 = n2250 & ~n5459 ;
  assign n5461 = n2254 & ~n5460 ;
  assign n5462 = n2258 & ~n5461 ;
  assign n5463 = n2262 & ~n5462 ;
  assign n5464 = n2266 & ~n5463 ;
  assign n5465 = n2270 & ~n5464 ;
  assign n5466 = n2274 & ~n5465 ;
  assign n5467 = n2278 & ~n5466 ;
  assign n5468 = n2282 & ~n5467 ;
  assign n5469 = n2286 & ~n5468 ;
  assign n5470 = n2290 & ~n5469 ;
  assign n5471 = n2836 & ~n5470 ;
  assign n5472 = n602 & ~n5471 ;
  assign n5473 = n606 & ~n5472 ;
  assign n5474 = n610 & ~n5473 ;
  assign n5475 = n614 & ~n5474 ;
  assign n5476 = n618 & ~n5475 ;
  assign n5477 = n622 & ~n5476 ;
  assign n5478 = n626 & ~n5477 ;
  assign n5479 = n630 & ~n5478 ;
  assign n5480 = n634 & ~n5479 ;
  assign n5481 = n638 & ~n5480 ;
  assign n5482 = n642 & ~n5481 ;
  assign n5483 = ~x148 & ~n644 ;
  assign n5484 = ~n5482 & n5483 ;
  assign n5487 = ~n5484 & ~x276 ;
  assign n5488 = ~n5486 & ~n5487 ;
  assign n5489 = n314 & ~n992 ;
  assign n5490 = n319 & ~n5489 ;
  assign n5491 = n323 & ~n5490 ;
  assign n5492 = n327 & ~n5491 ;
  assign n5493 = n331 & ~n5492 ;
  assign n5494 = n335 & ~n5493 ;
  assign n5495 = n339 & ~n5494 ;
  assign n5496 = n343 & ~n5495 ;
  assign n5497 = n347 & ~n5496 ;
  assign n5498 = n351 & ~n5497 ;
  assign n5499 = n355 & ~n5498 ;
  assign n5500 = n359 & ~n5499 ;
  assign n5501 = n363 & ~n5500 ;
  assign n5502 = n367 & ~n5501 ;
  assign n5503 = n371 & ~n5502 ;
  assign n5504 = n375 & ~n5503 ;
  assign n5505 = n379 & ~n5504 ;
  assign n5506 = n383 & ~n5505 ;
  assign n5507 = n387 & ~n5506 ;
  assign n5508 = n391 & ~n5507 ;
  assign n5509 = n395 & ~n5508 ;
  assign n5510 = n399 & ~n5509 ;
  assign n5511 = n403 & ~n5510 ;
  assign n5512 = n407 & ~n5511 ;
  assign n5513 = n411 & ~n5512 ;
  assign n5514 = n415 & ~n5513 ;
  assign n5515 = n419 & ~n5514 ;
  assign n5516 = n423 & ~n5515 ;
  assign n5517 = n427 & ~n5516 ;
  assign n5518 = n431 & ~n5517 ;
  assign n5519 = n435 & ~n5518 ;
  assign n5520 = n439 & ~n5519 ;
  assign n5521 = n443 & ~n5520 ;
  assign n5522 = n447 & ~n5521 ;
  assign n5523 = n451 & ~n5522 ;
  assign n5524 = n455 & ~n5523 ;
  assign n5525 = n459 & ~n5524 ;
  assign n5526 = n463 & ~n5525 ;
  assign n5527 = n467 & ~n5526 ;
  assign n5528 = n471 & ~n5527 ;
  assign n5529 = n475 & ~n5528 ;
  assign n5530 = n479 & ~n5529 ;
  assign n5531 = n483 & ~n5530 ;
  assign n5532 = n487 & ~n5531 ;
  assign n5533 = n491 & ~n5532 ;
  assign n5534 = n495 & ~n5533 ;
  assign n5535 = n499 & ~n5534 ;
  assign n5536 = n503 & ~n5535 ;
  assign n5537 = n507 & ~n5536 ;
  assign n5538 = n511 & ~n5537 ;
  assign n5539 = n515 & ~n5538 ;
  assign n5540 = n519 & ~n5539 ;
  assign n5541 = n523 & ~n5540 ;
  assign n5542 = n527 & ~n5541 ;
  assign n5543 = n531 & ~n5542 ;
  assign n5544 = n535 & ~n5543 ;
  assign n5545 = n539 & ~n5544 ;
  assign n5546 = n543 & ~n5545 ;
  assign n5547 = n547 & ~n5546 ;
  assign n5548 = n551 & ~n5547 ;
  assign n5549 = n555 & ~n5548 ;
  assign n5550 = n559 & ~n5549 ;
  assign n5551 = n563 & ~n5550 ;
  assign n5552 = n567 & ~n5551 ;
  assign n5553 = n571 & ~n5552 ;
  assign n5554 = n575 & ~n5553 ;
  assign n5555 = n579 & ~n5554 ;
  assign n5556 = n583 & ~n5555 ;
  assign n5557 = n587 & ~n5556 ;
  assign n5558 = n591 & ~n5557 ;
  assign n5559 = n2382 & ~n5558 ;
  assign n5560 = n2384 & ~n5559 ;
  assign n5561 = n2927 & ~n5560 ;
  assign n5562 = n945 & ~n5561 ;
  assign n5563 = n949 & ~n5562 ;
  assign n5564 = n953 & ~n5563 ;
  assign n5565 = n957 & ~n5564 ;
  assign n5566 = n961 & ~n5565 ;
  assign n5567 = n965 & ~n5566 ;
  assign n5568 = n969 & ~n5567 ;
  assign n5569 = n973 & ~n5568 ;
  assign n5570 = n977 & ~n5569 ;
  assign n5571 = n981 & ~n5570 ;
  assign n5572 = n985 & ~n5571 ;
  assign n5573 = x149 & ~n987 ;
  assign n5574 = ~n5572 & n5573 ;
  assign n5662 = n5574 & x277 ;
  assign n5575 = n653 & ~n1331 ;
  assign n5576 = n658 & ~n5575 ;
  assign n5577 = n662 & ~n5576 ;
  assign n5578 = n666 & ~n5577 ;
  assign n5579 = n670 & ~n5578 ;
  assign n5580 = n674 & ~n5579 ;
  assign n5581 = n678 & ~n5580 ;
  assign n5582 = n682 & ~n5581 ;
  assign n5583 = n686 & ~n5582 ;
  assign n5584 = n690 & ~n5583 ;
  assign n5585 = n694 & ~n5584 ;
  assign n5586 = n698 & ~n5585 ;
  assign n5587 = n702 & ~n5586 ;
  assign n5588 = n706 & ~n5587 ;
  assign n5589 = n710 & ~n5588 ;
  assign n5590 = n714 & ~n5589 ;
  assign n5591 = n718 & ~n5590 ;
  assign n5592 = n722 & ~n5591 ;
  assign n5593 = n726 & ~n5592 ;
  assign n5594 = n730 & ~n5593 ;
  assign n5595 = n734 & ~n5594 ;
  assign n5596 = n738 & ~n5595 ;
  assign n5597 = n742 & ~n5596 ;
  assign n5598 = n746 & ~n5597 ;
  assign n5599 = n750 & ~n5598 ;
  assign n5600 = n754 & ~n5599 ;
  assign n5601 = n758 & ~n5600 ;
  assign n5602 = n762 & ~n5601 ;
  assign n5603 = n766 & ~n5602 ;
  assign n5604 = n770 & ~n5603 ;
  assign n5605 = n774 & ~n5604 ;
  assign n5606 = n778 & ~n5605 ;
  assign n5607 = n782 & ~n5606 ;
  assign n5608 = n786 & ~n5607 ;
  assign n5609 = n790 & ~n5608 ;
  assign n5610 = n794 & ~n5609 ;
  assign n5611 = n798 & ~n5610 ;
  assign n5612 = n802 & ~n5611 ;
  assign n5613 = n806 & ~n5612 ;
  assign n5614 = n810 & ~n5613 ;
  assign n5615 = n814 & ~n5614 ;
  assign n5616 = n818 & ~n5615 ;
  assign n5617 = n822 & ~n5616 ;
  assign n5618 = n826 & ~n5617 ;
  assign n5619 = n830 & ~n5618 ;
  assign n5620 = n834 & ~n5619 ;
  assign n5621 = n838 & ~n5620 ;
  assign n5622 = n842 & ~n5621 ;
  assign n5623 = n846 & ~n5622 ;
  assign n5624 = n850 & ~n5623 ;
  assign n5625 = n854 & ~n5624 ;
  assign n5626 = n858 & ~n5625 ;
  assign n5627 = n862 & ~n5626 ;
  assign n5628 = n866 & ~n5627 ;
  assign n5629 = n870 & ~n5628 ;
  assign n5630 = n874 & ~n5629 ;
  assign n5631 = n878 & ~n5630 ;
  assign n5632 = n882 & ~n5631 ;
  assign n5633 = n886 & ~n5632 ;
  assign n5634 = n890 & ~n5633 ;
  assign n5635 = n894 & ~n5634 ;
  assign n5636 = n898 & ~n5635 ;
  assign n5637 = n902 & ~n5636 ;
  assign n5638 = n906 & ~n5637 ;
  assign n5639 = n910 & ~n5638 ;
  assign n5640 = n914 & ~n5639 ;
  assign n5641 = n918 & ~n5640 ;
  assign n5642 = n922 & ~n5641 ;
  assign n5643 = n926 & ~n5642 ;
  assign n5644 = n930 & ~n5643 ;
  assign n5645 = n2472 & ~n5644 ;
  assign n5646 = n2474 & ~n5645 ;
  assign n5647 = n3014 & ~n5646 ;
  assign n5648 = n1284 & ~n5647 ;
  assign n5649 = n1288 & ~n5648 ;
  assign n5650 = n1292 & ~n5649 ;
  assign n5651 = n1296 & ~n5650 ;
  assign n5652 = n1300 & ~n5651 ;
  assign n5653 = n1304 & ~n5652 ;
  assign n5654 = n1308 & ~n5653 ;
  assign n5655 = n1312 & ~n5654 ;
  assign n5656 = n1316 & ~n5655 ;
  assign n5657 = n1320 & ~n5656 ;
  assign n5658 = n1324 & ~n5657 ;
  assign n5659 = ~x149 & ~n1326 ;
  assign n5660 = ~n5658 & n5659 ;
  assign n5663 = ~n5660 & ~x277 ;
  assign n5664 = ~n5662 & ~n5663 ;
  assign n5665 = n996 & ~n1672 ;
  assign n5666 = n1001 & ~n5665 ;
  assign n5667 = n1005 & ~n5666 ;
  assign n5668 = n1009 & ~n5667 ;
  assign n5669 = n1013 & ~n5668 ;
  assign n5670 = n1017 & ~n5669 ;
  assign n5671 = n1021 & ~n5670 ;
  assign n5672 = n1025 & ~n5671 ;
  assign n5673 = n1029 & ~n5672 ;
  assign n5674 = n1033 & ~n5673 ;
  assign n5675 = n1037 & ~n5674 ;
  assign n5676 = n1041 & ~n5675 ;
  assign n5677 = n1045 & ~n5676 ;
  assign n5678 = n1049 & ~n5677 ;
  assign n5679 = n1053 & ~n5678 ;
  assign n5680 = n1057 & ~n5679 ;
  assign n5681 = n1061 & ~n5680 ;
  assign n5682 = n1065 & ~n5681 ;
  assign n5683 = n1069 & ~n5682 ;
  assign n5684 = n1073 & ~n5683 ;
  assign n5685 = n1077 & ~n5684 ;
  assign n5686 = n1081 & ~n5685 ;
  assign n5687 = n1085 & ~n5686 ;
  assign n5688 = n1089 & ~n5687 ;
  assign n5689 = n1093 & ~n5688 ;
  assign n5690 = n1097 & ~n5689 ;
  assign n5691 = n1101 & ~n5690 ;
  assign n5692 = n1105 & ~n5691 ;
  assign n5693 = n1109 & ~n5692 ;
  assign n5694 = n1113 & ~n5693 ;
  assign n5695 = n1117 & ~n5694 ;
  assign n5696 = n1121 & ~n5695 ;
  assign n5697 = n1125 & ~n5696 ;
  assign n5698 = n1129 & ~n5697 ;
  assign n5699 = n1133 & ~n5698 ;
  assign n5700 = n1137 & ~n5699 ;
  assign n5701 = n1141 & ~n5700 ;
  assign n5702 = n1145 & ~n5701 ;
  assign n5703 = n1149 & ~n5702 ;
  assign n5704 = n1153 & ~n5703 ;
  assign n5705 = n1157 & ~n5704 ;
  assign n5706 = n1161 & ~n5705 ;
  assign n5707 = n1165 & ~n5706 ;
  assign n5708 = n1169 & ~n5707 ;
  assign n5709 = n1173 & ~n5708 ;
  assign n5710 = n1177 & ~n5709 ;
  assign n5711 = n1181 & ~n5710 ;
  assign n5712 = n1185 & ~n5711 ;
  assign n5713 = n1189 & ~n5712 ;
  assign n5714 = n1193 & ~n5713 ;
  assign n5715 = n1197 & ~n5714 ;
  assign n5716 = n1201 & ~n5715 ;
  assign n5717 = n1205 & ~n5716 ;
  assign n5718 = n1209 & ~n5717 ;
  assign n5719 = n1213 & ~n5718 ;
  assign n5720 = n1217 & ~n5719 ;
  assign n5721 = n1221 & ~n5720 ;
  assign n5722 = n1225 & ~n5721 ;
  assign n5723 = n1229 & ~n5722 ;
  assign n5724 = n1233 & ~n5723 ;
  assign n5725 = n1237 & ~n5724 ;
  assign n5726 = n1241 & ~n5725 ;
  assign n5727 = n1245 & ~n5726 ;
  assign n5728 = n1249 & ~n5727 ;
  assign n5729 = n1253 & ~n5728 ;
  assign n5730 = n1257 & ~n5729 ;
  assign n5731 = n1261 & ~n5730 ;
  assign n5732 = n1265 & ~n5731 ;
  assign n5733 = n1269 & ~n5732 ;
  assign n5734 = n1273 & ~n5733 ;
  assign n5735 = n2566 & ~n5734 ;
  assign n5736 = n2568 & ~n5735 ;
  assign n5737 = n3105 & ~n5736 ;
  assign n5738 = n1625 & ~n5737 ;
  assign n5739 = n1629 & ~n5738 ;
  assign n5740 = n1633 & ~n5739 ;
  assign n5741 = n1637 & ~n5740 ;
  assign n5742 = n1641 & ~n5741 ;
  assign n5743 = n1645 & ~n5742 ;
  assign n5744 = n1649 & ~n5743 ;
  assign n5745 = n1653 & ~n5744 ;
  assign n5746 = n1657 & ~n5745 ;
  assign n5747 = n1661 & ~n5746 ;
  assign n5748 = n1665 & ~n5747 ;
  assign n5749 = x150 & ~n1667 ;
  assign n5750 = ~n5748 & n5749 ;
  assign n5838 = n5750 & x278 ;
  assign n5751 = n1335 & ~n2009 ;
  assign n5752 = n1340 & ~n5751 ;
  assign n5753 = n1344 & ~n5752 ;
  assign n5754 = n1348 & ~n5753 ;
  assign n5755 = n1352 & ~n5754 ;
  assign n5756 = n1356 & ~n5755 ;
  assign n5757 = n1360 & ~n5756 ;
  assign n5758 = n1364 & ~n5757 ;
  assign n5759 = n1368 & ~n5758 ;
  assign n5760 = n1372 & ~n5759 ;
  assign n5761 = n1376 & ~n5760 ;
  assign n5762 = n1380 & ~n5761 ;
  assign n5763 = n1384 & ~n5762 ;
  assign n5764 = n1388 & ~n5763 ;
  assign n5765 = n1392 & ~n5764 ;
  assign n5766 = n1396 & ~n5765 ;
  assign n5767 = n1400 & ~n5766 ;
  assign n5768 = n1404 & ~n5767 ;
  assign n5769 = n1408 & ~n5768 ;
  assign n5770 = n1412 & ~n5769 ;
  assign n5771 = n1416 & ~n5770 ;
  assign n5772 = n1420 & ~n5771 ;
  assign n5773 = n1424 & ~n5772 ;
  assign n5774 = n1428 & ~n5773 ;
  assign n5775 = n1432 & ~n5774 ;
  assign n5776 = n1436 & ~n5775 ;
  assign n5777 = n1440 & ~n5776 ;
  assign n5778 = n1444 & ~n5777 ;
  assign n5779 = n1448 & ~n5778 ;
  assign n5780 = n1452 & ~n5779 ;
  assign n5781 = n1456 & ~n5780 ;
  assign n5782 = n1460 & ~n5781 ;
  assign n5783 = n1464 & ~n5782 ;
  assign n5784 = n1468 & ~n5783 ;
  assign n5785 = n1472 & ~n5784 ;
  assign n5786 = n1476 & ~n5785 ;
  assign n5787 = n1480 & ~n5786 ;
  assign n5788 = n1484 & ~n5787 ;
  assign n5789 = n1488 & ~n5788 ;
  assign n5790 = n1492 & ~n5789 ;
  assign n5791 = n1496 & ~n5790 ;
  assign n5792 = n1500 & ~n5791 ;
  assign n5793 = n1504 & ~n5792 ;
  assign n5794 = n1508 & ~n5793 ;
  assign n5795 = n1512 & ~n5794 ;
  assign n5796 = n1516 & ~n5795 ;
  assign n5797 = n1520 & ~n5796 ;
  assign n5798 = n1524 & ~n5797 ;
  assign n5799 = n1528 & ~n5798 ;
  assign n5800 = n1532 & ~n5799 ;
  assign n5801 = n1536 & ~n5800 ;
  assign n5802 = n1540 & ~n5801 ;
  assign n5803 = n1544 & ~n5802 ;
  assign n5804 = n1548 & ~n5803 ;
  assign n5805 = n1552 & ~n5804 ;
  assign n5806 = n1556 & ~n5805 ;
  assign n5807 = n1560 & ~n5806 ;
  assign n5808 = n1564 & ~n5807 ;
  assign n5809 = n1568 & ~n5808 ;
  assign n5810 = n1572 & ~n5809 ;
  assign n5811 = n1576 & ~n5810 ;
  assign n5812 = n1580 & ~n5811 ;
  assign n5813 = n1584 & ~n5812 ;
  assign n5814 = n1588 & ~n5813 ;
  assign n5815 = n1592 & ~n5814 ;
  assign n5816 = n1596 & ~n5815 ;
  assign n5817 = n1600 & ~n5816 ;
  assign n5818 = n1604 & ~n5817 ;
  assign n5819 = n1608 & ~n5818 ;
  assign n5820 = n1612 & ~n5819 ;
  assign n5821 = n2656 & ~n5820 ;
  assign n5822 = n2658 & ~n5821 ;
  assign n5823 = n3192 & ~n5822 ;
  assign n5824 = n1962 & ~n5823 ;
  assign n5825 = n1966 & ~n5824 ;
  assign n5826 = n1970 & ~n5825 ;
  assign n5827 = n1974 & ~n5826 ;
  assign n5828 = n1978 & ~n5827 ;
  assign n5829 = n1982 & ~n5828 ;
  assign n5830 = n1986 & ~n5829 ;
  assign n5831 = n1990 & ~n5830 ;
  assign n5832 = n1994 & ~n5831 ;
  assign n5833 = n1998 & ~n5832 ;
  assign n5834 = n2002 & ~n5833 ;
  assign n5835 = ~x150 & ~n2004 ;
  assign n5836 = ~n5834 & n5835 ;
  assign n5839 = ~n5836 & ~x278 ;
  assign n5840 = ~n5838 & ~n5839 ;
  assign n5841 = ~n318 & n1676 ;
  assign n5842 = n1681 & ~n5841 ;
  assign n5843 = n1685 & ~n5842 ;
  assign n5844 = n1689 & ~n5843 ;
  assign n5845 = n1693 & ~n5844 ;
  assign n5846 = n1697 & ~n5845 ;
  assign n5847 = n1701 & ~n5846 ;
  assign n5848 = n1705 & ~n5847 ;
  assign n5849 = n1709 & ~n5848 ;
  assign n5850 = n1713 & ~n5849 ;
  assign n5851 = n1717 & ~n5850 ;
  assign n5852 = n1721 & ~n5851 ;
  assign n5853 = n1725 & ~n5852 ;
  assign n5854 = n1729 & ~n5853 ;
  assign n5855 = n1733 & ~n5854 ;
  assign n5856 = n1737 & ~n5855 ;
  assign n5857 = n1741 & ~n5856 ;
  assign n5858 = n1745 & ~n5857 ;
  assign n5859 = n1749 & ~n5858 ;
  assign n5860 = n1753 & ~n5859 ;
  assign n5861 = n1757 & ~n5860 ;
  assign n5862 = n1761 & ~n5861 ;
  assign n5863 = n1765 & ~n5862 ;
  assign n5864 = n1769 & ~n5863 ;
  assign n5865 = n1773 & ~n5864 ;
  assign n5866 = n1777 & ~n5865 ;
  assign n5867 = n1781 & ~n5866 ;
  assign n5868 = n1785 & ~n5867 ;
  assign n5869 = n1789 & ~n5868 ;
  assign n5870 = n1793 & ~n5869 ;
  assign n5871 = n1797 & ~n5870 ;
  assign n5872 = n1801 & ~n5871 ;
  assign n5873 = n1805 & ~n5872 ;
  assign n5874 = n1809 & ~n5873 ;
  assign n5875 = n1813 & ~n5874 ;
  assign n5876 = n1817 & ~n5875 ;
  assign n5877 = n1821 & ~n5876 ;
  assign n5878 = n1825 & ~n5877 ;
  assign n5879 = n1829 & ~n5878 ;
  assign n5880 = n1833 & ~n5879 ;
  assign n5881 = n1837 & ~n5880 ;
  assign n5882 = n1841 & ~n5881 ;
  assign n5883 = n1845 & ~n5882 ;
  assign n5884 = n1849 & ~n5883 ;
  assign n5885 = n1853 & ~n5884 ;
  assign n5886 = n1857 & ~n5885 ;
  assign n5887 = n1861 & ~n5886 ;
  assign n5888 = n1865 & ~n5887 ;
  assign n5889 = n1869 & ~n5888 ;
  assign n5890 = n1873 & ~n5889 ;
  assign n5891 = n1877 & ~n5890 ;
  assign n5892 = n1881 & ~n5891 ;
  assign n5893 = n1885 & ~n5892 ;
  assign n5894 = n1889 & ~n5893 ;
  assign n5895 = n1893 & ~n5894 ;
  assign n5896 = n1897 & ~n5895 ;
  assign n5897 = n1901 & ~n5896 ;
  assign n5898 = n1905 & ~n5897 ;
  assign n5899 = n1909 & ~n5898 ;
  assign n5900 = n1913 & ~n5899 ;
  assign n5901 = n1917 & ~n5900 ;
  assign n5902 = n1921 & ~n5901 ;
  assign n5903 = n1925 & ~n5902 ;
  assign n5904 = n1929 & ~n5903 ;
  assign n5905 = n1933 & ~n5904 ;
  assign n5906 = n1937 & ~n5905 ;
  assign n5907 = n1941 & ~n5906 ;
  assign n5908 = n1945 & ~n5907 ;
  assign n5909 = n1949 & ~n5908 ;
  assign n5910 = n1953 & ~n5909 ;
  assign n5911 = n2749 & ~n5910 ;
  assign n5912 = n263 & ~n5911 ;
  assign n5913 = n267 & ~n5912 ;
  assign n5914 = n271 & ~n5913 ;
  assign n5915 = n275 & ~n5914 ;
  assign n5916 = n279 & ~n5915 ;
  assign n5917 = n283 & ~n5916 ;
  assign n5918 = n287 & ~n5917 ;
  assign n5919 = n291 & ~n5918 ;
  assign n5920 = n295 & ~n5919 ;
  assign n5921 = n299 & ~n5920 ;
  assign n5922 = n303 & ~n5921 ;
  assign n5923 = n307 & ~n5922 ;
  assign n5924 = n311 & ~n5923 ;
  assign n5925 = x151 & ~n313 ;
  assign n5926 = ~n5924 & n5925 ;
  assign n6014 = n5926 & x279 ;
  assign n5927 = ~n657 & n2013 ;
  assign n5928 = n2018 & ~n5927 ;
  assign n5929 = n2022 & ~n5928 ;
  assign n5930 = n2026 & ~n5929 ;
  assign n5931 = n2030 & ~n5930 ;
  assign n5932 = n2034 & ~n5931 ;
  assign n5933 = n2038 & ~n5932 ;
  assign n5934 = n2042 & ~n5933 ;
  assign n5935 = n2046 & ~n5934 ;
  assign n5936 = n2050 & ~n5935 ;
  assign n5937 = n2054 & ~n5936 ;
  assign n5938 = n2058 & ~n5937 ;
  assign n5939 = n2062 & ~n5938 ;
  assign n5940 = n2066 & ~n5939 ;
  assign n5941 = n2070 & ~n5940 ;
  assign n5942 = n2074 & ~n5941 ;
  assign n5943 = n2078 & ~n5942 ;
  assign n5944 = n2082 & ~n5943 ;
  assign n5945 = n2086 & ~n5944 ;
  assign n5946 = n2090 & ~n5945 ;
  assign n5947 = n2094 & ~n5946 ;
  assign n5948 = n2098 & ~n5947 ;
  assign n5949 = n2102 & ~n5948 ;
  assign n5950 = n2106 & ~n5949 ;
  assign n5951 = n2110 & ~n5950 ;
  assign n5952 = n2114 & ~n5951 ;
  assign n5953 = n2118 & ~n5952 ;
  assign n5954 = n2122 & ~n5953 ;
  assign n5955 = n2126 & ~n5954 ;
  assign n5956 = n2130 & ~n5955 ;
  assign n5957 = n2134 & ~n5956 ;
  assign n5958 = n2138 & ~n5957 ;
  assign n5959 = n2142 & ~n5958 ;
  assign n5960 = n2146 & ~n5959 ;
  assign n5961 = n2150 & ~n5960 ;
  assign n5962 = n2154 & ~n5961 ;
  assign n5963 = n2158 & ~n5962 ;
  assign n5964 = n2162 & ~n5963 ;
  assign n5965 = n2166 & ~n5964 ;
  assign n5966 = n2170 & ~n5965 ;
  assign n5967 = n2174 & ~n5966 ;
  assign n5968 = n2178 & ~n5967 ;
  assign n5969 = n2182 & ~n5968 ;
  assign n5970 = n2186 & ~n5969 ;
  assign n5971 = n2190 & ~n5970 ;
  assign n5972 = n2194 & ~n5971 ;
  assign n5973 = n2198 & ~n5972 ;
  assign n5974 = n2202 & ~n5973 ;
  assign n5975 = n2206 & ~n5974 ;
  assign n5976 = n2210 & ~n5975 ;
  assign n5977 = n2214 & ~n5976 ;
  assign n5978 = n2218 & ~n5977 ;
  assign n5979 = n2222 & ~n5978 ;
  assign n5980 = n2226 & ~n5979 ;
  assign n5981 = n2230 & ~n5980 ;
  assign n5982 = n2234 & ~n5981 ;
  assign n5983 = n2238 & ~n5982 ;
  assign n5984 = n2242 & ~n5983 ;
  assign n5985 = n2246 & ~n5984 ;
  assign n5986 = n2250 & ~n5985 ;
  assign n5987 = n2254 & ~n5986 ;
  assign n5988 = n2258 & ~n5987 ;
  assign n5989 = n2262 & ~n5988 ;
  assign n5990 = n2266 & ~n5989 ;
  assign n5991 = n2270 & ~n5990 ;
  assign n5992 = n2274 & ~n5991 ;
  assign n5993 = n2278 & ~n5992 ;
  assign n5994 = n2282 & ~n5993 ;
  assign n5995 = n2286 & ~n5994 ;
  assign n5996 = n2290 & ~n5995 ;
  assign n5997 = n2836 & ~n5996 ;
  assign n5998 = n602 & ~n5997 ;
  assign n5999 = n606 & ~n5998 ;
  assign n6000 = n610 & ~n5999 ;
  assign n6001 = n614 & ~n6000 ;
  assign n6002 = n618 & ~n6001 ;
  assign n6003 = n622 & ~n6002 ;
  assign n6004 = n626 & ~n6003 ;
  assign n6005 = n630 & ~n6004 ;
  assign n6006 = n634 & ~n6005 ;
  assign n6007 = n638 & ~n6006 ;
  assign n6008 = n642 & ~n6007 ;
  assign n6009 = n646 & ~n6008 ;
  assign n6010 = n650 & ~n6009 ;
  assign n6011 = ~x151 & ~n652 ;
  assign n6012 = ~n6010 & n6011 ;
  assign n6015 = ~n6012 & ~x279 ;
  assign n6016 = ~n6014 & ~n6015 ;
  assign n6017 = n322 & ~n1000 ;
  assign n6018 = n327 & ~n6017 ;
  assign n6019 = n331 & ~n6018 ;
  assign n6020 = n335 & ~n6019 ;
  assign n6021 = n339 & ~n6020 ;
  assign n6022 = n343 & ~n6021 ;
  assign n6023 = n347 & ~n6022 ;
  assign n6024 = n351 & ~n6023 ;
  assign n6025 = n355 & ~n6024 ;
  assign n6026 = n359 & ~n6025 ;
  assign n6027 = n363 & ~n6026 ;
  assign n6028 = n367 & ~n6027 ;
  assign n6029 = n371 & ~n6028 ;
  assign n6030 = n375 & ~n6029 ;
  assign n6031 = n379 & ~n6030 ;
  assign n6032 = n383 & ~n6031 ;
  assign n6033 = n387 & ~n6032 ;
  assign n6034 = n391 & ~n6033 ;
  assign n6035 = n395 & ~n6034 ;
  assign n6036 = n399 & ~n6035 ;
  assign n6037 = n403 & ~n6036 ;
  assign n6038 = n407 & ~n6037 ;
  assign n6039 = n411 & ~n6038 ;
  assign n6040 = n415 & ~n6039 ;
  assign n6041 = n419 & ~n6040 ;
  assign n6042 = n423 & ~n6041 ;
  assign n6043 = n427 & ~n6042 ;
  assign n6044 = n431 & ~n6043 ;
  assign n6045 = n435 & ~n6044 ;
  assign n6046 = n439 & ~n6045 ;
  assign n6047 = n443 & ~n6046 ;
  assign n6048 = n447 & ~n6047 ;
  assign n6049 = n451 & ~n6048 ;
  assign n6050 = n455 & ~n6049 ;
  assign n6051 = n459 & ~n6050 ;
  assign n6052 = n463 & ~n6051 ;
  assign n6053 = n467 & ~n6052 ;
  assign n6054 = n471 & ~n6053 ;
  assign n6055 = n475 & ~n6054 ;
  assign n6056 = n479 & ~n6055 ;
  assign n6057 = n483 & ~n6056 ;
  assign n6058 = n487 & ~n6057 ;
  assign n6059 = n491 & ~n6058 ;
  assign n6060 = n495 & ~n6059 ;
  assign n6061 = n499 & ~n6060 ;
  assign n6062 = n503 & ~n6061 ;
  assign n6063 = n507 & ~n6062 ;
  assign n6064 = n511 & ~n6063 ;
  assign n6065 = n515 & ~n6064 ;
  assign n6066 = n519 & ~n6065 ;
  assign n6067 = n523 & ~n6066 ;
  assign n6068 = n527 & ~n6067 ;
  assign n6069 = n531 & ~n6068 ;
  assign n6070 = n535 & ~n6069 ;
  assign n6071 = n539 & ~n6070 ;
  assign n6072 = n543 & ~n6071 ;
  assign n6073 = n547 & ~n6072 ;
  assign n6074 = n551 & ~n6073 ;
  assign n6075 = n555 & ~n6074 ;
  assign n6076 = n559 & ~n6075 ;
  assign n6077 = n563 & ~n6076 ;
  assign n6078 = n567 & ~n6077 ;
  assign n6079 = n571 & ~n6078 ;
  assign n6080 = n575 & ~n6079 ;
  assign n6081 = n579 & ~n6080 ;
  assign n6082 = n583 & ~n6081 ;
  assign n6083 = n587 & ~n6082 ;
  assign n6084 = n591 & ~n6083 ;
  assign n6085 = n2382 & ~n6084 ;
  assign n6086 = n2384 & ~n6085 ;
  assign n6087 = n2927 & ~n6086 ;
  assign n6088 = n945 & ~n6087 ;
  assign n6089 = n949 & ~n6088 ;
  assign n6090 = n953 & ~n6089 ;
  assign n6091 = n957 & ~n6090 ;
  assign n6092 = n961 & ~n6091 ;
  assign n6093 = n965 & ~n6092 ;
  assign n6094 = n969 & ~n6093 ;
  assign n6095 = n973 & ~n6094 ;
  assign n6096 = n977 & ~n6095 ;
  assign n6097 = n981 & ~n6096 ;
  assign n6098 = n985 & ~n6097 ;
  assign n6099 = n989 & ~n6098 ;
  assign n6100 = n993 & ~n6099 ;
  assign n6101 = x152 & ~n995 ;
  assign n6102 = ~n6100 & n6101 ;
  assign n6190 = n6102 & x280 ;
  assign n6103 = n661 & ~n1339 ;
  assign n6104 = n666 & ~n6103 ;
  assign n6105 = n670 & ~n6104 ;
  assign n6106 = n674 & ~n6105 ;
  assign n6107 = n678 & ~n6106 ;
  assign n6108 = n682 & ~n6107 ;
  assign n6109 = n686 & ~n6108 ;
  assign n6110 = n690 & ~n6109 ;
  assign n6111 = n694 & ~n6110 ;
  assign n6112 = n698 & ~n6111 ;
  assign n6113 = n702 & ~n6112 ;
  assign n6114 = n706 & ~n6113 ;
  assign n6115 = n710 & ~n6114 ;
  assign n6116 = n714 & ~n6115 ;
  assign n6117 = n718 & ~n6116 ;
  assign n6118 = n722 & ~n6117 ;
  assign n6119 = n726 & ~n6118 ;
  assign n6120 = n730 & ~n6119 ;
  assign n6121 = n734 & ~n6120 ;
  assign n6122 = n738 & ~n6121 ;
  assign n6123 = n742 & ~n6122 ;
  assign n6124 = n746 & ~n6123 ;
  assign n6125 = n750 & ~n6124 ;
  assign n6126 = n754 & ~n6125 ;
  assign n6127 = n758 & ~n6126 ;
  assign n6128 = n762 & ~n6127 ;
  assign n6129 = n766 & ~n6128 ;
  assign n6130 = n770 & ~n6129 ;
  assign n6131 = n774 & ~n6130 ;
  assign n6132 = n778 & ~n6131 ;
  assign n6133 = n782 & ~n6132 ;
  assign n6134 = n786 & ~n6133 ;
  assign n6135 = n790 & ~n6134 ;
  assign n6136 = n794 & ~n6135 ;
  assign n6137 = n798 & ~n6136 ;
  assign n6138 = n802 & ~n6137 ;
  assign n6139 = n806 & ~n6138 ;
  assign n6140 = n810 & ~n6139 ;
  assign n6141 = n814 & ~n6140 ;
  assign n6142 = n818 & ~n6141 ;
  assign n6143 = n822 & ~n6142 ;
  assign n6144 = n826 & ~n6143 ;
  assign n6145 = n830 & ~n6144 ;
  assign n6146 = n834 & ~n6145 ;
  assign n6147 = n838 & ~n6146 ;
  assign n6148 = n842 & ~n6147 ;
  assign n6149 = n846 & ~n6148 ;
  assign n6150 = n850 & ~n6149 ;
  assign n6151 = n854 & ~n6150 ;
  assign n6152 = n858 & ~n6151 ;
  assign n6153 = n862 & ~n6152 ;
  assign n6154 = n866 & ~n6153 ;
  assign n6155 = n870 & ~n6154 ;
  assign n6156 = n874 & ~n6155 ;
  assign n6157 = n878 & ~n6156 ;
  assign n6158 = n882 & ~n6157 ;
  assign n6159 = n886 & ~n6158 ;
  assign n6160 = n890 & ~n6159 ;
  assign n6161 = n894 & ~n6160 ;
  assign n6162 = n898 & ~n6161 ;
  assign n6163 = n902 & ~n6162 ;
  assign n6164 = n906 & ~n6163 ;
  assign n6165 = n910 & ~n6164 ;
  assign n6166 = n914 & ~n6165 ;
  assign n6167 = n918 & ~n6166 ;
  assign n6168 = n922 & ~n6167 ;
  assign n6169 = n926 & ~n6168 ;
  assign n6170 = n930 & ~n6169 ;
  assign n6171 = n2472 & ~n6170 ;
  assign n6172 = n2474 & ~n6171 ;
  assign n6173 = n3014 & ~n6172 ;
  assign n6174 = n1284 & ~n6173 ;
  assign n6175 = n1288 & ~n6174 ;
  assign n6176 = n1292 & ~n6175 ;
  assign n6177 = n1296 & ~n6176 ;
  assign n6178 = n1300 & ~n6177 ;
  assign n6179 = n1304 & ~n6178 ;
  assign n6180 = n1308 & ~n6179 ;
  assign n6181 = n1312 & ~n6180 ;
  assign n6182 = n1316 & ~n6181 ;
  assign n6183 = n1320 & ~n6182 ;
  assign n6184 = n1324 & ~n6183 ;
  assign n6185 = n1328 & ~n6184 ;
  assign n6186 = n1332 & ~n6185 ;
  assign n6187 = ~x152 & ~n1334 ;
  assign n6188 = ~n6186 & n6187 ;
  assign n6191 = ~n6188 & ~x280 ;
  assign n6192 = ~n6190 & ~n6191 ;
  assign n6193 = n1004 & ~n1680 ;
  assign n6194 = n1009 & ~n6193 ;
  assign n6195 = n1013 & ~n6194 ;
  assign n6196 = n1017 & ~n6195 ;
  assign n6197 = n1021 & ~n6196 ;
  assign n6198 = n1025 & ~n6197 ;
  assign n6199 = n1029 & ~n6198 ;
  assign n6200 = n1033 & ~n6199 ;
  assign n6201 = n1037 & ~n6200 ;
  assign n6202 = n1041 & ~n6201 ;
  assign n6203 = n1045 & ~n6202 ;
  assign n6204 = n1049 & ~n6203 ;
  assign n6205 = n1053 & ~n6204 ;
  assign n6206 = n1057 & ~n6205 ;
  assign n6207 = n1061 & ~n6206 ;
  assign n6208 = n1065 & ~n6207 ;
  assign n6209 = n1069 & ~n6208 ;
  assign n6210 = n1073 & ~n6209 ;
  assign n6211 = n1077 & ~n6210 ;
  assign n6212 = n1081 & ~n6211 ;
  assign n6213 = n1085 & ~n6212 ;
  assign n6214 = n1089 & ~n6213 ;
  assign n6215 = n1093 & ~n6214 ;
  assign n6216 = n1097 & ~n6215 ;
  assign n6217 = n1101 & ~n6216 ;
  assign n6218 = n1105 & ~n6217 ;
  assign n6219 = n1109 & ~n6218 ;
  assign n6220 = n1113 & ~n6219 ;
  assign n6221 = n1117 & ~n6220 ;
  assign n6222 = n1121 & ~n6221 ;
  assign n6223 = n1125 & ~n6222 ;
  assign n6224 = n1129 & ~n6223 ;
  assign n6225 = n1133 & ~n6224 ;
  assign n6226 = n1137 & ~n6225 ;
  assign n6227 = n1141 & ~n6226 ;
  assign n6228 = n1145 & ~n6227 ;
  assign n6229 = n1149 & ~n6228 ;
  assign n6230 = n1153 & ~n6229 ;
  assign n6231 = n1157 & ~n6230 ;
  assign n6232 = n1161 & ~n6231 ;
  assign n6233 = n1165 & ~n6232 ;
  assign n6234 = n1169 & ~n6233 ;
  assign n6235 = n1173 & ~n6234 ;
  assign n6236 = n1177 & ~n6235 ;
  assign n6237 = n1181 & ~n6236 ;
  assign n6238 = n1185 & ~n6237 ;
  assign n6239 = n1189 & ~n6238 ;
  assign n6240 = n1193 & ~n6239 ;
  assign n6241 = n1197 & ~n6240 ;
  assign n6242 = n1201 & ~n6241 ;
  assign n6243 = n1205 & ~n6242 ;
  assign n6244 = n1209 & ~n6243 ;
  assign n6245 = n1213 & ~n6244 ;
  assign n6246 = n1217 & ~n6245 ;
  assign n6247 = n1221 & ~n6246 ;
  assign n6248 = n1225 & ~n6247 ;
  assign n6249 = n1229 & ~n6248 ;
  assign n6250 = n1233 & ~n6249 ;
  assign n6251 = n1237 & ~n6250 ;
  assign n6252 = n1241 & ~n6251 ;
  assign n6253 = n1245 & ~n6252 ;
  assign n6254 = n1249 & ~n6253 ;
  assign n6255 = n1253 & ~n6254 ;
  assign n6256 = n1257 & ~n6255 ;
  assign n6257 = n1261 & ~n6256 ;
  assign n6258 = n1265 & ~n6257 ;
  assign n6259 = n1269 & ~n6258 ;
  assign n6260 = n1273 & ~n6259 ;
  assign n6261 = n2566 & ~n6260 ;
  assign n6262 = n2568 & ~n6261 ;
  assign n6263 = n3105 & ~n6262 ;
  assign n6264 = n1625 & ~n6263 ;
  assign n6265 = n1629 & ~n6264 ;
  assign n6266 = n1633 & ~n6265 ;
  assign n6267 = n1637 & ~n6266 ;
  assign n6268 = n1641 & ~n6267 ;
  assign n6269 = n1645 & ~n6268 ;
  assign n6270 = n1649 & ~n6269 ;
  assign n6271 = n1653 & ~n6270 ;
  assign n6272 = n1657 & ~n6271 ;
  assign n6273 = n1661 & ~n6272 ;
  assign n6274 = n1665 & ~n6273 ;
  assign n6275 = n1669 & ~n6274 ;
  assign n6276 = n1673 & ~n6275 ;
  assign n6277 = x153 & ~n1675 ;
  assign n6278 = ~n6276 & n6277 ;
  assign n6366 = n6278 & x281 ;
  assign n6279 = n1343 & ~n2017 ;
  assign n6280 = n1348 & ~n6279 ;
  assign n6281 = n1352 & ~n6280 ;
  assign n6282 = n1356 & ~n6281 ;
  assign n6283 = n1360 & ~n6282 ;
  assign n6284 = n1364 & ~n6283 ;
  assign n6285 = n1368 & ~n6284 ;
  assign n6286 = n1372 & ~n6285 ;
  assign n6287 = n1376 & ~n6286 ;
  assign n6288 = n1380 & ~n6287 ;
  assign n6289 = n1384 & ~n6288 ;
  assign n6290 = n1388 & ~n6289 ;
  assign n6291 = n1392 & ~n6290 ;
  assign n6292 = n1396 & ~n6291 ;
  assign n6293 = n1400 & ~n6292 ;
  assign n6294 = n1404 & ~n6293 ;
  assign n6295 = n1408 & ~n6294 ;
  assign n6296 = n1412 & ~n6295 ;
  assign n6297 = n1416 & ~n6296 ;
  assign n6298 = n1420 & ~n6297 ;
  assign n6299 = n1424 & ~n6298 ;
  assign n6300 = n1428 & ~n6299 ;
  assign n6301 = n1432 & ~n6300 ;
  assign n6302 = n1436 & ~n6301 ;
  assign n6303 = n1440 & ~n6302 ;
  assign n6304 = n1444 & ~n6303 ;
  assign n6305 = n1448 & ~n6304 ;
  assign n6306 = n1452 & ~n6305 ;
  assign n6307 = n1456 & ~n6306 ;
  assign n6308 = n1460 & ~n6307 ;
  assign n6309 = n1464 & ~n6308 ;
  assign n6310 = n1468 & ~n6309 ;
  assign n6311 = n1472 & ~n6310 ;
  assign n6312 = n1476 & ~n6311 ;
  assign n6313 = n1480 & ~n6312 ;
  assign n6314 = n1484 & ~n6313 ;
  assign n6315 = n1488 & ~n6314 ;
  assign n6316 = n1492 & ~n6315 ;
  assign n6317 = n1496 & ~n6316 ;
  assign n6318 = n1500 & ~n6317 ;
  assign n6319 = n1504 & ~n6318 ;
  assign n6320 = n1508 & ~n6319 ;
  assign n6321 = n1512 & ~n6320 ;
  assign n6322 = n1516 & ~n6321 ;
  assign n6323 = n1520 & ~n6322 ;
  assign n6324 = n1524 & ~n6323 ;
  assign n6325 = n1528 & ~n6324 ;
  assign n6326 = n1532 & ~n6325 ;
  assign n6327 = n1536 & ~n6326 ;
  assign n6328 = n1540 & ~n6327 ;
  assign n6329 = n1544 & ~n6328 ;
  assign n6330 = n1548 & ~n6329 ;
  assign n6331 = n1552 & ~n6330 ;
  assign n6332 = n1556 & ~n6331 ;
  assign n6333 = n1560 & ~n6332 ;
  assign n6334 = n1564 & ~n6333 ;
  assign n6335 = n1568 & ~n6334 ;
  assign n6336 = n1572 & ~n6335 ;
  assign n6337 = n1576 & ~n6336 ;
  assign n6338 = n1580 & ~n6337 ;
  assign n6339 = n1584 & ~n6338 ;
  assign n6340 = n1588 & ~n6339 ;
  assign n6341 = n1592 & ~n6340 ;
  assign n6342 = n1596 & ~n6341 ;
  assign n6343 = n1600 & ~n6342 ;
  assign n6344 = n1604 & ~n6343 ;
  assign n6345 = n1608 & ~n6344 ;
  assign n6346 = n1612 & ~n6345 ;
  assign n6347 = n2656 & ~n6346 ;
  assign n6348 = n2658 & ~n6347 ;
  assign n6349 = n3192 & ~n6348 ;
  assign n6350 = n1962 & ~n6349 ;
  assign n6351 = n1966 & ~n6350 ;
  assign n6352 = n1970 & ~n6351 ;
  assign n6353 = n1974 & ~n6352 ;
  assign n6354 = n1978 & ~n6353 ;
  assign n6355 = n1982 & ~n6354 ;
  assign n6356 = n1986 & ~n6355 ;
  assign n6357 = n1990 & ~n6356 ;
  assign n6358 = n1994 & ~n6357 ;
  assign n6359 = n1998 & ~n6358 ;
  assign n6360 = n2002 & ~n6359 ;
  assign n6361 = n2006 & ~n6360 ;
  assign n6362 = n2010 & ~n6361 ;
  assign n6363 = ~x153 & ~n2012 ;
  assign n6364 = ~n6362 & n6363 ;
  assign n6367 = ~n6364 & ~x281 ;
  assign n6368 = ~n6366 & ~n6367 ;
  assign n6369 = ~n326 & n1684 ;
  assign n6370 = n1689 & ~n6369 ;
  assign n6371 = n1693 & ~n6370 ;
  assign n6372 = n1697 & ~n6371 ;
  assign n6373 = n1701 & ~n6372 ;
  assign n6374 = n1705 & ~n6373 ;
  assign n6375 = n1709 & ~n6374 ;
  assign n6376 = n1713 & ~n6375 ;
  assign n6377 = n1717 & ~n6376 ;
  assign n6378 = n1721 & ~n6377 ;
  assign n6379 = n1725 & ~n6378 ;
  assign n6380 = n1729 & ~n6379 ;
  assign n6381 = n1733 & ~n6380 ;
  assign n6382 = n1737 & ~n6381 ;
  assign n6383 = n1741 & ~n6382 ;
  assign n6384 = n1745 & ~n6383 ;
  assign n6385 = n1749 & ~n6384 ;
  assign n6386 = n1753 & ~n6385 ;
  assign n6387 = n1757 & ~n6386 ;
  assign n6388 = n1761 & ~n6387 ;
  assign n6389 = n1765 & ~n6388 ;
  assign n6390 = n1769 & ~n6389 ;
  assign n6391 = n1773 & ~n6390 ;
  assign n6392 = n1777 & ~n6391 ;
  assign n6393 = n1781 & ~n6392 ;
  assign n6394 = n1785 & ~n6393 ;
  assign n6395 = n1789 & ~n6394 ;
  assign n6396 = n1793 & ~n6395 ;
  assign n6397 = n1797 & ~n6396 ;
  assign n6398 = n1801 & ~n6397 ;
  assign n6399 = n1805 & ~n6398 ;
  assign n6400 = n1809 & ~n6399 ;
  assign n6401 = n1813 & ~n6400 ;
  assign n6402 = n1817 & ~n6401 ;
  assign n6403 = n1821 & ~n6402 ;
  assign n6404 = n1825 & ~n6403 ;
  assign n6405 = n1829 & ~n6404 ;
  assign n6406 = n1833 & ~n6405 ;
  assign n6407 = n1837 & ~n6406 ;
  assign n6408 = n1841 & ~n6407 ;
  assign n6409 = n1845 & ~n6408 ;
  assign n6410 = n1849 & ~n6409 ;
  assign n6411 = n1853 & ~n6410 ;
  assign n6412 = n1857 & ~n6411 ;
  assign n6413 = n1861 & ~n6412 ;
  assign n6414 = n1865 & ~n6413 ;
  assign n6415 = n1869 & ~n6414 ;
  assign n6416 = n1873 & ~n6415 ;
  assign n6417 = n1877 & ~n6416 ;
  assign n6418 = n1881 & ~n6417 ;
  assign n6419 = n1885 & ~n6418 ;
  assign n6420 = n1889 & ~n6419 ;
  assign n6421 = n1893 & ~n6420 ;
  assign n6422 = n1897 & ~n6421 ;
  assign n6423 = n1901 & ~n6422 ;
  assign n6424 = n1905 & ~n6423 ;
  assign n6425 = n1909 & ~n6424 ;
  assign n6426 = n1913 & ~n6425 ;
  assign n6427 = n1917 & ~n6426 ;
  assign n6428 = n1921 & ~n6427 ;
  assign n6429 = n1925 & ~n6428 ;
  assign n6430 = n1929 & ~n6429 ;
  assign n6431 = n1933 & ~n6430 ;
  assign n6432 = n1937 & ~n6431 ;
  assign n6433 = n1941 & ~n6432 ;
  assign n6434 = n1945 & ~n6433 ;
  assign n6435 = n1949 & ~n6434 ;
  assign n6436 = n1953 & ~n6435 ;
  assign n6437 = n2749 & ~n6436 ;
  assign n6438 = n263 & ~n6437 ;
  assign n6439 = n267 & ~n6438 ;
  assign n6440 = n271 & ~n6439 ;
  assign n6441 = n275 & ~n6440 ;
  assign n6442 = n279 & ~n6441 ;
  assign n6443 = n283 & ~n6442 ;
  assign n6444 = n287 & ~n6443 ;
  assign n6445 = n291 & ~n6444 ;
  assign n6446 = n295 & ~n6445 ;
  assign n6447 = n299 & ~n6446 ;
  assign n6448 = n303 & ~n6447 ;
  assign n6449 = n307 & ~n6448 ;
  assign n6450 = n311 & ~n6449 ;
  assign n6451 = n315 & ~n6450 ;
  assign n6452 = n319 & ~n6451 ;
  assign n6453 = x154 & ~n321 ;
  assign n6454 = ~n6452 & n6453 ;
  assign n6542 = n6454 & x282 ;
  assign n6455 = ~n665 & n2021 ;
  assign n6456 = n2026 & ~n6455 ;
  assign n6457 = n2030 & ~n6456 ;
  assign n6458 = n2034 & ~n6457 ;
  assign n6459 = n2038 & ~n6458 ;
  assign n6460 = n2042 & ~n6459 ;
  assign n6461 = n2046 & ~n6460 ;
  assign n6462 = n2050 & ~n6461 ;
  assign n6463 = n2054 & ~n6462 ;
  assign n6464 = n2058 & ~n6463 ;
  assign n6465 = n2062 & ~n6464 ;
  assign n6466 = n2066 & ~n6465 ;
  assign n6467 = n2070 & ~n6466 ;
  assign n6468 = n2074 & ~n6467 ;
  assign n6469 = n2078 & ~n6468 ;
  assign n6470 = n2082 & ~n6469 ;
  assign n6471 = n2086 & ~n6470 ;
  assign n6472 = n2090 & ~n6471 ;
  assign n6473 = n2094 & ~n6472 ;
  assign n6474 = n2098 & ~n6473 ;
  assign n6475 = n2102 & ~n6474 ;
  assign n6476 = n2106 & ~n6475 ;
  assign n6477 = n2110 & ~n6476 ;
  assign n6478 = n2114 & ~n6477 ;
  assign n6479 = n2118 & ~n6478 ;
  assign n6480 = n2122 & ~n6479 ;
  assign n6481 = n2126 & ~n6480 ;
  assign n6482 = n2130 & ~n6481 ;
  assign n6483 = n2134 & ~n6482 ;
  assign n6484 = n2138 & ~n6483 ;
  assign n6485 = n2142 & ~n6484 ;
  assign n6486 = n2146 & ~n6485 ;
  assign n6487 = n2150 & ~n6486 ;
  assign n6488 = n2154 & ~n6487 ;
  assign n6489 = n2158 & ~n6488 ;
  assign n6490 = n2162 & ~n6489 ;
  assign n6491 = n2166 & ~n6490 ;
  assign n6492 = n2170 & ~n6491 ;
  assign n6493 = n2174 & ~n6492 ;
  assign n6494 = n2178 & ~n6493 ;
  assign n6495 = n2182 & ~n6494 ;
  assign n6496 = n2186 & ~n6495 ;
  assign n6497 = n2190 & ~n6496 ;
  assign n6498 = n2194 & ~n6497 ;
  assign n6499 = n2198 & ~n6498 ;
  assign n6500 = n2202 & ~n6499 ;
  assign n6501 = n2206 & ~n6500 ;
  assign n6502 = n2210 & ~n6501 ;
  assign n6503 = n2214 & ~n6502 ;
  assign n6504 = n2218 & ~n6503 ;
  assign n6505 = n2222 & ~n6504 ;
  assign n6506 = n2226 & ~n6505 ;
  assign n6507 = n2230 & ~n6506 ;
  assign n6508 = n2234 & ~n6507 ;
  assign n6509 = n2238 & ~n6508 ;
  assign n6510 = n2242 & ~n6509 ;
  assign n6511 = n2246 & ~n6510 ;
  assign n6512 = n2250 & ~n6511 ;
  assign n6513 = n2254 & ~n6512 ;
  assign n6514 = n2258 & ~n6513 ;
  assign n6515 = n2262 & ~n6514 ;
  assign n6516 = n2266 & ~n6515 ;
  assign n6517 = n2270 & ~n6516 ;
  assign n6518 = n2274 & ~n6517 ;
  assign n6519 = n2278 & ~n6518 ;
  assign n6520 = n2282 & ~n6519 ;
  assign n6521 = n2286 & ~n6520 ;
  assign n6522 = n2290 & ~n6521 ;
  assign n6523 = n2836 & ~n6522 ;
  assign n6524 = n602 & ~n6523 ;
  assign n6525 = n606 & ~n6524 ;
  assign n6526 = n610 & ~n6525 ;
  assign n6527 = n614 & ~n6526 ;
  assign n6528 = n618 & ~n6527 ;
  assign n6529 = n622 & ~n6528 ;
  assign n6530 = n626 & ~n6529 ;
  assign n6531 = n630 & ~n6530 ;
  assign n6532 = n634 & ~n6531 ;
  assign n6533 = n638 & ~n6532 ;
  assign n6534 = n642 & ~n6533 ;
  assign n6535 = n646 & ~n6534 ;
  assign n6536 = n650 & ~n6535 ;
  assign n6537 = n654 & ~n6536 ;
  assign n6538 = n658 & ~n6537 ;
  assign n6539 = ~x154 & ~n660 ;
  assign n6540 = ~n6538 & n6539 ;
  assign n6543 = ~n6540 & ~x282 ;
  assign n6544 = ~n6542 & ~n6543 ;
  assign n6545 = n330 & ~n1008 ;
  assign n6546 = n335 & ~n6545 ;
  assign n6547 = n339 & ~n6546 ;
  assign n6548 = n343 & ~n6547 ;
  assign n6549 = n347 & ~n6548 ;
  assign n6550 = n351 & ~n6549 ;
  assign n6551 = n355 & ~n6550 ;
  assign n6552 = n359 & ~n6551 ;
  assign n6553 = n363 & ~n6552 ;
  assign n6554 = n367 & ~n6553 ;
  assign n6555 = n371 & ~n6554 ;
  assign n6556 = n375 & ~n6555 ;
  assign n6557 = n379 & ~n6556 ;
  assign n6558 = n383 & ~n6557 ;
  assign n6559 = n387 & ~n6558 ;
  assign n6560 = n391 & ~n6559 ;
  assign n6561 = n395 & ~n6560 ;
  assign n6562 = n399 & ~n6561 ;
  assign n6563 = n403 & ~n6562 ;
  assign n6564 = n407 & ~n6563 ;
  assign n6565 = n411 & ~n6564 ;
  assign n6566 = n415 & ~n6565 ;
  assign n6567 = n419 & ~n6566 ;
  assign n6568 = n423 & ~n6567 ;
  assign n6569 = n427 & ~n6568 ;
  assign n6570 = n431 & ~n6569 ;
  assign n6571 = n435 & ~n6570 ;
  assign n6572 = n439 & ~n6571 ;
  assign n6573 = n443 & ~n6572 ;
  assign n6574 = n447 & ~n6573 ;
  assign n6575 = n451 & ~n6574 ;
  assign n6576 = n455 & ~n6575 ;
  assign n6577 = n459 & ~n6576 ;
  assign n6578 = n463 & ~n6577 ;
  assign n6579 = n467 & ~n6578 ;
  assign n6580 = n471 & ~n6579 ;
  assign n6581 = n475 & ~n6580 ;
  assign n6582 = n479 & ~n6581 ;
  assign n6583 = n483 & ~n6582 ;
  assign n6584 = n487 & ~n6583 ;
  assign n6585 = n491 & ~n6584 ;
  assign n6586 = n495 & ~n6585 ;
  assign n6587 = n499 & ~n6586 ;
  assign n6588 = n503 & ~n6587 ;
  assign n6589 = n507 & ~n6588 ;
  assign n6590 = n511 & ~n6589 ;
  assign n6591 = n515 & ~n6590 ;
  assign n6592 = n519 & ~n6591 ;
  assign n6593 = n523 & ~n6592 ;
  assign n6594 = n527 & ~n6593 ;
  assign n6595 = n531 & ~n6594 ;
  assign n6596 = n535 & ~n6595 ;
  assign n6597 = n539 & ~n6596 ;
  assign n6598 = n543 & ~n6597 ;
  assign n6599 = n547 & ~n6598 ;
  assign n6600 = n551 & ~n6599 ;
  assign n6601 = n555 & ~n6600 ;
  assign n6602 = n559 & ~n6601 ;
  assign n6603 = n563 & ~n6602 ;
  assign n6604 = n567 & ~n6603 ;
  assign n6605 = n571 & ~n6604 ;
  assign n6606 = n575 & ~n6605 ;
  assign n6607 = n579 & ~n6606 ;
  assign n6608 = n583 & ~n6607 ;
  assign n6609 = n587 & ~n6608 ;
  assign n6610 = n591 & ~n6609 ;
  assign n6611 = n2382 & ~n6610 ;
  assign n6612 = n2384 & ~n6611 ;
  assign n6613 = n2927 & ~n6612 ;
  assign n6614 = n945 & ~n6613 ;
  assign n6615 = n949 & ~n6614 ;
  assign n6616 = n953 & ~n6615 ;
  assign n6617 = n957 & ~n6616 ;
  assign n6618 = n961 & ~n6617 ;
  assign n6619 = n965 & ~n6618 ;
  assign n6620 = n969 & ~n6619 ;
  assign n6621 = n973 & ~n6620 ;
  assign n6622 = n977 & ~n6621 ;
  assign n6623 = n981 & ~n6622 ;
  assign n6624 = n985 & ~n6623 ;
  assign n6625 = n989 & ~n6624 ;
  assign n6626 = n993 & ~n6625 ;
  assign n6627 = n997 & ~n6626 ;
  assign n6628 = n1001 & ~n6627 ;
  assign n6629 = x155 & ~n1003 ;
  assign n6630 = ~n6628 & n6629 ;
  assign n6718 = n6630 & x283 ;
  assign n6631 = n669 & ~n1347 ;
  assign n6632 = n674 & ~n6631 ;
  assign n6633 = n678 & ~n6632 ;
  assign n6634 = n682 & ~n6633 ;
  assign n6635 = n686 & ~n6634 ;
  assign n6636 = n690 & ~n6635 ;
  assign n6637 = n694 & ~n6636 ;
  assign n6638 = n698 & ~n6637 ;
  assign n6639 = n702 & ~n6638 ;
  assign n6640 = n706 & ~n6639 ;
  assign n6641 = n710 & ~n6640 ;
  assign n6642 = n714 & ~n6641 ;
  assign n6643 = n718 & ~n6642 ;
  assign n6644 = n722 & ~n6643 ;
  assign n6645 = n726 & ~n6644 ;
  assign n6646 = n730 & ~n6645 ;
  assign n6647 = n734 & ~n6646 ;
  assign n6648 = n738 & ~n6647 ;
  assign n6649 = n742 & ~n6648 ;
  assign n6650 = n746 & ~n6649 ;
  assign n6651 = n750 & ~n6650 ;
  assign n6652 = n754 & ~n6651 ;
  assign n6653 = n758 & ~n6652 ;
  assign n6654 = n762 & ~n6653 ;
  assign n6655 = n766 & ~n6654 ;
  assign n6656 = n770 & ~n6655 ;
  assign n6657 = n774 & ~n6656 ;
  assign n6658 = n778 & ~n6657 ;
  assign n6659 = n782 & ~n6658 ;
  assign n6660 = n786 & ~n6659 ;
  assign n6661 = n790 & ~n6660 ;
  assign n6662 = n794 & ~n6661 ;
  assign n6663 = n798 & ~n6662 ;
  assign n6664 = n802 & ~n6663 ;
  assign n6665 = n806 & ~n6664 ;
  assign n6666 = n810 & ~n6665 ;
  assign n6667 = n814 & ~n6666 ;
  assign n6668 = n818 & ~n6667 ;
  assign n6669 = n822 & ~n6668 ;
  assign n6670 = n826 & ~n6669 ;
  assign n6671 = n830 & ~n6670 ;
  assign n6672 = n834 & ~n6671 ;
  assign n6673 = n838 & ~n6672 ;
  assign n6674 = n842 & ~n6673 ;
  assign n6675 = n846 & ~n6674 ;
  assign n6676 = n850 & ~n6675 ;
  assign n6677 = n854 & ~n6676 ;
  assign n6678 = n858 & ~n6677 ;
  assign n6679 = n862 & ~n6678 ;
  assign n6680 = n866 & ~n6679 ;
  assign n6681 = n870 & ~n6680 ;
  assign n6682 = n874 & ~n6681 ;
  assign n6683 = n878 & ~n6682 ;
  assign n6684 = n882 & ~n6683 ;
  assign n6685 = n886 & ~n6684 ;
  assign n6686 = n890 & ~n6685 ;
  assign n6687 = n894 & ~n6686 ;
  assign n6688 = n898 & ~n6687 ;
  assign n6689 = n902 & ~n6688 ;
  assign n6690 = n906 & ~n6689 ;
  assign n6691 = n910 & ~n6690 ;
  assign n6692 = n914 & ~n6691 ;
  assign n6693 = n918 & ~n6692 ;
  assign n6694 = n922 & ~n6693 ;
  assign n6695 = n926 & ~n6694 ;
  assign n6696 = n930 & ~n6695 ;
  assign n6697 = n2472 & ~n6696 ;
  assign n6698 = n2474 & ~n6697 ;
  assign n6699 = n3014 & ~n6698 ;
  assign n6700 = n1284 & ~n6699 ;
  assign n6701 = n1288 & ~n6700 ;
  assign n6702 = n1292 & ~n6701 ;
  assign n6703 = n1296 & ~n6702 ;
  assign n6704 = n1300 & ~n6703 ;
  assign n6705 = n1304 & ~n6704 ;
  assign n6706 = n1308 & ~n6705 ;
  assign n6707 = n1312 & ~n6706 ;
  assign n6708 = n1316 & ~n6707 ;
  assign n6709 = n1320 & ~n6708 ;
  assign n6710 = n1324 & ~n6709 ;
  assign n6711 = n1328 & ~n6710 ;
  assign n6712 = n1332 & ~n6711 ;
  assign n6713 = n1336 & ~n6712 ;
  assign n6714 = n1340 & ~n6713 ;
  assign n6715 = ~x155 & ~n1342 ;
  assign n6716 = ~n6714 & n6715 ;
  assign n6719 = ~n6716 & ~x283 ;
  assign n6720 = ~n6718 & ~n6719 ;
  assign n6721 = n1012 & ~n1688 ;
  assign n6722 = n1017 & ~n6721 ;
  assign n6723 = n1021 & ~n6722 ;
  assign n6724 = n1025 & ~n6723 ;
  assign n6725 = n1029 & ~n6724 ;
  assign n6726 = n1033 & ~n6725 ;
  assign n6727 = n1037 & ~n6726 ;
  assign n6728 = n1041 & ~n6727 ;
  assign n6729 = n1045 & ~n6728 ;
  assign n6730 = n1049 & ~n6729 ;
  assign n6731 = n1053 & ~n6730 ;
  assign n6732 = n1057 & ~n6731 ;
  assign n6733 = n1061 & ~n6732 ;
  assign n6734 = n1065 & ~n6733 ;
  assign n6735 = n1069 & ~n6734 ;
  assign n6736 = n1073 & ~n6735 ;
  assign n6737 = n1077 & ~n6736 ;
  assign n6738 = n1081 & ~n6737 ;
  assign n6739 = n1085 & ~n6738 ;
  assign n6740 = n1089 & ~n6739 ;
  assign n6741 = n1093 & ~n6740 ;
  assign n6742 = n1097 & ~n6741 ;
  assign n6743 = n1101 & ~n6742 ;
  assign n6744 = n1105 & ~n6743 ;
  assign n6745 = n1109 & ~n6744 ;
  assign n6746 = n1113 & ~n6745 ;
  assign n6747 = n1117 & ~n6746 ;
  assign n6748 = n1121 & ~n6747 ;
  assign n6749 = n1125 & ~n6748 ;
  assign n6750 = n1129 & ~n6749 ;
  assign n6751 = n1133 & ~n6750 ;
  assign n6752 = n1137 & ~n6751 ;
  assign n6753 = n1141 & ~n6752 ;
  assign n6754 = n1145 & ~n6753 ;
  assign n6755 = n1149 & ~n6754 ;
  assign n6756 = n1153 & ~n6755 ;
  assign n6757 = n1157 & ~n6756 ;
  assign n6758 = n1161 & ~n6757 ;
  assign n6759 = n1165 & ~n6758 ;
  assign n6760 = n1169 & ~n6759 ;
  assign n6761 = n1173 & ~n6760 ;
  assign n6762 = n1177 & ~n6761 ;
  assign n6763 = n1181 & ~n6762 ;
  assign n6764 = n1185 & ~n6763 ;
  assign n6765 = n1189 & ~n6764 ;
  assign n6766 = n1193 & ~n6765 ;
  assign n6767 = n1197 & ~n6766 ;
  assign n6768 = n1201 & ~n6767 ;
  assign n6769 = n1205 & ~n6768 ;
  assign n6770 = n1209 & ~n6769 ;
  assign n6771 = n1213 & ~n6770 ;
  assign n6772 = n1217 & ~n6771 ;
  assign n6773 = n1221 & ~n6772 ;
  assign n6774 = n1225 & ~n6773 ;
  assign n6775 = n1229 & ~n6774 ;
  assign n6776 = n1233 & ~n6775 ;
  assign n6777 = n1237 & ~n6776 ;
  assign n6778 = n1241 & ~n6777 ;
  assign n6779 = n1245 & ~n6778 ;
  assign n6780 = n1249 & ~n6779 ;
  assign n6781 = n1253 & ~n6780 ;
  assign n6782 = n1257 & ~n6781 ;
  assign n6783 = n1261 & ~n6782 ;
  assign n6784 = n1265 & ~n6783 ;
  assign n6785 = n1269 & ~n6784 ;
  assign n6786 = n1273 & ~n6785 ;
  assign n6787 = n2566 & ~n6786 ;
  assign n6788 = n2568 & ~n6787 ;
  assign n6789 = n3105 & ~n6788 ;
  assign n6790 = n1625 & ~n6789 ;
  assign n6791 = n1629 & ~n6790 ;
  assign n6792 = n1633 & ~n6791 ;
  assign n6793 = n1637 & ~n6792 ;
  assign n6794 = n1641 & ~n6793 ;
  assign n6795 = n1645 & ~n6794 ;
  assign n6796 = n1649 & ~n6795 ;
  assign n6797 = n1653 & ~n6796 ;
  assign n6798 = n1657 & ~n6797 ;
  assign n6799 = n1661 & ~n6798 ;
  assign n6800 = n1665 & ~n6799 ;
  assign n6801 = n1669 & ~n6800 ;
  assign n6802 = n1673 & ~n6801 ;
  assign n6803 = n1677 & ~n6802 ;
  assign n6804 = n1681 & ~n6803 ;
  assign n6805 = x156 & ~n1683 ;
  assign n6806 = ~n6804 & n6805 ;
  assign n6894 = n6806 & x284 ;
  assign n6807 = n1351 & ~n2025 ;
  assign n6808 = n1356 & ~n6807 ;
  assign n6809 = n1360 & ~n6808 ;
  assign n6810 = n1364 & ~n6809 ;
  assign n6811 = n1368 & ~n6810 ;
  assign n6812 = n1372 & ~n6811 ;
  assign n6813 = n1376 & ~n6812 ;
  assign n6814 = n1380 & ~n6813 ;
  assign n6815 = n1384 & ~n6814 ;
  assign n6816 = n1388 & ~n6815 ;
  assign n6817 = n1392 & ~n6816 ;
  assign n6818 = n1396 & ~n6817 ;
  assign n6819 = n1400 & ~n6818 ;
  assign n6820 = n1404 & ~n6819 ;
  assign n6821 = n1408 & ~n6820 ;
  assign n6822 = n1412 & ~n6821 ;
  assign n6823 = n1416 & ~n6822 ;
  assign n6824 = n1420 & ~n6823 ;
  assign n6825 = n1424 & ~n6824 ;
  assign n6826 = n1428 & ~n6825 ;
  assign n6827 = n1432 & ~n6826 ;
  assign n6828 = n1436 & ~n6827 ;
  assign n6829 = n1440 & ~n6828 ;
  assign n6830 = n1444 & ~n6829 ;
  assign n6831 = n1448 & ~n6830 ;
  assign n6832 = n1452 & ~n6831 ;
  assign n6833 = n1456 & ~n6832 ;
  assign n6834 = n1460 & ~n6833 ;
  assign n6835 = n1464 & ~n6834 ;
  assign n6836 = n1468 & ~n6835 ;
  assign n6837 = n1472 & ~n6836 ;
  assign n6838 = n1476 & ~n6837 ;
  assign n6839 = n1480 & ~n6838 ;
  assign n6840 = n1484 & ~n6839 ;
  assign n6841 = n1488 & ~n6840 ;
  assign n6842 = n1492 & ~n6841 ;
  assign n6843 = n1496 & ~n6842 ;
  assign n6844 = n1500 & ~n6843 ;
  assign n6845 = n1504 & ~n6844 ;
  assign n6846 = n1508 & ~n6845 ;
  assign n6847 = n1512 & ~n6846 ;
  assign n6848 = n1516 & ~n6847 ;
  assign n6849 = n1520 & ~n6848 ;
  assign n6850 = n1524 & ~n6849 ;
  assign n6851 = n1528 & ~n6850 ;
  assign n6852 = n1532 & ~n6851 ;
  assign n6853 = n1536 & ~n6852 ;
  assign n6854 = n1540 & ~n6853 ;
  assign n6855 = n1544 & ~n6854 ;
  assign n6856 = n1548 & ~n6855 ;
  assign n6857 = n1552 & ~n6856 ;
  assign n6858 = n1556 & ~n6857 ;
  assign n6859 = n1560 & ~n6858 ;
  assign n6860 = n1564 & ~n6859 ;
  assign n6861 = n1568 & ~n6860 ;
  assign n6862 = n1572 & ~n6861 ;
  assign n6863 = n1576 & ~n6862 ;
  assign n6864 = n1580 & ~n6863 ;
  assign n6865 = n1584 & ~n6864 ;
  assign n6866 = n1588 & ~n6865 ;
  assign n6867 = n1592 & ~n6866 ;
  assign n6868 = n1596 & ~n6867 ;
  assign n6869 = n1600 & ~n6868 ;
  assign n6870 = n1604 & ~n6869 ;
  assign n6871 = n1608 & ~n6870 ;
  assign n6872 = n1612 & ~n6871 ;
  assign n6873 = n2656 & ~n6872 ;
  assign n6874 = n2658 & ~n6873 ;
  assign n6875 = n3192 & ~n6874 ;
  assign n6876 = n1962 & ~n6875 ;
  assign n6877 = n1966 & ~n6876 ;
  assign n6878 = n1970 & ~n6877 ;
  assign n6879 = n1974 & ~n6878 ;
  assign n6880 = n1978 & ~n6879 ;
  assign n6881 = n1982 & ~n6880 ;
  assign n6882 = n1986 & ~n6881 ;
  assign n6883 = n1990 & ~n6882 ;
  assign n6884 = n1994 & ~n6883 ;
  assign n6885 = n1998 & ~n6884 ;
  assign n6886 = n2002 & ~n6885 ;
  assign n6887 = n2006 & ~n6886 ;
  assign n6888 = n2010 & ~n6887 ;
  assign n6889 = n2014 & ~n6888 ;
  assign n6890 = n2018 & ~n6889 ;
  assign n6891 = ~x156 & ~n2020 ;
  assign n6892 = ~n6890 & n6891 ;
  assign n6895 = ~n6892 & ~x284 ;
  assign n6896 = ~n6894 & ~n6895 ;
  assign n6897 = ~n334 & n1692 ;
  assign n6898 = n1697 & ~n6897 ;
  assign n6899 = n1701 & ~n6898 ;
  assign n6900 = n1705 & ~n6899 ;
  assign n6901 = n1709 & ~n6900 ;
  assign n6902 = n1713 & ~n6901 ;
  assign n6903 = n1717 & ~n6902 ;
  assign n6904 = n1721 & ~n6903 ;
  assign n6905 = n1725 & ~n6904 ;
  assign n6906 = n1729 & ~n6905 ;
  assign n6907 = n1733 & ~n6906 ;
  assign n6908 = n1737 & ~n6907 ;
  assign n6909 = n1741 & ~n6908 ;
  assign n6910 = n1745 & ~n6909 ;
  assign n6911 = n1749 & ~n6910 ;
  assign n6912 = n1753 & ~n6911 ;
  assign n6913 = n1757 & ~n6912 ;
  assign n6914 = n1761 & ~n6913 ;
  assign n6915 = n1765 & ~n6914 ;
  assign n6916 = n1769 & ~n6915 ;
  assign n6917 = n1773 & ~n6916 ;
  assign n6918 = n1777 & ~n6917 ;
  assign n6919 = n1781 & ~n6918 ;
  assign n6920 = n1785 & ~n6919 ;
  assign n6921 = n1789 & ~n6920 ;
  assign n6922 = n1793 & ~n6921 ;
  assign n6923 = n1797 & ~n6922 ;
  assign n6924 = n1801 & ~n6923 ;
  assign n6925 = n1805 & ~n6924 ;
  assign n6926 = n1809 & ~n6925 ;
  assign n6927 = n1813 & ~n6926 ;
  assign n6928 = n1817 & ~n6927 ;
  assign n6929 = n1821 & ~n6928 ;
  assign n6930 = n1825 & ~n6929 ;
  assign n6931 = n1829 & ~n6930 ;
  assign n6932 = n1833 & ~n6931 ;
  assign n6933 = n1837 & ~n6932 ;
  assign n6934 = n1841 & ~n6933 ;
  assign n6935 = n1845 & ~n6934 ;
  assign n6936 = n1849 & ~n6935 ;
  assign n6937 = n1853 & ~n6936 ;
  assign n6938 = n1857 & ~n6937 ;
  assign n6939 = n1861 & ~n6938 ;
  assign n6940 = n1865 & ~n6939 ;
  assign n6941 = n1869 & ~n6940 ;
  assign n6942 = n1873 & ~n6941 ;
  assign n6943 = n1877 & ~n6942 ;
  assign n6944 = n1881 & ~n6943 ;
  assign n6945 = n1885 & ~n6944 ;
  assign n6946 = n1889 & ~n6945 ;
  assign n6947 = n1893 & ~n6946 ;
  assign n6948 = n1897 & ~n6947 ;
  assign n6949 = n1901 & ~n6948 ;
  assign n6950 = n1905 & ~n6949 ;
  assign n6951 = n1909 & ~n6950 ;
  assign n6952 = n1913 & ~n6951 ;
  assign n6953 = n1917 & ~n6952 ;
  assign n6954 = n1921 & ~n6953 ;
  assign n6955 = n1925 & ~n6954 ;
  assign n6956 = n1929 & ~n6955 ;
  assign n6957 = n1933 & ~n6956 ;
  assign n6958 = n1937 & ~n6957 ;
  assign n6959 = n1941 & ~n6958 ;
  assign n6960 = n1945 & ~n6959 ;
  assign n6961 = n1949 & ~n6960 ;
  assign n6962 = n1953 & ~n6961 ;
  assign n6963 = n2749 & ~n6962 ;
  assign n6964 = n263 & ~n6963 ;
  assign n6965 = n267 & ~n6964 ;
  assign n6966 = n271 & ~n6965 ;
  assign n6967 = n275 & ~n6966 ;
  assign n6968 = n279 & ~n6967 ;
  assign n6969 = n283 & ~n6968 ;
  assign n6970 = n287 & ~n6969 ;
  assign n6971 = n291 & ~n6970 ;
  assign n6972 = n295 & ~n6971 ;
  assign n6973 = n299 & ~n6972 ;
  assign n6974 = n303 & ~n6973 ;
  assign n6975 = n307 & ~n6974 ;
  assign n6976 = n311 & ~n6975 ;
  assign n6977 = n315 & ~n6976 ;
  assign n6978 = n319 & ~n6977 ;
  assign n6979 = n323 & ~n6978 ;
  assign n6980 = n327 & ~n6979 ;
  assign n6981 = x157 & ~n329 ;
  assign n6982 = ~n6980 & n6981 ;
  assign n7070 = n6982 & x285 ;
  assign n6983 = ~n673 & n2029 ;
  assign n6984 = n2034 & ~n6983 ;
  assign n6985 = n2038 & ~n6984 ;
  assign n6986 = n2042 & ~n6985 ;
  assign n6987 = n2046 & ~n6986 ;
  assign n6988 = n2050 & ~n6987 ;
  assign n6989 = n2054 & ~n6988 ;
  assign n6990 = n2058 & ~n6989 ;
  assign n6991 = n2062 & ~n6990 ;
  assign n6992 = n2066 & ~n6991 ;
  assign n6993 = n2070 & ~n6992 ;
  assign n6994 = n2074 & ~n6993 ;
  assign n6995 = n2078 & ~n6994 ;
  assign n6996 = n2082 & ~n6995 ;
  assign n6997 = n2086 & ~n6996 ;
  assign n6998 = n2090 & ~n6997 ;
  assign n6999 = n2094 & ~n6998 ;
  assign n7000 = n2098 & ~n6999 ;
  assign n7001 = n2102 & ~n7000 ;
  assign n7002 = n2106 & ~n7001 ;
  assign n7003 = n2110 & ~n7002 ;
  assign n7004 = n2114 & ~n7003 ;
  assign n7005 = n2118 & ~n7004 ;
  assign n7006 = n2122 & ~n7005 ;
  assign n7007 = n2126 & ~n7006 ;
  assign n7008 = n2130 & ~n7007 ;
  assign n7009 = n2134 & ~n7008 ;
  assign n7010 = n2138 & ~n7009 ;
  assign n7011 = n2142 & ~n7010 ;
  assign n7012 = n2146 & ~n7011 ;
  assign n7013 = n2150 & ~n7012 ;
  assign n7014 = n2154 & ~n7013 ;
  assign n7015 = n2158 & ~n7014 ;
  assign n7016 = n2162 & ~n7015 ;
  assign n7017 = n2166 & ~n7016 ;
  assign n7018 = n2170 & ~n7017 ;
  assign n7019 = n2174 & ~n7018 ;
  assign n7020 = n2178 & ~n7019 ;
  assign n7021 = n2182 & ~n7020 ;
  assign n7022 = n2186 & ~n7021 ;
  assign n7023 = n2190 & ~n7022 ;
  assign n7024 = n2194 & ~n7023 ;
  assign n7025 = n2198 & ~n7024 ;
  assign n7026 = n2202 & ~n7025 ;
  assign n7027 = n2206 & ~n7026 ;
  assign n7028 = n2210 & ~n7027 ;
  assign n7029 = n2214 & ~n7028 ;
  assign n7030 = n2218 & ~n7029 ;
  assign n7031 = n2222 & ~n7030 ;
  assign n7032 = n2226 & ~n7031 ;
  assign n7033 = n2230 & ~n7032 ;
  assign n7034 = n2234 & ~n7033 ;
  assign n7035 = n2238 & ~n7034 ;
  assign n7036 = n2242 & ~n7035 ;
  assign n7037 = n2246 & ~n7036 ;
  assign n7038 = n2250 & ~n7037 ;
  assign n7039 = n2254 & ~n7038 ;
  assign n7040 = n2258 & ~n7039 ;
  assign n7041 = n2262 & ~n7040 ;
  assign n7042 = n2266 & ~n7041 ;
  assign n7043 = n2270 & ~n7042 ;
  assign n7044 = n2274 & ~n7043 ;
  assign n7045 = n2278 & ~n7044 ;
  assign n7046 = n2282 & ~n7045 ;
  assign n7047 = n2286 & ~n7046 ;
  assign n7048 = n2290 & ~n7047 ;
  assign n7049 = n2836 & ~n7048 ;
  assign n7050 = n602 & ~n7049 ;
  assign n7051 = n606 & ~n7050 ;
  assign n7052 = n610 & ~n7051 ;
  assign n7053 = n614 & ~n7052 ;
  assign n7054 = n618 & ~n7053 ;
  assign n7055 = n622 & ~n7054 ;
  assign n7056 = n626 & ~n7055 ;
  assign n7057 = n630 & ~n7056 ;
  assign n7058 = n634 & ~n7057 ;
  assign n7059 = n638 & ~n7058 ;
  assign n7060 = n642 & ~n7059 ;
  assign n7061 = n646 & ~n7060 ;
  assign n7062 = n650 & ~n7061 ;
  assign n7063 = n654 & ~n7062 ;
  assign n7064 = n658 & ~n7063 ;
  assign n7065 = n662 & ~n7064 ;
  assign n7066 = n666 & ~n7065 ;
  assign n7067 = ~x157 & ~n668 ;
  assign n7068 = ~n7066 & n7067 ;
  assign n7071 = ~n7068 & ~x285 ;
  assign n7072 = ~n7070 & ~n7071 ;
  assign n7073 = n338 & ~n1016 ;
  assign n7074 = n343 & ~n7073 ;
  assign n7075 = n347 & ~n7074 ;
  assign n7076 = n351 & ~n7075 ;
  assign n7077 = n355 & ~n7076 ;
  assign n7078 = n359 & ~n7077 ;
  assign n7079 = n363 & ~n7078 ;
  assign n7080 = n367 & ~n7079 ;
  assign n7081 = n371 & ~n7080 ;
  assign n7082 = n375 & ~n7081 ;
  assign n7083 = n379 & ~n7082 ;
  assign n7084 = n383 & ~n7083 ;
  assign n7085 = n387 & ~n7084 ;
  assign n7086 = n391 & ~n7085 ;
  assign n7087 = n395 & ~n7086 ;
  assign n7088 = n399 & ~n7087 ;
  assign n7089 = n403 & ~n7088 ;
  assign n7090 = n407 & ~n7089 ;
  assign n7091 = n411 & ~n7090 ;
  assign n7092 = n415 & ~n7091 ;
  assign n7093 = n419 & ~n7092 ;
  assign n7094 = n423 & ~n7093 ;
  assign n7095 = n427 & ~n7094 ;
  assign n7096 = n431 & ~n7095 ;
  assign n7097 = n435 & ~n7096 ;
  assign n7098 = n439 & ~n7097 ;
  assign n7099 = n443 & ~n7098 ;
  assign n7100 = n447 & ~n7099 ;
  assign n7101 = n451 & ~n7100 ;
  assign n7102 = n455 & ~n7101 ;
  assign n7103 = n459 & ~n7102 ;
  assign n7104 = n463 & ~n7103 ;
  assign n7105 = n467 & ~n7104 ;
  assign n7106 = n471 & ~n7105 ;
  assign n7107 = n475 & ~n7106 ;
  assign n7108 = n479 & ~n7107 ;
  assign n7109 = n483 & ~n7108 ;
  assign n7110 = n487 & ~n7109 ;
  assign n7111 = n491 & ~n7110 ;
  assign n7112 = n495 & ~n7111 ;
  assign n7113 = n499 & ~n7112 ;
  assign n7114 = n503 & ~n7113 ;
  assign n7115 = n507 & ~n7114 ;
  assign n7116 = n511 & ~n7115 ;
  assign n7117 = n515 & ~n7116 ;
  assign n7118 = n519 & ~n7117 ;
  assign n7119 = n523 & ~n7118 ;
  assign n7120 = n527 & ~n7119 ;
  assign n7121 = n531 & ~n7120 ;
  assign n7122 = n535 & ~n7121 ;
  assign n7123 = n539 & ~n7122 ;
  assign n7124 = n543 & ~n7123 ;
  assign n7125 = n547 & ~n7124 ;
  assign n7126 = n551 & ~n7125 ;
  assign n7127 = n555 & ~n7126 ;
  assign n7128 = n559 & ~n7127 ;
  assign n7129 = n563 & ~n7128 ;
  assign n7130 = n567 & ~n7129 ;
  assign n7131 = n571 & ~n7130 ;
  assign n7132 = n575 & ~n7131 ;
  assign n7133 = n579 & ~n7132 ;
  assign n7134 = n583 & ~n7133 ;
  assign n7135 = n587 & ~n7134 ;
  assign n7136 = n591 & ~n7135 ;
  assign n7137 = n2382 & ~n7136 ;
  assign n7138 = n2384 & ~n7137 ;
  assign n7139 = n2927 & ~n7138 ;
  assign n7140 = n945 & ~n7139 ;
  assign n7141 = n949 & ~n7140 ;
  assign n7142 = n953 & ~n7141 ;
  assign n7143 = n957 & ~n7142 ;
  assign n7144 = n961 & ~n7143 ;
  assign n7145 = n965 & ~n7144 ;
  assign n7146 = n969 & ~n7145 ;
  assign n7147 = n973 & ~n7146 ;
  assign n7148 = n977 & ~n7147 ;
  assign n7149 = n981 & ~n7148 ;
  assign n7150 = n985 & ~n7149 ;
  assign n7151 = n989 & ~n7150 ;
  assign n7152 = n993 & ~n7151 ;
  assign n7153 = n997 & ~n7152 ;
  assign n7154 = n1001 & ~n7153 ;
  assign n7155 = n1005 & ~n7154 ;
  assign n7156 = n1009 & ~n7155 ;
  assign n7157 = x158 & ~n1011 ;
  assign n7158 = ~n7156 & n7157 ;
  assign n7246 = n7158 & x286 ;
  assign n7159 = n677 & ~n1355 ;
  assign n7160 = n682 & ~n7159 ;
  assign n7161 = n686 & ~n7160 ;
  assign n7162 = n690 & ~n7161 ;
  assign n7163 = n694 & ~n7162 ;
  assign n7164 = n698 & ~n7163 ;
  assign n7165 = n702 & ~n7164 ;
  assign n7166 = n706 & ~n7165 ;
  assign n7167 = n710 & ~n7166 ;
  assign n7168 = n714 & ~n7167 ;
  assign n7169 = n718 & ~n7168 ;
  assign n7170 = n722 & ~n7169 ;
  assign n7171 = n726 & ~n7170 ;
  assign n7172 = n730 & ~n7171 ;
  assign n7173 = n734 & ~n7172 ;
  assign n7174 = n738 & ~n7173 ;
  assign n7175 = n742 & ~n7174 ;
  assign n7176 = n746 & ~n7175 ;
  assign n7177 = n750 & ~n7176 ;
  assign n7178 = n754 & ~n7177 ;
  assign n7179 = n758 & ~n7178 ;
  assign n7180 = n762 & ~n7179 ;
  assign n7181 = n766 & ~n7180 ;
  assign n7182 = n770 & ~n7181 ;
  assign n7183 = n774 & ~n7182 ;
  assign n7184 = n778 & ~n7183 ;
  assign n7185 = n782 & ~n7184 ;
  assign n7186 = n786 & ~n7185 ;
  assign n7187 = n790 & ~n7186 ;
  assign n7188 = n794 & ~n7187 ;
  assign n7189 = n798 & ~n7188 ;
  assign n7190 = n802 & ~n7189 ;
  assign n7191 = n806 & ~n7190 ;
  assign n7192 = n810 & ~n7191 ;
  assign n7193 = n814 & ~n7192 ;
  assign n7194 = n818 & ~n7193 ;
  assign n7195 = n822 & ~n7194 ;
  assign n7196 = n826 & ~n7195 ;
  assign n7197 = n830 & ~n7196 ;
  assign n7198 = n834 & ~n7197 ;
  assign n7199 = n838 & ~n7198 ;
  assign n7200 = n842 & ~n7199 ;
  assign n7201 = n846 & ~n7200 ;
  assign n7202 = n850 & ~n7201 ;
  assign n7203 = n854 & ~n7202 ;
  assign n7204 = n858 & ~n7203 ;
  assign n7205 = n862 & ~n7204 ;
  assign n7206 = n866 & ~n7205 ;
  assign n7207 = n870 & ~n7206 ;
  assign n7208 = n874 & ~n7207 ;
  assign n7209 = n878 & ~n7208 ;
  assign n7210 = n882 & ~n7209 ;
  assign n7211 = n886 & ~n7210 ;
  assign n7212 = n890 & ~n7211 ;
  assign n7213 = n894 & ~n7212 ;
  assign n7214 = n898 & ~n7213 ;
  assign n7215 = n902 & ~n7214 ;
  assign n7216 = n906 & ~n7215 ;
  assign n7217 = n910 & ~n7216 ;
  assign n7218 = n914 & ~n7217 ;
  assign n7219 = n918 & ~n7218 ;
  assign n7220 = n922 & ~n7219 ;
  assign n7221 = n926 & ~n7220 ;
  assign n7222 = n930 & ~n7221 ;
  assign n7223 = n2472 & ~n7222 ;
  assign n7224 = n2474 & ~n7223 ;
  assign n7225 = n3014 & ~n7224 ;
  assign n7226 = n1284 & ~n7225 ;
  assign n7227 = n1288 & ~n7226 ;
  assign n7228 = n1292 & ~n7227 ;
  assign n7229 = n1296 & ~n7228 ;
  assign n7230 = n1300 & ~n7229 ;
  assign n7231 = n1304 & ~n7230 ;
  assign n7232 = n1308 & ~n7231 ;
  assign n7233 = n1312 & ~n7232 ;
  assign n7234 = n1316 & ~n7233 ;
  assign n7235 = n1320 & ~n7234 ;
  assign n7236 = n1324 & ~n7235 ;
  assign n7237 = n1328 & ~n7236 ;
  assign n7238 = n1332 & ~n7237 ;
  assign n7239 = n1336 & ~n7238 ;
  assign n7240 = n1340 & ~n7239 ;
  assign n7241 = n1344 & ~n7240 ;
  assign n7242 = n1348 & ~n7241 ;
  assign n7243 = ~x158 & ~n1350 ;
  assign n7244 = ~n7242 & n7243 ;
  assign n7247 = ~n7244 & ~x286 ;
  assign n7248 = ~n7246 & ~n7247 ;
  assign n7249 = n1020 & ~n1696 ;
  assign n7250 = n1025 & ~n7249 ;
  assign n7251 = n1029 & ~n7250 ;
  assign n7252 = n1033 & ~n7251 ;
  assign n7253 = n1037 & ~n7252 ;
  assign n7254 = n1041 & ~n7253 ;
  assign n7255 = n1045 & ~n7254 ;
  assign n7256 = n1049 & ~n7255 ;
  assign n7257 = n1053 & ~n7256 ;
  assign n7258 = n1057 & ~n7257 ;
  assign n7259 = n1061 & ~n7258 ;
  assign n7260 = n1065 & ~n7259 ;
  assign n7261 = n1069 & ~n7260 ;
  assign n7262 = n1073 & ~n7261 ;
  assign n7263 = n1077 & ~n7262 ;
  assign n7264 = n1081 & ~n7263 ;
  assign n7265 = n1085 & ~n7264 ;
  assign n7266 = n1089 & ~n7265 ;
  assign n7267 = n1093 & ~n7266 ;
  assign n7268 = n1097 & ~n7267 ;
  assign n7269 = n1101 & ~n7268 ;
  assign n7270 = n1105 & ~n7269 ;
  assign n7271 = n1109 & ~n7270 ;
  assign n7272 = n1113 & ~n7271 ;
  assign n7273 = n1117 & ~n7272 ;
  assign n7274 = n1121 & ~n7273 ;
  assign n7275 = n1125 & ~n7274 ;
  assign n7276 = n1129 & ~n7275 ;
  assign n7277 = n1133 & ~n7276 ;
  assign n7278 = n1137 & ~n7277 ;
  assign n7279 = n1141 & ~n7278 ;
  assign n7280 = n1145 & ~n7279 ;
  assign n7281 = n1149 & ~n7280 ;
  assign n7282 = n1153 & ~n7281 ;
  assign n7283 = n1157 & ~n7282 ;
  assign n7284 = n1161 & ~n7283 ;
  assign n7285 = n1165 & ~n7284 ;
  assign n7286 = n1169 & ~n7285 ;
  assign n7287 = n1173 & ~n7286 ;
  assign n7288 = n1177 & ~n7287 ;
  assign n7289 = n1181 & ~n7288 ;
  assign n7290 = n1185 & ~n7289 ;
  assign n7291 = n1189 & ~n7290 ;
  assign n7292 = n1193 & ~n7291 ;
  assign n7293 = n1197 & ~n7292 ;
  assign n7294 = n1201 & ~n7293 ;
  assign n7295 = n1205 & ~n7294 ;
  assign n7296 = n1209 & ~n7295 ;
  assign n7297 = n1213 & ~n7296 ;
  assign n7298 = n1217 & ~n7297 ;
  assign n7299 = n1221 & ~n7298 ;
  assign n7300 = n1225 & ~n7299 ;
  assign n7301 = n1229 & ~n7300 ;
  assign n7302 = n1233 & ~n7301 ;
  assign n7303 = n1237 & ~n7302 ;
  assign n7304 = n1241 & ~n7303 ;
  assign n7305 = n1245 & ~n7304 ;
  assign n7306 = n1249 & ~n7305 ;
  assign n7307 = n1253 & ~n7306 ;
  assign n7308 = n1257 & ~n7307 ;
  assign n7309 = n1261 & ~n7308 ;
  assign n7310 = n1265 & ~n7309 ;
  assign n7311 = n1269 & ~n7310 ;
  assign n7312 = n1273 & ~n7311 ;
  assign n7313 = n2566 & ~n7312 ;
  assign n7314 = n2568 & ~n7313 ;
  assign n7315 = n3105 & ~n7314 ;
  assign n7316 = n1625 & ~n7315 ;
  assign n7317 = n1629 & ~n7316 ;
  assign n7318 = n1633 & ~n7317 ;
  assign n7319 = n1637 & ~n7318 ;
  assign n7320 = n1641 & ~n7319 ;
  assign n7321 = n1645 & ~n7320 ;
  assign n7322 = n1649 & ~n7321 ;
  assign n7323 = n1653 & ~n7322 ;
  assign n7324 = n1657 & ~n7323 ;
  assign n7325 = n1661 & ~n7324 ;
  assign n7326 = n1665 & ~n7325 ;
  assign n7327 = n1669 & ~n7326 ;
  assign n7328 = n1673 & ~n7327 ;
  assign n7329 = n1677 & ~n7328 ;
  assign n7330 = n1681 & ~n7329 ;
  assign n7331 = n1685 & ~n7330 ;
  assign n7332 = n1689 & ~n7331 ;
  assign n7333 = x159 & ~n1691 ;
  assign n7334 = ~n7332 & n7333 ;
  assign n7422 = n7334 & x287 ;
  assign n7335 = n1359 & ~n2033 ;
  assign n7336 = n1364 & ~n7335 ;
  assign n7337 = n1368 & ~n7336 ;
  assign n7338 = n1372 & ~n7337 ;
  assign n7339 = n1376 & ~n7338 ;
  assign n7340 = n1380 & ~n7339 ;
  assign n7341 = n1384 & ~n7340 ;
  assign n7342 = n1388 & ~n7341 ;
  assign n7343 = n1392 & ~n7342 ;
  assign n7344 = n1396 & ~n7343 ;
  assign n7345 = n1400 & ~n7344 ;
  assign n7346 = n1404 & ~n7345 ;
  assign n7347 = n1408 & ~n7346 ;
  assign n7348 = n1412 & ~n7347 ;
  assign n7349 = n1416 & ~n7348 ;
  assign n7350 = n1420 & ~n7349 ;
  assign n7351 = n1424 & ~n7350 ;
  assign n7352 = n1428 & ~n7351 ;
  assign n7353 = n1432 & ~n7352 ;
  assign n7354 = n1436 & ~n7353 ;
  assign n7355 = n1440 & ~n7354 ;
  assign n7356 = n1444 & ~n7355 ;
  assign n7357 = n1448 & ~n7356 ;
  assign n7358 = n1452 & ~n7357 ;
  assign n7359 = n1456 & ~n7358 ;
  assign n7360 = n1460 & ~n7359 ;
  assign n7361 = n1464 & ~n7360 ;
  assign n7362 = n1468 & ~n7361 ;
  assign n7363 = n1472 & ~n7362 ;
  assign n7364 = n1476 & ~n7363 ;
  assign n7365 = n1480 & ~n7364 ;
  assign n7366 = n1484 & ~n7365 ;
  assign n7367 = n1488 & ~n7366 ;
  assign n7368 = n1492 & ~n7367 ;
  assign n7369 = n1496 & ~n7368 ;
  assign n7370 = n1500 & ~n7369 ;
  assign n7371 = n1504 & ~n7370 ;
  assign n7372 = n1508 & ~n7371 ;
  assign n7373 = n1512 & ~n7372 ;
  assign n7374 = n1516 & ~n7373 ;
  assign n7375 = n1520 & ~n7374 ;
  assign n7376 = n1524 & ~n7375 ;
  assign n7377 = n1528 & ~n7376 ;
  assign n7378 = n1532 & ~n7377 ;
  assign n7379 = n1536 & ~n7378 ;
  assign n7380 = n1540 & ~n7379 ;
  assign n7381 = n1544 & ~n7380 ;
  assign n7382 = n1548 & ~n7381 ;
  assign n7383 = n1552 & ~n7382 ;
  assign n7384 = n1556 & ~n7383 ;
  assign n7385 = n1560 & ~n7384 ;
  assign n7386 = n1564 & ~n7385 ;
  assign n7387 = n1568 & ~n7386 ;
  assign n7388 = n1572 & ~n7387 ;
  assign n7389 = n1576 & ~n7388 ;
  assign n7390 = n1580 & ~n7389 ;
  assign n7391 = n1584 & ~n7390 ;
  assign n7392 = n1588 & ~n7391 ;
  assign n7393 = n1592 & ~n7392 ;
  assign n7394 = n1596 & ~n7393 ;
  assign n7395 = n1600 & ~n7394 ;
  assign n7396 = n1604 & ~n7395 ;
  assign n7397 = n1608 & ~n7396 ;
  assign n7398 = n1612 & ~n7397 ;
  assign n7399 = n2656 & ~n7398 ;
  assign n7400 = n2658 & ~n7399 ;
  assign n7401 = n3192 & ~n7400 ;
  assign n7402 = n1962 & ~n7401 ;
  assign n7403 = n1966 & ~n7402 ;
  assign n7404 = n1970 & ~n7403 ;
  assign n7405 = n1974 & ~n7404 ;
  assign n7406 = n1978 & ~n7405 ;
  assign n7407 = n1982 & ~n7406 ;
  assign n7408 = n1986 & ~n7407 ;
  assign n7409 = n1990 & ~n7408 ;
  assign n7410 = n1994 & ~n7409 ;
  assign n7411 = n1998 & ~n7410 ;
  assign n7412 = n2002 & ~n7411 ;
  assign n7413 = n2006 & ~n7412 ;
  assign n7414 = n2010 & ~n7413 ;
  assign n7415 = n2014 & ~n7414 ;
  assign n7416 = n2018 & ~n7415 ;
  assign n7417 = n2022 & ~n7416 ;
  assign n7418 = n2026 & ~n7417 ;
  assign n7419 = ~x159 & ~n2028 ;
  assign n7420 = ~n7418 & n7419 ;
  assign n7423 = ~n7420 & ~x287 ;
  assign n7424 = ~n7422 & ~n7423 ;
  assign n7425 = ~n342 & n1700 ;
  assign n7426 = n1705 & ~n7425 ;
  assign n7427 = n1709 & ~n7426 ;
  assign n7428 = n1713 & ~n7427 ;
  assign n7429 = n1717 & ~n7428 ;
  assign n7430 = n1721 & ~n7429 ;
  assign n7431 = n1725 & ~n7430 ;
  assign n7432 = n1729 & ~n7431 ;
  assign n7433 = n1733 & ~n7432 ;
  assign n7434 = n1737 & ~n7433 ;
  assign n7435 = n1741 & ~n7434 ;
  assign n7436 = n1745 & ~n7435 ;
  assign n7437 = n1749 & ~n7436 ;
  assign n7438 = n1753 & ~n7437 ;
  assign n7439 = n1757 & ~n7438 ;
  assign n7440 = n1761 & ~n7439 ;
  assign n7441 = n1765 & ~n7440 ;
  assign n7442 = n1769 & ~n7441 ;
  assign n7443 = n1773 & ~n7442 ;
  assign n7444 = n1777 & ~n7443 ;
  assign n7445 = n1781 & ~n7444 ;
  assign n7446 = n1785 & ~n7445 ;
  assign n7447 = n1789 & ~n7446 ;
  assign n7448 = n1793 & ~n7447 ;
  assign n7449 = n1797 & ~n7448 ;
  assign n7450 = n1801 & ~n7449 ;
  assign n7451 = n1805 & ~n7450 ;
  assign n7452 = n1809 & ~n7451 ;
  assign n7453 = n1813 & ~n7452 ;
  assign n7454 = n1817 & ~n7453 ;
  assign n7455 = n1821 & ~n7454 ;
  assign n7456 = n1825 & ~n7455 ;
  assign n7457 = n1829 & ~n7456 ;
  assign n7458 = n1833 & ~n7457 ;
  assign n7459 = n1837 & ~n7458 ;
  assign n7460 = n1841 & ~n7459 ;
  assign n7461 = n1845 & ~n7460 ;
  assign n7462 = n1849 & ~n7461 ;
  assign n7463 = n1853 & ~n7462 ;
  assign n7464 = n1857 & ~n7463 ;
  assign n7465 = n1861 & ~n7464 ;
  assign n7466 = n1865 & ~n7465 ;
  assign n7467 = n1869 & ~n7466 ;
  assign n7468 = n1873 & ~n7467 ;
  assign n7469 = n1877 & ~n7468 ;
  assign n7470 = n1881 & ~n7469 ;
  assign n7471 = n1885 & ~n7470 ;
  assign n7472 = n1889 & ~n7471 ;
  assign n7473 = n1893 & ~n7472 ;
  assign n7474 = n1897 & ~n7473 ;
  assign n7475 = n1901 & ~n7474 ;
  assign n7476 = n1905 & ~n7475 ;
  assign n7477 = n1909 & ~n7476 ;
  assign n7478 = n1913 & ~n7477 ;
  assign n7479 = n1917 & ~n7478 ;
  assign n7480 = n1921 & ~n7479 ;
  assign n7481 = n1925 & ~n7480 ;
  assign n7482 = n1929 & ~n7481 ;
  assign n7483 = n1933 & ~n7482 ;
  assign n7484 = n1937 & ~n7483 ;
  assign n7485 = n1941 & ~n7484 ;
  assign n7486 = n1945 & ~n7485 ;
  assign n7487 = n1949 & ~n7486 ;
  assign n7488 = n1953 & ~n7487 ;
  assign n7489 = n2749 & ~n7488 ;
  assign n7490 = n263 & ~n7489 ;
  assign n7491 = n267 & ~n7490 ;
  assign n7492 = n271 & ~n7491 ;
  assign n7493 = n275 & ~n7492 ;
  assign n7494 = n279 & ~n7493 ;
  assign n7495 = n283 & ~n7494 ;
  assign n7496 = n287 & ~n7495 ;
  assign n7497 = n291 & ~n7496 ;
  assign n7498 = n295 & ~n7497 ;
  assign n7499 = n299 & ~n7498 ;
  assign n7500 = n303 & ~n7499 ;
  assign n7501 = n307 & ~n7500 ;
  assign n7502 = n311 & ~n7501 ;
  assign n7503 = n315 & ~n7502 ;
  assign n7504 = n319 & ~n7503 ;
  assign n7505 = n323 & ~n7504 ;
  assign n7506 = n327 & ~n7505 ;
  assign n7507 = n331 & ~n7506 ;
  assign n7508 = n335 & ~n7507 ;
  assign n7509 = x160 & ~n337 ;
  assign n7510 = ~n7508 & n7509 ;
  assign n7598 = n7510 & x288 ;
  assign n7511 = ~n681 & n2037 ;
  assign n7512 = n2042 & ~n7511 ;
  assign n7513 = n2046 & ~n7512 ;
  assign n7514 = n2050 & ~n7513 ;
  assign n7515 = n2054 & ~n7514 ;
  assign n7516 = n2058 & ~n7515 ;
  assign n7517 = n2062 & ~n7516 ;
  assign n7518 = n2066 & ~n7517 ;
  assign n7519 = n2070 & ~n7518 ;
  assign n7520 = n2074 & ~n7519 ;
  assign n7521 = n2078 & ~n7520 ;
  assign n7522 = n2082 & ~n7521 ;
  assign n7523 = n2086 & ~n7522 ;
  assign n7524 = n2090 & ~n7523 ;
  assign n7525 = n2094 & ~n7524 ;
  assign n7526 = n2098 & ~n7525 ;
  assign n7527 = n2102 & ~n7526 ;
  assign n7528 = n2106 & ~n7527 ;
  assign n7529 = n2110 & ~n7528 ;
  assign n7530 = n2114 & ~n7529 ;
  assign n7531 = n2118 & ~n7530 ;
  assign n7532 = n2122 & ~n7531 ;
  assign n7533 = n2126 & ~n7532 ;
  assign n7534 = n2130 & ~n7533 ;
  assign n7535 = n2134 & ~n7534 ;
  assign n7536 = n2138 & ~n7535 ;
  assign n7537 = n2142 & ~n7536 ;
  assign n7538 = n2146 & ~n7537 ;
  assign n7539 = n2150 & ~n7538 ;
  assign n7540 = n2154 & ~n7539 ;
  assign n7541 = n2158 & ~n7540 ;
  assign n7542 = n2162 & ~n7541 ;
  assign n7543 = n2166 & ~n7542 ;
  assign n7544 = n2170 & ~n7543 ;
  assign n7545 = n2174 & ~n7544 ;
  assign n7546 = n2178 & ~n7545 ;
  assign n7547 = n2182 & ~n7546 ;
  assign n7548 = n2186 & ~n7547 ;
  assign n7549 = n2190 & ~n7548 ;
  assign n7550 = n2194 & ~n7549 ;
  assign n7551 = n2198 & ~n7550 ;
  assign n7552 = n2202 & ~n7551 ;
  assign n7553 = n2206 & ~n7552 ;
  assign n7554 = n2210 & ~n7553 ;
  assign n7555 = n2214 & ~n7554 ;
  assign n7556 = n2218 & ~n7555 ;
  assign n7557 = n2222 & ~n7556 ;
  assign n7558 = n2226 & ~n7557 ;
  assign n7559 = n2230 & ~n7558 ;
  assign n7560 = n2234 & ~n7559 ;
  assign n7561 = n2238 & ~n7560 ;
  assign n7562 = n2242 & ~n7561 ;
  assign n7563 = n2246 & ~n7562 ;
  assign n7564 = n2250 & ~n7563 ;
  assign n7565 = n2254 & ~n7564 ;
  assign n7566 = n2258 & ~n7565 ;
  assign n7567 = n2262 & ~n7566 ;
  assign n7568 = n2266 & ~n7567 ;
  assign n7569 = n2270 & ~n7568 ;
  assign n7570 = n2274 & ~n7569 ;
  assign n7571 = n2278 & ~n7570 ;
  assign n7572 = n2282 & ~n7571 ;
  assign n7573 = n2286 & ~n7572 ;
  assign n7574 = n2290 & ~n7573 ;
  assign n7575 = n2836 & ~n7574 ;
  assign n7576 = n602 & ~n7575 ;
  assign n7577 = n606 & ~n7576 ;
  assign n7578 = n610 & ~n7577 ;
  assign n7579 = n614 & ~n7578 ;
  assign n7580 = n618 & ~n7579 ;
  assign n7581 = n622 & ~n7580 ;
  assign n7582 = n626 & ~n7581 ;
  assign n7583 = n630 & ~n7582 ;
  assign n7584 = n634 & ~n7583 ;
  assign n7585 = n638 & ~n7584 ;
  assign n7586 = n642 & ~n7585 ;
  assign n7587 = n646 & ~n7586 ;
  assign n7588 = n650 & ~n7587 ;
  assign n7589 = n654 & ~n7588 ;
  assign n7590 = n658 & ~n7589 ;
  assign n7591 = n662 & ~n7590 ;
  assign n7592 = n666 & ~n7591 ;
  assign n7593 = n670 & ~n7592 ;
  assign n7594 = n674 & ~n7593 ;
  assign n7595 = ~x160 & ~n676 ;
  assign n7596 = ~n7594 & n7595 ;
  assign n7599 = ~n7596 & ~x288 ;
  assign n7600 = ~n7598 & ~n7599 ;
  assign n7601 = n346 & ~n1024 ;
  assign n7602 = n351 & ~n7601 ;
  assign n7603 = n355 & ~n7602 ;
  assign n7604 = n359 & ~n7603 ;
  assign n7605 = n363 & ~n7604 ;
  assign n7606 = n367 & ~n7605 ;
  assign n7607 = n371 & ~n7606 ;
  assign n7608 = n375 & ~n7607 ;
  assign n7609 = n379 & ~n7608 ;
  assign n7610 = n383 & ~n7609 ;
  assign n7611 = n387 & ~n7610 ;
  assign n7612 = n391 & ~n7611 ;
  assign n7613 = n395 & ~n7612 ;
  assign n7614 = n399 & ~n7613 ;
  assign n7615 = n403 & ~n7614 ;
  assign n7616 = n407 & ~n7615 ;
  assign n7617 = n411 & ~n7616 ;
  assign n7618 = n415 & ~n7617 ;
  assign n7619 = n419 & ~n7618 ;
  assign n7620 = n423 & ~n7619 ;
  assign n7621 = n427 & ~n7620 ;
  assign n7622 = n431 & ~n7621 ;
  assign n7623 = n435 & ~n7622 ;
  assign n7624 = n439 & ~n7623 ;
  assign n7625 = n443 & ~n7624 ;
  assign n7626 = n447 & ~n7625 ;
  assign n7627 = n451 & ~n7626 ;
  assign n7628 = n455 & ~n7627 ;
  assign n7629 = n459 & ~n7628 ;
  assign n7630 = n463 & ~n7629 ;
  assign n7631 = n467 & ~n7630 ;
  assign n7632 = n471 & ~n7631 ;
  assign n7633 = n475 & ~n7632 ;
  assign n7634 = n479 & ~n7633 ;
  assign n7635 = n483 & ~n7634 ;
  assign n7636 = n487 & ~n7635 ;
  assign n7637 = n491 & ~n7636 ;
  assign n7638 = n495 & ~n7637 ;
  assign n7639 = n499 & ~n7638 ;
  assign n7640 = n503 & ~n7639 ;
  assign n7641 = n507 & ~n7640 ;
  assign n7642 = n511 & ~n7641 ;
  assign n7643 = n515 & ~n7642 ;
  assign n7644 = n519 & ~n7643 ;
  assign n7645 = n523 & ~n7644 ;
  assign n7646 = n527 & ~n7645 ;
  assign n7647 = n531 & ~n7646 ;
  assign n7648 = n535 & ~n7647 ;
  assign n7649 = n539 & ~n7648 ;
  assign n7650 = n543 & ~n7649 ;
  assign n7651 = n547 & ~n7650 ;
  assign n7652 = n551 & ~n7651 ;
  assign n7653 = n555 & ~n7652 ;
  assign n7654 = n559 & ~n7653 ;
  assign n7655 = n563 & ~n7654 ;
  assign n7656 = n567 & ~n7655 ;
  assign n7657 = n571 & ~n7656 ;
  assign n7658 = n575 & ~n7657 ;
  assign n7659 = n579 & ~n7658 ;
  assign n7660 = n583 & ~n7659 ;
  assign n7661 = n587 & ~n7660 ;
  assign n7662 = n591 & ~n7661 ;
  assign n7663 = n2382 & ~n7662 ;
  assign n7664 = n2384 & ~n7663 ;
  assign n7665 = n2927 & ~n7664 ;
  assign n7666 = n945 & ~n7665 ;
  assign n7667 = n949 & ~n7666 ;
  assign n7668 = n953 & ~n7667 ;
  assign n7669 = n957 & ~n7668 ;
  assign n7670 = n961 & ~n7669 ;
  assign n7671 = n965 & ~n7670 ;
  assign n7672 = n969 & ~n7671 ;
  assign n7673 = n973 & ~n7672 ;
  assign n7674 = n977 & ~n7673 ;
  assign n7675 = n981 & ~n7674 ;
  assign n7676 = n985 & ~n7675 ;
  assign n7677 = n989 & ~n7676 ;
  assign n7678 = n993 & ~n7677 ;
  assign n7679 = n997 & ~n7678 ;
  assign n7680 = n1001 & ~n7679 ;
  assign n7681 = n1005 & ~n7680 ;
  assign n7682 = n1009 & ~n7681 ;
  assign n7683 = n1013 & ~n7682 ;
  assign n7684 = n1017 & ~n7683 ;
  assign n7685 = x161 & ~n1019 ;
  assign n7686 = ~n7684 & n7685 ;
  assign n7774 = n7686 & x289 ;
  assign n7687 = n685 & ~n1363 ;
  assign n7688 = n690 & ~n7687 ;
  assign n7689 = n694 & ~n7688 ;
  assign n7690 = n698 & ~n7689 ;
  assign n7691 = n702 & ~n7690 ;
  assign n7692 = n706 & ~n7691 ;
  assign n7693 = n710 & ~n7692 ;
  assign n7694 = n714 & ~n7693 ;
  assign n7695 = n718 & ~n7694 ;
  assign n7696 = n722 & ~n7695 ;
  assign n7697 = n726 & ~n7696 ;
  assign n7698 = n730 & ~n7697 ;
  assign n7699 = n734 & ~n7698 ;
  assign n7700 = n738 & ~n7699 ;
  assign n7701 = n742 & ~n7700 ;
  assign n7702 = n746 & ~n7701 ;
  assign n7703 = n750 & ~n7702 ;
  assign n7704 = n754 & ~n7703 ;
  assign n7705 = n758 & ~n7704 ;
  assign n7706 = n762 & ~n7705 ;
  assign n7707 = n766 & ~n7706 ;
  assign n7708 = n770 & ~n7707 ;
  assign n7709 = n774 & ~n7708 ;
  assign n7710 = n778 & ~n7709 ;
  assign n7711 = n782 & ~n7710 ;
  assign n7712 = n786 & ~n7711 ;
  assign n7713 = n790 & ~n7712 ;
  assign n7714 = n794 & ~n7713 ;
  assign n7715 = n798 & ~n7714 ;
  assign n7716 = n802 & ~n7715 ;
  assign n7717 = n806 & ~n7716 ;
  assign n7718 = n810 & ~n7717 ;
  assign n7719 = n814 & ~n7718 ;
  assign n7720 = n818 & ~n7719 ;
  assign n7721 = n822 & ~n7720 ;
  assign n7722 = n826 & ~n7721 ;
  assign n7723 = n830 & ~n7722 ;
  assign n7724 = n834 & ~n7723 ;
  assign n7725 = n838 & ~n7724 ;
  assign n7726 = n842 & ~n7725 ;
  assign n7727 = n846 & ~n7726 ;
  assign n7728 = n850 & ~n7727 ;
  assign n7729 = n854 & ~n7728 ;
  assign n7730 = n858 & ~n7729 ;
  assign n7731 = n862 & ~n7730 ;
  assign n7732 = n866 & ~n7731 ;
  assign n7733 = n870 & ~n7732 ;
  assign n7734 = n874 & ~n7733 ;
  assign n7735 = n878 & ~n7734 ;
  assign n7736 = n882 & ~n7735 ;
  assign n7737 = n886 & ~n7736 ;
  assign n7738 = n890 & ~n7737 ;
  assign n7739 = n894 & ~n7738 ;
  assign n7740 = n898 & ~n7739 ;
  assign n7741 = n902 & ~n7740 ;
  assign n7742 = n906 & ~n7741 ;
  assign n7743 = n910 & ~n7742 ;
  assign n7744 = n914 & ~n7743 ;
  assign n7745 = n918 & ~n7744 ;
  assign n7746 = n922 & ~n7745 ;
  assign n7747 = n926 & ~n7746 ;
  assign n7748 = n930 & ~n7747 ;
  assign n7749 = n2472 & ~n7748 ;
  assign n7750 = n2474 & ~n7749 ;
  assign n7751 = n3014 & ~n7750 ;
  assign n7752 = n1284 & ~n7751 ;
  assign n7753 = n1288 & ~n7752 ;
  assign n7754 = n1292 & ~n7753 ;
  assign n7755 = n1296 & ~n7754 ;
  assign n7756 = n1300 & ~n7755 ;
  assign n7757 = n1304 & ~n7756 ;
  assign n7758 = n1308 & ~n7757 ;
  assign n7759 = n1312 & ~n7758 ;
  assign n7760 = n1316 & ~n7759 ;
  assign n7761 = n1320 & ~n7760 ;
  assign n7762 = n1324 & ~n7761 ;
  assign n7763 = n1328 & ~n7762 ;
  assign n7764 = n1332 & ~n7763 ;
  assign n7765 = n1336 & ~n7764 ;
  assign n7766 = n1340 & ~n7765 ;
  assign n7767 = n1344 & ~n7766 ;
  assign n7768 = n1348 & ~n7767 ;
  assign n7769 = n1352 & ~n7768 ;
  assign n7770 = n1356 & ~n7769 ;
  assign n7771 = ~x161 & ~n1358 ;
  assign n7772 = ~n7770 & n7771 ;
  assign n7775 = ~n7772 & ~x289 ;
  assign n7776 = ~n7774 & ~n7775 ;
  assign n7777 = n1028 & ~n1704 ;
  assign n7778 = n1033 & ~n7777 ;
  assign n7779 = n1037 & ~n7778 ;
  assign n7780 = n1041 & ~n7779 ;
  assign n7781 = n1045 & ~n7780 ;
  assign n7782 = n1049 & ~n7781 ;
  assign n7783 = n1053 & ~n7782 ;
  assign n7784 = n1057 & ~n7783 ;
  assign n7785 = n1061 & ~n7784 ;
  assign n7786 = n1065 & ~n7785 ;
  assign n7787 = n1069 & ~n7786 ;
  assign n7788 = n1073 & ~n7787 ;
  assign n7789 = n1077 & ~n7788 ;
  assign n7790 = n1081 & ~n7789 ;
  assign n7791 = n1085 & ~n7790 ;
  assign n7792 = n1089 & ~n7791 ;
  assign n7793 = n1093 & ~n7792 ;
  assign n7794 = n1097 & ~n7793 ;
  assign n7795 = n1101 & ~n7794 ;
  assign n7796 = n1105 & ~n7795 ;
  assign n7797 = n1109 & ~n7796 ;
  assign n7798 = n1113 & ~n7797 ;
  assign n7799 = n1117 & ~n7798 ;
  assign n7800 = n1121 & ~n7799 ;
  assign n7801 = n1125 & ~n7800 ;
  assign n7802 = n1129 & ~n7801 ;
  assign n7803 = n1133 & ~n7802 ;
  assign n7804 = n1137 & ~n7803 ;
  assign n7805 = n1141 & ~n7804 ;
  assign n7806 = n1145 & ~n7805 ;
  assign n7807 = n1149 & ~n7806 ;
  assign n7808 = n1153 & ~n7807 ;
  assign n7809 = n1157 & ~n7808 ;
  assign n7810 = n1161 & ~n7809 ;
  assign n7811 = n1165 & ~n7810 ;
  assign n7812 = n1169 & ~n7811 ;
  assign n7813 = n1173 & ~n7812 ;
  assign n7814 = n1177 & ~n7813 ;
  assign n7815 = n1181 & ~n7814 ;
  assign n7816 = n1185 & ~n7815 ;
  assign n7817 = n1189 & ~n7816 ;
  assign n7818 = n1193 & ~n7817 ;
  assign n7819 = n1197 & ~n7818 ;
  assign n7820 = n1201 & ~n7819 ;
  assign n7821 = n1205 & ~n7820 ;
  assign n7822 = n1209 & ~n7821 ;
  assign n7823 = n1213 & ~n7822 ;
  assign n7824 = n1217 & ~n7823 ;
  assign n7825 = n1221 & ~n7824 ;
  assign n7826 = n1225 & ~n7825 ;
  assign n7827 = n1229 & ~n7826 ;
  assign n7828 = n1233 & ~n7827 ;
  assign n7829 = n1237 & ~n7828 ;
  assign n7830 = n1241 & ~n7829 ;
  assign n7831 = n1245 & ~n7830 ;
  assign n7832 = n1249 & ~n7831 ;
  assign n7833 = n1253 & ~n7832 ;
  assign n7834 = n1257 & ~n7833 ;
  assign n7835 = n1261 & ~n7834 ;
  assign n7836 = n1265 & ~n7835 ;
  assign n7837 = n1269 & ~n7836 ;
  assign n7838 = n1273 & ~n7837 ;
  assign n7839 = n2566 & ~n7838 ;
  assign n7840 = n2568 & ~n7839 ;
  assign n7841 = n3105 & ~n7840 ;
  assign n7842 = n1625 & ~n7841 ;
  assign n7843 = n1629 & ~n7842 ;
  assign n7844 = n1633 & ~n7843 ;
  assign n7845 = n1637 & ~n7844 ;
  assign n7846 = n1641 & ~n7845 ;
  assign n7847 = n1645 & ~n7846 ;
  assign n7848 = n1649 & ~n7847 ;
  assign n7849 = n1653 & ~n7848 ;
  assign n7850 = n1657 & ~n7849 ;
  assign n7851 = n1661 & ~n7850 ;
  assign n7852 = n1665 & ~n7851 ;
  assign n7853 = n1669 & ~n7852 ;
  assign n7854 = n1673 & ~n7853 ;
  assign n7855 = n1677 & ~n7854 ;
  assign n7856 = n1681 & ~n7855 ;
  assign n7857 = n1685 & ~n7856 ;
  assign n7858 = n1689 & ~n7857 ;
  assign n7859 = n1693 & ~n7858 ;
  assign n7860 = n1697 & ~n7859 ;
  assign n7861 = x162 & ~n1699 ;
  assign n7862 = ~n7860 & n7861 ;
  assign n7950 = n7862 & x290 ;
  assign n7863 = n1367 & ~n2041 ;
  assign n7864 = n1372 & ~n7863 ;
  assign n7865 = n1376 & ~n7864 ;
  assign n7866 = n1380 & ~n7865 ;
  assign n7867 = n1384 & ~n7866 ;
  assign n7868 = n1388 & ~n7867 ;
  assign n7869 = n1392 & ~n7868 ;
  assign n7870 = n1396 & ~n7869 ;
  assign n7871 = n1400 & ~n7870 ;
  assign n7872 = n1404 & ~n7871 ;
  assign n7873 = n1408 & ~n7872 ;
  assign n7874 = n1412 & ~n7873 ;
  assign n7875 = n1416 & ~n7874 ;
  assign n7876 = n1420 & ~n7875 ;
  assign n7877 = n1424 & ~n7876 ;
  assign n7878 = n1428 & ~n7877 ;
  assign n7879 = n1432 & ~n7878 ;
  assign n7880 = n1436 & ~n7879 ;
  assign n7881 = n1440 & ~n7880 ;
  assign n7882 = n1444 & ~n7881 ;
  assign n7883 = n1448 & ~n7882 ;
  assign n7884 = n1452 & ~n7883 ;
  assign n7885 = n1456 & ~n7884 ;
  assign n7886 = n1460 & ~n7885 ;
  assign n7887 = n1464 & ~n7886 ;
  assign n7888 = n1468 & ~n7887 ;
  assign n7889 = n1472 & ~n7888 ;
  assign n7890 = n1476 & ~n7889 ;
  assign n7891 = n1480 & ~n7890 ;
  assign n7892 = n1484 & ~n7891 ;
  assign n7893 = n1488 & ~n7892 ;
  assign n7894 = n1492 & ~n7893 ;
  assign n7895 = n1496 & ~n7894 ;
  assign n7896 = n1500 & ~n7895 ;
  assign n7897 = n1504 & ~n7896 ;
  assign n7898 = n1508 & ~n7897 ;
  assign n7899 = n1512 & ~n7898 ;
  assign n7900 = n1516 & ~n7899 ;
  assign n7901 = n1520 & ~n7900 ;
  assign n7902 = n1524 & ~n7901 ;
  assign n7903 = n1528 & ~n7902 ;
  assign n7904 = n1532 & ~n7903 ;
  assign n7905 = n1536 & ~n7904 ;
  assign n7906 = n1540 & ~n7905 ;
  assign n7907 = n1544 & ~n7906 ;
  assign n7908 = n1548 & ~n7907 ;
  assign n7909 = n1552 & ~n7908 ;
  assign n7910 = n1556 & ~n7909 ;
  assign n7911 = n1560 & ~n7910 ;
  assign n7912 = n1564 & ~n7911 ;
  assign n7913 = n1568 & ~n7912 ;
  assign n7914 = n1572 & ~n7913 ;
  assign n7915 = n1576 & ~n7914 ;
  assign n7916 = n1580 & ~n7915 ;
  assign n7917 = n1584 & ~n7916 ;
  assign n7918 = n1588 & ~n7917 ;
  assign n7919 = n1592 & ~n7918 ;
  assign n7920 = n1596 & ~n7919 ;
  assign n7921 = n1600 & ~n7920 ;
  assign n7922 = n1604 & ~n7921 ;
  assign n7923 = n1608 & ~n7922 ;
  assign n7924 = n1612 & ~n7923 ;
  assign n7925 = n2656 & ~n7924 ;
  assign n7926 = n2658 & ~n7925 ;
  assign n7927 = n3192 & ~n7926 ;
  assign n7928 = n1962 & ~n7927 ;
  assign n7929 = n1966 & ~n7928 ;
  assign n7930 = n1970 & ~n7929 ;
  assign n7931 = n1974 & ~n7930 ;
  assign n7932 = n1978 & ~n7931 ;
  assign n7933 = n1982 & ~n7932 ;
  assign n7934 = n1986 & ~n7933 ;
  assign n7935 = n1990 & ~n7934 ;
  assign n7936 = n1994 & ~n7935 ;
  assign n7937 = n1998 & ~n7936 ;
  assign n7938 = n2002 & ~n7937 ;
  assign n7939 = n2006 & ~n7938 ;
  assign n7940 = n2010 & ~n7939 ;
  assign n7941 = n2014 & ~n7940 ;
  assign n7942 = n2018 & ~n7941 ;
  assign n7943 = n2022 & ~n7942 ;
  assign n7944 = n2026 & ~n7943 ;
  assign n7945 = n2030 & ~n7944 ;
  assign n7946 = n2034 & ~n7945 ;
  assign n7947 = ~x162 & ~n2036 ;
  assign n7948 = ~n7946 & n7947 ;
  assign n7951 = ~n7948 & ~x290 ;
  assign n7952 = ~n7950 & ~n7951 ;
  assign n7953 = ~n350 & n1708 ;
  assign n7954 = n1713 & ~n7953 ;
  assign n7955 = n1717 & ~n7954 ;
  assign n7956 = n1721 & ~n7955 ;
  assign n7957 = n1725 & ~n7956 ;
  assign n7958 = n1729 & ~n7957 ;
  assign n7959 = n1733 & ~n7958 ;
  assign n7960 = n1737 & ~n7959 ;
  assign n7961 = n1741 & ~n7960 ;
  assign n7962 = n1745 & ~n7961 ;
  assign n7963 = n1749 & ~n7962 ;
  assign n7964 = n1753 & ~n7963 ;
  assign n7965 = n1757 & ~n7964 ;
  assign n7966 = n1761 & ~n7965 ;
  assign n7967 = n1765 & ~n7966 ;
  assign n7968 = n1769 & ~n7967 ;
  assign n7969 = n1773 & ~n7968 ;
  assign n7970 = n1777 & ~n7969 ;
  assign n7971 = n1781 & ~n7970 ;
  assign n7972 = n1785 & ~n7971 ;
  assign n7973 = n1789 & ~n7972 ;
  assign n7974 = n1793 & ~n7973 ;
  assign n7975 = n1797 & ~n7974 ;
  assign n7976 = n1801 & ~n7975 ;
  assign n7977 = n1805 & ~n7976 ;
  assign n7978 = n1809 & ~n7977 ;
  assign n7979 = n1813 & ~n7978 ;
  assign n7980 = n1817 & ~n7979 ;
  assign n7981 = n1821 & ~n7980 ;
  assign n7982 = n1825 & ~n7981 ;
  assign n7983 = n1829 & ~n7982 ;
  assign n7984 = n1833 & ~n7983 ;
  assign n7985 = n1837 & ~n7984 ;
  assign n7986 = n1841 & ~n7985 ;
  assign n7987 = n1845 & ~n7986 ;
  assign n7988 = n1849 & ~n7987 ;
  assign n7989 = n1853 & ~n7988 ;
  assign n7990 = n1857 & ~n7989 ;
  assign n7991 = n1861 & ~n7990 ;
  assign n7992 = n1865 & ~n7991 ;
  assign n7993 = n1869 & ~n7992 ;
  assign n7994 = n1873 & ~n7993 ;
  assign n7995 = n1877 & ~n7994 ;
  assign n7996 = n1881 & ~n7995 ;
  assign n7997 = n1885 & ~n7996 ;
  assign n7998 = n1889 & ~n7997 ;
  assign n7999 = n1893 & ~n7998 ;
  assign n8000 = n1897 & ~n7999 ;
  assign n8001 = n1901 & ~n8000 ;
  assign n8002 = n1905 & ~n8001 ;
  assign n8003 = n1909 & ~n8002 ;
  assign n8004 = n1913 & ~n8003 ;
  assign n8005 = n1917 & ~n8004 ;
  assign n8006 = n1921 & ~n8005 ;
  assign n8007 = n1925 & ~n8006 ;
  assign n8008 = n1929 & ~n8007 ;
  assign n8009 = n1933 & ~n8008 ;
  assign n8010 = n1937 & ~n8009 ;
  assign n8011 = n1941 & ~n8010 ;
  assign n8012 = n1945 & ~n8011 ;
  assign n8013 = n1949 & ~n8012 ;
  assign n8014 = n1953 & ~n8013 ;
  assign n8015 = n2749 & ~n8014 ;
  assign n8016 = n263 & ~n8015 ;
  assign n8017 = n267 & ~n8016 ;
  assign n8018 = n271 & ~n8017 ;
  assign n8019 = n275 & ~n8018 ;
  assign n8020 = n279 & ~n8019 ;
  assign n8021 = n283 & ~n8020 ;
  assign n8022 = n287 & ~n8021 ;
  assign n8023 = n291 & ~n8022 ;
  assign n8024 = n295 & ~n8023 ;
  assign n8025 = n299 & ~n8024 ;
  assign n8026 = n303 & ~n8025 ;
  assign n8027 = n307 & ~n8026 ;
  assign n8028 = n311 & ~n8027 ;
  assign n8029 = n315 & ~n8028 ;
  assign n8030 = n319 & ~n8029 ;
  assign n8031 = n323 & ~n8030 ;
  assign n8032 = n327 & ~n8031 ;
  assign n8033 = n331 & ~n8032 ;
  assign n8034 = n335 & ~n8033 ;
  assign n8035 = n339 & ~n8034 ;
  assign n8036 = n343 & ~n8035 ;
  assign n8037 = x163 & ~n345 ;
  assign n8038 = ~n8036 & n8037 ;
  assign n8126 = n8038 & x291 ;
  assign n8039 = ~n689 & n2045 ;
  assign n8040 = n2050 & ~n8039 ;
  assign n8041 = n2054 & ~n8040 ;
  assign n8042 = n2058 & ~n8041 ;
  assign n8043 = n2062 & ~n8042 ;
  assign n8044 = n2066 & ~n8043 ;
  assign n8045 = n2070 & ~n8044 ;
  assign n8046 = n2074 & ~n8045 ;
  assign n8047 = n2078 & ~n8046 ;
  assign n8048 = n2082 & ~n8047 ;
  assign n8049 = n2086 & ~n8048 ;
  assign n8050 = n2090 & ~n8049 ;
  assign n8051 = n2094 & ~n8050 ;
  assign n8052 = n2098 & ~n8051 ;
  assign n8053 = n2102 & ~n8052 ;
  assign n8054 = n2106 & ~n8053 ;
  assign n8055 = n2110 & ~n8054 ;
  assign n8056 = n2114 & ~n8055 ;
  assign n8057 = n2118 & ~n8056 ;
  assign n8058 = n2122 & ~n8057 ;
  assign n8059 = n2126 & ~n8058 ;
  assign n8060 = n2130 & ~n8059 ;
  assign n8061 = n2134 & ~n8060 ;
  assign n8062 = n2138 & ~n8061 ;
  assign n8063 = n2142 & ~n8062 ;
  assign n8064 = n2146 & ~n8063 ;
  assign n8065 = n2150 & ~n8064 ;
  assign n8066 = n2154 & ~n8065 ;
  assign n8067 = n2158 & ~n8066 ;
  assign n8068 = n2162 & ~n8067 ;
  assign n8069 = n2166 & ~n8068 ;
  assign n8070 = n2170 & ~n8069 ;
  assign n8071 = n2174 & ~n8070 ;
  assign n8072 = n2178 & ~n8071 ;
  assign n8073 = n2182 & ~n8072 ;
  assign n8074 = n2186 & ~n8073 ;
  assign n8075 = n2190 & ~n8074 ;
  assign n8076 = n2194 & ~n8075 ;
  assign n8077 = n2198 & ~n8076 ;
  assign n8078 = n2202 & ~n8077 ;
  assign n8079 = n2206 & ~n8078 ;
  assign n8080 = n2210 & ~n8079 ;
  assign n8081 = n2214 & ~n8080 ;
  assign n8082 = n2218 & ~n8081 ;
  assign n8083 = n2222 & ~n8082 ;
  assign n8084 = n2226 & ~n8083 ;
  assign n8085 = n2230 & ~n8084 ;
  assign n8086 = n2234 & ~n8085 ;
  assign n8087 = n2238 & ~n8086 ;
  assign n8088 = n2242 & ~n8087 ;
  assign n8089 = n2246 & ~n8088 ;
  assign n8090 = n2250 & ~n8089 ;
  assign n8091 = n2254 & ~n8090 ;
  assign n8092 = n2258 & ~n8091 ;
  assign n8093 = n2262 & ~n8092 ;
  assign n8094 = n2266 & ~n8093 ;
  assign n8095 = n2270 & ~n8094 ;
  assign n8096 = n2274 & ~n8095 ;
  assign n8097 = n2278 & ~n8096 ;
  assign n8098 = n2282 & ~n8097 ;
  assign n8099 = n2286 & ~n8098 ;
  assign n8100 = n2290 & ~n8099 ;
  assign n8101 = n2836 & ~n8100 ;
  assign n8102 = n602 & ~n8101 ;
  assign n8103 = n606 & ~n8102 ;
  assign n8104 = n610 & ~n8103 ;
  assign n8105 = n614 & ~n8104 ;
  assign n8106 = n618 & ~n8105 ;
  assign n8107 = n622 & ~n8106 ;
  assign n8108 = n626 & ~n8107 ;
  assign n8109 = n630 & ~n8108 ;
  assign n8110 = n634 & ~n8109 ;
  assign n8111 = n638 & ~n8110 ;
  assign n8112 = n642 & ~n8111 ;
  assign n8113 = n646 & ~n8112 ;
  assign n8114 = n650 & ~n8113 ;
  assign n8115 = n654 & ~n8114 ;
  assign n8116 = n658 & ~n8115 ;
  assign n8117 = n662 & ~n8116 ;
  assign n8118 = n666 & ~n8117 ;
  assign n8119 = n670 & ~n8118 ;
  assign n8120 = n674 & ~n8119 ;
  assign n8121 = n678 & ~n8120 ;
  assign n8122 = n682 & ~n8121 ;
  assign n8123 = ~x163 & ~n684 ;
  assign n8124 = ~n8122 & n8123 ;
  assign n8127 = ~n8124 & ~x291 ;
  assign n8128 = ~n8126 & ~n8127 ;
  assign n8129 = n354 & ~n1032 ;
  assign n8130 = n359 & ~n8129 ;
  assign n8131 = n363 & ~n8130 ;
  assign n8132 = n367 & ~n8131 ;
  assign n8133 = n371 & ~n8132 ;
  assign n8134 = n375 & ~n8133 ;
  assign n8135 = n379 & ~n8134 ;
  assign n8136 = n383 & ~n8135 ;
  assign n8137 = n387 & ~n8136 ;
  assign n8138 = n391 & ~n8137 ;
  assign n8139 = n395 & ~n8138 ;
  assign n8140 = n399 & ~n8139 ;
  assign n8141 = n403 & ~n8140 ;
  assign n8142 = n407 & ~n8141 ;
  assign n8143 = n411 & ~n8142 ;
  assign n8144 = n415 & ~n8143 ;
  assign n8145 = n419 & ~n8144 ;
  assign n8146 = n423 & ~n8145 ;
  assign n8147 = n427 & ~n8146 ;
  assign n8148 = n431 & ~n8147 ;
  assign n8149 = n435 & ~n8148 ;
  assign n8150 = n439 & ~n8149 ;
  assign n8151 = n443 & ~n8150 ;
  assign n8152 = n447 & ~n8151 ;
  assign n8153 = n451 & ~n8152 ;
  assign n8154 = n455 & ~n8153 ;
  assign n8155 = n459 & ~n8154 ;
  assign n8156 = n463 & ~n8155 ;
  assign n8157 = n467 & ~n8156 ;
  assign n8158 = n471 & ~n8157 ;
  assign n8159 = n475 & ~n8158 ;
  assign n8160 = n479 & ~n8159 ;
  assign n8161 = n483 & ~n8160 ;
  assign n8162 = n487 & ~n8161 ;
  assign n8163 = n491 & ~n8162 ;
  assign n8164 = n495 & ~n8163 ;
  assign n8165 = n499 & ~n8164 ;
  assign n8166 = n503 & ~n8165 ;
  assign n8167 = n507 & ~n8166 ;
  assign n8168 = n511 & ~n8167 ;
  assign n8169 = n515 & ~n8168 ;
  assign n8170 = n519 & ~n8169 ;
  assign n8171 = n523 & ~n8170 ;
  assign n8172 = n527 & ~n8171 ;
  assign n8173 = n531 & ~n8172 ;
  assign n8174 = n535 & ~n8173 ;
  assign n8175 = n539 & ~n8174 ;
  assign n8176 = n543 & ~n8175 ;
  assign n8177 = n547 & ~n8176 ;
  assign n8178 = n551 & ~n8177 ;
  assign n8179 = n555 & ~n8178 ;
  assign n8180 = n559 & ~n8179 ;
  assign n8181 = n563 & ~n8180 ;
  assign n8182 = n567 & ~n8181 ;
  assign n8183 = n571 & ~n8182 ;
  assign n8184 = n575 & ~n8183 ;
  assign n8185 = n579 & ~n8184 ;
  assign n8186 = n583 & ~n8185 ;
  assign n8187 = n587 & ~n8186 ;
  assign n8188 = n591 & ~n8187 ;
  assign n8189 = n2382 & ~n8188 ;
  assign n8190 = n2384 & ~n8189 ;
  assign n8191 = n2927 & ~n8190 ;
  assign n8192 = n945 & ~n8191 ;
  assign n8193 = n949 & ~n8192 ;
  assign n8194 = n953 & ~n8193 ;
  assign n8195 = n957 & ~n8194 ;
  assign n8196 = n961 & ~n8195 ;
  assign n8197 = n965 & ~n8196 ;
  assign n8198 = n969 & ~n8197 ;
  assign n8199 = n973 & ~n8198 ;
  assign n8200 = n977 & ~n8199 ;
  assign n8201 = n981 & ~n8200 ;
  assign n8202 = n985 & ~n8201 ;
  assign n8203 = n989 & ~n8202 ;
  assign n8204 = n993 & ~n8203 ;
  assign n8205 = n997 & ~n8204 ;
  assign n8206 = n1001 & ~n8205 ;
  assign n8207 = n1005 & ~n8206 ;
  assign n8208 = n1009 & ~n8207 ;
  assign n8209 = n1013 & ~n8208 ;
  assign n8210 = n1017 & ~n8209 ;
  assign n8211 = n1021 & ~n8210 ;
  assign n8212 = n1025 & ~n8211 ;
  assign n8213 = x164 & ~n1027 ;
  assign n8214 = ~n8212 & n8213 ;
  assign n8302 = n8214 & x292 ;
  assign n8215 = n693 & ~n1371 ;
  assign n8216 = n698 & ~n8215 ;
  assign n8217 = n702 & ~n8216 ;
  assign n8218 = n706 & ~n8217 ;
  assign n8219 = n710 & ~n8218 ;
  assign n8220 = n714 & ~n8219 ;
  assign n8221 = n718 & ~n8220 ;
  assign n8222 = n722 & ~n8221 ;
  assign n8223 = n726 & ~n8222 ;
  assign n8224 = n730 & ~n8223 ;
  assign n8225 = n734 & ~n8224 ;
  assign n8226 = n738 & ~n8225 ;
  assign n8227 = n742 & ~n8226 ;
  assign n8228 = n746 & ~n8227 ;
  assign n8229 = n750 & ~n8228 ;
  assign n8230 = n754 & ~n8229 ;
  assign n8231 = n758 & ~n8230 ;
  assign n8232 = n762 & ~n8231 ;
  assign n8233 = n766 & ~n8232 ;
  assign n8234 = n770 & ~n8233 ;
  assign n8235 = n774 & ~n8234 ;
  assign n8236 = n778 & ~n8235 ;
  assign n8237 = n782 & ~n8236 ;
  assign n8238 = n786 & ~n8237 ;
  assign n8239 = n790 & ~n8238 ;
  assign n8240 = n794 & ~n8239 ;
  assign n8241 = n798 & ~n8240 ;
  assign n8242 = n802 & ~n8241 ;
  assign n8243 = n806 & ~n8242 ;
  assign n8244 = n810 & ~n8243 ;
  assign n8245 = n814 & ~n8244 ;
  assign n8246 = n818 & ~n8245 ;
  assign n8247 = n822 & ~n8246 ;
  assign n8248 = n826 & ~n8247 ;
  assign n8249 = n830 & ~n8248 ;
  assign n8250 = n834 & ~n8249 ;
  assign n8251 = n838 & ~n8250 ;
  assign n8252 = n842 & ~n8251 ;
  assign n8253 = n846 & ~n8252 ;
  assign n8254 = n850 & ~n8253 ;
  assign n8255 = n854 & ~n8254 ;
  assign n8256 = n858 & ~n8255 ;
  assign n8257 = n862 & ~n8256 ;
  assign n8258 = n866 & ~n8257 ;
  assign n8259 = n870 & ~n8258 ;
  assign n8260 = n874 & ~n8259 ;
  assign n8261 = n878 & ~n8260 ;
  assign n8262 = n882 & ~n8261 ;
  assign n8263 = n886 & ~n8262 ;
  assign n8264 = n890 & ~n8263 ;
  assign n8265 = n894 & ~n8264 ;
  assign n8266 = n898 & ~n8265 ;
  assign n8267 = n902 & ~n8266 ;
  assign n8268 = n906 & ~n8267 ;
  assign n8269 = n910 & ~n8268 ;
  assign n8270 = n914 & ~n8269 ;
  assign n8271 = n918 & ~n8270 ;
  assign n8272 = n922 & ~n8271 ;
  assign n8273 = n926 & ~n8272 ;
  assign n8274 = n930 & ~n8273 ;
  assign n8275 = n2472 & ~n8274 ;
  assign n8276 = n2474 & ~n8275 ;
  assign n8277 = n3014 & ~n8276 ;
  assign n8278 = n1284 & ~n8277 ;
  assign n8279 = n1288 & ~n8278 ;
  assign n8280 = n1292 & ~n8279 ;
  assign n8281 = n1296 & ~n8280 ;
  assign n8282 = n1300 & ~n8281 ;
  assign n8283 = n1304 & ~n8282 ;
  assign n8284 = n1308 & ~n8283 ;
  assign n8285 = n1312 & ~n8284 ;
  assign n8286 = n1316 & ~n8285 ;
  assign n8287 = n1320 & ~n8286 ;
  assign n8288 = n1324 & ~n8287 ;
  assign n8289 = n1328 & ~n8288 ;
  assign n8290 = n1332 & ~n8289 ;
  assign n8291 = n1336 & ~n8290 ;
  assign n8292 = n1340 & ~n8291 ;
  assign n8293 = n1344 & ~n8292 ;
  assign n8294 = n1348 & ~n8293 ;
  assign n8295 = n1352 & ~n8294 ;
  assign n8296 = n1356 & ~n8295 ;
  assign n8297 = n1360 & ~n8296 ;
  assign n8298 = n1364 & ~n8297 ;
  assign n8299 = ~x164 & ~n1366 ;
  assign n8300 = ~n8298 & n8299 ;
  assign n8303 = ~n8300 & ~x292 ;
  assign n8304 = ~n8302 & ~n8303 ;
  assign n8305 = n1036 & ~n1712 ;
  assign n8306 = n1041 & ~n8305 ;
  assign n8307 = n1045 & ~n8306 ;
  assign n8308 = n1049 & ~n8307 ;
  assign n8309 = n1053 & ~n8308 ;
  assign n8310 = n1057 & ~n8309 ;
  assign n8311 = n1061 & ~n8310 ;
  assign n8312 = n1065 & ~n8311 ;
  assign n8313 = n1069 & ~n8312 ;
  assign n8314 = n1073 & ~n8313 ;
  assign n8315 = n1077 & ~n8314 ;
  assign n8316 = n1081 & ~n8315 ;
  assign n8317 = n1085 & ~n8316 ;
  assign n8318 = n1089 & ~n8317 ;
  assign n8319 = n1093 & ~n8318 ;
  assign n8320 = n1097 & ~n8319 ;
  assign n8321 = n1101 & ~n8320 ;
  assign n8322 = n1105 & ~n8321 ;
  assign n8323 = n1109 & ~n8322 ;
  assign n8324 = n1113 & ~n8323 ;
  assign n8325 = n1117 & ~n8324 ;
  assign n8326 = n1121 & ~n8325 ;
  assign n8327 = n1125 & ~n8326 ;
  assign n8328 = n1129 & ~n8327 ;
  assign n8329 = n1133 & ~n8328 ;
  assign n8330 = n1137 & ~n8329 ;
  assign n8331 = n1141 & ~n8330 ;
  assign n8332 = n1145 & ~n8331 ;
  assign n8333 = n1149 & ~n8332 ;
  assign n8334 = n1153 & ~n8333 ;
  assign n8335 = n1157 & ~n8334 ;
  assign n8336 = n1161 & ~n8335 ;
  assign n8337 = n1165 & ~n8336 ;
  assign n8338 = n1169 & ~n8337 ;
  assign n8339 = n1173 & ~n8338 ;
  assign n8340 = n1177 & ~n8339 ;
  assign n8341 = n1181 & ~n8340 ;
  assign n8342 = n1185 & ~n8341 ;
  assign n8343 = n1189 & ~n8342 ;
  assign n8344 = n1193 & ~n8343 ;
  assign n8345 = n1197 & ~n8344 ;
  assign n8346 = n1201 & ~n8345 ;
  assign n8347 = n1205 & ~n8346 ;
  assign n8348 = n1209 & ~n8347 ;
  assign n8349 = n1213 & ~n8348 ;
  assign n8350 = n1217 & ~n8349 ;
  assign n8351 = n1221 & ~n8350 ;
  assign n8352 = n1225 & ~n8351 ;
  assign n8353 = n1229 & ~n8352 ;
  assign n8354 = n1233 & ~n8353 ;
  assign n8355 = n1237 & ~n8354 ;
  assign n8356 = n1241 & ~n8355 ;
  assign n8357 = n1245 & ~n8356 ;
  assign n8358 = n1249 & ~n8357 ;
  assign n8359 = n1253 & ~n8358 ;
  assign n8360 = n1257 & ~n8359 ;
  assign n8361 = n1261 & ~n8360 ;
  assign n8362 = n1265 & ~n8361 ;
  assign n8363 = n1269 & ~n8362 ;
  assign n8364 = n1273 & ~n8363 ;
  assign n8365 = n2566 & ~n8364 ;
  assign n8366 = n2568 & ~n8365 ;
  assign n8367 = n3105 & ~n8366 ;
  assign n8368 = n1625 & ~n8367 ;
  assign n8369 = n1629 & ~n8368 ;
  assign n8370 = n1633 & ~n8369 ;
  assign n8371 = n1637 & ~n8370 ;
  assign n8372 = n1641 & ~n8371 ;
  assign n8373 = n1645 & ~n8372 ;
  assign n8374 = n1649 & ~n8373 ;
  assign n8375 = n1653 & ~n8374 ;
  assign n8376 = n1657 & ~n8375 ;
  assign n8377 = n1661 & ~n8376 ;
  assign n8378 = n1665 & ~n8377 ;
  assign n8379 = n1669 & ~n8378 ;
  assign n8380 = n1673 & ~n8379 ;
  assign n8381 = n1677 & ~n8380 ;
  assign n8382 = n1681 & ~n8381 ;
  assign n8383 = n1685 & ~n8382 ;
  assign n8384 = n1689 & ~n8383 ;
  assign n8385 = n1693 & ~n8384 ;
  assign n8386 = n1697 & ~n8385 ;
  assign n8387 = n1701 & ~n8386 ;
  assign n8388 = n1705 & ~n8387 ;
  assign n8389 = x165 & ~n1707 ;
  assign n8390 = ~n8388 & n8389 ;
  assign n8478 = n8390 & x293 ;
  assign n8391 = n1375 & ~n2049 ;
  assign n8392 = n1380 & ~n8391 ;
  assign n8393 = n1384 & ~n8392 ;
  assign n8394 = n1388 & ~n8393 ;
  assign n8395 = n1392 & ~n8394 ;
  assign n8396 = n1396 & ~n8395 ;
  assign n8397 = n1400 & ~n8396 ;
  assign n8398 = n1404 & ~n8397 ;
  assign n8399 = n1408 & ~n8398 ;
  assign n8400 = n1412 & ~n8399 ;
  assign n8401 = n1416 & ~n8400 ;
  assign n8402 = n1420 & ~n8401 ;
  assign n8403 = n1424 & ~n8402 ;
  assign n8404 = n1428 & ~n8403 ;
  assign n8405 = n1432 & ~n8404 ;
  assign n8406 = n1436 & ~n8405 ;
  assign n8407 = n1440 & ~n8406 ;
  assign n8408 = n1444 & ~n8407 ;
  assign n8409 = n1448 & ~n8408 ;
  assign n8410 = n1452 & ~n8409 ;
  assign n8411 = n1456 & ~n8410 ;
  assign n8412 = n1460 & ~n8411 ;
  assign n8413 = n1464 & ~n8412 ;
  assign n8414 = n1468 & ~n8413 ;
  assign n8415 = n1472 & ~n8414 ;
  assign n8416 = n1476 & ~n8415 ;
  assign n8417 = n1480 & ~n8416 ;
  assign n8418 = n1484 & ~n8417 ;
  assign n8419 = n1488 & ~n8418 ;
  assign n8420 = n1492 & ~n8419 ;
  assign n8421 = n1496 & ~n8420 ;
  assign n8422 = n1500 & ~n8421 ;
  assign n8423 = n1504 & ~n8422 ;
  assign n8424 = n1508 & ~n8423 ;
  assign n8425 = n1512 & ~n8424 ;
  assign n8426 = n1516 & ~n8425 ;
  assign n8427 = n1520 & ~n8426 ;
  assign n8428 = n1524 & ~n8427 ;
  assign n8429 = n1528 & ~n8428 ;
  assign n8430 = n1532 & ~n8429 ;
  assign n8431 = n1536 & ~n8430 ;
  assign n8432 = n1540 & ~n8431 ;
  assign n8433 = n1544 & ~n8432 ;
  assign n8434 = n1548 & ~n8433 ;
  assign n8435 = n1552 & ~n8434 ;
  assign n8436 = n1556 & ~n8435 ;
  assign n8437 = n1560 & ~n8436 ;
  assign n8438 = n1564 & ~n8437 ;
  assign n8439 = n1568 & ~n8438 ;
  assign n8440 = n1572 & ~n8439 ;
  assign n8441 = n1576 & ~n8440 ;
  assign n8442 = n1580 & ~n8441 ;
  assign n8443 = n1584 & ~n8442 ;
  assign n8444 = n1588 & ~n8443 ;
  assign n8445 = n1592 & ~n8444 ;
  assign n8446 = n1596 & ~n8445 ;
  assign n8447 = n1600 & ~n8446 ;
  assign n8448 = n1604 & ~n8447 ;
  assign n8449 = n1608 & ~n8448 ;
  assign n8450 = n1612 & ~n8449 ;
  assign n8451 = n2656 & ~n8450 ;
  assign n8452 = n2658 & ~n8451 ;
  assign n8453 = n3192 & ~n8452 ;
  assign n8454 = n1962 & ~n8453 ;
  assign n8455 = n1966 & ~n8454 ;
  assign n8456 = n1970 & ~n8455 ;
  assign n8457 = n1974 & ~n8456 ;
  assign n8458 = n1978 & ~n8457 ;
  assign n8459 = n1982 & ~n8458 ;
  assign n8460 = n1986 & ~n8459 ;
  assign n8461 = n1990 & ~n8460 ;
  assign n8462 = n1994 & ~n8461 ;
  assign n8463 = n1998 & ~n8462 ;
  assign n8464 = n2002 & ~n8463 ;
  assign n8465 = n2006 & ~n8464 ;
  assign n8466 = n2010 & ~n8465 ;
  assign n8467 = n2014 & ~n8466 ;
  assign n8468 = n2018 & ~n8467 ;
  assign n8469 = n2022 & ~n8468 ;
  assign n8470 = n2026 & ~n8469 ;
  assign n8471 = n2030 & ~n8470 ;
  assign n8472 = n2034 & ~n8471 ;
  assign n8473 = n2038 & ~n8472 ;
  assign n8474 = n2042 & ~n8473 ;
  assign n8475 = ~x165 & ~n2044 ;
  assign n8476 = ~n8474 & n8475 ;
  assign n8479 = ~n8476 & ~x293 ;
  assign n8480 = ~n8478 & ~n8479 ;
  assign n8481 = ~n358 & n1716 ;
  assign n8482 = n1721 & ~n8481 ;
  assign n8483 = n1725 & ~n8482 ;
  assign n8484 = n1729 & ~n8483 ;
  assign n8485 = n1733 & ~n8484 ;
  assign n8486 = n1737 & ~n8485 ;
  assign n8487 = n1741 & ~n8486 ;
  assign n8488 = n1745 & ~n8487 ;
  assign n8489 = n1749 & ~n8488 ;
  assign n8490 = n1753 & ~n8489 ;
  assign n8491 = n1757 & ~n8490 ;
  assign n8492 = n1761 & ~n8491 ;
  assign n8493 = n1765 & ~n8492 ;
  assign n8494 = n1769 & ~n8493 ;
  assign n8495 = n1773 & ~n8494 ;
  assign n8496 = n1777 & ~n8495 ;
  assign n8497 = n1781 & ~n8496 ;
  assign n8498 = n1785 & ~n8497 ;
  assign n8499 = n1789 & ~n8498 ;
  assign n8500 = n1793 & ~n8499 ;
  assign n8501 = n1797 & ~n8500 ;
  assign n8502 = n1801 & ~n8501 ;
  assign n8503 = n1805 & ~n8502 ;
  assign n8504 = n1809 & ~n8503 ;
  assign n8505 = n1813 & ~n8504 ;
  assign n8506 = n1817 & ~n8505 ;
  assign n8507 = n1821 & ~n8506 ;
  assign n8508 = n1825 & ~n8507 ;
  assign n8509 = n1829 & ~n8508 ;
  assign n8510 = n1833 & ~n8509 ;
  assign n8511 = n1837 & ~n8510 ;
  assign n8512 = n1841 & ~n8511 ;
  assign n8513 = n1845 & ~n8512 ;
  assign n8514 = n1849 & ~n8513 ;
  assign n8515 = n1853 & ~n8514 ;
  assign n8516 = n1857 & ~n8515 ;
  assign n8517 = n1861 & ~n8516 ;
  assign n8518 = n1865 & ~n8517 ;
  assign n8519 = n1869 & ~n8518 ;
  assign n8520 = n1873 & ~n8519 ;
  assign n8521 = n1877 & ~n8520 ;
  assign n8522 = n1881 & ~n8521 ;
  assign n8523 = n1885 & ~n8522 ;
  assign n8524 = n1889 & ~n8523 ;
  assign n8525 = n1893 & ~n8524 ;
  assign n8526 = n1897 & ~n8525 ;
  assign n8527 = n1901 & ~n8526 ;
  assign n8528 = n1905 & ~n8527 ;
  assign n8529 = n1909 & ~n8528 ;
  assign n8530 = n1913 & ~n8529 ;
  assign n8531 = n1917 & ~n8530 ;
  assign n8532 = n1921 & ~n8531 ;
  assign n8533 = n1925 & ~n8532 ;
  assign n8534 = n1929 & ~n8533 ;
  assign n8535 = n1933 & ~n8534 ;
  assign n8536 = n1937 & ~n8535 ;
  assign n8537 = n1941 & ~n8536 ;
  assign n8538 = n1945 & ~n8537 ;
  assign n8539 = n1949 & ~n8538 ;
  assign n8540 = n1953 & ~n8539 ;
  assign n8541 = n2749 & ~n8540 ;
  assign n8542 = n263 & ~n8541 ;
  assign n8543 = n267 & ~n8542 ;
  assign n8544 = n271 & ~n8543 ;
  assign n8545 = n275 & ~n8544 ;
  assign n8546 = n279 & ~n8545 ;
  assign n8547 = n283 & ~n8546 ;
  assign n8548 = n287 & ~n8547 ;
  assign n8549 = n291 & ~n8548 ;
  assign n8550 = n295 & ~n8549 ;
  assign n8551 = n299 & ~n8550 ;
  assign n8552 = n303 & ~n8551 ;
  assign n8553 = n307 & ~n8552 ;
  assign n8554 = n311 & ~n8553 ;
  assign n8555 = n315 & ~n8554 ;
  assign n8556 = n319 & ~n8555 ;
  assign n8557 = n323 & ~n8556 ;
  assign n8558 = n327 & ~n8557 ;
  assign n8559 = n331 & ~n8558 ;
  assign n8560 = n335 & ~n8559 ;
  assign n8561 = n339 & ~n8560 ;
  assign n8562 = n343 & ~n8561 ;
  assign n8563 = n347 & ~n8562 ;
  assign n8564 = n351 & ~n8563 ;
  assign n8565 = x166 & ~n353 ;
  assign n8566 = ~n8564 & n8565 ;
  assign n8654 = n8566 & x294 ;
  assign n8567 = ~n697 & n2053 ;
  assign n8568 = n2058 & ~n8567 ;
  assign n8569 = n2062 & ~n8568 ;
  assign n8570 = n2066 & ~n8569 ;
  assign n8571 = n2070 & ~n8570 ;
  assign n8572 = n2074 & ~n8571 ;
  assign n8573 = n2078 & ~n8572 ;
  assign n8574 = n2082 & ~n8573 ;
  assign n8575 = n2086 & ~n8574 ;
  assign n8576 = n2090 & ~n8575 ;
  assign n8577 = n2094 & ~n8576 ;
  assign n8578 = n2098 & ~n8577 ;
  assign n8579 = n2102 & ~n8578 ;
  assign n8580 = n2106 & ~n8579 ;
  assign n8581 = n2110 & ~n8580 ;
  assign n8582 = n2114 & ~n8581 ;
  assign n8583 = n2118 & ~n8582 ;
  assign n8584 = n2122 & ~n8583 ;
  assign n8585 = n2126 & ~n8584 ;
  assign n8586 = n2130 & ~n8585 ;
  assign n8587 = n2134 & ~n8586 ;
  assign n8588 = n2138 & ~n8587 ;
  assign n8589 = n2142 & ~n8588 ;
  assign n8590 = n2146 & ~n8589 ;
  assign n8591 = n2150 & ~n8590 ;
  assign n8592 = n2154 & ~n8591 ;
  assign n8593 = n2158 & ~n8592 ;
  assign n8594 = n2162 & ~n8593 ;
  assign n8595 = n2166 & ~n8594 ;
  assign n8596 = n2170 & ~n8595 ;
  assign n8597 = n2174 & ~n8596 ;
  assign n8598 = n2178 & ~n8597 ;
  assign n8599 = n2182 & ~n8598 ;
  assign n8600 = n2186 & ~n8599 ;
  assign n8601 = n2190 & ~n8600 ;
  assign n8602 = n2194 & ~n8601 ;
  assign n8603 = n2198 & ~n8602 ;
  assign n8604 = n2202 & ~n8603 ;
  assign n8605 = n2206 & ~n8604 ;
  assign n8606 = n2210 & ~n8605 ;
  assign n8607 = n2214 & ~n8606 ;
  assign n8608 = n2218 & ~n8607 ;
  assign n8609 = n2222 & ~n8608 ;
  assign n8610 = n2226 & ~n8609 ;
  assign n8611 = n2230 & ~n8610 ;
  assign n8612 = n2234 & ~n8611 ;
  assign n8613 = n2238 & ~n8612 ;
  assign n8614 = n2242 & ~n8613 ;
  assign n8615 = n2246 & ~n8614 ;
  assign n8616 = n2250 & ~n8615 ;
  assign n8617 = n2254 & ~n8616 ;
  assign n8618 = n2258 & ~n8617 ;
  assign n8619 = n2262 & ~n8618 ;
  assign n8620 = n2266 & ~n8619 ;
  assign n8621 = n2270 & ~n8620 ;
  assign n8622 = n2274 & ~n8621 ;
  assign n8623 = n2278 & ~n8622 ;
  assign n8624 = n2282 & ~n8623 ;
  assign n8625 = n2286 & ~n8624 ;
  assign n8626 = n2290 & ~n8625 ;
  assign n8627 = n2836 & ~n8626 ;
  assign n8628 = n602 & ~n8627 ;
  assign n8629 = n606 & ~n8628 ;
  assign n8630 = n610 & ~n8629 ;
  assign n8631 = n614 & ~n8630 ;
  assign n8632 = n618 & ~n8631 ;
  assign n8633 = n622 & ~n8632 ;
  assign n8634 = n626 & ~n8633 ;
  assign n8635 = n630 & ~n8634 ;
  assign n8636 = n634 & ~n8635 ;
  assign n8637 = n638 & ~n8636 ;
  assign n8638 = n642 & ~n8637 ;
  assign n8639 = n646 & ~n8638 ;
  assign n8640 = n650 & ~n8639 ;
  assign n8641 = n654 & ~n8640 ;
  assign n8642 = n658 & ~n8641 ;
  assign n8643 = n662 & ~n8642 ;
  assign n8644 = n666 & ~n8643 ;
  assign n8645 = n670 & ~n8644 ;
  assign n8646 = n674 & ~n8645 ;
  assign n8647 = n678 & ~n8646 ;
  assign n8648 = n682 & ~n8647 ;
  assign n8649 = n686 & ~n8648 ;
  assign n8650 = n690 & ~n8649 ;
  assign n8651 = ~x166 & ~n692 ;
  assign n8652 = ~n8650 & n8651 ;
  assign n8655 = ~n8652 & ~x294 ;
  assign n8656 = ~n8654 & ~n8655 ;
  assign n8657 = n362 & ~n1040 ;
  assign n8658 = n367 & ~n8657 ;
  assign n8659 = n371 & ~n8658 ;
  assign n8660 = n375 & ~n8659 ;
  assign n8661 = n379 & ~n8660 ;
  assign n8662 = n383 & ~n8661 ;
  assign n8663 = n387 & ~n8662 ;
  assign n8664 = n391 & ~n8663 ;
  assign n8665 = n395 & ~n8664 ;
  assign n8666 = n399 & ~n8665 ;
  assign n8667 = n403 & ~n8666 ;
  assign n8668 = n407 & ~n8667 ;
  assign n8669 = n411 & ~n8668 ;
  assign n8670 = n415 & ~n8669 ;
  assign n8671 = n419 & ~n8670 ;
  assign n8672 = n423 & ~n8671 ;
  assign n8673 = n427 & ~n8672 ;
  assign n8674 = n431 & ~n8673 ;
  assign n8675 = n435 & ~n8674 ;
  assign n8676 = n439 & ~n8675 ;
  assign n8677 = n443 & ~n8676 ;
  assign n8678 = n447 & ~n8677 ;
  assign n8679 = n451 & ~n8678 ;
  assign n8680 = n455 & ~n8679 ;
  assign n8681 = n459 & ~n8680 ;
  assign n8682 = n463 & ~n8681 ;
  assign n8683 = n467 & ~n8682 ;
  assign n8684 = n471 & ~n8683 ;
  assign n8685 = n475 & ~n8684 ;
  assign n8686 = n479 & ~n8685 ;
  assign n8687 = n483 & ~n8686 ;
  assign n8688 = n487 & ~n8687 ;
  assign n8689 = n491 & ~n8688 ;
  assign n8690 = n495 & ~n8689 ;
  assign n8691 = n499 & ~n8690 ;
  assign n8692 = n503 & ~n8691 ;
  assign n8693 = n507 & ~n8692 ;
  assign n8694 = n511 & ~n8693 ;
  assign n8695 = n515 & ~n8694 ;
  assign n8696 = n519 & ~n8695 ;
  assign n8697 = n523 & ~n8696 ;
  assign n8698 = n527 & ~n8697 ;
  assign n8699 = n531 & ~n8698 ;
  assign n8700 = n535 & ~n8699 ;
  assign n8701 = n539 & ~n8700 ;
  assign n8702 = n543 & ~n8701 ;
  assign n8703 = n547 & ~n8702 ;
  assign n8704 = n551 & ~n8703 ;
  assign n8705 = n555 & ~n8704 ;
  assign n8706 = n559 & ~n8705 ;
  assign n8707 = n563 & ~n8706 ;
  assign n8708 = n567 & ~n8707 ;
  assign n8709 = n571 & ~n8708 ;
  assign n8710 = n575 & ~n8709 ;
  assign n8711 = n579 & ~n8710 ;
  assign n8712 = n583 & ~n8711 ;
  assign n8713 = n587 & ~n8712 ;
  assign n8714 = n591 & ~n8713 ;
  assign n8715 = n2382 & ~n8714 ;
  assign n8716 = n2384 & ~n8715 ;
  assign n8717 = n2927 & ~n8716 ;
  assign n8718 = n945 & ~n8717 ;
  assign n8719 = n949 & ~n8718 ;
  assign n8720 = n953 & ~n8719 ;
  assign n8721 = n957 & ~n8720 ;
  assign n8722 = n961 & ~n8721 ;
  assign n8723 = n965 & ~n8722 ;
  assign n8724 = n969 & ~n8723 ;
  assign n8725 = n973 & ~n8724 ;
  assign n8726 = n977 & ~n8725 ;
  assign n8727 = n981 & ~n8726 ;
  assign n8728 = n985 & ~n8727 ;
  assign n8729 = n989 & ~n8728 ;
  assign n8730 = n993 & ~n8729 ;
  assign n8731 = n997 & ~n8730 ;
  assign n8732 = n1001 & ~n8731 ;
  assign n8733 = n1005 & ~n8732 ;
  assign n8734 = n1009 & ~n8733 ;
  assign n8735 = n1013 & ~n8734 ;
  assign n8736 = n1017 & ~n8735 ;
  assign n8737 = n1021 & ~n8736 ;
  assign n8738 = n1025 & ~n8737 ;
  assign n8739 = n1029 & ~n8738 ;
  assign n8740 = n1033 & ~n8739 ;
  assign n8741 = x167 & ~n1035 ;
  assign n8742 = ~n8740 & n8741 ;
  assign n8830 = n8742 & x295 ;
  assign n8743 = n701 & ~n1379 ;
  assign n8744 = n706 & ~n8743 ;
  assign n8745 = n710 & ~n8744 ;
  assign n8746 = n714 & ~n8745 ;
  assign n8747 = n718 & ~n8746 ;
  assign n8748 = n722 & ~n8747 ;
  assign n8749 = n726 & ~n8748 ;
  assign n8750 = n730 & ~n8749 ;
  assign n8751 = n734 & ~n8750 ;
  assign n8752 = n738 & ~n8751 ;
  assign n8753 = n742 & ~n8752 ;
  assign n8754 = n746 & ~n8753 ;
  assign n8755 = n750 & ~n8754 ;
  assign n8756 = n754 & ~n8755 ;
  assign n8757 = n758 & ~n8756 ;
  assign n8758 = n762 & ~n8757 ;
  assign n8759 = n766 & ~n8758 ;
  assign n8760 = n770 & ~n8759 ;
  assign n8761 = n774 & ~n8760 ;
  assign n8762 = n778 & ~n8761 ;
  assign n8763 = n782 & ~n8762 ;
  assign n8764 = n786 & ~n8763 ;
  assign n8765 = n790 & ~n8764 ;
  assign n8766 = n794 & ~n8765 ;
  assign n8767 = n798 & ~n8766 ;
  assign n8768 = n802 & ~n8767 ;
  assign n8769 = n806 & ~n8768 ;
  assign n8770 = n810 & ~n8769 ;
  assign n8771 = n814 & ~n8770 ;
  assign n8772 = n818 & ~n8771 ;
  assign n8773 = n822 & ~n8772 ;
  assign n8774 = n826 & ~n8773 ;
  assign n8775 = n830 & ~n8774 ;
  assign n8776 = n834 & ~n8775 ;
  assign n8777 = n838 & ~n8776 ;
  assign n8778 = n842 & ~n8777 ;
  assign n8779 = n846 & ~n8778 ;
  assign n8780 = n850 & ~n8779 ;
  assign n8781 = n854 & ~n8780 ;
  assign n8782 = n858 & ~n8781 ;
  assign n8783 = n862 & ~n8782 ;
  assign n8784 = n866 & ~n8783 ;
  assign n8785 = n870 & ~n8784 ;
  assign n8786 = n874 & ~n8785 ;
  assign n8787 = n878 & ~n8786 ;
  assign n8788 = n882 & ~n8787 ;
  assign n8789 = n886 & ~n8788 ;
  assign n8790 = n890 & ~n8789 ;
  assign n8791 = n894 & ~n8790 ;
  assign n8792 = n898 & ~n8791 ;
  assign n8793 = n902 & ~n8792 ;
  assign n8794 = n906 & ~n8793 ;
  assign n8795 = n910 & ~n8794 ;
  assign n8796 = n914 & ~n8795 ;
  assign n8797 = n918 & ~n8796 ;
  assign n8798 = n922 & ~n8797 ;
  assign n8799 = n926 & ~n8798 ;
  assign n8800 = n930 & ~n8799 ;
  assign n8801 = n2472 & ~n8800 ;
  assign n8802 = n2474 & ~n8801 ;
  assign n8803 = n3014 & ~n8802 ;
  assign n8804 = n1284 & ~n8803 ;
  assign n8805 = n1288 & ~n8804 ;
  assign n8806 = n1292 & ~n8805 ;
  assign n8807 = n1296 & ~n8806 ;
  assign n8808 = n1300 & ~n8807 ;
  assign n8809 = n1304 & ~n8808 ;
  assign n8810 = n1308 & ~n8809 ;
  assign n8811 = n1312 & ~n8810 ;
  assign n8812 = n1316 & ~n8811 ;
  assign n8813 = n1320 & ~n8812 ;
  assign n8814 = n1324 & ~n8813 ;
  assign n8815 = n1328 & ~n8814 ;
  assign n8816 = n1332 & ~n8815 ;
  assign n8817 = n1336 & ~n8816 ;
  assign n8818 = n1340 & ~n8817 ;
  assign n8819 = n1344 & ~n8818 ;
  assign n8820 = n1348 & ~n8819 ;
  assign n8821 = n1352 & ~n8820 ;
  assign n8822 = n1356 & ~n8821 ;
  assign n8823 = n1360 & ~n8822 ;
  assign n8824 = n1364 & ~n8823 ;
  assign n8825 = n1368 & ~n8824 ;
  assign n8826 = n1372 & ~n8825 ;
  assign n8827 = ~x167 & ~n1374 ;
  assign n8828 = ~n8826 & n8827 ;
  assign n8831 = ~n8828 & ~x295 ;
  assign n8832 = ~n8830 & ~n8831 ;
  assign n8833 = n1044 & ~n1720 ;
  assign n8834 = n1049 & ~n8833 ;
  assign n8835 = n1053 & ~n8834 ;
  assign n8836 = n1057 & ~n8835 ;
  assign n8837 = n1061 & ~n8836 ;
  assign n8838 = n1065 & ~n8837 ;
  assign n8839 = n1069 & ~n8838 ;
  assign n8840 = n1073 & ~n8839 ;
  assign n8841 = n1077 & ~n8840 ;
  assign n8842 = n1081 & ~n8841 ;
  assign n8843 = n1085 & ~n8842 ;
  assign n8844 = n1089 & ~n8843 ;
  assign n8845 = n1093 & ~n8844 ;
  assign n8846 = n1097 & ~n8845 ;
  assign n8847 = n1101 & ~n8846 ;
  assign n8848 = n1105 & ~n8847 ;
  assign n8849 = n1109 & ~n8848 ;
  assign n8850 = n1113 & ~n8849 ;
  assign n8851 = n1117 & ~n8850 ;
  assign n8852 = n1121 & ~n8851 ;
  assign n8853 = n1125 & ~n8852 ;
  assign n8854 = n1129 & ~n8853 ;
  assign n8855 = n1133 & ~n8854 ;
  assign n8856 = n1137 & ~n8855 ;
  assign n8857 = n1141 & ~n8856 ;
  assign n8858 = n1145 & ~n8857 ;
  assign n8859 = n1149 & ~n8858 ;
  assign n8860 = n1153 & ~n8859 ;
  assign n8861 = n1157 & ~n8860 ;
  assign n8862 = n1161 & ~n8861 ;
  assign n8863 = n1165 & ~n8862 ;
  assign n8864 = n1169 & ~n8863 ;
  assign n8865 = n1173 & ~n8864 ;
  assign n8866 = n1177 & ~n8865 ;
  assign n8867 = n1181 & ~n8866 ;
  assign n8868 = n1185 & ~n8867 ;
  assign n8869 = n1189 & ~n8868 ;
  assign n8870 = n1193 & ~n8869 ;
  assign n8871 = n1197 & ~n8870 ;
  assign n8872 = n1201 & ~n8871 ;
  assign n8873 = n1205 & ~n8872 ;
  assign n8874 = n1209 & ~n8873 ;
  assign n8875 = n1213 & ~n8874 ;
  assign n8876 = n1217 & ~n8875 ;
  assign n8877 = n1221 & ~n8876 ;
  assign n8878 = n1225 & ~n8877 ;
  assign n8879 = n1229 & ~n8878 ;
  assign n8880 = n1233 & ~n8879 ;
  assign n8881 = n1237 & ~n8880 ;
  assign n8882 = n1241 & ~n8881 ;
  assign n8883 = n1245 & ~n8882 ;
  assign n8884 = n1249 & ~n8883 ;
  assign n8885 = n1253 & ~n8884 ;
  assign n8886 = n1257 & ~n8885 ;
  assign n8887 = n1261 & ~n8886 ;
  assign n8888 = n1265 & ~n8887 ;
  assign n8889 = n1269 & ~n8888 ;
  assign n8890 = n1273 & ~n8889 ;
  assign n8891 = n2566 & ~n8890 ;
  assign n8892 = n2568 & ~n8891 ;
  assign n8893 = n3105 & ~n8892 ;
  assign n8894 = n1625 & ~n8893 ;
  assign n8895 = n1629 & ~n8894 ;
  assign n8896 = n1633 & ~n8895 ;
  assign n8897 = n1637 & ~n8896 ;
  assign n8898 = n1641 & ~n8897 ;
  assign n8899 = n1645 & ~n8898 ;
  assign n8900 = n1649 & ~n8899 ;
  assign n8901 = n1653 & ~n8900 ;
  assign n8902 = n1657 & ~n8901 ;
  assign n8903 = n1661 & ~n8902 ;
  assign n8904 = n1665 & ~n8903 ;
  assign n8905 = n1669 & ~n8904 ;
  assign n8906 = n1673 & ~n8905 ;
  assign n8907 = n1677 & ~n8906 ;
  assign n8908 = n1681 & ~n8907 ;
  assign n8909 = n1685 & ~n8908 ;
  assign n8910 = n1689 & ~n8909 ;
  assign n8911 = n1693 & ~n8910 ;
  assign n8912 = n1697 & ~n8911 ;
  assign n8913 = n1701 & ~n8912 ;
  assign n8914 = n1705 & ~n8913 ;
  assign n8915 = n1709 & ~n8914 ;
  assign n8916 = n1713 & ~n8915 ;
  assign n8917 = x168 & ~n1715 ;
  assign n8918 = ~n8916 & n8917 ;
  assign n9006 = n8918 & x296 ;
  assign n8919 = n1383 & ~n2057 ;
  assign n8920 = n1388 & ~n8919 ;
  assign n8921 = n1392 & ~n8920 ;
  assign n8922 = n1396 & ~n8921 ;
  assign n8923 = n1400 & ~n8922 ;
  assign n8924 = n1404 & ~n8923 ;
  assign n8925 = n1408 & ~n8924 ;
  assign n8926 = n1412 & ~n8925 ;
  assign n8927 = n1416 & ~n8926 ;
  assign n8928 = n1420 & ~n8927 ;
  assign n8929 = n1424 & ~n8928 ;
  assign n8930 = n1428 & ~n8929 ;
  assign n8931 = n1432 & ~n8930 ;
  assign n8932 = n1436 & ~n8931 ;
  assign n8933 = n1440 & ~n8932 ;
  assign n8934 = n1444 & ~n8933 ;
  assign n8935 = n1448 & ~n8934 ;
  assign n8936 = n1452 & ~n8935 ;
  assign n8937 = n1456 & ~n8936 ;
  assign n8938 = n1460 & ~n8937 ;
  assign n8939 = n1464 & ~n8938 ;
  assign n8940 = n1468 & ~n8939 ;
  assign n8941 = n1472 & ~n8940 ;
  assign n8942 = n1476 & ~n8941 ;
  assign n8943 = n1480 & ~n8942 ;
  assign n8944 = n1484 & ~n8943 ;
  assign n8945 = n1488 & ~n8944 ;
  assign n8946 = n1492 & ~n8945 ;
  assign n8947 = n1496 & ~n8946 ;
  assign n8948 = n1500 & ~n8947 ;
  assign n8949 = n1504 & ~n8948 ;
  assign n8950 = n1508 & ~n8949 ;
  assign n8951 = n1512 & ~n8950 ;
  assign n8952 = n1516 & ~n8951 ;
  assign n8953 = n1520 & ~n8952 ;
  assign n8954 = n1524 & ~n8953 ;
  assign n8955 = n1528 & ~n8954 ;
  assign n8956 = n1532 & ~n8955 ;
  assign n8957 = n1536 & ~n8956 ;
  assign n8958 = n1540 & ~n8957 ;
  assign n8959 = n1544 & ~n8958 ;
  assign n8960 = n1548 & ~n8959 ;
  assign n8961 = n1552 & ~n8960 ;
  assign n8962 = n1556 & ~n8961 ;
  assign n8963 = n1560 & ~n8962 ;
  assign n8964 = n1564 & ~n8963 ;
  assign n8965 = n1568 & ~n8964 ;
  assign n8966 = n1572 & ~n8965 ;
  assign n8967 = n1576 & ~n8966 ;
  assign n8968 = n1580 & ~n8967 ;
  assign n8969 = n1584 & ~n8968 ;
  assign n8970 = n1588 & ~n8969 ;
  assign n8971 = n1592 & ~n8970 ;
  assign n8972 = n1596 & ~n8971 ;
  assign n8973 = n1600 & ~n8972 ;
  assign n8974 = n1604 & ~n8973 ;
  assign n8975 = n1608 & ~n8974 ;
  assign n8976 = n1612 & ~n8975 ;
  assign n8977 = n2656 & ~n8976 ;
  assign n8978 = n2658 & ~n8977 ;
  assign n8979 = n3192 & ~n8978 ;
  assign n8980 = n1962 & ~n8979 ;
  assign n8981 = n1966 & ~n8980 ;
  assign n8982 = n1970 & ~n8981 ;
  assign n8983 = n1974 & ~n8982 ;
  assign n8984 = n1978 & ~n8983 ;
  assign n8985 = n1982 & ~n8984 ;
  assign n8986 = n1986 & ~n8985 ;
  assign n8987 = n1990 & ~n8986 ;
  assign n8988 = n1994 & ~n8987 ;
  assign n8989 = n1998 & ~n8988 ;
  assign n8990 = n2002 & ~n8989 ;
  assign n8991 = n2006 & ~n8990 ;
  assign n8992 = n2010 & ~n8991 ;
  assign n8993 = n2014 & ~n8992 ;
  assign n8994 = n2018 & ~n8993 ;
  assign n8995 = n2022 & ~n8994 ;
  assign n8996 = n2026 & ~n8995 ;
  assign n8997 = n2030 & ~n8996 ;
  assign n8998 = n2034 & ~n8997 ;
  assign n8999 = n2038 & ~n8998 ;
  assign n9000 = n2042 & ~n8999 ;
  assign n9001 = n2046 & ~n9000 ;
  assign n9002 = n2050 & ~n9001 ;
  assign n9003 = ~x168 & ~n2052 ;
  assign n9004 = ~n9002 & n9003 ;
  assign n9007 = ~n9004 & ~x296 ;
  assign n9008 = ~n9006 & ~n9007 ;
  assign n9009 = ~n366 & n1724 ;
  assign n9010 = n1729 & ~n9009 ;
  assign n9011 = n1733 & ~n9010 ;
  assign n9012 = n1737 & ~n9011 ;
  assign n9013 = n1741 & ~n9012 ;
  assign n9014 = n1745 & ~n9013 ;
  assign n9015 = n1749 & ~n9014 ;
  assign n9016 = n1753 & ~n9015 ;
  assign n9017 = n1757 & ~n9016 ;
  assign n9018 = n1761 & ~n9017 ;
  assign n9019 = n1765 & ~n9018 ;
  assign n9020 = n1769 & ~n9019 ;
  assign n9021 = n1773 & ~n9020 ;
  assign n9022 = n1777 & ~n9021 ;
  assign n9023 = n1781 & ~n9022 ;
  assign n9024 = n1785 & ~n9023 ;
  assign n9025 = n1789 & ~n9024 ;
  assign n9026 = n1793 & ~n9025 ;
  assign n9027 = n1797 & ~n9026 ;
  assign n9028 = n1801 & ~n9027 ;
  assign n9029 = n1805 & ~n9028 ;
  assign n9030 = n1809 & ~n9029 ;
  assign n9031 = n1813 & ~n9030 ;
  assign n9032 = n1817 & ~n9031 ;
  assign n9033 = n1821 & ~n9032 ;
  assign n9034 = n1825 & ~n9033 ;
  assign n9035 = n1829 & ~n9034 ;
  assign n9036 = n1833 & ~n9035 ;
  assign n9037 = n1837 & ~n9036 ;
  assign n9038 = n1841 & ~n9037 ;
  assign n9039 = n1845 & ~n9038 ;
  assign n9040 = n1849 & ~n9039 ;
  assign n9041 = n1853 & ~n9040 ;
  assign n9042 = n1857 & ~n9041 ;
  assign n9043 = n1861 & ~n9042 ;
  assign n9044 = n1865 & ~n9043 ;
  assign n9045 = n1869 & ~n9044 ;
  assign n9046 = n1873 & ~n9045 ;
  assign n9047 = n1877 & ~n9046 ;
  assign n9048 = n1881 & ~n9047 ;
  assign n9049 = n1885 & ~n9048 ;
  assign n9050 = n1889 & ~n9049 ;
  assign n9051 = n1893 & ~n9050 ;
  assign n9052 = n1897 & ~n9051 ;
  assign n9053 = n1901 & ~n9052 ;
  assign n9054 = n1905 & ~n9053 ;
  assign n9055 = n1909 & ~n9054 ;
  assign n9056 = n1913 & ~n9055 ;
  assign n9057 = n1917 & ~n9056 ;
  assign n9058 = n1921 & ~n9057 ;
  assign n9059 = n1925 & ~n9058 ;
  assign n9060 = n1929 & ~n9059 ;
  assign n9061 = n1933 & ~n9060 ;
  assign n9062 = n1937 & ~n9061 ;
  assign n9063 = n1941 & ~n9062 ;
  assign n9064 = n1945 & ~n9063 ;
  assign n9065 = n1949 & ~n9064 ;
  assign n9066 = n1953 & ~n9065 ;
  assign n9067 = n2749 & ~n9066 ;
  assign n9068 = n263 & ~n9067 ;
  assign n9069 = n267 & ~n9068 ;
  assign n9070 = n271 & ~n9069 ;
  assign n9071 = n275 & ~n9070 ;
  assign n9072 = n279 & ~n9071 ;
  assign n9073 = n283 & ~n9072 ;
  assign n9074 = n287 & ~n9073 ;
  assign n9075 = n291 & ~n9074 ;
  assign n9076 = n295 & ~n9075 ;
  assign n9077 = n299 & ~n9076 ;
  assign n9078 = n303 & ~n9077 ;
  assign n9079 = n307 & ~n9078 ;
  assign n9080 = n311 & ~n9079 ;
  assign n9081 = n315 & ~n9080 ;
  assign n9082 = n319 & ~n9081 ;
  assign n9083 = n323 & ~n9082 ;
  assign n9084 = n327 & ~n9083 ;
  assign n9085 = n331 & ~n9084 ;
  assign n9086 = n335 & ~n9085 ;
  assign n9087 = n339 & ~n9086 ;
  assign n9088 = n343 & ~n9087 ;
  assign n9089 = n347 & ~n9088 ;
  assign n9090 = n351 & ~n9089 ;
  assign n9091 = n355 & ~n9090 ;
  assign n9092 = n359 & ~n9091 ;
  assign n9093 = x169 & ~n361 ;
  assign n9094 = ~n9092 & n9093 ;
  assign n9182 = n9094 & x297 ;
  assign n9095 = ~n705 & n2061 ;
  assign n9096 = n2066 & ~n9095 ;
  assign n9097 = n2070 & ~n9096 ;
  assign n9098 = n2074 & ~n9097 ;
  assign n9099 = n2078 & ~n9098 ;
  assign n9100 = n2082 & ~n9099 ;
  assign n9101 = n2086 & ~n9100 ;
  assign n9102 = n2090 & ~n9101 ;
  assign n9103 = n2094 & ~n9102 ;
  assign n9104 = n2098 & ~n9103 ;
  assign n9105 = n2102 & ~n9104 ;
  assign n9106 = n2106 & ~n9105 ;
  assign n9107 = n2110 & ~n9106 ;
  assign n9108 = n2114 & ~n9107 ;
  assign n9109 = n2118 & ~n9108 ;
  assign n9110 = n2122 & ~n9109 ;
  assign n9111 = n2126 & ~n9110 ;
  assign n9112 = n2130 & ~n9111 ;
  assign n9113 = n2134 & ~n9112 ;
  assign n9114 = n2138 & ~n9113 ;
  assign n9115 = n2142 & ~n9114 ;
  assign n9116 = n2146 & ~n9115 ;
  assign n9117 = n2150 & ~n9116 ;
  assign n9118 = n2154 & ~n9117 ;
  assign n9119 = n2158 & ~n9118 ;
  assign n9120 = n2162 & ~n9119 ;
  assign n9121 = n2166 & ~n9120 ;
  assign n9122 = n2170 & ~n9121 ;
  assign n9123 = n2174 & ~n9122 ;
  assign n9124 = n2178 & ~n9123 ;
  assign n9125 = n2182 & ~n9124 ;
  assign n9126 = n2186 & ~n9125 ;
  assign n9127 = n2190 & ~n9126 ;
  assign n9128 = n2194 & ~n9127 ;
  assign n9129 = n2198 & ~n9128 ;
  assign n9130 = n2202 & ~n9129 ;
  assign n9131 = n2206 & ~n9130 ;
  assign n9132 = n2210 & ~n9131 ;
  assign n9133 = n2214 & ~n9132 ;
  assign n9134 = n2218 & ~n9133 ;
  assign n9135 = n2222 & ~n9134 ;
  assign n9136 = n2226 & ~n9135 ;
  assign n9137 = n2230 & ~n9136 ;
  assign n9138 = n2234 & ~n9137 ;
  assign n9139 = n2238 & ~n9138 ;
  assign n9140 = n2242 & ~n9139 ;
  assign n9141 = n2246 & ~n9140 ;
  assign n9142 = n2250 & ~n9141 ;
  assign n9143 = n2254 & ~n9142 ;
  assign n9144 = n2258 & ~n9143 ;
  assign n9145 = n2262 & ~n9144 ;
  assign n9146 = n2266 & ~n9145 ;
  assign n9147 = n2270 & ~n9146 ;
  assign n9148 = n2274 & ~n9147 ;
  assign n9149 = n2278 & ~n9148 ;
  assign n9150 = n2282 & ~n9149 ;
  assign n9151 = n2286 & ~n9150 ;
  assign n9152 = n2290 & ~n9151 ;
  assign n9153 = n2836 & ~n9152 ;
  assign n9154 = n602 & ~n9153 ;
  assign n9155 = n606 & ~n9154 ;
  assign n9156 = n610 & ~n9155 ;
  assign n9157 = n614 & ~n9156 ;
  assign n9158 = n618 & ~n9157 ;
  assign n9159 = n622 & ~n9158 ;
  assign n9160 = n626 & ~n9159 ;
  assign n9161 = n630 & ~n9160 ;
  assign n9162 = n634 & ~n9161 ;
  assign n9163 = n638 & ~n9162 ;
  assign n9164 = n642 & ~n9163 ;
  assign n9165 = n646 & ~n9164 ;
  assign n9166 = n650 & ~n9165 ;
  assign n9167 = n654 & ~n9166 ;
  assign n9168 = n658 & ~n9167 ;
  assign n9169 = n662 & ~n9168 ;
  assign n9170 = n666 & ~n9169 ;
  assign n9171 = n670 & ~n9170 ;
  assign n9172 = n674 & ~n9171 ;
  assign n9173 = n678 & ~n9172 ;
  assign n9174 = n682 & ~n9173 ;
  assign n9175 = n686 & ~n9174 ;
  assign n9176 = n690 & ~n9175 ;
  assign n9177 = n694 & ~n9176 ;
  assign n9178 = n698 & ~n9177 ;
  assign n9179 = ~x169 & ~n700 ;
  assign n9180 = ~n9178 & n9179 ;
  assign n9183 = ~n9180 & ~x297 ;
  assign n9184 = ~n9182 & ~n9183 ;
  assign n9185 = n370 & ~n1048 ;
  assign n9186 = n375 & ~n9185 ;
  assign n9187 = n379 & ~n9186 ;
  assign n9188 = n383 & ~n9187 ;
  assign n9189 = n387 & ~n9188 ;
  assign n9190 = n391 & ~n9189 ;
  assign n9191 = n395 & ~n9190 ;
  assign n9192 = n399 & ~n9191 ;
  assign n9193 = n403 & ~n9192 ;
  assign n9194 = n407 & ~n9193 ;
  assign n9195 = n411 & ~n9194 ;
  assign n9196 = n415 & ~n9195 ;
  assign n9197 = n419 & ~n9196 ;
  assign n9198 = n423 & ~n9197 ;
  assign n9199 = n427 & ~n9198 ;
  assign n9200 = n431 & ~n9199 ;
  assign n9201 = n435 & ~n9200 ;
  assign n9202 = n439 & ~n9201 ;
  assign n9203 = n443 & ~n9202 ;
  assign n9204 = n447 & ~n9203 ;
  assign n9205 = n451 & ~n9204 ;
  assign n9206 = n455 & ~n9205 ;
  assign n9207 = n459 & ~n9206 ;
  assign n9208 = n463 & ~n9207 ;
  assign n9209 = n467 & ~n9208 ;
  assign n9210 = n471 & ~n9209 ;
  assign n9211 = n475 & ~n9210 ;
  assign n9212 = n479 & ~n9211 ;
  assign n9213 = n483 & ~n9212 ;
  assign n9214 = n487 & ~n9213 ;
  assign n9215 = n491 & ~n9214 ;
  assign n9216 = n495 & ~n9215 ;
  assign n9217 = n499 & ~n9216 ;
  assign n9218 = n503 & ~n9217 ;
  assign n9219 = n507 & ~n9218 ;
  assign n9220 = n511 & ~n9219 ;
  assign n9221 = n515 & ~n9220 ;
  assign n9222 = n519 & ~n9221 ;
  assign n9223 = n523 & ~n9222 ;
  assign n9224 = n527 & ~n9223 ;
  assign n9225 = n531 & ~n9224 ;
  assign n9226 = n535 & ~n9225 ;
  assign n9227 = n539 & ~n9226 ;
  assign n9228 = n543 & ~n9227 ;
  assign n9229 = n547 & ~n9228 ;
  assign n9230 = n551 & ~n9229 ;
  assign n9231 = n555 & ~n9230 ;
  assign n9232 = n559 & ~n9231 ;
  assign n9233 = n563 & ~n9232 ;
  assign n9234 = n567 & ~n9233 ;
  assign n9235 = n571 & ~n9234 ;
  assign n9236 = n575 & ~n9235 ;
  assign n9237 = n579 & ~n9236 ;
  assign n9238 = n583 & ~n9237 ;
  assign n9239 = n587 & ~n9238 ;
  assign n9240 = n591 & ~n9239 ;
  assign n9241 = n2382 & ~n9240 ;
  assign n9242 = n2384 & ~n9241 ;
  assign n9243 = n2927 & ~n9242 ;
  assign n9244 = n945 & ~n9243 ;
  assign n9245 = n949 & ~n9244 ;
  assign n9246 = n953 & ~n9245 ;
  assign n9247 = n957 & ~n9246 ;
  assign n9248 = n961 & ~n9247 ;
  assign n9249 = n965 & ~n9248 ;
  assign n9250 = n969 & ~n9249 ;
  assign n9251 = n973 & ~n9250 ;
  assign n9252 = n977 & ~n9251 ;
  assign n9253 = n981 & ~n9252 ;
  assign n9254 = n985 & ~n9253 ;
  assign n9255 = n989 & ~n9254 ;
  assign n9256 = n993 & ~n9255 ;
  assign n9257 = n997 & ~n9256 ;
  assign n9258 = n1001 & ~n9257 ;
  assign n9259 = n1005 & ~n9258 ;
  assign n9260 = n1009 & ~n9259 ;
  assign n9261 = n1013 & ~n9260 ;
  assign n9262 = n1017 & ~n9261 ;
  assign n9263 = n1021 & ~n9262 ;
  assign n9264 = n1025 & ~n9263 ;
  assign n9265 = n1029 & ~n9264 ;
  assign n9266 = n1033 & ~n9265 ;
  assign n9267 = n1037 & ~n9266 ;
  assign n9268 = n1041 & ~n9267 ;
  assign n9269 = x170 & ~n1043 ;
  assign n9270 = ~n9268 & n9269 ;
  assign n9358 = n9270 & x298 ;
  assign n9271 = n709 & ~n1387 ;
  assign n9272 = n714 & ~n9271 ;
  assign n9273 = n718 & ~n9272 ;
  assign n9274 = n722 & ~n9273 ;
  assign n9275 = n726 & ~n9274 ;
  assign n9276 = n730 & ~n9275 ;
  assign n9277 = n734 & ~n9276 ;
  assign n9278 = n738 & ~n9277 ;
  assign n9279 = n742 & ~n9278 ;
  assign n9280 = n746 & ~n9279 ;
  assign n9281 = n750 & ~n9280 ;
  assign n9282 = n754 & ~n9281 ;
  assign n9283 = n758 & ~n9282 ;
  assign n9284 = n762 & ~n9283 ;
  assign n9285 = n766 & ~n9284 ;
  assign n9286 = n770 & ~n9285 ;
  assign n9287 = n774 & ~n9286 ;
  assign n9288 = n778 & ~n9287 ;
  assign n9289 = n782 & ~n9288 ;
  assign n9290 = n786 & ~n9289 ;
  assign n9291 = n790 & ~n9290 ;
  assign n9292 = n794 & ~n9291 ;
  assign n9293 = n798 & ~n9292 ;
  assign n9294 = n802 & ~n9293 ;
  assign n9295 = n806 & ~n9294 ;
  assign n9296 = n810 & ~n9295 ;
  assign n9297 = n814 & ~n9296 ;
  assign n9298 = n818 & ~n9297 ;
  assign n9299 = n822 & ~n9298 ;
  assign n9300 = n826 & ~n9299 ;
  assign n9301 = n830 & ~n9300 ;
  assign n9302 = n834 & ~n9301 ;
  assign n9303 = n838 & ~n9302 ;
  assign n9304 = n842 & ~n9303 ;
  assign n9305 = n846 & ~n9304 ;
  assign n9306 = n850 & ~n9305 ;
  assign n9307 = n854 & ~n9306 ;
  assign n9308 = n858 & ~n9307 ;
  assign n9309 = n862 & ~n9308 ;
  assign n9310 = n866 & ~n9309 ;
  assign n9311 = n870 & ~n9310 ;
  assign n9312 = n874 & ~n9311 ;
  assign n9313 = n878 & ~n9312 ;
  assign n9314 = n882 & ~n9313 ;
  assign n9315 = n886 & ~n9314 ;
  assign n9316 = n890 & ~n9315 ;
  assign n9317 = n894 & ~n9316 ;
  assign n9318 = n898 & ~n9317 ;
  assign n9319 = n902 & ~n9318 ;
  assign n9320 = n906 & ~n9319 ;
  assign n9321 = n910 & ~n9320 ;
  assign n9322 = n914 & ~n9321 ;
  assign n9323 = n918 & ~n9322 ;
  assign n9324 = n922 & ~n9323 ;
  assign n9325 = n926 & ~n9324 ;
  assign n9326 = n930 & ~n9325 ;
  assign n9327 = n2472 & ~n9326 ;
  assign n9328 = n2474 & ~n9327 ;
  assign n9329 = n3014 & ~n9328 ;
  assign n9330 = n1284 & ~n9329 ;
  assign n9331 = n1288 & ~n9330 ;
  assign n9332 = n1292 & ~n9331 ;
  assign n9333 = n1296 & ~n9332 ;
  assign n9334 = n1300 & ~n9333 ;
  assign n9335 = n1304 & ~n9334 ;
  assign n9336 = n1308 & ~n9335 ;
  assign n9337 = n1312 & ~n9336 ;
  assign n9338 = n1316 & ~n9337 ;
  assign n9339 = n1320 & ~n9338 ;
  assign n9340 = n1324 & ~n9339 ;
  assign n9341 = n1328 & ~n9340 ;
  assign n9342 = n1332 & ~n9341 ;
  assign n9343 = n1336 & ~n9342 ;
  assign n9344 = n1340 & ~n9343 ;
  assign n9345 = n1344 & ~n9344 ;
  assign n9346 = n1348 & ~n9345 ;
  assign n9347 = n1352 & ~n9346 ;
  assign n9348 = n1356 & ~n9347 ;
  assign n9349 = n1360 & ~n9348 ;
  assign n9350 = n1364 & ~n9349 ;
  assign n9351 = n1368 & ~n9350 ;
  assign n9352 = n1372 & ~n9351 ;
  assign n9353 = n1376 & ~n9352 ;
  assign n9354 = n1380 & ~n9353 ;
  assign n9355 = ~x170 & ~n1382 ;
  assign n9356 = ~n9354 & n9355 ;
  assign n9359 = ~n9356 & ~x298 ;
  assign n9360 = ~n9358 & ~n9359 ;
  assign n9361 = n1052 & ~n1728 ;
  assign n9362 = n1057 & ~n9361 ;
  assign n9363 = n1061 & ~n9362 ;
  assign n9364 = n1065 & ~n9363 ;
  assign n9365 = n1069 & ~n9364 ;
  assign n9366 = n1073 & ~n9365 ;
  assign n9367 = n1077 & ~n9366 ;
  assign n9368 = n1081 & ~n9367 ;
  assign n9369 = n1085 & ~n9368 ;
  assign n9370 = n1089 & ~n9369 ;
  assign n9371 = n1093 & ~n9370 ;
  assign n9372 = n1097 & ~n9371 ;
  assign n9373 = n1101 & ~n9372 ;
  assign n9374 = n1105 & ~n9373 ;
  assign n9375 = n1109 & ~n9374 ;
  assign n9376 = n1113 & ~n9375 ;
  assign n9377 = n1117 & ~n9376 ;
  assign n9378 = n1121 & ~n9377 ;
  assign n9379 = n1125 & ~n9378 ;
  assign n9380 = n1129 & ~n9379 ;
  assign n9381 = n1133 & ~n9380 ;
  assign n9382 = n1137 & ~n9381 ;
  assign n9383 = n1141 & ~n9382 ;
  assign n9384 = n1145 & ~n9383 ;
  assign n9385 = n1149 & ~n9384 ;
  assign n9386 = n1153 & ~n9385 ;
  assign n9387 = n1157 & ~n9386 ;
  assign n9388 = n1161 & ~n9387 ;
  assign n9389 = n1165 & ~n9388 ;
  assign n9390 = n1169 & ~n9389 ;
  assign n9391 = n1173 & ~n9390 ;
  assign n9392 = n1177 & ~n9391 ;
  assign n9393 = n1181 & ~n9392 ;
  assign n9394 = n1185 & ~n9393 ;
  assign n9395 = n1189 & ~n9394 ;
  assign n9396 = n1193 & ~n9395 ;
  assign n9397 = n1197 & ~n9396 ;
  assign n9398 = n1201 & ~n9397 ;
  assign n9399 = n1205 & ~n9398 ;
  assign n9400 = n1209 & ~n9399 ;
  assign n9401 = n1213 & ~n9400 ;
  assign n9402 = n1217 & ~n9401 ;
  assign n9403 = n1221 & ~n9402 ;
  assign n9404 = n1225 & ~n9403 ;
  assign n9405 = n1229 & ~n9404 ;
  assign n9406 = n1233 & ~n9405 ;
  assign n9407 = n1237 & ~n9406 ;
  assign n9408 = n1241 & ~n9407 ;
  assign n9409 = n1245 & ~n9408 ;
  assign n9410 = n1249 & ~n9409 ;
  assign n9411 = n1253 & ~n9410 ;
  assign n9412 = n1257 & ~n9411 ;
  assign n9413 = n1261 & ~n9412 ;
  assign n9414 = n1265 & ~n9413 ;
  assign n9415 = n1269 & ~n9414 ;
  assign n9416 = n1273 & ~n9415 ;
  assign n9417 = n2566 & ~n9416 ;
  assign n9418 = n2568 & ~n9417 ;
  assign n9419 = n3105 & ~n9418 ;
  assign n9420 = n1625 & ~n9419 ;
  assign n9421 = n1629 & ~n9420 ;
  assign n9422 = n1633 & ~n9421 ;
  assign n9423 = n1637 & ~n9422 ;
  assign n9424 = n1641 & ~n9423 ;
  assign n9425 = n1645 & ~n9424 ;
  assign n9426 = n1649 & ~n9425 ;
  assign n9427 = n1653 & ~n9426 ;
  assign n9428 = n1657 & ~n9427 ;
  assign n9429 = n1661 & ~n9428 ;
  assign n9430 = n1665 & ~n9429 ;
  assign n9431 = n1669 & ~n9430 ;
  assign n9432 = n1673 & ~n9431 ;
  assign n9433 = n1677 & ~n9432 ;
  assign n9434 = n1681 & ~n9433 ;
  assign n9435 = n1685 & ~n9434 ;
  assign n9436 = n1689 & ~n9435 ;
  assign n9437 = n1693 & ~n9436 ;
  assign n9438 = n1697 & ~n9437 ;
  assign n9439 = n1701 & ~n9438 ;
  assign n9440 = n1705 & ~n9439 ;
  assign n9441 = n1709 & ~n9440 ;
  assign n9442 = n1713 & ~n9441 ;
  assign n9443 = n1717 & ~n9442 ;
  assign n9444 = n1721 & ~n9443 ;
  assign n9445 = x171 & ~n1723 ;
  assign n9446 = ~n9444 & n9445 ;
  assign n9534 = n9446 & x299 ;
  assign n9447 = n1391 & ~n2065 ;
  assign n9448 = n1396 & ~n9447 ;
  assign n9449 = n1400 & ~n9448 ;
  assign n9450 = n1404 & ~n9449 ;
  assign n9451 = n1408 & ~n9450 ;
  assign n9452 = n1412 & ~n9451 ;
  assign n9453 = n1416 & ~n9452 ;
  assign n9454 = n1420 & ~n9453 ;
  assign n9455 = n1424 & ~n9454 ;
  assign n9456 = n1428 & ~n9455 ;
  assign n9457 = n1432 & ~n9456 ;
  assign n9458 = n1436 & ~n9457 ;
  assign n9459 = n1440 & ~n9458 ;
  assign n9460 = n1444 & ~n9459 ;
  assign n9461 = n1448 & ~n9460 ;
  assign n9462 = n1452 & ~n9461 ;
  assign n9463 = n1456 & ~n9462 ;
  assign n9464 = n1460 & ~n9463 ;
  assign n9465 = n1464 & ~n9464 ;
  assign n9466 = n1468 & ~n9465 ;
  assign n9467 = n1472 & ~n9466 ;
  assign n9468 = n1476 & ~n9467 ;
  assign n9469 = n1480 & ~n9468 ;
  assign n9470 = n1484 & ~n9469 ;
  assign n9471 = n1488 & ~n9470 ;
  assign n9472 = n1492 & ~n9471 ;
  assign n9473 = n1496 & ~n9472 ;
  assign n9474 = n1500 & ~n9473 ;
  assign n9475 = n1504 & ~n9474 ;
  assign n9476 = n1508 & ~n9475 ;
  assign n9477 = n1512 & ~n9476 ;
  assign n9478 = n1516 & ~n9477 ;
  assign n9479 = n1520 & ~n9478 ;
  assign n9480 = n1524 & ~n9479 ;
  assign n9481 = n1528 & ~n9480 ;
  assign n9482 = n1532 & ~n9481 ;
  assign n9483 = n1536 & ~n9482 ;
  assign n9484 = n1540 & ~n9483 ;
  assign n9485 = n1544 & ~n9484 ;
  assign n9486 = n1548 & ~n9485 ;
  assign n9487 = n1552 & ~n9486 ;
  assign n9488 = n1556 & ~n9487 ;
  assign n9489 = n1560 & ~n9488 ;
  assign n9490 = n1564 & ~n9489 ;
  assign n9491 = n1568 & ~n9490 ;
  assign n9492 = n1572 & ~n9491 ;
  assign n9493 = n1576 & ~n9492 ;
  assign n9494 = n1580 & ~n9493 ;
  assign n9495 = n1584 & ~n9494 ;
  assign n9496 = n1588 & ~n9495 ;
  assign n9497 = n1592 & ~n9496 ;
  assign n9498 = n1596 & ~n9497 ;
  assign n9499 = n1600 & ~n9498 ;
  assign n9500 = n1604 & ~n9499 ;
  assign n9501 = n1608 & ~n9500 ;
  assign n9502 = n1612 & ~n9501 ;
  assign n9503 = n2656 & ~n9502 ;
  assign n9504 = n2658 & ~n9503 ;
  assign n9505 = n3192 & ~n9504 ;
  assign n9506 = n1962 & ~n9505 ;
  assign n9507 = n1966 & ~n9506 ;
  assign n9508 = n1970 & ~n9507 ;
  assign n9509 = n1974 & ~n9508 ;
  assign n9510 = n1978 & ~n9509 ;
  assign n9511 = n1982 & ~n9510 ;
  assign n9512 = n1986 & ~n9511 ;
  assign n9513 = n1990 & ~n9512 ;
  assign n9514 = n1994 & ~n9513 ;
  assign n9515 = n1998 & ~n9514 ;
  assign n9516 = n2002 & ~n9515 ;
  assign n9517 = n2006 & ~n9516 ;
  assign n9518 = n2010 & ~n9517 ;
  assign n9519 = n2014 & ~n9518 ;
  assign n9520 = n2018 & ~n9519 ;
  assign n9521 = n2022 & ~n9520 ;
  assign n9522 = n2026 & ~n9521 ;
  assign n9523 = n2030 & ~n9522 ;
  assign n9524 = n2034 & ~n9523 ;
  assign n9525 = n2038 & ~n9524 ;
  assign n9526 = n2042 & ~n9525 ;
  assign n9527 = n2046 & ~n9526 ;
  assign n9528 = n2050 & ~n9527 ;
  assign n9529 = n2054 & ~n9528 ;
  assign n9530 = n2058 & ~n9529 ;
  assign n9531 = ~x171 & ~n2060 ;
  assign n9532 = ~n9530 & n9531 ;
  assign n9535 = ~n9532 & ~x299 ;
  assign n9536 = ~n9534 & ~n9535 ;
  assign n9537 = ~n374 & n1732 ;
  assign n9538 = n1737 & ~n9537 ;
  assign n9539 = n1741 & ~n9538 ;
  assign n9540 = n1745 & ~n9539 ;
  assign n9541 = n1749 & ~n9540 ;
  assign n9542 = n1753 & ~n9541 ;
  assign n9543 = n1757 & ~n9542 ;
  assign n9544 = n1761 & ~n9543 ;
  assign n9545 = n1765 & ~n9544 ;
  assign n9546 = n1769 & ~n9545 ;
  assign n9547 = n1773 & ~n9546 ;
  assign n9548 = n1777 & ~n9547 ;
  assign n9549 = n1781 & ~n9548 ;
  assign n9550 = n1785 & ~n9549 ;
  assign n9551 = n1789 & ~n9550 ;
  assign n9552 = n1793 & ~n9551 ;
  assign n9553 = n1797 & ~n9552 ;
  assign n9554 = n1801 & ~n9553 ;
  assign n9555 = n1805 & ~n9554 ;
  assign n9556 = n1809 & ~n9555 ;
  assign n9557 = n1813 & ~n9556 ;
  assign n9558 = n1817 & ~n9557 ;
  assign n9559 = n1821 & ~n9558 ;
  assign n9560 = n1825 & ~n9559 ;
  assign n9561 = n1829 & ~n9560 ;
  assign n9562 = n1833 & ~n9561 ;
  assign n9563 = n1837 & ~n9562 ;
  assign n9564 = n1841 & ~n9563 ;
  assign n9565 = n1845 & ~n9564 ;
  assign n9566 = n1849 & ~n9565 ;
  assign n9567 = n1853 & ~n9566 ;
  assign n9568 = n1857 & ~n9567 ;
  assign n9569 = n1861 & ~n9568 ;
  assign n9570 = n1865 & ~n9569 ;
  assign n9571 = n1869 & ~n9570 ;
  assign n9572 = n1873 & ~n9571 ;
  assign n9573 = n1877 & ~n9572 ;
  assign n9574 = n1881 & ~n9573 ;
  assign n9575 = n1885 & ~n9574 ;
  assign n9576 = n1889 & ~n9575 ;
  assign n9577 = n1893 & ~n9576 ;
  assign n9578 = n1897 & ~n9577 ;
  assign n9579 = n1901 & ~n9578 ;
  assign n9580 = n1905 & ~n9579 ;
  assign n9581 = n1909 & ~n9580 ;
  assign n9582 = n1913 & ~n9581 ;
  assign n9583 = n1917 & ~n9582 ;
  assign n9584 = n1921 & ~n9583 ;
  assign n9585 = n1925 & ~n9584 ;
  assign n9586 = n1929 & ~n9585 ;
  assign n9587 = n1933 & ~n9586 ;
  assign n9588 = n1937 & ~n9587 ;
  assign n9589 = n1941 & ~n9588 ;
  assign n9590 = n1945 & ~n9589 ;
  assign n9591 = n1949 & ~n9590 ;
  assign n9592 = n1953 & ~n9591 ;
  assign n9593 = n2749 & ~n9592 ;
  assign n9594 = n263 & ~n9593 ;
  assign n9595 = n267 & ~n9594 ;
  assign n9596 = n271 & ~n9595 ;
  assign n9597 = n275 & ~n9596 ;
  assign n9598 = n279 & ~n9597 ;
  assign n9599 = n283 & ~n9598 ;
  assign n9600 = n287 & ~n9599 ;
  assign n9601 = n291 & ~n9600 ;
  assign n9602 = n295 & ~n9601 ;
  assign n9603 = n299 & ~n9602 ;
  assign n9604 = n303 & ~n9603 ;
  assign n9605 = n307 & ~n9604 ;
  assign n9606 = n311 & ~n9605 ;
  assign n9607 = n315 & ~n9606 ;
  assign n9608 = n319 & ~n9607 ;
  assign n9609 = n323 & ~n9608 ;
  assign n9610 = n327 & ~n9609 ;
  assign n9611 = n331 & ~n9610 ;
  assign n9612 = n335 & ~n9611 ;
  assign n9613 = n339 & ~n9612 ;
  assign n9614 = n343 & ~n9613 ;
  assign n9615 = n347 & ~n9614 ;
  assign n9616 = n351 & ~n9615 ;
  assign n9617 = n355 & ~n9616 ;
  assign n9618 = n359 & ~n9617 ;
  assign n9619 = n363 & ~n9618 ;
  assign n9620 = n367 & ~n9619 ;
  assign n9621 = x172 & ~n369 ;
  assign n9622 = ~n9620 & n9621 ;
  assign n9710 = n9622 & x300 ;
  assign n9623 = ~n713 & n2069 ;
  assign n9624 = n2074 & ~n9623 ;
  assign n9625 = n2078 & ~n9624 ;
  assign n9626 = n2082 & ~n9625 ;
  assign n9627 = n2086 & ~n9626 ;
  assign n9628 = n2090 & ~n9627 ;
  assign n9629 = n2094 & ~n9628 ;
  assign n9630 = n2098 & ~n9629 ;
  assign n9631 = n2102 & ~n9630 ;
  assign n9632 = n2106 & ~n9631 ;
  assign n9633 = n2110 & ~n9632 ;
  assign n9634 = n2114 & ~n9633 ;
  assign n9635 = n2118 & ~n9634 ;
  assign n9636 = n2122 & ~n9635 ;
  assign n9637 = n2126 & ~n9636 ;
  assign n9638 = n2130 & ~n9637 ;
  assign n9639 = n2134 & ~n9638 ;
  assign n9640 = n2138 & ~n9639 ;
  assign n9641 = n2142 & ~n9640 ;
  assign n9642 = n2146 & ~n9641 ;
  assign n9643 = n2150 & ~n9642 ;
  assign n9644 = n2154 & ~n9643 ;
  assign n9645 = n2158 & ~n9644 ;
  assign n9646 = n2162 & ~n9645 ;
  assign n9647 = n2166 & ~n9646 ;
  assign n9648 = n2170 & ~n9647 ;
  assign n9649 = n2174 & ~n9648 ;
  assign n9650 = n2178 & ~n9649 ;
  assign n9651 = n2182 & ~n9650 ;
  assign n9652 = n2186 & ~n9651 ;
  assign n9653 = n2190 & ~n9652 ;
  assign n9654 = n2194 & ~n9653 ;
  assign n9655 = n2198 & ~n9654 ;
  assign n9656 = n2202 & ~n9655 ;
  assign n9657 = n2206 & ~n9656 ;
  assign n9658 = n2210 & ~n9657 ;
  assign n9659 = n2214 & ~n9658 ;
  assign n9660 = n2218 & ~n9659 ;
  assign n9661 = n2222 & ~n9660 ;
  assign n9662 = n2226 & ~n9661 ;
  assign n9663 = n2230 & ~n9662 ;
  assign n9664 = n2234 & ~n9663 ;
  assign n9665 = n2238 & ~n9664 ;
  assign n9666 = n2242 & ~n9665 ;
  assign n9667 = n2246 & ~n9666 ;
  assign n9668 = n2250 & ~n9667 ;
  assign n9669 = n2254 & ~n9668 ;
  assign n9670 = n2258 & ~n9669 ;
  assign n9671 = n2262 & ~n9670 ;
  assign n9672 = n2266 & ~n9671 ;
  assign n9673 = n2270 & ~n9672 ;
  assign n9674 = n2274 & ~n9673 ;
  assign n9675 = n2278 & ~n9674 ;
  assign n9676 = n2282 & ~n9675 ;
  assign n9677 = n2286 & ~n9676 ;
  assign n9678 = n2290 & ~n9677 ;
  assign n9679 = n2836 & ~n9678 ;
  assign n9680 = n602 & ~n9679 ;
  assign n9681 = n606 & ~n9680 ;
  assign n9682 = n610 & ~n9681 ;
  assign n9683 = n614 & ~n9682 ;
  assign n9684 = n618 & ~n9683 ;
  assign n9685 = n622 & ~n9684 ;
  assign n9686 = n626 & ~n9685 ;
  assign n9687 = n630 & ~n9686 ;
  assign n9688 = n634 & ~n9687 ;
  assign n9689 = n638 & ~n9688 ;
  assign n9690 = n642 & ~n9689 ;
  assign n9691 = n646 & ~n9690 ;
  assign n9692 = n650 & ~n9691 ;
  assign n9693 = n654 & ~n9692 ;
  assign n9694 = n658 & ~n9693 ;
  assign n9695 = n662 & ~n9694 ;
  assign n9696 = n666 & ~n9695 ;
  assign n9697 = n670 & ~n9696 ;
  assign n9698 = n674 & ~n9697 ;
  assign n9699 = n678 & ~n9698 ;
  assign n9700 = n682 & ~n9699 ;
  assign n9701 = n686 & ~n9700 ;
  assign n9702 = n690 & ~n9701 ;
  assign n9703 = n694 & ~n9702 ;
  assign n9704 = n698 & ~n9703 ;
  assign n9705 = n702 & ~n9704 ;
  assign n9706 = n706 & ~n9705 ;
  assign n9707 = ~x172 & ~n708 ;
  assign n9708 = ~n9706 & n9707 ;
  assign n9711 = ~n9708 & ~x300 ;
  assign n9712 = ~n9710 & ~n9711 ;
  assign n9713 = n378 & ~n1056 ;
  assign n9714 = n383 & ~n9713 ;
  assign n9715 = n387 & ~n9714 ;
  assign n9716 = n391 & ~n9715 ;
  assign n9717 = n395 & ~n9716 ;
  assign n9718 = n399 & ~n9717 ;
  assign n9719 = n403 & ~n9718 ;
  assign n9720 = n407 & ~n9719 ;
  assign n9721 = n411 & ~n9720 ;
  assign n9722 = n415 & ~n9721 ;
  assign n9723 = n419 & ~n9722 ;
  assign n9724 = n423 & ~n9723 ;
  assign n9725 = n427 & ~n9724 ;
  assign n9726 = n431 & ~n9725 ;
  assign n9727 = n435 & ~n9726 ;
  assign n9728 = n439 & ~n9727 ;
  assign n9729 = n443 & ~n9728 ;
  assign n9730 = n447 & ~n9729 ;
  assign n9731 = n451 & ~n9730 ;
  assign n9732 = n455 & ~n9731 ;
  assign n9733 = n459 & ~n9732 ;
  assign n9734 = n463 & ~n9733 ;
  assign n9735 = n467 & ~n9734 ;
  assign n9736 = n471 & ~n9735 ;
  assign n9737 = n475 & ~n9736 ;
  assign n9738 = n479 & ~n9737 ;
  assign n9739 = n483 & ~n9738 ;
  assign n9740 = n487 & ~n9739 ;
  assign n9741 = n491 & ~n9740 ;
  assign n9742 = n495 & ~n9741 ;
  assign n9743 = n499 & ~n9742 ;
  assign n9744 = n503 & ~n9743 ;
  assign n9745 = n507 & ~n9744 ;
  assign n9746 = n511 & ~n9745 ;
  assign n9747 = n515 & ~n9746 ;
  assign n9748 = n519 & ~n9747 ;
  assign n9749 = n523 & ~n9748 ;
  assign n9750 = n527 & ~n9749 ;
  assign n9751 = n531 & ~n9750 ;
  assign n9752 = n535 & ~n9751 ;
  assign n9753 = n539 & ~n9752 ;
  assign n9754 = n543 & ~n9753 ;
  assign n9755 = n547 & ~n9754 ;
  assign n9756 = n551 & ~n9755 ;
  assign n9757 = n555 & ~n9756 ;
  assign n9758 = n559 & ~n9757 ;
  assign n9759 = n563 & ~n9758 ;
  assign n9760 = n567 & ~n9759 ;
  assign n9761 = n571 & ~n9760 ;
  assign n9762 = n575 & ~n9761 ;
  assign n9763 = n579 & ~n9762 ;
  assign n9764 = n583 & ~n9763 ;
  assign n9765 = n587 & ~n9764 ;
  assign n9766 = n591 & ~n9765 ;
  assign n9767 = n2382 & ~n9766 ;
  assign n9768 = n2384 & ~n9767 ;
  assign n9769 = n2927 & ~n9768 ;
  assign n9770 = n945 & ~n9769 ;
  assign n9771 = n949 & ~n9770 ;
  assign n9772 = n953 & ~n9771 ;
  assign n9773 = n957 & ~n9772 ;
  assign n9774 = n961 & ~n9773 ;
  assign n9775 = n965 & ~n9774 ;
  assign n9776 = n969 & ~n9775 ;
  assign n9777 = n973 & ~n9776 ;
  assign n9778 = n977 & ~n9777 ;
  assign n9779 = n981 & ~n9778 ;
  assign n9780 = n985 & ~n9779 ;
  assign n9781 = n989 & ~n9780 ;
  assign n9782 = n993 & ~n9781 ;
  assign n9783 = n997 & ~n9782 ;
  assign n9784 = n1001 & ~n9783 ;
  assign n9785 = n1005 & ~n9784 ;
  assign n9786 = n1009 & ~n9785 ;
  assign n9787 = n1013 & ~n9786 ;
  assign n9788 = n1017 & ~n9787 ;
  assign n9789 = n1021 & ~n9788 ;
  assign n9790 = n1025 & ~n9789 ;
  assign n9791 = n1029 & ~n9790 ;
  assign n9792 = n1033 & ~n9791 ;
  assign n9793 = n1037 & ~n9792 ;
  assign n9794 = n1041 & ~n9793 ;
  assign n9795 = n1045 & ~n9794 ;
  assign n9796 = n1049 & ~n9795 ;
  assign n9797 = x173 & ~n1051 ;
  assign n9798 = ~n9796 & n9797 ;
  assign n9886 = n9798 & x301 ;
  assign n9799 = n717 & ~n1395 ;
  assign n9800 = n722 & ~n9799 ;
  assign n9801 = n726 & ~n9800 ;
  assign n9802 = n730 & ~n9801 ;
  assign n9803 = n734 & ~n9802 ;
  assign n9804 = n738 & ~n9803 ;
  assign n9805 = n742 & ~n9804 ;
  assign n9806 = n746 & ~n9805 ;
  assign n9807 = n750 & ~n9806 ;
  assign n9808 = n754 & ~n9807 ;
  assign n9809 = n758 & ~n9808 ;
  assign n9810 = n762 & ~n9809 ;
  assign n9811 = n766 & ~n9810 ;
  assign n9812 = n770 & ~n9811 ;
  assign n9813 = n774 & ~n9812 ;
  assign n9814 = n778 & ~n9813 ;
  assign n9815 = n782 & ~n9814 ;
  assign n9816 = n786 & ~n9815 ;
  assign n9817 = n790 & ~n9816 ;
  assign n9818 = n794 & ~n9817 ;
  assign n9819 = n798 & ~n9818 ;
  assign n9820 = n802 & ~n9819 ;
  assign n9821 = n806 & ~n9820 ;
  assign n9822 = n810 & ~n9821 ;
  assign n9823 = n814 & ~n9822 ;
  assign n9824 = n818 & ~n9823 ;
  assign n9825 = n822 & ~n9824 ;
  assign n9826 = n826 & ~n9825 ;
  assign n9827 = n830 & ~n9826 ;
  assign n9828 = n834 & ~n9827 ;
  assign n9829 = n838 & ~n9828 ;
  assign n9830 = n842 & ~n9829 ;
  assign n9831 = n846 & ~n9830 ;
  assign n9832 = n850 & ~n9831 ;
  assign n9833 = n854 & ~n9832 ;
  assign n9834 = n858 & ~n9833 ;
  assign n9835 = n862 & ~n9834 ;
  assign n9836 = n866 & ~n9835 ;
  assign n9837 = n870 & ~n9836 ;
  assign n9838 = n874 & ~n9837 ;
  assign n9839 = n878 & ~n9838 ;
  assign n9840 = n882 & ~n9839 ;
  assign n9841 = n886 & ~n9840 ;
  assign n9842 = n890 & ~n9841 ;
  assign n9843 = n894 & ~n9842 ;
  assign n9844 = n898 & ~n9843 ;
  assign n9845 = n902 & ~n9844 ;
  assign n9846 = n906 & ~n9845 ;
  assign n9847 = n910 & ~n9846 ;
  assign n9848 = n914 & ~n9847 ;
  assign n9849 = n918 & ~n9848 ;
  assign n9850 = n922 & ~n9849 ;
  assign n9851 = n926 & ~n9850 ;
  assign n9852 = n930 & ~n9851 ;
  assign n9853 = n2472 & ~n9852 ;
  assign n9854 = n2474 & ~n9853 ;
  assign n9855 = n3014 & ~n9854 ;
  assign n9856 = n1284 & ~n9855 ;
  assign n9857 = n1288 & ~n9856 ;
  assign n9858 = n1292 & ~n9857 ;
  assign n9859 = n1296 & ~n9858 ;
  assign n9860 = n1300 & ~n9859 ;
  assign n9861 = n1304 & ~n9860 ;
  assign n9862 = n1308 & ~n9861 ;
  assign n9863 = n1312 & ~n9862 ;
  assign n9864 = n1316 & ~n9863 ;
  assign n9865 = n1320 & ~n9864 ;
  assign n9866 = n1324 & ~n9865 ;
  assign n9867 = n1328 & ~n9866 ;
  assign n9868 = n1332 & ~n9867 ;
  assign n9869 = n1336 & ~n9868 ;
  assign n9870 = n1340 & ~n9869 ;
  assign n9871 = n1344 & ~n9870 ;
  assign n9872 = n1348 & ~n9871 ;
  assign n9873 = n1352 & ~n9872 ;
  assign n9874 = n1356 & ~n9873 ;
  assign n9875 = n1360 & ~n9874 ;
  assign n9876 = n1364 & ~n9875 ;
  assign n9877 = n1368 & ~n9876 ;
  assign n9878 = n1372 & ~n9877 ;
  assign n9879 = n1376 & ~n9878 ;
  assign n9880 = n1380 & ~n9879 ;
  assign n9881 = n1384 & ~n9880 ;
  assign n9882 = n1388 & ~n9881 ;
  assign n9883 = ~x173 & ~n1390 ;
  assign n9884 = ~n9882 & n9883 ;
  assign n9887 = ~n9884 & ~x301 ;
  assign n9888 = ~n9886 & ~n9887 ;
  assign n9889 = n1060 & ~n1736 ;
  assign n9890 = n1065 & ~n9889 ;
  assign n9891 = n1069 & ~n9890 ;
  assign n9892 = n1073 & ~n9891 ;
  assign n9893 = n1077 & ~n9892 ;
  assign n9894 = n1081 & ~n9893 ;
  assign n9895 = n1085 & ~n9894 ;
  assign n9896 = n1089 & ~n9895 ;
  assign n9897 = n1093 & ~n9896 ;
  assign n9898 = n1097 & ~n9897 ;
  assign n9899 = n1101 & ~n9898 ;
  assign n9900 = n1105 & ~n9899 ;
  assign n9901 = n1109 & ~n9900 ;
  assign n9902 = n1113 & ~n9901 ;
  assign n9903 = n1117 & ~n9902 ;
  assign n9904 = n1121 & ~n9903 ;
  assign n9905 = n1125 & ~n9904 ;
  assign n9906 = n1129 & ~n9905 ;
  assign n9907 = n1133 & ~n9906 ;
  assign n9908 = n1137 & ~n9907 ;
  assign n9909 = n1141 & ~n9908 ;
  assign n9910 = n1145 & ~n9909 ;
  assign n9911 = n1149 & ~n9910 ;
  assign n9912 = n1153 & ~n9911 ;
  assign n9913 = n1157 & ~n9912 ;
  assign n9914 = n1161 & ~n9913 ;
  assign n9915 = n1165 & ~n9914 ;
  assign n9916 = n1169 & ~n9915 ;
  assign n9917 = n1173 & ~n9916 ;
  assign n9918 = n1177 & ~n9917 ;
  assign n9919 = n1181 & ~n9918 ;
  assign n9920 = n1185 & ~n9919 ;
  assign n9921 = n1189 & ~n9920 ;
  assign n9922 = n1193 & ~n9921 ;
  assign n9923 = n1197 & ~n9922 ;
  assign n9924 = n1201 & ~n9923 ;
  assign n9925 = n1205 & ~n9924 ;
  assign n9926 = n1209 & ~n9925 ;
  assign n9927 = n1213 & ~n9926 ;
  assign n9928 = n1217 & ~n9927 ;
  assign n9929 = n1221 & ~n9928 ;
  assign n9930 = n1225 & ~n9929 ;
  assign n9931 = n1229 & ~n9930 ;
  assign n9932 = n1233 & ~n9931 ;
  assign n9933 = n1237 & ~n9932 ;
  assign n9934 = n1241 & ~n9933 ;
  assign n9935 = n1245 & ~n9934 ;
  assign n9936 = n1249 & ~n9935 ;
  assign n9937 = n1253 & ~n9936 ;
  assign n9938 = n1257 & ~n9937 ;
  assign n9939 = n1261 & ~n9938 ;
  assign n9940 = n1265 & ~n9939 ;
  assign n9941 = n1269 & ~n9940 ;
  assign n9942 = n1273 & ~n9941 ;
  assign n9943 = n2566 & ~n9942 ;
  assign n9944 = n2568 & ~n9943 ;
  assign n9945 = n3105 & ~n9944 ;
  assign n9946 = n1625 & ~n9945 ;
  assign n9947 = n1629 & ~n9946 ;
  assign n9948 = n1633 & ~n9947 ;
  assign n9949 = n1637 & ~n9948 ;
  assign n9950 = n1641 & ~n9949 ;
  assign n9951 = n1645 & ~n9950 ;
  assign n9952 = n1649 & ~n9951 ;
  assign n9953 = n1653 & ~n9952 ;
  assign n9954 = n1657 & ~n9953 ;
  assign n9955 = n1661 & ~n9954 ;
  assign n9956 = n1665 & ~n9955 ;
  assign n9957 = n1669 & ~n9956 ;
  assign n9958 = n1673 & ~n9957 ;
  assign n9959 = n1677 & ~n9958 ;
  assign n9960 = n1681 & ~n9959 ;
  assign n9961 = n1685 & ~n9960 ;
  assign n9962 = n1689 & ~n9961 ;
  assign n9963 = n1693 & ~n9962 ;
  assign n9964 = n1697 & ~n9963 ;
  assign n9965 = n1701 & ~n9964 ;
  assign n9966 = n1705 & ~n9965 ;
  assign n9967 = n1709 & ~n9966 ;
  assign n9968 = n1713 & ~n9967 ;
  assign n9969 = n1717 & ~n9968 ;
  assign n9970 = n1721 & ~n9969 ;
  assign n9971 = n1725 & ~n9970 ;
  assign n9972 = n1729 & ~n9971 ;
  assign n9973 = x174 & ~n1731 ;
  assign n9974 = ~n9972 & n9973 ;
  assign n10062 = n9974 & x302 ;
  assign n9975 = n1399 & ~n2073 ;
  assign n9976 = n1404 & ~n9975 ;
  assign n9977 = n1408 & ~n9976 ;
  assign n9978 = n1412 & ~n9977 ;
  assign n9979 = n1416 & ~n9978 ;
  assign n9980 = n1420 & ~n9979 ;
  assign n9981 = n1424 & ~n9980 ;
  assign n9982 = n1428 & ~n9981 ;
  assign n9983 = n1432 & ~n9982 ;
  assign n9984 = n1436 & ~n9983 ;
  assign n9985 = n1440 & ~n9984 ;
  assign n9986 = n1444 & ~n9985 ;
  assign n9987 = n1448 & ~n9986 ;
  assign n9988 = n1452 & ~n9987 ;
  assign n9989 = n1456 & ~n9988 ;
  assign n9990 = n1460 & ~n9989 ;
  assign n9991 = n1464 & ~n9990 ;
  assign n9992 = n1468 & ~n9991 ;
  assign n9993 = n1472 & ~n9992 ;
  assign n9994 = n1476 & ~n9993 ;
  assign n9995 = n1480 & ~n9994 ;
  assign n9996 = n1484 & ~n9995 ;
  assign n9997 = n1488 & ~n9996 ;
  assign n9998 = n1492 & ~n9997 ;
  assign n9999 = n1496 & ~n9998 ;
  assign n10000 = n1500 & ~n9999 ;
  assign n10001 = n1504 & ~n10000 ;
  assign n10002 = n1508 & ~n10001 ;
  assign n10003 = n1512 & ~n10002 ;
  assign n10004 = n1516 & ~n10003 ;
  assign n10005 = n1520 & ~n10004 ;
  assign n10006 = n1524 & ~n10005 ;
  assign n10007 = n1528 & ~n10006 ;
  assign n10008 = n1532 & ~n10007 ;
  assign n10009 = n1536 & ~n10008 ;
  assign n10010 = n1540 & ~n10009 ;
  assign n10011 = n1544 & ~n10010 ;
  assign n10012 = n1548 & ~n10011 ;
  assign n10013 = n1552 & ~n10012 ;
  assign n10014 = n1556 & ~n10013 ;
  assign n10015 = n1560 & ~n10014 ;
  assign n10016 = n1564 & ~n10015 ;
  assign n10017 = n1568 & ~n10016 ;
  assign n10018 = n1572 & ~n10017 ;
  assign n10019 = n1576 & ~n10018 ;
  assign n10020 = n1580 & ~n10019 ;
  assign n10021 = n1584 & ~n10020 ;
  assign n10022 = n1588 & ~n10021 ;
  assign n10023 = n1592 & ~n10022 ;
  assign n10024 = n1596 & ~n10023 ;
  assign n10025 = n1600 & ~n10024 ;
  assign n10026 = n1604 & ~n10025 ;
  assign n10027 = n1608 & ~n10026 ;
  assign n10028 = n1612 & ~n10027 ;
  assign n10029 = n2656 & ~n10028 ;
  assign n10030 = n2658 & ~n10029 ;
  assign n10031 = n3192 & ~n10030 ;
  assign n10032 = n1962 & ~n10031 ;
  assign n10033 = n1966 & ~n10032 ;
  assign n10034 = n1970 & ~n10033 ;
  assign n10035 = n1974 & ~n10034 ;
  assign n10036 = n1978 & ~n10035 ;
  assign n10037 = n1982 & ~n10036 ;
  assign n10038 = n1986 & ~n10037 ;
  assign n10039 = n1990 & ~n10038 ;
  assign n10040 = n1994 & ~n10039 ;
  assign n10041 = n1998 & ~n10040 ;
  assign n10042 = n2002 & ~n10041 ;
  assign n10043 = n2006 & ~n10042 ;
  assign n10044 = n2010 & ~n10043 ;
  assign n10045 = n2014 & ~n10044 ;
  assign n10046 = n2018 & ~n10045 ;
  assign n10047 = n2022 & ~n10046 ;
  assign n10048 = n2026 & ~n10047 ;
  assign n10049 = n2030 & ~n10048 ;
  assign n10050 = n2034 & ~n10049 ;
  assign n10051 = n2038 & ~n10050 ;
  assign n10052 = n2042 & ~n10051 ;
  assign n10053 = n2046 & ~n10052 ;
  assign n10054 = n2050 & ~n10053 ;
  assign n10055 = n2054 & ~n10054 ;
  assign n10056 = n2058 & ~n10055 ;
  assign n10057 = n2062 & ~n10056 ;
  assign n10058 = n2066 & ~n10057 ;
  assign n10059 = ~x174 & ~n2068 ;
  assign n10060 = ~n10058 & n10059 ;
  assign n10063 = ~n10060 & ~x302 ;
  assign n10064 = ~n10062 & ~n10063 ;
  assign n10065 = ~n382 & n1740 ;
  assign n10066 = n1745 & ~n10065 ;
  assign n10067 = n1749 & ~n10066 ;
  assign n10068 = n1753 & ~n10067 ;
  assign n10069 = n1757 & ~n10068 ;
  assign n10070 = n1761 & ~n10069 ;
  assign n10071 = n1765 & ~n10070 ;
  assign n10072 = n1769 & ~n10071 ;
  assign n10073 = n1773 & ~n10072 ;
  assign n10074 = n1777 & ~n10073 ;
  assign n10075 = n1781 & ~n10074 ;
  assign n10076 = n1785 & ~n10075 ;
  assign n10077 = n1789 & ~n10076 ;
  assign n10078 = n1793 & ~n10077 ;
  assign n10079 = n1797 & ~n10078 ;
  assign n10080 = n1801 & ~n10079 ;
  assign n10081 = n1805 & ~n10080 ;
  assign n10082 = n1809 & ~n10081 ;
  assign n10083 = n1813 & ~n10082 ;
  assign n10084 = n1817 & ~n10083 ;
  assign n10085 = n1821 & ~n10084 ;
  assign n10086 = n1825 & ~n10085 ;
  assign n10087 = n1829 & ~n10086 ;
  assign n10088 = n1833 & ~n10087 ;
  assign n10089 = n1837 & ~n10088 ;
  assign n10090 = n1841 & ~n10089 ;
  assign n10091 = n1845 & ~n10090 ;
  assign n10092 = n1849 & ~n10091 ;
  assign n10093 = n1853 & ~n10092 ;
  assign n10094 = n1857 & ~n10093 ;
  assign n10095 = n1861 & ~n10094 ;
  assign n10096 = n1865 & ~n10095 ;
  assign n10097 = n1869 & ~n10096 ;
  assign n10098 = n1873 & ~n10097 ;
  assign n10099 = n1877 & ~n10098 ;
  assign n10100 = n1881 & ~n10099 ;
  assign n10101 = n1885 & ~n10100 ;
  assign n10102 = n1889 & ~n10101 ;
  assign n10103 = n1893 & ~n10102 ;
  assign n10104 = n1897 & ~n10103 ;
  assign n10105 = n1901 & ~n10104 ;
  assign n10106 = n1905 & ~n10105 ;
  assign n10107 = n1909 & ~n10106 ;
  assign n10108 = n1913 & ~n10107 ;
  assign n10109 = n1917 & ~n10108 ;
  assign n10110 = n1921 & ~n10109 ;
  assign n10111 = n1925 & ~n10110 ;
  assign n10112 = n1929 & ~n10111 ;
  assign n10113 = n1933 & ~n10112 ;
  assign n10114 = n1937 & ~n10113 ;
  assign n10115 = n1941 & ~n10114 ;
  assign n10116 = n1945 & ~n10115 ;
  assign n10117 = n1949 & ~n10116 ;
  assign n10118 = n1953 & ~n10117 ;
  assign n10119 = n2749 & ~n10118 ;
  assign n10120 = n263 & ~n10119 ;
  assign n10121 = n267 & ~n10120 ;
  assign n10122 = n271 & ~n10121 ;
  assign n10123 = n275 & ~n10122 ;
  assign n10124 = n279 & ~n10123 ;
  assign n10125 = n283 & ~n10124 ;
  assign n10126 = n287 & ~n10125 ;
  assign n10127 = n291 & ~n10126 ;
  assign n10128 = n295 & ~n10127 ;
  assign n10129 = n299 & ~n10128 ;
  assign n10130 = n303 & ~n10129 ;
  assign n10131 = n307 & ~n10130 ;
  assign n10132 = n311 & ~n10131 ;
  assign n10133 = n315 & ~n10132 ;
  assign n10134 = n319 & ~n10133 ;
  assign n10135 = n323 & ~n10134 ;
  assign n10136 = n327 & ~n10135 ;
  assign n10137 = n331 & ~n10136 ;
  assign n10138 = n335 & ~n10137 ;
  assign n10139 = n339 & ~n10138 ;
  assign n10140 = n343 & ~n10139 ;
  assign n10141 = n347 & ~n10140 ;
  assign n10142 = n351 & ~n10141 ;
  assign n10143 = n355 & ~n10142 ;
  assign n10144 = n359 & ~n10143 ;
  assign n10145 = n363 & ~n10144 ;
  assign n10146 = n367 & ~n10145 ;
  assign n10147 = n371 & ~n10146 ;
  assign n10148 = n375 & ~n10147 ;
  assign n10149 = x175 & ~n377 ;
  assign n10150 = ~n10148 & n10149 ;
  assign n10238 = n10150 & x303 ;
  assign n10151 = ~n721 & n2077 ;
  assign n10152 = n2082 & ~n10151 ;
  assign n10153 = n2086 & ~n10152 ;
  assign n10154 = n2090 & ~n10153 ;
  assign n10155 = n2094 & ~n10154 ;
  assign n10156 = n2098 & ~n10155 ;
  assign n10157 = n2102 & ~n10156 ;
  assign n10158 = n2106 & ~n10157 ;
  assign n10159 = n2110 & ~n10158 ;
  assign n10160 = n2114 & ~n10159 ;
  assign n10161 = n2118 & ~n10160 ;
  assign n10162 = n2122 & ~n10161 ;
  assign n10163 = n2126 & ~n10162 ;
  assign n10164 = n2130 & ~n10163 ;
  assign n10165 = n2134 & ~n10164 ;
  assign n10166 = n2138 & ~n10165 ;
  assign n10167 = n2142 & ~n10166 ;
  assign n10168 = n2146 & ~n10167 ;
  assign n10169 = n2150 & ~n10168 ;
  assign n10170 = n2154 & ~n10169 ;
  assign n10171 = n2158 & ~n10170 ;
  assign n10172 = n2162 & ~n10171 ;
  assign n10173 = n2166 & ~n10172 ;
  assign n10174 = n2170 & ~n10173 ;
  assign n10175 = n2174 & ~n10174 ;
  assign n10176 = n2178 & ~n10175 ;
  assign n10177 = n2182 & ~n10176 ;
  assign n10178 = n2186 & ~n10177 ;
  assign n10179 = n2190 & ~n10178 ;
  assign n10180 = n2194 & ~n10179 ;
  assign n10181 = n2198 & ~n10180 ;
  assign n10182 = n2202 & ~n10181 ;
  assign n10183 = n2206 & ~n10182 ;
  assign n10184 = n2210 & ~n10183 ;
  assign n10185 = n2214 & ~n10184 ;
  assign n10186 = n2218 & ~n10185 ;
  assign n10187 = n2222 & ~n10186 ;
  assign n10188 = n2226 & ~n10187 ;
  assign n10189 = n2230 & ~n10188 ;
  assign n10190 = n2234 & ~n10189 ;
  assign n10191 = n2238 & ~n10190 ;
  assign n10192 = n2242 & ~n10191 ;
  assign n10193 = n2246 & ~n10192 ;
  assign n10194 = n2250 & ~n10193 ;
  assign n10195 = n2254 & ~n10194 ;
  assign n10196 = n2258 & ~n10195 ;
  assign n10197 = n2262 & ~n10196 ;
  assign n10198 = n2266 & ~n10197 ;
  assign n10199 = n2270 & ~n10198 ;
  assign n10200 = n2274 & ~n10199 ;
  assign n10201 = n2278 & ~n10200 ;
  assign n10202 = n2282 & ~n10201 ;
  assign n10203 = n2286 & ~n10202 ;
  assign n10204 = n2290 & ~n10203 ;
  assign n10205 = n2836 & ~n10204 ;
  assign n10206 = n602 & ~n10205 ;
  assign n10207 = n606 & ~n10206 ;
  assign n10208 = n610 & ~n10207 ;
  assign n10209 = n614 & ~n10208 ;
  assign n10210 = n618 & ~n10209 ;
  assign n10211 = n622 & ~n10210 ;
  assign n10212 = n626 & ~n10211 ;
  assign n10213 = n630 & ~n10212 ;
  assign n10214 = n634 & ~n10213 ;
  assign n10215 = n638 & ~n10214 ;
  assign n10216 = n642 & ~n10215 ;
  assign n10217 = n646 & ~n10216 ;
  assign n10218 = n650 & ~n10217 ;
  assign n10219 = n654 & ~n10218 ;
  assign n10220 = n658 & ~n10219 ;
  assign n10221 = n662 & ~n10220 ;
  assign n10222 = n666 & ~n10221 ;
  assign n10223 = n670 & ~n10222 ;
  assign n10224 = n674 & ~n10223 ;
  assign n10225 = n678 & ~n10224 ;
  assign n10226 = n682 & ~n10225 ;
  assign n10227 = n686 & ~n10226 ;
  assign n10228 = n690 & ~n10227 ;
  assign n10229 = n694 & ~n10228 ;
  assign n10230 = n698 & ~n10229 ;
  assign n10231 = n702 & ~n10230 ;
  assign n10232 = n706 & ~n10231 ;
  assign n10233 = n710 & ~n10232 ;
  assign n10234 = n714 & ~n10233 ;
  assign n10235 = ~x175 & ~n716 ;
  assign n10236 = ~n10234 & n10235 ;
  assign n10239 = ~n10236 & ~x303 ;
  assign n10240 = ~n10238 & ~n10239 ;
  assign n10241 = n386 & ~n1064 ;
  assign n10242 = n391 & ~n10241 ;
  assign n10243 = n395 & ~n10242 ;
  assign n10244 = n399 & ~n10243 ;
  assign n10245 = n403 & ~n10244 ;
  assign n10246 = n407 & ~n10245 ;
  assign n10247 = n411 & ~n10246 ;
  assign n10248 = n415 & ~n10247 ;
  assign n10249 = n419 & ~n10248 ;
  assign n10250 = n423 & ~n10249 ;
  assign n10251 = n427 & ~n10250 ;
  assign n10252 = n431 & ~n10251 ;
  assign n10253 = n435 & ~n10252 ;
  assign n10254 = n439 & ~n10253 ;
  assign n10255 = n443 & ~n10254 ;
  assign n10256 = n447 & ~n10255 ;
  assign n10257 = n451 & ~n10256 ;
  assign n10258 = n455 & ~n10257 ;
  assign n10259 = n459 & ~n10258 ;
  assign n10260 = n463 & ~n10259 ;
  assign n10261 = n467 & ~n10260 ;
  assign n10262 = n471 & ~n10261 ;
  assign n10263 = n475 & ~n10262 ;
  assign n10264 = n479 & ~n10263 ;
  assign n10265 = n483 & ~n10264 ;
  assign n10266 = n487 & ~n10265 ;
  assign n10267 = n491 & ~n10266 ;
  assign n10268 = n495 & ~n10267 ;
  assign n10269 = n499 & ~n10268 ;
  assign n10270 = n503 & ~n10269 ;
  assign n10271 = n507 & ~n10270 ;
  assign n10272 = n511 & ~n10271 ;
  assign n10273 = n515 & ~n10272 ;
  assign n10274 = n519 & ~n10273 ;
  assign n10275 = n523 & ~n10274 ;
  assign n10276 = n527 & ~n10275 ;
  assign n10277 = n531 & ~n10276 ;
  assign n10278 = n535 & ~n10277 ;
  assign n10279 = n539 & ~n10278 ;
  assign n10280 = n543 & ~n10279 ;
  assign n10281 = n547 & ~n10280 ;
  assign n10282 = n551 & ~n10281 ;
  assign n10283 = n555 & ~n10282 ;
  assign n10284 = n559 & ~n10283 ;
  assign n10285 = n563 & ~n10284 ;
  assign n10286 = n567 & ~n10285 ;
  assign n10287 = n571 & ~n10286 ;
  assign n10288 = n575 & ~n10287 ;
  assign n10289 = n579 & ~n10288 ;
  assign n10290 = n583 & ~n10289 ;
  assign n10291 = n587 & ~n10290 ;
  assign n10292 = n591 & ~n10291 ;
  assign n10293 = n2382 & ~n10292 ;
  assign n10294 = n2384 & ~n10293 ;
  assign n10295 = n2927 & ~n10294 ;
  assign n10296 = n945 & ~n10295 ;
  assign n10297 = n949 & ~n10296 ;
  assign n10298 = n953 & ~n10297 ;
  assign n10299 = n957 & ~n10298 ;
  assign n10300 = n961 & ~n10299 ;
  assign n10301 = n965 & ~n10300 ;
  assign n10302 = n969 & ~n10301 ;
  assign n10303 = n973 & ~n10302 ;
  assign n10304 = n977 & ~n10303 ;
  assign n10305 = n981 & ~n10304 ;
  assign n10306 = n985 & ~n10305 ;
  assign n10307 = n989 & ~n10306 ;
  assign n10308 = n993 & ~n10307 ;
  assign n10309 = n997 & ~n10308 ;
  assign n10310 = n1001 & ~n10309 ;
  assign n10311 = n1005 & ~n10310 ;
  assign n10312 = n1009 & ~n10311 ;
  assign n10313 = n1013 & ~n10312 ;
  assign n10314 = n1017 & ~n10313 ;
  assign n10315 = n1021 & ~n10314 ;
  assign n10316 = n1025 & ~n10315 ;
  assign n10317 = n1029 & ~n10316 ;
  assign n10318 = n1033 & ~n10317 ;
  assign n10319 = n1037 & ~n10318 ;
  assign n10320 = n1041 & ~n10319 ;
  assign n10321 = n1045 & ~n10320 ;
  assign n10322 = n1049 & ~n10321 ;
  assign n10323 = n1053 & ~n10322 ;
  assign n10324 = n1057 & ~n10323 ;
  assign n10325 = x176 & ~n1059 ;
  assign n10326 = ~n10324 & n10325 ;
  assign n10414 = n10326 & x304 ;
  assign n10327 = n725 & ~n1403 ;
  assign n10328 = n730 & ~n10327 ;
  assign n10329 = n734 & ~n10328 ;
  assign n10330 = n738 & ~n10329 ;
  assign n10331 = n742 & ~n10330 ;
  assign n10332 = n746 & ~n10331 ;
  assign n10333 = n750 & ~n10332 ;
  assign n10334 = n754 & ~n10333 ;
  assign n10335 = n758 & ~n10334 ;
  assign n10336 = n762 & ~n10335 ;
  assign n10337 = n766 & ~n10336 ;
  assign n10338 = n770 & ~n10337 ;
  assign n10339 = n774 & ~n10338 ;
  assign n10340 = n778 & ~n10339 ;
  assign n10341 = n782 & ~n10340 ;
  assign n10342 = n786 & ~n10341 ;
  assign n10343 = n790 & ~n10342 ;
  assign n10344 = n794 & ~n10343 ;
  assign n10345 = n798 & ~n10344 ;
  assign n10346 = n802 & ~n10345 ;
  assign n10347 = n806 & ~n10346 ;
  assign n10348 = n810 & ~n10347 ;
  assign n10349 = n814 & ~n10348 ;
  assign n10350 = n818 & ~n10349 ;
  assign n10351 = n822 & ~n10350 ;
  assign n10352 = n826 & ~n10351 ;
  assign n10353 = n830 & ~n10352 ;
  assign n10354 = n834 & ~n10353 ;
  assign n10355 = n838 & ~n10354 ;
  assign n10356 = n842 & ~n10355 ;
  assign n10357 = n846 & ~n10356 ;
  assign n10358 = n850 & ~n10357 ;
  assign n10359 = n854 & ~n10358 ;
  assign n10360 = n858 & ~n10359 ;
  assign n10361 = n862 & ~n10360 ;
  assign n10362 = n866 & ~n10361 ;
  assign n10363 = n870 & ~n10362 ;
  assign n10364 = n874 & ~n10363 ;
  assign n10365 = n878 & ~n10364 ;
  assign n10366 = n882 & ~n10365 ;
  assign n10367 = n886 & ~n10366 ;
  assign n10368 = n890 & ~n10367 ;
  assign n10369 = n894 & ~n10368 ;
  assign n10370 = n898 & ~n10369 ;
  assign n10371 = n902 & ~n10370 ;
  assign n10372 = n906 & ~n10371 ;
  assign n10373 = n910 & ~n10372 ;
  assign n10374 = n914 & ~n10373 ;
  assign n10375 = n918 & ~n10374 ;
  assign n10376 = n922 & ~n10375 ;
  assign n10377 = n926 & ~n10376 ;
  assign n10378 = n930 & ~n10377 ;
  assign n10379 = n2472 & ~n10378 ;
  assign n10380 = n2474 & ~n10379 ;
  assign n10381 = n3014 & ~n10380 ;
  assign n10382 = n1284 & ~n10381 ;
  assign n10383 = n1288 & ~n10382 ;
  assign n10384 = n1292 & ~n10383 ;
  assign n10385 = n1296 & ~n10384 ;
  assign n10386 = n1300 & ~n10385 ;
  assign n10387 = n1304 & ~n10386 ;
  assign n10388 = n1308 & ~n10387 ;
  assign n10389 = n1312 & ~n10388 ;
  assign n10390 = n1316 & ~n10389 ;
  assign n10391 = n1320 & ~n10390 ;
  assign n10392 = n1324 & ~n10391 ;
  assign n10393 = n1328 & ~n10392 ;
  assign n10394 = n1332 & ~n10393 ;
  assign n10395 = n1336 & ~n10394 ;
  assign n10396 = n1340 & ~n10395 ;
  assign n10397 = n1344 & ~n10396 ;
  assign n10398 = n1348 & ~n10397 ;
  assign n10399 = n1352 & ~n10398 ;
  assign n10400 = n1356 & ~n10399 ;
  assign n10401 = n1360 & ~n10400 ;
  assign n10402 = n1364 & ~n10401 ;
  assign n10403 = n1368 & ~n10402 ;
  assign n10404 = n1372 & ~n10403 ;
  assign n10405 = n1376 & ~n10404 ;
  assign n10406 = n1380 & ~n10405 ;
  assign n10407 = n1384 & ~n10406 ;
  assign n10408 = n1388 & ~n10407 ;
  assign n10409 = n1392 & ~n10408 ;
  assign n10410 = n1396 & ~n10409 ;
  assign n10411 = ~x176 & ~n1398 ;
  assign n10412 = ~n10410 & n10411 ;
  assign n10415 = ~n10412 & ~x304 ;
  assign n10416 = ~n10414 & ~n10415 ;
  assign n10417 = n1068 & ~n1744 ;
  assign n10418 = n1073 & ~n10417 ;
  assign n10419 = n1077 & ~n10418 ;
  assign n10420 = n1081 & ~n10419 ;
  assign n10421 = n1085 & ~n10420 ;
  assign n10422 = n1089 & ~n10421 ;
  assign n10423 = n1093 & ~n10422 ;
  assign n10424 = n1097 & ~n10423 ;
  assign n10425 = n1101 & ~n10424 ;
  assign n10426 = n1105 & ~n10425 ;
  assign n10427 = n1109 & ~n10426 ;
  assign n10428 = n1113 & ~n10427 ;
  assign n10429 = n1117 & ~n10428 ;
  assign n10430 = n1121 & ~n10429 ;
  assign n10431 = n1125 & ~n10430 ;
  assign n10432 = n1129 & ~n10431 ;
  assign n10433 = n1133 & ~n10432 ;
  assign n10434 = n1137 & ~n10433 ;
  assign n10435 = n1141 & ~n10434 ;
  assign n10436 = n1145 & ~n10435 ;
  assign n10437 = n1149 & ~n10436 ;
  assign n10438 = n1153 & ~n10437 ;
  assign n10439 = n1157 & ~n10438 ;
  assign n10440 = n1161 & ~n10439 ;
  assign n10441 = n1165 & ~n10440 ;
  assign n10442 = n1169 & ~n10441 ;
  assign n10443 = n1173 & ~n10442 ;
  assign n10444 = n1177 & ~n10443 ;
  assign n10445 = n1181 & ~n10444 ;
  assign n10446 = n1185 & ~n10445 ;
  assign n10447 = n1189 & ~n10446 ;
  assign n10448 = n1193 & ~n10447 ;
  assign n10449 = n1197 & ~n10448 ;
  assign n10450 = n1201 & ~n10449 ;
  assign n10451 = n1205 & ~n10450 ;
  assign n10452 = n1209 & ~n10451 ;
  assign n10453 = n1213 & ~n10452 ;
  assign n10454 = n1217 & ~n10453 ;
  assign n10455 = n1221 & ~n10454 ;
  assign n10456 = n1225 & ~n10455 ;
  assign n10457 = n1229 & ~n10456 ;
  assign n10458 = n1233 & ~n10457 ;
  assign n10459 = n1237 & ~n10458 ;
  assign n10460 = n1241 & ~n10459 ;
  assign n10461 = n1245 & ~n10460 ;
  assign n10462 = n1249 & ~n10461 ;
  assign n10463 = n1253 & ~n10462 ;
  assign n10464 = n1257 & ~n10463 ;
  assign n10465 = n1261 & ~n10464 ;
  assign n10466 = n1265 & ~n10465 ;
  assign n10467 = n1269 & ~n10466 ;
  assign n10468 = n1273 & ~n10467 ;
  assign n10469 = n2566 & ~n10468 ;
  assign n10470 = n2568 & ~n10469 ;
  assign n10471 = n3105 & ~n10470 ;
  assign n10472 = n1625 & ~n10471 ;
  assign n10473 = n1629 & ~n10472 ;
  assign n10474 = n1633 & ~n10473 ;
  assign n10475 = n1637 & ~n10474 ;
  assign n10476 = n1641 & ~n10475 ;
  assign n10477 = n1645 & ~n10476 ;
  assign n10478 = n1649 & ~n10477 ;
  assign n10479 = n1653 & ~n10478 ;
  assign n10480 = n1657 & ~n10479 ;
  assign n10481 = n1661 & ~n10480 ;
  assign n10482 = n1665 & ~n10481 ;
  assign n10483 = n1669 & ~n10482 ;
  assign n10484 = n1673 & ~n10483 ;
  assign n10485 = n1677 & ~n10484 ;
  assign n10486 = n1681 & ~n10485 ;
  assign n10487 = n1685 & ~n10486 ;
  assign n10488 = n1689 & ~n10487 ;
  assign n10489 = n1693 & ~n10488 ;
  assign n10490 = n1697 & ~n10489 ;
  assign n10491 = n1701 & ~n10490 ;
  assign n10492 = n1705 & ~n10491 ;
  assign n10493 = n1709 & ~n10492 ;
  assign n10494 = n1713 & ~n10493 ;
  assign n10495 = n1717 & ~n10494 ;
  assign n10496 = n1721 & ~n10495 ;
  assign n10497 = n1725 & ~n10496 ;
  assign n10498 = n1729 & ~n10497 ;
  assign n10499 = n1733 & ~n10498 ;
  assign n10500 = n1737 & ~n10499 ;
  assign n10501 = x177 & ~n1739 ;
  assign n10502 = ~n10500 & n10501 ;
  assign n10590 = n10502 & x305 ;
  assign n10503 = n1407 & ~n2081 ;
  assign n10504 = n1412 & ~n10503 ;
  assign n10505 = n1416 & ~n10504 ;
  assign n10506 = n1420 & ~n10505 ;
  assign n10507 = n1424 & ~n10506 ;
  assign n10508 = n1428 & ~n10507 ;
  assign n10509 = n1432 & ~n10508 ;
  assign n10510 = n1436 & ~n10509 ;
  assign n10511 = n1440 & ~n10510 ;
  assign n10512 = n1444 & ~n10511 ;
  assign n10513 = n1448 & ~n10512 ;
  assign n10514 = n1452 & ~n10513 ;
  assign n10515 = n1456 & ~n10514 ;
  assign n10516 = n1460 & ~n10515 ;
  assign n10517 = n1464 & ~n10516 ;
  assign n10518 = n1468 & ~n10517 ;
  assign n10519 = n1472 & ~n10518 ;
  assign n10520 = n1476 & ~n10519 ;
  assign n10521 = n1480 & ~n10520 ;
  assign n10522 = n1484 & ~n10521 ;
  assign n10523 = n1488 & ~n10522 ;
  assign n10524 = n1492 & ~n10523 ;
  assign n10525 = n1496 & ~n10524 ;
  assign n10526 = n1500 & ~n10525 ;
  assign n10527 = n1504 & ~n10526 ;
  assign n10528 = n1508 & ~n10527 ;
  assign n10529 = n1512 & ~n10528 ;
  assign n10530 = n1516 & ~n10529 ;
  assign n10531 = n1520 & ~n10530 ;
  assign n10532 = n1524 & ~n10531 ;
  assign n10533 = n1528 & ~n10532 ;
  assign n10534 = n1532 & ~n10533 ;
  assign n10535 = n1536 & ~n10534 ;
  assign n10536 = n1540 & ~n10535 ;
  assign n10537 = n1544 & ~n10536 ;
  assign n10538 = n1548 & ~n10537 ;
  assign n10539 = n1552 & ~n10538 ;
  assign n10540 = n1556 & ~n10539 ;
  assign n10541 = n1560 & ~n10540 ;
  assign n10542 = n1564 & ~n10541 ;
  assign n10543 = n1568 & ~n10542 ;
  assign n10544 = n1572 & ~n10543 ;
  assign n10545 = n1576 & ~n10544 ;
  assign n10546 = n1580 & ~n10545 ;
  assign n10547 = n1584 & ~n10546 ;
  assign n10548 = n1588 & ~n10547 ;
  assign n10549 = n1592 & ~n10548 ;
  assign n10550 = n1596 & ~n10549 ;
  assign n10551 = n1600 & ~n10550 ;
  assign n10552 = n1604 & ~n10551 ;
  assign n10553 = n1608 & ~n10552 ;
  assign n10554 = n1612 & ~n10553 ;
  assign n10555 = n2656 & ~n10554 ;
  assign n10556 = n2658 & ~n10555 ;
  assign n10557 = n3192 & ~n10556 ;
  assign n10558 = n1962 & ~n10557 ;
  assign n10559 = n1966 & ~n10558 ;
  assign n10560 = n1970 & ~n10559 ;
  assign n10561 = n1974 & ~n10560 ;
  assign n10562 = n1978 & ~n10561 ;
  assign n10563 = n1982 & ~n10562 ;
  assign n10564 = n1986 & ~n10563 ;
  assign n10565 = n1990 & ~n10564 ;
  assign n10566 = n1994 & ~n10565 ;
  assign n10567 = n1998 & ~n10566 ;
  assign n10568 = n2002 & ~n10567 ;
  assign n10569 = n2006 & ~n10568 ;
  assign n10570 = n2010 & ~n10569 ;
  assign n10571 = n2014 & ~n10570 ;
  assign n10572 = n2018 & ~n10571 ;
  assign n10573 = n2022 & ~n10572 ;
  assign n10574 = n2026 & ~n10573 ;
  assign n10575 = n2030 & ~n10574 ;
  assign n10576 = n2034 & ~n10575 ;
  assign n10577 = n2038 & ~n10576 ;
  assign n10578 = n2042 & ~n10577 ;
  assign n10579 = n2046 & ~n10578 ;
  assign n10580 = n2050 & ~n10579 ;
  assign n10581 = n2054 & ~n10580 ;
  assign n10582 = n2058 & ~n10581 ;
  assign n10583 = n2062 & ~n10582 ;
  assign n10584 = n2066 & ~n10583 ;
  assign n10585 = n2070 & ~n10584 ;
  assign n10586 = n2074 & ~n10585 ;
  assign n10587 = ~x177 & ~n2076 ;
  assign n10588 = ~n10586 & n10587 ;
  assign n10591 = ~n10588 & ~x305 ;
  assign n10592 = ~n10590 & ~n10591 ;
  assign n10593 = ~n390 & n1748 ;
  assign n10594 = n1753 & ~n10593 ;
  assign n10595 = n1757 & ~n10594 ;
  assign n10596 = n1761 & ~n10595 ;
  assign n10597 = n1765 & ~n10596 ;
  assign n10598 = n1769 & ~n10597 ;
  assign n10599 = n1773 & ~n10598 ;
  assign n10600 = n1777 & ~n10599 ;
  assign n10601 = n1781 & ~n10600 ;
  assign n10602 = n1785 & ~n10601 ;
  assign n10603 = n1789 & ~n10602 ;
  assign n10604 = n1793 & ~n10603 ;
  assign n10605 = n1797 & ~n10604 ;
  assign n10606 = n1801 & ~n10605 ;
  assign n10607 = n1805 & ~n10606 ;
  assign n10608 = n1809 & ~n10607 ;
  assign n10609 = n1813 & ~n10608 ;
  assign n10610 = n1817 & ~n10609 ;
  assign n10611 = n1821 & ~n10610 ;
  assign n10612 = n1825 & ~n10611 ;
  assign n10613 = n1829 & ~n10612 ;
  assign n10614 = n1833 & ~n10613 ;
  assign n10615 = n1837 & ~n10614 ;
  assign n10616 = n1841 & ~n10615 ;
  assign n10617 = n1845 & ~n10616 ;
  assign n10618 = n1849 & ~n10617 ;
  assign n10619 = n1853 & ~n10618 ;
  assign n10620 = n1857 & ~n10619 ;
  assign n10621 = n1861 & ~n10620 ;
  assign n10622 = n1865 & ~n10621 ;
  assign n10623 = n1869 & ~n10622 ;
  assign n10624 = n1873 & ~n10623 ;
  assign n10625 = n1877 & ~n10624 ;
  assign n10626 = n1881 & ~n10625 ;
  assign n10627 = n1885 & ~n10626 ;
  assign n10628 = n1889 & ~n10627 ;
  assign n10629 = n1893 & ~n10628 ;
  assign n10630 = n1897 & ~n10629 ;
  assign n10631 = n1901 & ~n10630 ;
  assign n10632 = n1905 & ~n10631 ;
  assign n10633 = n1909 & ~n10632 ;
  assign n10634 = n1913 & ~n10633 ;
  assign n10635 = n1917 & ~n10634 ;
  assign n10636 = n1921 & ~n10635 ;
  assign n10637 = n1925 & ~n10636 ;
  assign n10638 = n1929 & ~n10637 ;
  assign n10639 = n1933 & ~n10638 ;
  assign n10640 = n1937 & ~n10639 ;
  assign n10641 = n1941 & ~n10640 ;
  assign n10642 = n1945 & ~n10641 ;
  assign n10643 = n1949 & ~n10642 ;
  assign n10644 = n1953 & ~n10643 ;
  assign n10645 = n2749 & ~n10644 ;
  assign n10646 = n263 & ~n10645 ;
  assign n10647 = n267 & ~n10646 ;
  assign n10648 = n271 & ~n10647 ;
  assign n10649 = n275 & ~n10648 ;
  assign n10650 = n279 & ~n10649 ;
  assign n10651 = n283 & ~n10650 ;
  assign n10652 = n287 & ~n10651 ;
  assign n10653 = n291 & ~n10652 ;
  assign n10654 = n295 & ~n10653 ;
  assign n10655 = n299 & ~n10654 ;
  assign n10656 = n303 & ~n10655 ;
  assign n10657 = n307 & ~n10656 ;
  assign n10658 = n311 & ~n10657 ;
  assign n10659 = n315 & ~n10658 ;
  assign n10660 = n319 & ~n10659 ;
  assign n10661 = n323 & ~n10660 ;
  assign n10662 = n327 & ~n10661 ;
  assign n10663 = n331 & ~n10662 ;
  assign n10664 = n335 & ~n10663 ;
  assign n10665 = n339 & ~n10664 ;
  assign n10666 = n343 & ~n10665 ;
  assign n10667 = n347 & ~n10666 ;
  assign n10668 = n351 & ~n10667 ;
  assign n10669 = n355 & ~n10668 ;
  assign n10670 = n359 & ~n10669 ;
  assign n10671 = n363 & ~n10670 ;
  assign n10672 = n367 & ~n10671 ;
  assign n10673 = n371 & ~n10672 ;
  assign n10674 = n375 & ~n10673 ;
  assign n10675 = n379 & ~n10674 ;
  assign n10676 = n383 & ~n10675 ;
  assign n10677 = x178 & ~n385 ;
  assign n10678 = ~n10676 & n10677 ;
  assign n10766 = n10678 & x306 ;
  assign n10679 = ~n729 & n2085 ;
  assign n10680 = n2090 & ~n10679 ;
  assign n10681 = n2094 & ~n10680 ;
  assign n10682 = n2098 & ~n10681 ;
  assign n10683 = n2102 & ~n10682 ;
  assign n10684 = n2106 & ~n10683 ;
  assign n10685 = n2110 & ~n10684 ;
  assign n10686 = n2114 & ~n10685 ;
  assign n10687 = n2118 & ~n10686 ;
  assign n10688 = n2122 & ~n10687 ;
  assign n10689 = n2126 & ~n10688 ;
  assign n10690 = n2130 & ~n10689 ;
  assign n10691 = n2134 & ~n10690 ;
  assign n10692 = n2138 & ~n10691 ;
  assign n10693 = n2142 & ~n10692 ;
  assign n10694 = n2146 & ~n10693 ;
  assign n10695 = n2150 & ~n10694 ;
  assign n10696 = n2154 & ~n10695 ;
  assign n10697 = n2158 & ~n10696 ;
  assign n10698 = n2162 & ~n10697 ;
  assign n10699 = n2166 & ~n10698 ;
  assign n10700 = n2170 & ~n10699 ;
  assign n10701 = n2174 & ~n10700 ;
  assign n10702 = n2178 & ~n10701 ;
  assign n10703 = n2182 & ~n10702 ;
  assign n10704 = n2186 & ~n10703 ;
  assign n10705 = n2190 & ~n10704 ;
  assign n10706 = n2194 & ~n10705 ;
  assign n10707 = n2198 & ~n10706 ;
  assign n10708 = n2202 & ~n10707 ;
  assign n10709 = n2206 & ~n10708 ;
  assign n10710 = n2210 & ~n10709 ;
  assign n10711 = n2214 & ~n10710 ;
  assign n10712 = n2218 & ~n10711 ;
  assign n10713 = n2222 & ~n10712 ;
  assign n10714 = n2226 & ~n10713 ;
  assign n10715 = n2230 & ~n10714 ;
  assign n10716 = n2234 & ~n10715 ;
  assign n10717 = n2238 & ~n10716 ;
  assign n10718 = n2242 & ~n10717 ;
  assign n10719 = n2246 & ~n10718 ;
  assign n10720 = n2250 & ~n10719 ;
  assign n10721 = n2254 & ~n10720 ;
  assign n10722 = n2258 & ~n10721 ;
  assign n10723 = n2262 & ~n10722 ;
  assign n10724 = n2266 & ~n10723 ;
  assign n10725 = n2270 & ~n10724 ;
  assign n10726 = n2274 & ~n10725 ;
  assign n10727 = n2278 & ~n10726 ;
  assign n10728 = n2282 & ~n10727 ;
  assign n10729 = n2286 & ~n10728 ;
  assign n10730 = n2290 & ~n10729 ;
  assign n10731 = n2836 & ~n10730 ;
  assign n10732 = n602 & ~n10731 ;
  assign n10733 = n606 & ~n10732 ;
  assign n10734 = n610 & ~n10733 ;
  assign n10735 = n614 & ~n10734 ;
  assign n10736 = n618 & ~n10735 ;
  assign n10737 = n622 & ~n10736 ;
  assign n10738 = n626 & ~n10737 ;
  assign n10739 = n630 & ~n10738 ;
  assign n10740 = n634 & ~n10739 ;
  assign n10741 = n638 & ~n10740 ;
  assign n10742 = n642 & ~n10741 ;
  assign n10743 = n646 & ~n10742 ;
  assign n10744 = n650 & ~n10743 ;
  assign n10745 = n654 & ~n10744 ;
  assign n10746 = n658 & ~n10745 ;
  assign n10747 = n662 & ~n10746 ;
  assign n10748 = n666 & ~n10747 ;
  assign n10749 = n670 & ~n10748 ;
  assign n10750 = n674 & ~n10749 ;
  assign n10751 = n678 & ~n10750 ;
  assign n10752 = n682 & ~n10751 ;
  assign n10753 = n686 & ~n10752 ;
  assign n10754 = n690 & ~n10753 ;
  assign n10755 = n694 & ~n10754 ;
  assign n10756 = n698 & ~n10755 ;
  assign n10757 = n702 & ~n10756 ;
  assign n10758 = n706 & ~n10757 ;
  assign n10759 = n710 & ~n10758 ;
  assign n10760 = n714 & ~n10759 ;
  assign n10761 = n718 & ~n10760 ;
  assign n10762 = n722 & ~n10761 ;
  assign n10763 = ~x178 & ~n724 ;
  assign n10764 = ~n10762 & n10763 ;
  assign n10767 = ~n10764 & ~x306 ;
  assign n10768 = ~n10766 & ~n10767 ;
  assign n10769 = n394 & ~n1072 ;
  assign n10770 = n399 & ~n10769 ;
  assign n10771 = n403 & ~n10770 ;
  assign n10772 = n407 & ~n10771 ;
  assign n10773 = n411 & ~n10772 ;
  assign n10774 = n415 & ~n10773 ;
  assign n10775 = n419 & ~n10774 ;
  assign n10776 = n423 & ~n10775 ;
  assign n10777 = n427 & ~n10776 ;
  assign n10778 = n431 & ~n10777 ;
  assign n10779 = n435 & ~n10778 ;
  assign n10780 = n439 & ~n10779 ;
  assign n10781 = n443 & ~n10780 ;
  assign n10782 = n447 & ~n10781 ;
  assign n10783 = n451 & ~n10782 ;
  assign n10784 = n455 & ~n10783 ;
  assign n10785 = n459 & ~n10784 ;
  assign n10786 = n463 & ~n10785 ;
  assign n10787 = n467 & ~n10786 ;
  assign n10788 = n471 & ~n10787 ;
  assign n10789 = n475 & ~n10788 ;
  assign n10790 = n479 & ~n10789 ;
  assign n10791 = n483 & ~n10790 ;
  assign n10792 = n487 & ~n10791 ;
  assign n10793 = n491 & ~n10792 ;
  assign n10794 = n495 & ~n10793 ;
  assign n10795 = n499 & ~n10794 ;
  assign n10796 = n503 & ~n10795 ;
  assign n10797 = n507 & ~n10796 ;
  assign n10798 = n511 & ~n10797 ;
  assign n10799 = n515 & ~n10798 ;
  assign n10800 = n519 & ~n10799 ;
  assign n10801 = n523 & ~n10800 ;
  assign n10802 = n527 & ~n10801 ;
  assign n10803 = n531 & ~n10802 ;
  assign n10804 = n535 & ~n10803 ;
  assign n10805 = n539 & ~n10804 ;
  assign n10806 = n543 & ~n10805 ;
  assign n10807 = n547 & ~n10806 ;
  assign n10808 = n551 & ~n10807 ;
  assign n10809 = n555 & ~n10808 ;
  assign n10810 = n559 & ~n10809 ;
  assign n10811 = n563 & ~n10810 ;
  assign n10812 = n567 & ~n10811 ;
  assign n10813 = n571 & ~n10812 ;
  assign n10814 = n575 & ~n10813 ;
  assign n10815 = n579 & ~n10814 ;
  assign n10816 = n583 & ~n10815 ;
  assign n10817 = n587 & ~n10816 ;
  assign n10818 = n591 & ~n10817 ;
  assign n10819 = n2382 & ~n10818 ;
  assign n10820 = n2384 & ~n10819 ;
  assign n10821 = n2927 & ~n10820 ;
  assign n10822 = n945 & ~n10821 ;
  assign n10823 = n949 & ~n10822 ;
  assign n10824 = n953 & ~n10823 ;
  assign n10825 = n957 & ~n10824 ;
  assign n10826 = n961 & ~n10825 ;
  assign n10827 = n965 & ~n10826 ;
  assign n10828 = n969 & ~n10827 ;
  assign n10829 = n973 & ~n10828 ;
  assign n10830 = n977 & ~n10829 ;
  assign n10831 = n981 & ~n10830 ;
  assign n10832 = n985 & ~n10831 ;
  assign n10833 = n989 & ~n10832 ;
  assign n10834 = n993 & ~n10833 ;
  assign n10835 = n997 & ~n10834 ;
  assign n10836 = n1001 & ~n10835 ;
  assign n10837 = n1005 & ~n10836 ;
  assign n10838 = n1009 & ~n10837 ;
  assign n10839 = n1013 & ~n10838 ;
  assign n10840 = n1017 & ~n10839 ;
  assign n10841 = n1021 & ~n10840 ;
  assign n10842 = n1025 & ~n10841 ;
  assign n10843 = n1029 & ~n10842 ;
  assign n10844 = n1033 & ~n10843 ;
  assign n10845 = n1037 & ~n10844 ;
  assign n10846 = n1041 & ~n10845 ;
  assign n10847 = n1045 & ~n10846 ;
  assign n10848 = n1049 & ~n10847 ;
  assign n10849 = n1053 & ~n10848 ;
  assign n10850 = n1057 & ~n10849 ;
  assign n10851 = n1061 & ~n10850 ;
  assign n10852 = n1065 & ~n10851 ;
  assign n10853 = x179 & ~n1067 ;
  assign n10854 = ~n10852 & n10853 ;
  assign n10942 = n10854 & x307 ;
  assign n10855 = n733 & ~n1411 ;
  assign n10856 = n738 & ~n10855 ;
  assign n10857 = n742 & ~n10856 ;
  assign n10858 = n746 & ~n10857 ;
  assign n10859 = n750 & ~n10858 ;
  assign n10860 = n754 & ~n10859 ;
  assign n10861 = n758 & ~n10860 ;
  assign n10862 = n762 & ~n10861 ;
  assign n10863 = n766 & ~n10862 ;
  assign n10864 = n770 & ~n10863 ;
  assign n10865 = n774 & ~n10864 ;
  assign n10866 = n778 & ~n10865 ;
  assign n10867 = n782 & ~n10866 ;
  assign n10868 = n786 & ~n10867 ;
  assign n10869 = n790 & ~n10868 ;
  assign n10870 = n794 & ~n10869 ;
  assign n10871 = n798 & ~n10870 ;
  assign n10872 = n802 & ~n10871 ;
  assign n10873 = n806 & ~n10872 ;
  assign n10874 = n810 & ~n10873 ;
  assign n10875 = n814 & ~n10874 ;
  assign n10876 = n818 & ~n10875 ;
  assign n10877 = n822 & ~n10876 ;
  assign n10878 = n826 & ~n10877 ;
  assign n10879 = n830 & ~n10878 ;
  assign n10880 = n834 & ~n10879 ;
  assign n10881 = n838 & ~n10880 ;
  assign n10882 = n842 & ~n10881 ;
  assign n10883 = n846 & ~n10882 ;
  assign n10884 = n850 & ~n10883 ;
  assign n10885 = n854 & ~n10884 ;
  assign n10886 = n858 & ~n10885 ;
  assign n10887 = n862 & ~n10886 ;
  assign n10888 = n866 & ~n10887 ;
  assign n10889 = n870 & ~n10888 ;
  assign n10890 = n874 & ~n10889 ;
  assign n10891 = n878 & ~n10890 ;
  assign n10892 = n882 & ~n10891 ;
  assign n10893 = n886 & ~n10892 ;
  assign n10894 = n890 & ~n10893 ;
  assign n10895 = n894 & ~n10894 ;
  assign n10896 = n898 & ~n10895 ;
  assign n10897 = n902 & ~n10896 ;
  assign n10898 = n906 & ~n10897 ;
  assign n10899 = n910 & ~n10898 ;
  assign n10900 = n914 & ~n10899 ;
  assign n10901 = n918 & ~n10900 ;
  assign n10902 = n922 & ~n10901 ;
  assign n10903 = n926 & ~n10902 ;
  assign n10904 = n930 & ~n10903 ;
  assign n10905 = n2472 & ~n10904 ;
  assign n10906 = n2474 & ~n10905 ;
  assign n10907 = n3014 & ~n10906 ;
  assign n10908 = n1284 & ~n10907 ;
  assign n10909 = n1288 & ~n10908 ;
  assign n10910 = n1292 & ~n10909 ;
  assign n10911 = n1296 & ~n10910 ;
  assign n10912 = n1300 & ~n10911 ;
  assign n10913 = n1304 & ~n10912 ;
  assign n10914 = n1308 & ~n10913 ;
  assign n10915 = n1312 & ~n10914 ;
  assign n10916 = n1316 & ~n10915 ;
  assign n10917 = n1320 & ~n10916 ;
  assign n10918 = n1324 & ~n10917 ;
  assign n10919 = n1328 & ~n10918 ;
  assign n10920 = n1332 & ~n10919 ;
  assign n10921 = n1336 & ~n10920 ;
  assign n10922 = n1340 & ~n10921 ;
  assign n10923 = n1344 & ~n10922 ;
  assign n10924 = n1348 & ~n10923 ;
  assign n10925 = n1352 & ~n10924 ;
  assign n10926 = n1356 & ~n10925 ;
  assign n10927 = n1360 & ~n10926 ;
  assign n10928 = n1364 & ~n10927 ;
  assign n10929 = n1368 & ~n10928 ;
  assign n10930 = n1372 & ~n10929 ;
  assign n10931 = n1376 & ~n10930 ;
  assign n10932 = n1380 & ~n10931 ;
  assign n10933 = n1384 & ~n10932 ;
  assign n10934 = n1388 & ~n10933 ;
  assign n10935 = n1392 & ~n10934 ;
  assign n10936 = n1396 & ~n10935 ;
  assign n10937 = n1400 & ~n10936 ;
  assign n10938 = n1404 & ~n10937 ;
  assign n10939 = ~x179 & ~n1406 ;
  assign n10940 = ~n10938 & n10939 ;
  assign n10943 = ~n10940 & ~x307 ;
  assign n10944 = ~n10942 & ~n10943 ;
  assign n10945 = n1076 & ~n1752 ;
  assign n10946 = n1081 & ~n10945 ;
  assign n10947 = n1085 & ~n10946 ;
  assign n10948 = n1089 & ~n10947 ;
  assign n10949 = n1093 & ~n10948 ;
  assign n10950 = n1097 & ~n10949 ;
  assign n10951 = n1101 & ~n10950 ;
  assign n10952 = n1105 & ~n10951 ;
  assign n10953 = n1109 & ~n10952 ;
  assign n10954 = n1113 & ~n10953 ;
  assign n10955 = n1117 & ~n10954 ;
  assign n10956 = n1121 & ~n10955 ;
  assign n10957 = n1125 & ~n10956 ;
  assign n10958 = n1129 & ~n10957 ;
  assign n10959 = n1133 & ~n10958 ;
  assign n10960 = n1137 & ~n10959 ;
  assign n10961 = n1141 & ~n10960 ;
  assign n10962 = n1145 & ~n10961 ;
  assign n10963 = n1149 & ~n10962 ;
  assign n10964 = n1153 & ~n10963 ;
  assign n10965 = n1157 & ~n10964 ;
  assign n10966 = n1161 & ~n10965 ;
  assign n10967 = n1165 & ~n10966 ;
  assign n10968 = n1169 & ~n10967 ;
  assign n10969 = n1173 & ~n10968 ;
  assign n10970 = n1177 & ~n10969 ;
  assign n10971 = n1181 & ~n10970 ;
  assign n10972 = n1185 & ~n10971 ;
  assign n10973 = n1189 & ~n10972 ;
  assign n10974 = n1193 & ~n10973 ;
  assign n10975 = n1197 & ~n10974 ;
  assign n10976 = n1201 & ~n10975 ;
  assign n10977 = n1205 & ~n10976 ;
  assign n10978 = n1209 & ~n10977 ;
  assign n10979 = n1213 & ~n10978 ;
  assign n10980 = n1217 & ~n10979 ;
  assign n10981 = n1221 & ~n10980 ;
  assign n10982 = n1225 & ~n10981 ;
  assign n10983 = n1229 & ~n10982 ;
  assign n10984 = n1233 & ~n10983 ;
  assign n10985 = n1237 & ~n10984 ;
  assign n10986 = n1241 & ~n10985 ;
  assign n10987 = n1245 & ~n10986 ;
  assign n10988 = n1249 & ~n10987 ;
  assign n10989 = n1253 & ~n10988 ;
  assign n10990 = n1257 & ~n10989 ;
  assign n10991 = n1261 & ~n10990 ;
  assign n10992 = n1265 & ~n10991 ;
  assign n10993 = n1269 & ~n10992 ;
  assign n10994 = n1273 & ~n10993 ;
  assign n10995 = n2566 & ~n10994 ;
  assign n10996 = n2568 & ~n10995 ;
  assign n10997 = n3105 & ~n10996 ;
  assign n10998 = n1625 & ~n10997 ;
  assign n10999 = n1629 & ~n10998 ;
  assign n11000 = n1633 & ~n10999 ;
  assign n11001 = n1637 & ~n11000 ;
  assign n11002 = n1641 & ~n11001 ;
  assign n11003 = n1645 & ~n11002 ;
  assign n11004 = n1649 & ~n11003 ;
  assign n11005 = n1653 & ~n11004 ;
  assign n11006 = n1657 & ~n11005 ;
  assign n11007 = n1661 & ~n11006 ;
  assign n11008 = n1665 & ~n11007 ;
  assign n11009 = n1669 & ~n11008 ;
  assign n11010 = n1673 & ~n11009 ;
  assign n11011 = n1677 & ~n11010 ;
  assign n11012 = n1681 & ~n11011 ;
  assign n11013 = n1685 & ~n11012 ;
  assign n11014 = n1689 & ~n11013 ;
  assign n11015 = n1693 & ~n11014 ;
  assign n11016 = n1697 & ~n11015 ;
  assign n11017 = n1701 & ~n11016 ;
  assign n11018 = n1705 & ~n11017 ;
  assign n11019 = n1709 & ~n11018 ;
  assign n11020 = n1713 & ~n11019 ;
  assign n11021 = n1717 & ~n11020 ;
  assign n11022 = n1721 & ~n11021 ;
  assign n11023 = n1725 & ~n11022 ;
  assign n11024 = n1729 & ~n11023 ;
  assign n11025 = n1733 & ~n11024 ;
  assign n11026 = n1737 & ~n11025 ;
  assign n11027 = n1741 & ~n11026 ;
  assign n11028 = n1745 & ~n11027 ;
  assign n11029 = x180 & ~n1747 ;
  assign n11030 = ~n11028 & n11029 ;
  assign n11118 = n11030 & x308 ;
  assign n11031 = n1415 & ~n2089 ;
  assign n11032 = n1420 & ~n11031 ;
  assign n11033 = n1424 & ~n11032 ;
  assign n11034 = n1428 & ~n11033 ;
  assign n11035 = n1432 & ~n11034 ;
  assign n11036 = n1436 & ~n11035 ;
  assign n11037 = n1440 & ~n11036 ;
  assign n11038 = n1444 & ~n11037 ;
  assign n11039 = n1448 & ~n11038 ;
  assign n11040 = n1452 & ~n11039 ;
  assign n11041 = n1456 & ~n11040 ;
  assign n11042 = n1460 & ~n11041 ;
  assign n11043 = n1464 & ~n11042 ;
  assign n11044 = n1468 & ~n11043 ;
  assign n11045 = n1472 & ~n11044 ;
  assign n11046 = n1476 & ~n11045 ;
  assign n11047 = n1480 & ~n11046 ;
  assign n11048 = n1484 & ~n11047 ;
  assign n11049 = n1488 & ~n11048 ;
  assign n11050 = n1492 & ~n11049 ;
  assign n11051 = n1496 & ~n11050 ;
  assign n11052 = n1500 & ~n11051 ;
  assign n11053 = n1504 & ~n11052 ;
  assign n11054 = n1508 & ~n11053 ;
  assign n11055 = n1512 & ~n11054 ;
  assign n11056 = n1516 & ~n11055 ;
  assign n11057 = n1520 & ~n11056 ;
  assign n11058 = n1524 & ~n11057 ;
  assign n11059 = n1528 & ~n11058 ;
  assign n11060 = n1532 & ~n11059 ;
  assign n11061 = n1536 & ~n11060 ;
  assign n11062 = n1540 & ~n11061 ;
  assign n11063 = n1544 & ~n11062 ;
  assign n11064 = n1548 & ~n11063 ;
  assign n11065 = n1552 & ~n11064 ;
  assign n11066 = n1556 & ~n11065 ;
  assign n11067 = n1560 & ~n11066 ;
  assign n11068 = n1564 & ~n11067 ;
  assign n11069 = n1568 & ~n11068 ;
  assign n11070 = n1572 & ~n11069 ;
  assign n11071 = n1576 & ~n11070 ;
  assign n11072 = n1580 & ~n11071 ;
  assign n11073 = n1584 & ~n11072 ;
  assign n11074 = n1588 & ~n11073 ;
  assign n11075 = n1592 & ~n11074 ;
  assign n11076 = n1596 & ~n11075 ;
  assign n11077 = n1600 & ~n11076 ;
  assign n11078 = n1604 & ~n11077 ;
  assign n11079 = n1608 & ~n11078 ;
  assign n11080 = n1612 & ~n11079 ;
  assign n11081 = n2656 & ~n11080 ;
  assign n11082 = n2658 & ~n11081 ;
  assign n11083 = n3192 & ~n11082 ;
  assign n11084 = n1962 & ~n11083 ;
  assign n11085 = n1966 & ~n11084 ;
  assign n11086 = n1970 & ~n11085 ;
  assign n11087 = n1974 & ~n11086 ;
  assign n11088 = n1978 & ~n11087 ;
  assign n11089 = n1982 & ~n11088 ;
  assign n11090 = n1986 & ~n11089 ;
  assign n11091 = n1990 & ~n11090 ;
  assign n11092 = n1994 & ~n11091 ;
  assign n11093 = n1998 & ~n11092 ;
  assign n11094 = n2002 & ~n11093 ;
  assign n11095 = n2006 & ~n11094 ;
  assign n11096 = n2010 & ~n11095 ;
  assign n11097 = n2014 & ~n11096 ;
  assign n11098 = n2018 & ~n11097 ;
  assign n11099 = n2022 & ~n11098 ;
  assign n11100 = n2026 & ~n11099 ;
  assign n11101 = n2030 & ~n11100 ;
  assign n11102 = n2034 & ~n11101 ;
  assign n11103 = n2038 & ~n11102 ;
  assign n11104 = n2042 & ~n11103 ;
  assign n11105 = n2046 & ~n11104 ;
  assign n11106 = n2050 & ~n11105 ;
  assign n11107 = n2054 & ~n11106 ;
  assign n11108 = n2058 & ~n11107 ;
  assign n11109 = n2062 & ~n11108 ;
  assign n11110 = n2066 & ~n11109 ;
  assign n11111 = n2070 & ~n11110 ;
  assign n11112 = n2074 & ~n11111 ;
  assign n11113 = n2078 & ~n11112 ;
  assign n11114 = n2082 & ~n11113 ;
  assign n11115 = ~x180 & ~n2084 ;
  assign n11116 = ~n11114 & n11115 ;
  assign n11119 = ~n11116 & ~x308 ;
  assign n11120 = ~n11118 & ~n11119 ;
  assign n11121 = ~n398 & n1756 ;
  assign n11122 = n1761 & ~n11121 ;
  assign n11123 = n1765 & ~n11122 ;
  assign n11124 = n1769 & ~n11123 ;
  assign n11125 = n1773 & ~n11124 ;
  assign n11126 = n1777 & ~n11125 ;
  assign n11127 = n1781 & ~n11126 ;
  assign n11128 = n1785 & ~n11127 ;
  assign n11129 = n1789 & ~n11128 ;
  assign n11130 = n1793 & ~n11129 ;
  assign n11131 = n1797 & ~n11130 ;
  assign n11132 = n1801 & ~n11131 ;
  assign n11133 = n1805 & ~n11132 ;
  assign n11134 = n1809 & ~n11133 ;
  assign n11135 = n1813 & ~n11134 ;
  assign n11136 = n1817 & ~n11135 ;
  assign n11137 = n1821 & ~n11136 ;
  assign n11138 = n1825 & ~n11137 ;
  assign n11139 = n1829 & ~n11138 ;
  assign n11140 = n1833 & ~n11139 ;
  assign n11141 = n1837 & ~n11140 ;
  assign n11142 = n1841 & ~n11141 ;
  assign n11143 = n1845 & ~n11142 ;
  assign n11144 = n1849 & ~n11143 ;
  assign n11145 = n1853 & ~n11144 ;
  assign n11146 = n1857 & ~n11145 ;
  assign n11147 = n1861 & ~n11146 ;
  assign n11148 = n1865 & ~n11147 ;
  assign n11149 = n1869 & ~n11148 ;
  assign n11150 = n1873 & ~n11149 ;
  assign n11151 = n1877 & ~n11150 ;
  assign n11152 = n1881 & ~n11151 ;
  assign n11153 = n1885 & ~n11152 ;
  assign n11154 = n1889 & ~n11153 ;
  assign n11155 = n1893 & ~n11154 ;
  assign n11156 = n1897 & ~n11155 ;
  assign n11157 = n1901 & ~n11156 ;
  assign n11158 = n1905 & ~n11157 ;
  assign n11159 = n1909 & ~n11158 ;
  assign n11160 = n1913 & ~n11159 ;
  assign n11161 = n1917 & ~n11160 ;
  assign n11162 = n1921 & ~n11161 ;
  assign n11163 = n1925 & ~n11162 ;
  assign n11164 = n1929 & ~n11163 ;
  assign n11165 = n1933 & ~n11164 ;
  assign n11166 = n1937 & ~n11165 ;
  assign n11167 = n1941 & ~n11166 ;
  assign n11168 = n1945 & ~n11167 ;
  assign n11169 = n1949 & ~n11168 ;
  assign n11170 = n1953 & ~n11169 ;
  assign n11171 = n2749 & ~n11170 ;
  assign n11172 = n263 & ~n11171 ;
  assign n11173 = n267 & ~n11172 ;
  assign n11174 = n271 & ~n11173 ;
  assign n11175 = n275 & ~n11174 ;
  assign n11176 = n279 & ~n11175 ;
  assign n11177 = n283 & ~n11176 ;
  assign n11178 = n287 & ~n11177 ;
  assign n11179 = n291 & ~n11178 ;
  assign n11180 = n295 & ~n11179 ;
  assign n11181 = n299 & ~n11180 ;
  assign n11182 = n303 & ~n11181 ;
  assign n11183 = n307 & ~n11182 ;
  assign n11184 = n311 & ~n11183 ;
  assign n11185 = n315 & ~n11184 ;
  assign n11186 = n319 & ~n11185 ;
  assign n11187 = n323 & ~n11186 ;
  assign n11188 = n327 & ~n11187 ;
  assign n11189 = n331 & ~n11188 ;
  assign n11190 = n335 & ~n11189 ;
  assign n11191 = n339 & ~n11190 ;
  assign n11192 = n343 & ~n11191 ;
  assign n11193 = n347 & ~n11192 ;
  assign n11194 = n351 & ~n11193 ;
  assign n11195 = n355 & ~n11194 ;
  assign n11196 = n359 & ~n11195 ;
  assign n11197 = n363 & ~n11196 ;
  assign n11198 = n367 & ~n11197 ;
  assign n11199 = n371 & ~n11198 ;
  assign n11200 = n375 & ~n11199 ;
  assign n11201 = n379 & ~n11200 ;
  assign n11202 = n383 & ~n11201 ;
  assign n11203 = n387 & ~n11202 ;
  assign n11204 = n391 & ~n11203 ;
  assign n11205 = x181 & ~n393 ;
  assign n11206 = ~n11204 & n11205 ;
  assign n11294 = n11206 & x309 ;
  assign n11207 = ~n737 & n2093 ;
  assign n11208 = n2098 & ~n11207 ;
  assign n11209 = n2102 & ~n11208 ;
  assign n11210 = n2106 & ~n11209 ;
  assign n11211 = n2110 & ~n11210 ;
  assign n11212 = n2114 & ~n11211 ;
  assign n11213 = n2118 & ~n11212 ;
  assign n11214 = n2122 & ~n11213 ;
  assign n11215 = n2126 & ~n11214 ;
  assign n11216 = n2130 & ~n11215 ;
  assign n11217 = n2134 & ~n11216 ;
  assign n11218 = n2138 & ~n11217 ;
  assign n11219 = n2142 & ~n11218 ;
  assign n11220 = n2146 & ~n11219 ;
  assign n11221 = n2150 & ~n11220 ;
  assign n11222 = n2154 & ~n11221 ;
  assign n11223 = n2158 & ~n11222 ;
  assign n11224 = n2162 & ~n11223 ;
  assign n11225 = n2166 & ~n11224 ;
  assign n11226 = n2170 & ~n11225 ;
  assign n11227 = n2174 & ~n11226 ;
  assign n11228 = n2178 & ~n11227 ;
  assign n11229 = n2182 & ~n11228 ;
  assign n11230 = n2186 & ~n11229 ;
  assign n11231 = n2190 & ~n11230 ;
  assign n11232 = n2194 & ~n11231 ;
  assign n11233 = n2198 & ~n11232 ;
  assign n11234 = n2202 & ~n11233 ;
  assign n11235 = n2206 & ~n11234 ;
  assign n11236 = n2210 & ~n11235 ;
  assign n11237 = n2214 & ~n11236 ;
  assign n11238 = n2218 & ~n11237 ;
  assign n11239 = n2222 & ~n11238 ;
  assign n11240 = n2226 & ~n11239 ;
  assign n11241 = n2230 & ~n11240 ;
  assign n11242 = n2234 & ~n11241 ;
  assign n11243 = n2238 & ~n11242 ;
  assign n11244 = n2242 & ~n11243 ;
  assign n11245 = n2246 & ~n11244 ;
  assign n11246 = n2250 & ~n11245 ;
  assign n11247 = n2254 & ~n11246 ;
  assign n11248 = n2258 & ~n11247 ;
  assign n11249 = n2262 & ~n11248 ;
  assign n11250 = n2266 & ~n11249 ;
  assign n11251 = n2270 & ~n11250 ;
  assign n11252 = n2274 & ~n11251 ;
  assign n11253 = n2278 & ~n11252 ;
  assign n11254 = n2282 & ~n11253 ;
  assign n11255 = n2286 & ~n11254 ;
  assign n11256 = n2290 & ~n11255 ;
  assign n11257 = n2836 & ~n11256 ;
  assign n11258 = n602 & ~n11257 ;
  assign n11259 = n606 & ~n11258 ;
  assign n11260 = n610 & ~n11259 ;
  assign n11261 = n614 & ~n11260 ;
  assign n11262 = n618 & ~n11261 ;
  assign n11263 = n622 & ~n11262 ;
  assign n11264 = n626 & ~n11263 ;
  assign n11265 = n630 & ~n11264 ;
  assign n11266 = n634 & ~n11265 ;
  assign n11267 = n638 & ~n11266 ;
  assign n11268 = n642 & ~n11267 ;
  assign n11269 = n646 & ~n11268 ;
  assign n11270 = n650 & ~n11269 ;
  assign n11271 = n654 & ~n11270 ;
  assign n11272 = n658 & ~n11271 ;
  assign n11273 = n662 & ~n11272 ;
  assign n11274 = n666 & ~n11273 ;
  assign n11275 = n670 & ~n11274 ;
  assign n11276 = n674 & ~n11275 ;
  assign n11277 = n678 & ~n11276 ;
  assign n11278 = n682 & ~n11277 ;
  assign n11279 = n686 & ~n11278 ;
  assign n11280 = n690 & ~n11279 ;
  assign n11281 = n694 & ~n11280 ;
  assign n11282 = n698 & ~n11281 ;
  assign n11283 = n702 & ~n11282 ;
  assign n11284 = n706 & ~n11283 ;
  assign n11285 = n710 & ~n11284 ;
  assign n11286 = n714 & ~n11285 ;
  assign n11287 = n718 & ~n11286 ;
  assign n11288 = n722 & ~n11287 ;
  assign n11289 = n726 & ~n11288 ;
  assign n11290 = n730 & ~n11289 ;
  assign n11291 = ~x181 & ~n732 ;
  assign n11292 = ~n11290 & n11291 ;
  assign n11295 = ~n11292 & ~x309 ;
  assign n11296 = ~n11294 & ~n11295 ;
  assign n11297 = n402 & ~n1080 ;
  assign n11298 = n407 & ~n11297 ;
  assign n11299 = n411 & ~n11298 ;
  assign n11300 = n415 & ~n11299 ;
  assign n11301 = n419 & ~n11300 ;
  assign n11302 = n423 & ~n11301 ;
  assign n11303 = n427 & ~n11302 ;
  assign n11304 = n431 & ~n11303 ;
  assign n11305 = n435 & ~n11304 ;
  assign n11306 = n439 & ~n11305 ;
  assign n11307 = n443 & ~n11306 ;
  assign n11308 = n447 & ~n11307 ;
  assign n11309 = n451 & ~n11308 ;
  assign n11310 = n455 & ~n11309 ;
  assign n11311 = n459 & ~n11310 ;
  assign n11312 = n463 & ~n11311 ;
  assign n11313 = n467 & ~n11312 ;
  assign n11314 = n471 & ~n11313 ;
  assign n11315 = n475 & ~n11314 ;
  assign n11316 = n479 & ~n11315 ;
  assign n11317 = n483 & ~n11316 ;
  assign n11318 = n487 & ~n11317 ;
  assign n11319 = n491 & ~n11318 ;
  assign n11320 = n495 & ~n11319 ;
  assign n11321 = n499 & ~n11320 ;
  assign n11322 = n503 & ~n11321 ;
  assign n11323 = n507 & ~n11322 ;
  assign n11324 = n511 & ~n11323 ;
  assign n11325 = n515 & ~n11324 ;
  assign n11326 = n519 & ~n11325 ;
  assign n11327 = n523 & ~n11326 ;
  assign n11328 = n527 & ~n11327 ;
  assign n11329 = n531 & ~n11328 ;
  assign n11330 = n535 & ~n11329 ;
  assign n11331 = n539 & ~n11330 ;
  assign n11332 = n543 & ~n11331 ;
  assign n11333 = n547 & ~n11332 ;
  assign n11334 = n551 & ~n11333 ;
  assign n11335 = n555 & ~n11334 ;
  assign n11336 = n559 & ~n11335 ;
  assign n11337 = n563 & ~n11336 ;
  assign n11338 = n567 & ~n11337 ;
  assign n11339 = n571 & ~n11338 ;
  assign n11340 = n575 & ~n11339 ;
  assign n11341 = n579 & ~n11340 ;
  assign n11342 = n583 & ~n11341 ;
  assign n11343 = n587 & ~n11342 ;
  assign n11344 = n591 & ~n11343 ;
  assign n11345 = n2382 & ~n11344 ;
  assign n11346 = n2384 & ~n11345 ;
  assign n11347 = n2927 & ~n11346 ;
  assign n11348 = n945 & ~n11347 ;
  assign n11349 = n949 & ~n11348 ;
  assign n11350 = n953 & ~n11349 ;
  assign n11351 = n957 & ~n11350 ;
  assign n11352 = n961 & ~n11351 ;
  assign n11353 = n965 & ~n11352 ;
  assign n11354 = n969 & ~n11353 ;
  assign n11355 = n973 & ~n11354 ;
  assign n11356 = n977 & ~n11355 ;
  assign n11357 = n981 & ~n11356 ;
  assign n11358 = n985 & ~n11357 ;
  assign n11359 = n989 & ~n11358 ;
  assign n11360 = n993 & ~n11359 ;
  assign n11361 = n997 & ~n11360 ;
  assign n11362 = n1001 & ~n11361 ;
  assign n11363 = n1005 & ~n11362 ;
  assign n11364 = n1009 & ~n11363 ;
  assign n11365 = n1013 & ~n11364 ;
  assign n11366 = n1017 & ~n11365 ;
  assign n11367 = n1021 & ~n11366 ;
  assign n11368 = n1025 & ~n11367 ;
  assign n11369 = n1029 & ~n11368 ;
  assign n11370 = n1033 & ~n11369 ;
  assign n11371 = n1037 & ~n11370 ;
  assign n11372 = n1041 & ~n11371 ;
  assign n11373 = n1045 & ~n11372 ;
  assign n11374 = n1049 & ~n11373 ;
  assign n11375 = n1053 & ~n11374 ;
  assign n11376 = n1057 & ~n11375 ;
  assign n11377 = n1061 & ~n11376 ;
  assign n11378 = n1065 & ~n11377 ;
  assign n11379 = n1069 & ~n11378 ;
  assign n11380 = n1073 & ~n11379 ;
  assign n11381 = x182 & ~n1075 ;
  assign n11382 = ~n11380 & n11381 ;
  assign n11470 = n11382 & x310 ;
  assign n11383 = n741 & ~n1419 ;
  assign n11384 = n746 & ~n11383 ;
  assign n11385 = n750 & ~n11384 ;
  assign n11386 = n754 & ~n11385 ;
  assign n11387 = n758 & ~n11386 ;
  assign n11388 = n762 & ~n11387 ;
  assign n11389 = n766 & ~n11388 ;
  assign n11390 = n770 & ~n11389 ;
  assign n11391 = n774 & ~n11390 ;
  assign n11392 = n778 & ~n11391 ;
  assign n11393 = n782 & ~n11392 ;
  assign n11394 = n786 & ~n11393 ;
  assign n11395 = n790 & ~n11394 ;
  assign n11396 = n794 & ~n11395 ;
  assign n11397 = n798 & ~n11396 ;
  assign n11398 = n802 & ~n11397 ;
  assign n11399 = n806 & ~n11398 ;
  assign n11400 = n810 & ~n11399 ;
  assign n11401 = n814 & ~n11400 ;
  assign n11402 = n818 & ~n11401 ;
  assign n11403 = n822 & ~n11402 ;
  assign n11404 = n826 & ~n11403 ;
  assign n11405 = n830 & ~n11404 ;
  assign n11406 = n834 & ~n11405 ;
  assign n11407 = n838 & ~n11406 ;
  assign n11408 = n842 & ~n11407 ;
  assign n11409 = n846 & ~n11408 ;
  assign n11410 = n850 & ~n11409 ;
  assign n11411 = n854 & ~n11410 ;
  assign n11412 = n858 & ~n11411 ;
  assign n11413 = n862 & ~n11412 ;
  assign n11414 = n866 & ~n11413 ;
  assign n11415 = n870 & ~n11414 ;
  assign n11416 = n874 & ~n11415 ;
  assign n11417 = n878 & ~n11416 ;
  assign n11418 = n882 & ~n11417 ;
  assign n11419 = n886 & ~n11418 ;
  assign n11420 = n890 & ~n11419 ;
  assign n11421 = n894 & ~n11420 ;
  assign n11422 = n898 & ~n11421 ;
  assign n11423 = n902 & ~n11422 ;
  assign n11424 = n906 & ~n11423 ;
  assign n11425 = n910 & ~n11424 ;
  assign n11426 = n914 & ~n11425 ;
  assign n11427 = n918 & ~n11426 ;
  assign n11428 = n922 & ~n11427 ;
  assign n11429 = n926 & ~n11428 ;
  assign n11430 = n930 & ~n11429 ;
  assign n11431 = n2472 & ~n11430 ;
  assign n11432 = n2474 & ~n11431 ;
  assign n11433 = n3014 & ~n11432 ;
  assign n11434 = n1284 & ~n11433 ;
  assign n11435 = n1288 & ~n11434 ;
  assign n11436 = n1292 & ~n11435 ;
  assign n11437 = n1296 & ~n11436 ;
  assign n11438 = n1300 & ~n11437 ;
  assign n11439 = n1304 & ~n11438 ;
  assign n11440 = n1308 & ~n11439 ;
  assign n11441 = n1312 & ~n11440 ;
  assign n11442 = n1316 & ~n11441 ;
  assign n11443 = n1320 & ~n11442 ;
  assign n11444 = n1324 & ~n11443 ;
  assign n11445 = n1328 & ~n11444 ;
  assign n11446 = n1332 & ~n11445 ;
  assign n11447 = n1336 & ~n11446 ;
  assign n11448 = n1340 & ~n11447 ;
  assign n11449 = n1344 & ~n11448 ;
  assign n11450 = n1348 & ~n11449 ;
  assign n11451 = n1352 & ~n11450 ;
  assign n11452 = n1356 & ~n11451 ;
  assign n11453 = n1360 & ~n11452 ;
  assign n11454 = n1364 & ~n11453 ;
  assign n11455 = n1368 & ~n11454 ;
  assign n11456 = n1372 & ~n11455 ;
  assign n11457 = n1376 & ~n11456 ;
  assign n11458 = n1380 & ~n11457 ;
  assign n11459 = n1384 & ~n11458 ;
  assign n11460 = n1388 & ~n11459 ;
  assign n11461 = n1392 & ~n11460 ;
  assign n11462 = n1396 & ~n11461 ;
  assign n11463 = n1400 & ~n11462 ;
  assign n11464 = n1404 & ~n11463 ;
  assign n11465 = n1408 & ~n11464 ;
  assign n11466 = n1412 & ~n11465 ;
  assign n11467 = ~x182 & ~n1414 ;
  assign n11468 = ~n11466 & n11467 ;
  assign n11471 = ~n11468 & ~x310 ;
  assign n11472 = ~n11470 & ~n11471 ;
  assign n11473 = n1084 & ~n1760 ;
  assign n11474 = n1089 & ~n11473 ;
  assign n11475 = n1093 & ~n11474 ;
  assign n11476 = n1097 & ~n11475 ;
  assign n11477 = n1101 & ~n11476 ;
  assign n11478 = n1105 & ~n11477 ;
  assign n11479 = n1109 & ~n11478 ;
  assign n11480 = n1113 & ~n11479 ;
  assign n11481 = n1117 & ~n11480 ;
  assign n11482 = n1121 & ~n11481 ;
  assign n11483 = n1125 & ~n11482 ;
  assign n11484 = n1129 & ~n11483 ;
  assign n11485 = n1133 & ~n11484 ;
  assign n11486 = n1137 & ~n11485 ;
  assign n11487 = n1141 & ~n11486 ;
  assign n11488 = n1145 & ~n11487 ;
  assign n11489 = n1149 & ~n11488 ;
  assign n11490 = n1153 & ~n11489 ;
  assign n11491 = n1157 & ~n11490 ;
  assign n11492 = n1161 & ~n11491 ;
  assign n11493 = n1165 & ~n11492 ;
  assign n11494 = n1169 & ~n11493 ;
  assign n11495 = n1173 & ~n11494 ;
  assign n11496 = n1177 & ~n11495 ;
  assign n11497 = n1181 & ~n11496 ;
  assign n11498 = n1185 & ~n11497 ;
  assign n11499 = n1189 & ~n11498 ;
  assign n11500 = n1193 & ~n11499 ;
  assign n11501 = n1197 & ~n11500 ;
  assign n11502 = n1201 & ~n11501 ;
  assign n11503 = n1205 & ~n11502 ;
  assign n11504 = n1209 & ~n11503 ;
  assign n11505 = n1213 & ~n11504 ;
  assign n11506 = n1217 & ~n11505 ;
  assign n11507 = n1221 & ~n11506 ;
  assign n11508 = n1225 & ~n11507 ;
  assign n11509 = n1229 & ~n11508 ;
  assign n11510 = n1233 & ~n11509 ;
  assign n11511 = n1237 & ~n11510 ;
  assign n11512 = n1241 & ~n11511 ;
  assign n11513 = n1245 & ~n11512 ;
  assign n11514 = n1249 & ~n11513 ;
  assign n11515 = n1253 & ~n11514 ;
  assign n11516 = n1257 & ~n11515 ;
  assign n11517 = n1261 & ~n11516 ;
  assign n11518 = n1265 & ~n11517 ;
  assign n11519 = n1269 & ~n11518 ;
  assign n11520 = n1273 & ~n11519 ;
  assign n11521 = n2566 & ~n11520 ;
  assign n11522 = n2568 & ~n11521 ;
  assign n11523 = n3105 & ~n11522 ;
  assign n11524 = n1625 & ~n11523 ;
  assign n11525 = n1629 & ~n11524 ;
  assign n11526 = n1633 & ~n11525 ;
  assign n11527 = n1637 & ~n11526 ;
  assign n11528 = n1641 & ~n11527 ;
  assign n11529 = n1645 & ~n11528 ;
  assign n11530 = n1649 & ~n11529 ;
  assign n11531 = n1653 & ~n11530 ;
  assign n11532 = n1657 & ~n11531 ;
  assign n11533 = n1661 & ~n11532 ;
  assign n11534 = n1665 & ~n11533 ;
  assign n11535 = n1669 & ~n11534 ;
  assign n11536 = n1673 & ~n11535 ;
  assign n11537 = n1677 & ~n11536 ;
  assign n11538 = n1681 & ~n11537 ;
  assign n11539 = n1685 & ~n11538 ;
  assign n11540 = n1689 & ~n11539 ;
  assign n11541 = n1693 & ~n11540 ;
  assign n11542 = n1697 & ~n11541 ;
  assign n11543 = n1701 & ~n11542 ;
  assign n11544 = n1705 & ~n11543 ;
  assign n11545 = n1709 & ~n11544 ;
  assign n11546 = n1713 & ~n11545 ;
  assign n11547 = n1717 & ~n11546 ;
  assign n11548 = n1721 & ~n11547 ;
  assign n11549 = n1725 & ~n11548 ;
  assign n11550 = n1729 & ~n11549 ;
  assign n11551 = n1733 & ~n11550 ;
  assign n11552 = n1737 & ~n11551 ;
  assign n11553 = n1741 & ~n11552 ;
  assign n11554 = n1745 & ~n11553 ;
  assign n11555 = n1749 & ~n11554 ;
  assign n11556 = n1753 & ~n11555 ;
  assign n11557 = x183 & ~n1755 ;
  assign n11558 = ~n11556 & n11557 ;
  assign n11646 = n11558 & x311 ;
  assign n11559 = n1423 & ~n2097 ;
  assign n11560 = n1428 & ~n11559 ;
  assign n11561 = n1432 & ~n11560 ;
  assign n11562 = n1436 & ~n11561 ;
  assign n11563 = n1440 & ~n11562 ;
  assign n11564 = n1444 & ~n11563 ;
  assign n11565 = n1448 & ~n11564 ;
  assign n11566 = n1452 & ~n11565 ;
  assign n11567 = n1456 & ~n11566 ;
  assign n11568 = n1460 & ~n11567 ;
  assign n11569 = n1464 & ~n11568 ;
  assign n11570 = n1468 & ~n11569 ;
  assign n11571 = n1472 & ~n11570 ;
  assign n11572 = n1476 & ~n11571 ;
  assign n11573 = n1480 & ~n11572 ;
  assign n11574 = n1484 & ~n11573 ;
  assign n11575 = n1488 & ~n11574 ;
  assign n11576 = n1492 & ~n11575 ;
  assign n11577 = n1496 & ~n11576 ;
  assign n11578 = n1500 & ~n11577 ;
  assign n11579 = n1504 & ~n11578 ;
  assign n11580 = n1508 & ~n11579 ;
  assign n11581 = n1512 & ~n11580 ;
  assign n11582 = n1516 & ~n11581 ;
  assign n11583 = n1520 & ~n11582 ;
  assign n11584 = n1524 & ~n11583 ;
  assign n11585 = n1528 & ~n11584 ;
  assign n11586 = n1532 & ~n11585 ;
  assign n11587 = n1536 & ~n11586 ;
  assign n11588 = n1540 & ~n11587 ;
  assign n11589 = n1544 & ~n11588 ;
  assign n11590 = n1548 & ~n11589 ;
  assign n11591 = n1552 & ~n11590 ;
  assign n11592 = n1556 & ~n11591 ;
  assign n11593 = n1560 & ~n11592 ;
  assign n11594 = n1564 & ~n11593 ;
  assign n11595 = n1568 & ~n11594 ;
  assign n11596 = n1572 & ~n11595 ;
  assign n11597 = n1576 & ~n11596 ;
  assign n11598 = n1580 & ~n11597 ;
  assign n11599 = n1584 & ~n11598 ;
  assign n11600 = n1588 & ~n11599 ;
  assign n11601 = n1592 & ~n11600 ;
  assign n11602 = n1596 & ~n11601 ;
  assign n11603 = n1600 & ~n11602 ;
  assign n11604 = n1604 & ~n11603 ;
  assign n11605 = n1608 & ~n11604 ;
  assign n11606 = n1612 & ~n11605 ;
  assign n11607 = n2656 & ~n11606 ;
  assign n11608 = n2658 & ~n11607 ;
  assign n11609 = n3192 & ~n11608 ;
  assign n11610 = n1962 & ~n11609 ;
  assign n11611 = n1966 & ~n11610 ;
  assign n11612 = n1970 & ~n11611 ;
  assign n11613 = n1974 & ~n11612 ;
  assign n11614 = n1978 & ~n11613 ;
  assign n11615 = n1982 & ~n11614 ;
  assign n11616 = n1986 & ~n11615 ;
  assign n11617 = n1990 & ~n11616 ;
  assign n11618 = n1994 & ~n11617 ;
  assign n11619 = n1998 & ~n11618 ;
  assign n11620 = n2002 & ~n11619 ;
  assign n11621 = n2006 & ~n11620 ;
  assign n11622 = n2010 & ~n11621 ;
  assign n11623 = n2014 & ~n11622 ;
  assign n11624 = n2018 & ~n11623 ;
  assign n11625 = n2022 & ~n11624 ;
  assign n11626 = n2026 & ~n11625 ;
  assign n11627 = n2030 & ~n11626 ;
  assign n11628 = n2034 & ~n11627 ;
  assign n11629 = n2038 & ~n11628 ;
  assign n11630 = n2042 & ~n11629 ;
  assign n11631 = n2046 & ~n11630 ;
  assign n11632 = n2050 & ~n11631 ;
  assign n11633 = n2054 & ~n11632 ;
  assign n11634 = n2058 & ~n11633 ;
  assign n11635 = n2062 & ~n11634 ;
  assign n11636 = n2066 & ~n11635 ;
  assign n11637 = n2070 & ~n11636 ;
  assign n11638 = n2074 & ~n11637 ;
  assign n11639 = n2078 & ~n11638 ;
  assign n11640 = n2082 & ~n11639 ;
  assign n11641 = n2086 & ~n11640 ;
  assign n11642 = n2090 & ~n11641 ;
  assign n11643 = ~x183 & ~n2092 ;
  assign n11644 = ~n11642 & n11643 ;
  assign n11647 = ~n11644 & ~x311 ;
  assign n11648 = ~n11646 & ~n11647 ;
  assign n11649 = ~n406 & n1764 ;
  assign n11650 = n1769 & ~n11649 ;
  assign n11651 = n1773 & ~n11650 ;
  assign n11652 = n1777 & ~n11651 ;
  assign n11653 = n1781 & ~n11652 ;
  assign n11654 = n1785 & ~n11653 ;
  assign n11655 = n1789 & ~n11654 ;
  assign n11656 = n1793 & ~n11655 ;
  assign n11657 = n1797 & ~n11656 ;
  assign n11658 = n1801 & ~n11657 ;
  assign n11659 = n1805 & ~n11658 ;
  assign n11660 = n1809 & ~n11659 ;
  assign n11661 = n1813 & ~n11660 ;
  assign n11662 = n1817 & ~n11661 ;
  assign n11663 = n1821 & ~n11662 ;
  assign n11664 = n1825 & ~n11663 ;
  assign n11665 = n1829 & ~n11664 ;
  assign n11666 = n1833 & ~n11665 ;
  assign n11667 = n1837 & ~n11666 ;
  assign n11668 = n1841 & ~n11667 ;
  assign n11669 = n1845 & ~n11668 ;
  assign n11670 = n1849 & ~n11669 ;
  assign n11671 = n1853 & ~n11670 ;
  assign n11672 = n1857 & ~n11671 ;
  assign n11673 = n1861 & ~n11672 ;
  assign n11674 = n1865 & ~n11673 ;
  assign n11675 = n1869 & ~n11674 ;
  assign n11676 = n1873 & ~n11675 ;
  assign n11677 = n1877 & ~n11676 ;
  assign n11678 = n1881 & ~n11677 ;
  assign n11679 = n1885 & ~n11678 ;
  assign n11680 = n1889 & ~n11679 ;
  assign n11681 = n1893 & ~n11680 ;
  assign n11682 = n1897 & ~n11681 ;
  assign n11683 = n1901 & ~n11682 ;
  assign n11684 = n1905 & ~n11683 ;
  assign n11685 = n1909 & ~n11684 ;
  assign n11686 = n1913 & ~n11685 ;
  assign n11687 = n1917 & ~n11686 ;
  assign n11688 = n1921 & ~n11687 ;
  assign n11689 = n1925 & ~n11688 ;
  assign n11690 = n1929 & ~n11689 ;
  assign n11691 = n1933 & ~n11690 ;
  assign n11692 = n1937 & ~n11691 ;
  assign n11693 = n1941 & ~n11692 ;
  assign n11694 = n1945 & ~n11693 ;
  assign n11695 = n1949 & ~n11694 ;
  assign n11696 = n1953 & ~n11695 ;
  assign n11697 = n2749 & ~n11696 ;
  assign n11698 = n263 & ~n11697 ;
  assign n11699 = n267 & ~n11698 ;
  assign n11700 = n271 & ~n11699 ;
  assign n11701 = n275 & ~n11700 ;
  assign n11702 = n279 & ~n11701 ;
  assign n11703 = n283 & ~n11702 ;
  assign n11704 = n287 & ~n11703 ;
  assign n11705 = n291 & ~n11704 ;
  assign n11706 = n295 & ~n11705 ;
  assign n11707 = n299 & ~n11706 ;
  assign n11708 = n303 & ~n11707 ;
  assign n11709 = n307 & ~n11708 ;
  assign n11710 = n311 & ~n11709 ;
  assign n11711 = n315 & ~n11710 ;
  assign n11712 = n319 & ~n11711 ;
  assign n11713 = n323 & ~n11712 ;
  assign n11714 = n327 & ~n11713 ;
  assign n11715 = n331 & ~n11714 ;
  assign n11716 = n335 & ~n11715 ;
  assign n11717 = n339 & ~n11716 ;
  assign n11718 = n343 & ~n11717 ;
  assign n11719 = n347 & ~n11718 ;
  assign n11720 = n351 & ~n11719 ;
  assign n11721 = n355 & ~n11720 ;
  assign n11722 = n359 & ~n11721 ;
  assign n11723 = n363 & ~n11722 ;
  assign n11724 = n367 & ~n11723 ;
  assign n11725 = n371 & ~n11724 ;
  assign n11726 = n375 & ~n11725 ;
  assign n11727 = n379 & ~n11726 ;
  assign n11728 = n383 & ~n11727 ;
  assign n11729 = n387 & ~n11728 ;
  assign n11730 = n391 & ~n11729 ;
  assign n11731 = n395 & ~n11730 ;
  assign n11732 = n399 & ~n11731 ;
  assign n11733 = x184 & ~n401 ;
  assign n11734 = ~n11732 & n11733 ;
  assign n11822 = n11734 & x312 ;
  assign n11735 = ~n745 & n2101 ;
  assign n11736 = n2106 & ~n11735 ;
  assign n11737 = n2110 & ~n11736 ;
  assign n11738 = n2114 & ~n11737 ;
  assign n11739 = n2118 & ~n11738 ;
  assign n11740 = n2122 & ~n11739 ;
  assign n11741 = n2126 & ~n11740 ;
  assign n11742 = n2130 & ~n11741 ;
  assign n11743 = n2134 & ~n11742 ;
  assign n11744 = n2138 & ~n11743 ;
  assign n11745 = n2142 & ~n11744 ;
  assign n11746 = n2146 & ~n11745 ;
  assign n11747 = n2150 & ~n11746 ;
  assign n11748 = n2154 & ~n11747 ;
  assign n11749 = n2158 & ~n11748 ;
  assign n11750 = n2162 & ~n11749 ;
  assign n11751 = n2166 & ~n11750 ;
  assign n11752 = n2170 & ~n11751 ;
  assign n11753 = n2174 & ~n11752 ;
  assign n11754 = n2178 & ~n11753 ;
  assign n11755 = n2182 & ~n11754 ;
  assign n11756 = n2186 & ~n11755 ;
  assign n11757 = n2190 & ~n11756 ;
  assign n11758 = n2194 & ~n11757 ;
  assign n11759 = n2198 & ~n11758 ;
  assign n11760 = n2202 & ~n11759 ;
  assign n11761 = n2206 & ~n11760 ;
  assign n11762 = n2210 & ~n11761 ;
  assign n11763 = n2214 & ~n11762 ;
  assign n11764 = n2218 & ~n11763 ;
  assign n11765 = n2222 & ~n11764 ;
  assign n11766 = n2226 & ~n11765 ;
  assign n11767 = n2230 & ~n11766 ;
  assign n11768 = n2234 & ~n11767 ;
  assign n11769 = n2238 & ~n11768 ;
  assign n11770 = n2242 & ~n11769 ;
  assign n11771 = n2246 & ~n11770 ;
  assign n11772 = n2250 & ~n11771 ;
  assign n11773 = n2254 & ~n11772 ;
  assign n11774 = n2258 & ~n11773 ;
  assign n11775 = n2262 & ~n11774 ;
  assign n11776 = n2266 & ~n11775 ;
  assign n11777 = n2270 & ~n11776 ;
  assign n11778 = n2274 & ~n11777 ;
  assign n11779 = n2278 & ~n11778 ;
  assign n11780 = n2282 & ~n11779 ;
  assign n11781 = n2286 & ~n11780 ;
  assign n11782 = n2290 & ~n11781 ;
  assign n11783 = n2836 & ~n11782 ;
  assign n11784 = n602 & ~n11783 ;
  assign n11785 = n606 & ~n11784 ;
  assign n11786 = n610 & ~n11785 ;
  assign n11787 = n614 & ~n11786 ;
  assign n11788 = n618 & ~n11787 ;
  assign n11789 = n622 & ~n11788 ;
  assign n11790 = n626 & ~n11789 ;
  assign n11791 = n630 & ~n11790 ;
  assign n11792 = n634 & ~n11791 ;
  assign n11793 = n638 & ~n11792 ;
  assign n11794 = n642 & ~n11793 ;
  assign n11795 = n646 & ~n11794 ;
  assign n11796 = n650 & ~n11795 ;
  assign n11797 = n654 & ~n11796 ;
  assign n11798 = n658 & ~n11797 ;
  assign n11799 = n662 & ~n11798 ;
  assign n11800 = n666 & ~n11799 ;
  assign n11801 = n670 & ~n11800 ;
  assign n11802 = n674 & ~n11801 ;
  assign n11803 = n678 & ~n11802 ;
  assign n11804 = n682 & ~n11803 ;
  assign n11805 = n686 & ~n11804 ;
  assign n11806 = n690 & ~n11805 ;
  assign n11807 = n694 & ~n11806 ;
  assign n11808 = n698 & ~n11807 ;
  assign n11809 = n702 & ~n11808 ;
  assign n11810 = n706 & ~n11809 ;
  assign n11811 = n710 & ~n11810 ;
  assign n11812 = n714 & ~n11811 ;
  assign n11813 = n718 & ~n11812 ;
  assign n11814 = n722 & ~n11813 ;
  assign n11815 = n726 & ~n11814 ;
  assign n11816 = n730 & ~n11815 ;
  assign n11817 = n734 & ~n11816 ;
  assign n11818 = n738 & ~n11817 ;
  assign n11819 = ~x184 & ~n740 ;
  assign n11820 = ~n11818 & n11819 ;
  assign n11823 = ~n11820 & ~x312 ;
  assign n11824 = ~n11822 & ~n11823 ;
  assign n11825 = n410 & ~n1088 ;
  assign n11826 = n415 & ~n11825 ;
  assign n11827 = n419 & ~n11826 ;
  assign n11828 = n423 & ~n11827 ;
  assign n11829 = n427 & ~n11828 ;
  assign n11830 = n431 & ~n11829 ;
  assign n11831 = n435 & ~n11830 ;
  assign n11832 = n439 & ~n11831 ;
  assign n11833 = n443 & ~n11832 ;
  assign n11834 = n447 & ~n11833 ;
  assign n11835 = n451 & ~n11834 ;
  assign n11836 = n455 & ~n11835 ;
  assign n11837 = n459 & ~n11836 ;
  assign n11838 = n463 & ~n11837 ;
  assign n11839 = n467 & ~n11838 ;
  assign n11840 = n471 & ~n11839 ;
  assign n11841 = n475 & ~n11840 ;
  assign n11842 = n479 & ~n11841 ;
  assign n11843 = n483 & ~n11842 ;
  assign n11844 = n487 & ~n11843 ;
  assign n11845 = n491 & ~n11844 ;
  assign n11846 = n495 & ~n11845 ;
  assign n11847 = n499 & ~n11846 ;
  assign n11848 = n503 & ~n11847 ;
  assign n11849 = n507 & ~n11848 ;
  assign n11850 = n511 & ~n11849 ;
  assign n11851 = n515 & ~n11850 ;
  assign n11852 = n519 & ~n11851 ;
  assign n11853 = n523 & ~n11852 ;
  assign n11854 = n527 & ~n11853 ;
  assign n11855 = n531 & ~n11854 ;
  assign n11856 = n535 & ~n11855 ;
  assign n11857 = n539 & ~n11856 ;
  assign n11858 = n543 & ~n11857 ;
  assign n11859 = n547 & ~n11858 ;
  assign n11860 = n551 & ~n11859 ;
  assign n11861 = n555 & ~n11860 ;
  assign n11862 = n559 & ~n11861 ;
  assign n11863 = n563 & ~n11862 ;
  assign n11864 = n567 & ~n11863 ;
  assign n11865 = n571 & ~n11864 ;
  assign n11866 = n575 & ~n11865 ;
  assign n11867 = n579 & ~n11866 ;
  assign n11868 = n583 & ~n11867 ;
  assign n11869 = n587 & ~n11868 ;
  assign n11870 = n591 & ~n11869 ;
  assign n11871 = n2382 & ~n11870 ;
  assign n11872 = n2384 & ~n11871 ;
  assign n11873 = n2927 & ~n11872 ;
  assign n11874 = n945 & ~n11873 ;
  assign n11875 = n949 & ~n11874 ;
  assign n11876 = n953 & ~n11875 ;
  assign n11877 = n957 & ~n11876 ;
  assign n11878 = n961 & ~n11877 ;
  assign n11879 = n965 & ~n11878 ;
  assign n11880 = n969 & ~n11879 ;
  assign n11881 = n973 & ~n11880 ;
  assign n11882 = n977 & ~n11881 ;
  assign n11883 = n981 & ~n11882 ;
  assign n11884 = n985 & ~n11883 ;
  assign n11885 = n989 & ~n11884 ;
  assign n11886 = n993 & ~n11885 ;
  assign n11887 = n997 & ~n11886 ;
  assign n11888 = n1001 & ~n11887 ;
  assign n11889 = n1005 & ~n11888 ;
  assign n11890 = n1009 & ~n11889 ;
  assign n11891 = n1013 & ~n11890 ;
  assign n11892 = n1017 & ~n11891 ;
  assign n11893 = n1021 & ~n11892 ;
  assign n11894 = n1025 & ~n11893 ;
  assign n11895 = n1029 & ~n11894 ;
  assign n11896 = n1033 & ~n11895 ;
  assign n11897 = n1037 & ~n11896 ;
  assign n11898 = n1041 & ~n11897 ;
  assign n11899 = n1045 & ~n11898 ;
  assign n11900 = n1049 & ~n11899 ;
  assign n11901 = n1053 & ~n11900 ;
  assign n11902 = n1057 & ~n11901 ;
  assign n11903 = n1061 & ~n11902 ;
  assign n11904 = n1065 & ~n11903 ;
  assign n11905 = n1069 & ~n11904 ;
  assign n11906 = n1073 & ~n11905 ;
  assign n11907 = n1077 & ~n11906 ;
  assign n11908 = n1081 & ~n11907 ;
  assign n11909 = x185 & ~n1083 ;
  assign n11910 = ~n11908 & n11909 ;
  assign n11998 = n11910 & x313 ;
  assign n11911 = n749 & ~n1427 ;
  assign n11912 = n754 & ~n11911 ;
  assign n11913 = n758 & ~n11912 ;
  assign n11914 = n762 & ~n11913 ;
  assign n11915 = n766 & ~n11914 ;
  assign n11916 = n770 & ~n11915 ;
  assign n11917 = n774 & ~n11916 ;
  assign n11918 = n778 & ~n11917 ;
  assign n11919 = n782 & ~n11918 ;
  assign n11920 = n786 & ~n11919 ;
  assign n11921 = n790 & ~n11920 ;
  assign n11922 = n794 & ~n11921 ;
  assign n11923 = n798 & ~n11922 ;
  assign n11924 = n802 & ~n11923 ;
  assign n11925 = n806 & ~n11924 ;
  assign n11926 = n810 & ~n11925 ;
  assign n11927 = n814 & ~n11926 ;
  assign n11928 = n818 & ~n11927 ;
  assign n11929 = n822 & ~n11928 ;
  assign n11930 = n826 & ~n11929 ;
  assign n11931 = n830 & ~n11930 ;
  assign n11932 = n834 & ~n11931 ;
  assign n11933 = n838 & ~n11932 ;
  assign n11934 = n842 & ~n11933 ;
  assign n11935 = n846 & ~n11934 ;
  assign n11936 = n850 & ~n11935 ;
  assign n11937 = n854 & ~n11936 ;
  assign n11938 = n858 & ~n11937 ;
  assign n11939 = n862 & ~n11938 ;
  assign n11940 = n866 & ~n11939 ;
  assign n11941 = n870 & ~n11940 ;
  assign n11942 = n874 & ~n11941 ;
  assign n11943 = n878 & ~n11942 ;
  assign n11944 = n882 & ~n11943 ;
  assign n11945 = n886 & ~n11944 ;
  assign n11946 = n890 & ~n11945 ;
  assign n11947 = n894 & ~n11946 ;
  assign n11948 = n898 & ~n11947 ;
  assign n11949 = n902 & ~n11948 ;
  assign n11950 = n906 & ~n11949 ;
  assign n11951 = n910 & ~n11950 ;
  assign n11952 = n914 & ~n11951 ;
  assign n11953 = n918 & ~n11952 ;
  assign n11954 = n922 & ~n11953 ;
  assign n11955 = n926 & ~n11954 ;
  assign n11956 = n930 & ~n11955 ;
  assign n11957 = n2472 & ~n11956 ;
  assign n11958 = n2474 & ~n11957 ;
  assign n11959 = n3014 & ~n11958 ;
  assign n11960 = n1284 & ~n11959 ;
  assign n11961 = n1288 & ~n11960 ;
  assign n11962 = n1292 & ~n11961 ;
  assign n11963 = n1296 & ~n11962 ;
  assign n11964 = n1300 & ~n11963 ;
  assign n11965 = n1304 & ~n11964 ;
  assign n11966 = n1308 & ~n11965 ;
  assign n11967 = n1312 & ~n11966 ;
  assign n11968 = n1316 & ~n11967 ;
  assign n11969 = n1320 & ~n11968 ;
  assign n11970 = n1324 & ~n11969 ;
  assign n11971 = n1328 & ~n11970 ;
  assign n11972 = n1332 & ~n11971 ;
  assign n11973 = n1336 & ~n11972 ;
  assign n11974 = n1340 & ~n11973 ;
  assign n11975 = n1344 & ~n11974 ;
  assign n11976 = n1348 & ~n11975 ;
  assign n11977 = n1352 & ~n11976 ;
  assign n11978 = n1356 & ~n11977 ;
  assign n11979 = n1360 & ~n11978 ;
  assign n11980 = n1364 & ~n11979 ;
  assign n11981 = n1368 & ~n11980 ;
  assign n11982 = n1372 & ~n11981 ;
  assign n11983 = n1376 & ~n11982 ;
  assign n11984 = n1380 & ~n11983 ;
  assign n11985 = n1384 & ~n11984 ;
  assign n11986 = n1388 & ~n11985 ;
  assign n11987 = n1392 & ~n11986 ;
  assign n11988 = n1396 & ~n11987 ;
  assign n11989 = n1400 & ~n11988 ;
  assign n11990 = n1404 & ~n11989 ;
  assign n11991 = n1408 & ~n11990 ;
  assign n11992 = n1412 & ~n11991 ;
  assign n11993 = n1416 & ~n11992 ;
  assign n11994 = n1420 & ~n11993 ;
  assign n11995 = ~x185 & ~n1422 ;
  assign n11996 = ~n11994 & n11995 ;
  assign n11999 = ~n11996 & ~x313 ;
  assign n12000 = ~n11998 & ~n11999 ;
  assign n12001 = n1092 & ~n1768 ;
  assign n12002 = n1097 & ~n12001 ;
  assign n12003 = n1101 & ~n12002 ;
  assign n12004 = n1105 & ~n12003 ;
  assign n12005 = n1109 & ~n12004 ;
  assign n12006 = n1113 & ~n12005 ;
  assign n12007 = n1117 & ~n12006 ;
  assign n12008 = n1121 & ~n12007 ;
  assign n12009 = n1125 & ~n12008 ;
  assign n12010 = n1129 & ~n12009 ;
  assign n12011 = n1133 & ~n12010 ;
  assign n12012 = n1137 & ~n12011 ;
  assign n12013 = n1141 & ~n12012 ;
  assign n12014 = n1145 & ~n12013 ;
  assign n12015 = n1149 & ~n12014 ;
  assign n12016 = n1153 & ~n12015 ;
  assign n12017 = n1157 & ~n12016 ;
  assign n12018 = n1161 & ~n12017 ;
  assign n12019 = n1165 & ~n12018 ;
  assign n12020 = n1169 & ~n12019 ;
  assign n12021 = n1173 & ~n12020 ;
  assign n12022 = n1177 & ~n12021 ;
  assign n12023 = n1181 & ~n12022 ;
  assign n12024 = n1185 & ~n12023 ;
  assign n12025 = n1189 & ~n12024 ;
  assign n12026 = n1193 & ~n12025 ;
  assign n12027 = n1197 & ~n12026 ;
  assign n12028 = n1201 & ~n12027 ;
  assign n12029 = n1205 & ~n12028 ;
  assign n12030 = n1209 & ~n12029 ;
  assign n12031 = n1213 & ~n12030 ;
  assign n12032 = n1217 & ~n12031 ;
  assign n12033 = n1221 & ~n12032 ;
  assign n12034 = n1225 & ~n12033 ;
  assign n12035 = n1229 & ~n12034 ;
  assign n12036 = n1233 & ~n12035 ;
  assign n12037 = n1237 & ~n12036 ;
  assign n12038 = n1241 & ~n12037 ;
  assign n12039 = n1245 & ~n12038 ;
  assign n12040 = n1249 & ~n12039 ;
  assign n12041 = n1253 & ~n12040 ;
  assign n12042 = n1257 & ~n12041 ;
  assign n12043 = n1261 & ~n12042 ;
  assign n12044 = n1265 & ~n12043 ;
  assign n12045 = n1269 & ~n12044 ;
  assign n12046 = n1273 & ~n12045 ;
  assign n12047 = n2566 & ~n12046 ;
  assign n12048 = n2568 & ~n12047 ;
  assign n12049 = n3105 & ~n12048 ;
  assign n12050 = n1625 & ~n12049 ;
  assign n12051 = n1629 & ~n12050 ;
  assign n12052 = n1633 & ~n12051 ;
  assign n12053 = n1637 & ~n12052 ;
  assign n12054 = n1641 & ~n12053 ;
  assign n12055 = n1645 & ~n12054 ;
  assign n12056 = n1649 & ~n12055 ;
  assign n12057 = n1653 & ~n12056 ;
  assign n12058 = n1657 & ~n12057 ;
  assign n12059 = n1661 & ~n12058 ;
  assign n12060 = n1665 & ~n12059 ;
  assign n12061 = n1669 & ~n12060 ;
  assign n12062 = n1673 & ~n12061 ;
  assign n12063 = n1677 & ~n12062 ;
  assign n12064 = n1681 & ~n12063 ;
  assign n12065 = n1685 & ~n12064 ;
  assign n12066 = n1689 & ~n12065 ;
  assign n12067 = n1693 & ~n12066 ;
  assign n12068 = n1697 & ~n12067 ;
  assign n12069 = n1701 & ~n12068 ;
  assign n12070 = n1705 & ~n12069 ;
  assign n12071 = n1709 & ~n12070 ;
  assign n12072 = n1713 & ~n12071 ;
  assign n12073 = n1717 & ~n12072 ;
  assign n12074 = n1721 & ~n12073 ;
  assign n12075 = n1725 & ~n12074 ;
  assign n12076 = n1729 & ~n12075 ;
  assign n12077 = n1733 & ~n12076 ;
  assign n12078 = n1737 & ~n12077 ;
  assign n12079 = n1741 & ~n12078 ;
  assign n12080 = n1745 & ~n12079 ;
  assign n12081 = n1749 & ~n12080 ;
  assign n12082 = n1753 & ~n12081 ;
  assign n12083 = n1757 & ~n12082 ;
  assign n12084 = n1761 & ~n12083 ;
  assign n12085 = x186 & ~n1763 ;
  assign n12086 = ~n12084 & n12085 ;
  assign n12174 = n12086 & x314 ;
  assign n12087 = n1431 & ~n2105 ;
  assign n12088 = n1436 & ~n12087 ;
  assign n12089 = n1440 & ~n12088 ;
  assign n12090 = n1444 & ~n12089 ;
  assign n12091 = n1448 & ~n12090 ;
  assign n12092 = n1452 & ~n12091 ;
  assign n12093 = n1456 & ~n12092 ;
  assign n12094 = n1460 & ~n12093 ;
  assign n12095 = n1464 & ~n12094 ;
  assign n12096 = n1468 & ~n12095 ;
  assign n12097 = n1472 & ~n12096 ;
  assign n12098 = n1476 & ~n12097 ;
  assign n12099 = n1480 & ~n12098 ;
  assign n12100 = n1484 & ~n12099 ;
  assign n12101 = n1488 & ~n12100 ;
  assign n12102 = n1492 & ~n12101 ;
  assign n12103 = n1496 & ~n12102 ;
  assign n12104 = n1500 & ~n12103 ;
  assign n12105 = n1504 & ~n12104 ;
  assign n12106 = n1508 & ~n12105 ;
  assign n12107 = n1512 & ~n12106 ;
  assign n12108 = n1516 & ~n12107 ;
  assign n12109 = n1520 & ~n12108 ;
  assign n12110 = n1524 & ~n12109 ;
  assign n12111 = n1528 & ~n12110 ;
  assign n12112 = n1532 & ~n12111 ;
  assign n12113 = n1536 & ~n12112 ;
  assign n12114 = n1540 & ~n12113 ;
  assign n12115 = n1544 & ~n12114 ;
  assign n12116 = n1548 & ~n12115 ;
  assign n12117 = n1552 & ~n12116 ;
  assign n12118 = n1556 & ~n12117 ;
  assign n12119 = n1560 & ~n12118 ;
  assign n12120 = n1564 & ~n12119 ;
  assign n12121 = n1568 & ~n12120 ;
  assign n12122 = n1572 & ~n12121 ;
  assign n12123 = n1576 & ~n12122 ;
  assign n12124 = n1580 & ~n12123 ;
  assign n12125 = n1584 & ~n12124 ;
  assign n12126 = n1588 & ~n12125 ;
  assign n12127 = n1592 & ~n12126 ;
  assign n12128 = n1596 & ~n12127 ;
  assign n12129 = n1600 & ~n12128 ;
  assign n12130 = n1604 & ~n12129 ;
  assign n12131 = n1608 & ~n12130 ;
  assign n12132 = n1612 & ~n12131 ;
  assign n12133 = n2656 & ~n12132 ;
  assign n12134 = n2658 & ~n12133 ;
  assign n12135 = n3192 & ~n12134 ;
  assign n12136 = n1962 & ~n12135 ;
  assign n12137 = n1966 & ~n12136 ;
  assign n12138 = n1970 & ~n12137 ;
  assign n12139 = n1974 & ~n12138 ;
  assign n12140 = n1978 & ~n12139 ;
  assign n12141 = n1982 & ~n12140 ;
  assign n12142 = n1986 & ~n12141 ;
  assign n12143 = n1990 & ~n12142 ;
  assign n12144 = n1994 & ~n12143 ;
  assign n12145 = n1998 & ~n12144 ;
  assign n12146 = n2002 & ~n12145 ;
  assign n12147 = n2006 & ~n12146 ;
  assign n12148 = n2010 & ~n12147 ;
  assign n12149 = n2014 & ~n12148 ;
  assign n12150 = n2018 & ~n12149 ;
  assign n12151 = n2022 & ~n12150 ;
  assign n12152 = n2026 & ~n12151 ;
  assign n12153 = n2030 & ~n12152 ;
  assign n12154 = n2034 & ~n12153 ;
  assign n12155 = n2038 & ~n12154 ;
  assign n12156 = n2042 & ~n12155 ;
  assign n12157 = n2046 & ~n12156 ;
  assign n12158 = n2050 & ~n12157 ;
  assign n12159 = n2054 & ~n12158 ;
  assign n12160 = n2058 & ~n12159 ;
  assign n12161 = n2062 & ~n12160 ;
  assign n12162 = n2066 & ~n12161 ;
  assign n12163 = n2070 & ~n12162 ;
  assign n12164 = n2074 & ~n12163 ;
  assign n12165 = n2078 & ~n12164 ;
  assign n12166 = n2082 & ~n12165 ;
  assign n12167 = n2086 & ~n12166 ;
  assign n12168 = n2090 & ~n12167 ;
  assign n12169 = n2094 & ~n12168 ;
  assign n12170 = n2098 & ~n12169 ;
  assign n12171 = ~x186 & ~n2100 ;
  assign n12172 = ~n12170 & n12171 ;
  assign n12175 = ~n12172 & ~x314 ;
  assign n12176 = ~n12174 & ~n12175 ;
  assign n12177 = ~n414 & n1772 ;
  assign n12178 = n1777 & ~n12177 ;
  assign n12179 = n1781 & ~n12178 ;
  assign n12180 = n1785 & ~n12179 ;
  assign n12181 = n1789 & ~n12180 ;
  assign n12182 = n1793 & ~n12181 ;
  assign n12183 = n1797 & ~n12182 ;
  assign n12184 = n1801 & ~n12183 ;
  assign n12185 = n1805 & ~n12184 ;
  assign n12186 = n1809 & ~n12185 ;
  assign n12187 = n1813 & ~n12186 ;
  assign n12188 = n1817 & ~n12187 ;
  assign n12189 = n1821 & ~n12188 ;
  assign n12190 = n1825 & ~n12189 ;
  assign n12191 = n1829 & ~n12190 ;
  assign n12192 = n1833 & ~n12191 ;
  assign n12193 = n1837 & ~n12192 ;
  assign n12194 = n1841 & ~n12193 ;
  assign n12195 = n1845 & ~n12194 ;
  assign n12196 = n1849 & ~n12195 ;
  assign n12197 = n1853 & ~n12196 ;
  assign n12198 = n1857 & ~n12197 ;
  assign n12199 = n1861 & ~n12198 ;
  assign n12200 = n1865 & ~n12199 ;
  assign n12201 = n1869 & ~n12200 ;
  assign n12202 = n1873 & ~n12201 ;
  assign n12203 = n1877 & ~n12202 ;
  assign n12204 = n1881 & ~n12203 ;
  assign n12205 = n1885 & ~n12204 ;
  assign n12206 = n1889 & ~n12205 ;
  assign n12207 = n1893 & ~n12206 ;
  assign n12208 = n1897 & ~n12207 ;
  assign n12209 = n1901 & ~n12208 ;
  assign n12210 = n1905 & ~n12209 ;
  assign n12211 = n1909 & ~n12210 ;
  assign n12212 = n1913 & ~n12211 ;
  assign n12213 = n1917 & ~n12212 ;
  assign n12214 = n1921 & ~n12213 ;
  assign n12215 = n1925 & ~n12214 ;
  assign n12216 = n1929 & ~n12215 ;
  assign n12217 = n1933 & ~n12216 ;
  assign n12218 = n1937 & ~n12217 ;
  assign n12219 = n1941 & ~n12218 ;
  assign n12220 = n1945 & ~n12219 ;
  assign n12221 = n1949 & ~n12220 ;
  assign n12222 = n1953 & ~n12221 ;
  assign n12223 = n2749 & ~n12222 ;
  assign n12224 = n263 & ~n12223 ;
  assign n12225 = n267 & ~n12224 ;
  assign n12226 = n271 & ~n12225 ;
  assign n12227 = n275 & ~n12226 ;
  assign n12228 = n279 & ~n12227 ;
  assign n12229 = n283 & ~n12228 ;
  assign n12230 = n287 & ~n12229 ;
  assign n12231 = n291 & ~n12230 ;
  assign n12232 = n295 & ~n12231 ;
  assign n12233 = n299 & ~n12232 ;
  assign n12234 = n303 & ~n12233 ;
  assign n12235 = n307 & ~n12234 ;
  assign n12236 = n311 & ~n12235 ;
  assign n12237 = n315 & ~n12236 ;
  assign n12238 = n319 & ~n12237 ;
  assign n12239 = n323 & ~n12238 ;
  assign n12240 = n327 & ~n12239 ;
  assign n12241 = n331 & ~n12240 ;
  assign n12242 = n335 & ~n12241 ;
  assign n12243 = n339 & ~n12242 ;
  assign n12244 = n343 & ~n12243 ;
  assign n12245 = n347 & ~n12244 ;
  assign n12246 = n351 & ~n12245 ;
  assign n12247 = n355 & ~n12246 ;
  assign n12248 = n359 & ~n12247 ;
  assign n12249 = n363 & ~n12248 ;
  assign n12250 = n367 & ~n12249 ;
  assign n12251 = n371 & ~n12250 ;
  assign n12252 = n375 & ~n12251 ;
  assign n12253 = n379 & ~n12252 ;
  assign n12254 = n383 & ~n12253 ;
  assign n12255 = n387 & ~n12254 ;
  assign n12256 = n391 & ~n12255 ;
  assign n12257 = n395 & ~n12256 ;
  assign n12258 = n399 & ~n12257 ;
  assign n12259 = n403 & ~n12258 ;
  assign n12260 = n407 & ~n12259 ;
  assign n12261 = x187 & ~n409 ;
  assign n12262 = ~n12260 & n12261 ;
  assign n12350 = n12262 & x315 ;
  assign n12263 = ~n753 & n2109 ;
  assign n12264 = n2114 & ~n12263 ;
  assign n12265 = n2118 & ~n12264 ;
  assign n12266 = n2122 & ~n12265 ;
  assign n12267 = n2126 & ~n12266 ;
  assign n12268 = n2130 & ~n12267 ;
  assign n12269 = n2134 & ~n12268 ;
  assign n12270 = n2138 & ~n12269 ;
  assign n12271 = n2142 & ~n12270 ;
  assign n12272 = n2146 & ~n12271 ;
  assign n12273 = n2150 & ~n12272 ;
  assign n12274 = n2154 & ~n12273 ;
  assign n12275 = n2158 & ~n12274 ;
  assign n12276 = n2162 & ~n12275 ;
  assign n12277 = n2166 & ~n12276 ;
  assign n12278 = n2170 & ~n12277 ;
  assign n12279 = n2174 & ~n12278 ;
  assign n12280 = n2178 & ~n12279 ;
  assign n12281 = n2182 & ~n12280 ;
  assign n12282 = n2186 & ~n12281 ;
  assign n12283 = n2190 & ~n12282 ;
  assign n12284 = n2194 & ~n12283 ;
  assign n12285 = n2198 & ~n12284 ;
  assign n12286 = n2202 & ~n12285 ;
  assign n12287 = n2206 & ~n12286 ;
  assign n12288 = n2210 & ~n12287 ;
  assign n12289 = n2214 & ~n12288 ;
  assign n12290 = n2218 & ~n12289 ;
  assign n12291 = n2222 & ~n12290 ;
  assign n12292 = n2226 & ~n12291 ;
  assign n12293 = n2230 & ~n12292 ;
  assign n12294 = n2234 & ~n12293 ;
  assign n12295 = n2238 & ~n12294 ;
  assign n12296 = n2242 & ~n12295 ;
  assign n12297 = n2246 & ~n12296 ;
  assign n12298 = n2250 & ~n12297 ;
  assign n12299 = n2254 & ~n12298 ;
  assign n12300 = n2258 & ~n12299 ;
  assign n12301 = n2262 & ~n12300 ;
  assign n12302 = n2266 & ~n12301 ;
  assign n12303 = n2270 & ~n12302 ;
  assign n12304 = n2274 & ~n12303 ;
  assign n12305 = n2278 & ~n12304 ;
  assign n12306 = n2282 & ~n12305 ;
  assign n12307 = n2286 & ~n12306 ;
  assign n12308 = n2290 & ~n12307 ;
  assign n12309 = n2836 & ~n12308 ;
  assign n12310 = n602 & ~n12309 ;
  assign n12311 = n606 & ~n12310 ;
  assign n12312 = n610 & ~n12311 ;
  assign n12313 = n614 & ~n12312 ;
  assign n12314 = n618 & ~n12313 ;
  assign n12315 = n622 & ~n12314 ;
  assign n12316 = n626 & ~n12315 ;
  assign n12317 = n630 & ~n12316 ;
  assign n12318 = n634 & ~n12317 ;
  assign n12319 = n638 & ~n12318 ;
  assign n12320 = n642 & ~n12319 ;
  assign n12321 = n646 & ~n12320 ;
  assign n12322 = n650 & ~n12321 ;
  assign n12323 = n654 & ~n12322 ;
  assign n12324 = n658 & ~n12323 ;
  assign n12325 = n662 & ~n12324 ;
  assign n12326 = n666 & ~n12325 ;
  assign n12327 = n670 & ~n12326 ;
  assign n12328 = n674 & ~n12327 ;
  assign n12329 = n678 & ~n12328 ;
  assign n12330 = n682 & ~n12329 ;
  assign n12331 = n686 & ~n12330 ;
  assign n12332 = n690 & ~n12331 ;
  assign n12333 = n694 & ~n12332 ;
  assign n12334 = n698 & ~n12333 ;
  assign n12335 = n702 & ~n12334 ;
  assign n12336 = n706 & ~n12335 ;
  assign n12337 = n710 & ~n12336 ;
  assign n12338 = n714 & ~n12337 ;
  assign n12339 = n718 & ~n12338 ;
  assign n12340 = n722 & ~n12339 ;
  assign n12341 = n726 & ~n12340 ;
  assign n12342 = n730 & ~n12341 ;
  assign n12343 = n734 & ~n12342 ;
  assign n12344 = n738 & ~n12343 ;
  assign n12345 = n742 & ~n12344 ;
  assign n12346 = n746 & ~n12345 ;
  assign n12347 = ~x187 & ~n748 ;
  assign n12348 = ~n12346 & n12347 ;
  assign n12351 = ~n12348 & ~x315 ;
  assign n12352 = ~n12350 & ~n12351 ;
  assign n12353 = n418 & ~n1096 ;
  assign n12354 = n423 & ~n12353 ;
  assign n12355 = n427 & ~n12354 ;
  assign n12356 = n431 & ~n12355 ;
  assign n12357 = n435 & ~n12356 ;
  assign n12358 = n439 & ~n12357 ;
  assign n12359 = n443 & ~n12358 ;
  assign n12360 = n447 & ~n12359 ;
  assign n12361 = n451 & ~n12360 ;
  assign n12362 = n455 & ~n12361 ;
  assign n12363 = n459 & ~n12362 ;
  assign n12364 = n463 & ~n12363 ;
  assign n12365 = n467 & ~n12364 ;
  assign n12366 = n471 & ~n12365 ;
  assign n12367 = n475 & ~n12366 ;
  assign n12368 = n479 & ~n12367 ;
  assign n12369 = n483 & ~n12368 ;
  assign n12370 = n487 & ~n12369 ;
  assign n12371 = n491 & ~n12370 ;
  assign n12372 = n495 & ~n12371 ;
  assign n12373 = n499 & ~n12372 ;
  assign n12374 = n503 & ~n12373 ;
  assign n12375 = n507 & ~n12374 ;
  assign n12376 = n511 & ~n12375 ;
  assign n12377 = n515 & ~n12376 ;
  assign n12378 = n519 & ~n12377 ;
  assign n12379 = n523 & ~n12378 ;
  assign n12380 = n527 & ~n12379 ;
  assign n12381 = n531 & ~n12380 ;
  assign n12382 = n535 & ~n12381 ;
  assign n12383 = n539 & ~n12382 ;
  assign n12384 = n543 & ~n12383 ;
  assign n12385 = n547 & ~n12384 ;
  assign n12386 = n551 & ~n12385 ;
  assign n12387 = n555 & ~n12386 ;
  assign n12388 = n559 & ~n12387 ;
  assign n12389 = n563 & ~n12388 ;
  assign n12390 = n567 & ~n12389 ;
  assign n12391 = n571 & ~n12390 ;
  assign n12392 = n575 & ~n12391 ;
  assign n12393 = n579 & ~n12392 ;
  assign n12394 = n583 & ~n12393 ;
  assign n12395 = n587 & ~n12394 ;
  assign n12396 = n591 & ~n12395 ;
  assign n12397 = n2382 & ~n12396 ;
  assign n12398 = n2384 & ~n12397 ;
  assign n12399 = n2927 & ~n12398 ;
  assign n12400 = n945 & ~n12399 ;
  assign n12401 = n949 & ~n12400 ;
  assign n12402 = n953 & ~n12401 ;
  assign n12403 = n957 & ~n12402 ;
  assign n12404 = n961 & ~n12403 ;
  assign n12405 = n965 & ~n12404 ;
  assign n12406 = n969 & ~n12405 ;
  assign n12407 = n973 & ~n12406 ;
  assign n12408 = n977 & ~n12407 ;
  assign n12409 = n981 & ~n12408 ;
  assign n12410 = n985 & ~n12409 ;
  assign n12411 = n989 & ~n12410 ;
  assign n12412 = n993 & ~n12411 ;
  assign n12413 = n997 & ~n12412 ;
  assign n12414 = n1001 & ~n12413 ;
  assign n12415 = n1005 & ~n12414 ;
  assign n12416 = n1009 & ~n12415 ;
  assign n12417 = n1013 & ~n12416 ;
  assign n12418 = n1017 & ~n12417 ;
  assign n12419 = n1021 & ~n12418 ;
  assign n12420 = n1025 & ~n12419 ;
  assign n12421 = n1029 & ~n12420 ;
  assign n12422 = n1033 & ~n12421 ;
  assign n12423 = n1037 & ~n12422 ;
  assign n12424 = n1041 & ~n12423 ;
  assign n12425 = n1045 & ~n12424 ;
  assign n12426 = n1049 & ~n12425 ;
  assign n12427 = n1053 & ~n12426 ;
  assign n12428 = n1057 & ~n12427 ;
  assign n12429 = n1061 & ~n12428 ;
  assign n12430 = n1065 & ~n12429 ;
  assign n12431 = n1069 & ~n12430 ;
  assign n12432 = n1073 & ~n12431 ;
  assign n12433 = n1077 & ~n12432 ;
  assign n12434 = n1081 & ~n12433 ;
  assign n12435 = n1085 & ~n12434 ;
  assign n12436 = n1089 & ~n12435 ;
  assign n12437 = x188 & ~n1091 ;
  assign n12438 = ~n12436 & n12437 ;
  assign n12526 = n12438 & x316 ;
  assign n12439 = n757 & ~n1435 ;
  assign n12440 = n762 & ~n12439 ;
  assign n12441 = n766 & ~n12440 ;
  assign n12442 = n770 & ~n12441 ;
  assign n12443 = n774 & ~n12442 ;
  assign n12444 = n778 & ~n12443 ;
  assign n12445 = n782 & ~n12444 ;
  assign n12446 = n786 & ~n12445 ;
  assign n12447 = n790 & ~n12446 ;
  assign n12448 = n794 & ~n12447 ;
  assign n12449 = n798 & ~n12448 ;
  assign n12450 = n802 & ~n12449 ;
  assign n12451 = n806 & ~n12450 ;
  assign n12452 = n810 & ~n12451 ;
  assign n12453 = n814 & ~n12452 ;
  assign n12454 = n818 & ~n12453 ;
  assign n12455 = n822 & ~n12454 ;
  assign n12456 = n826 & ~n12455 ;
  assign n12457 = n830 & ~n12456 ;
  assign n12458 = n834 & ~n12457 ;
  assign n12459 = n838 & ~n12458 ;
  assign n12460 = n842 & ~n12459 ;
  assign n12461 = n846 & ~n12460 ;
  assign n12462 = n850 & ~n12461 ;
  assign n12463 = n854 & ~n12462 ;
  assign n12464 = n858 & ~n12463 ;
  assign n12465 = n862 & ~n12464 ;
  assign n12466 = n866 & ~n12465 ;
  assign n12467 = n870 & ~n12466 ;
  assign n12468 = n874 & ~n12467 ;
  assign n12469 = n878 & ~n12468 ;
  assign n12470 = n882 & ~n12469 ;
  assign n12471 = n886 & ~n12470 ;
  assign n12472 = n890 & ~n12471 ;
  assign n12473 = n894 & ~n12472 ;
  assign n12474 = n898 & ~n12473 ;
  assign n12475 = n902 & ~n12474 ;
  assign n12476 = n906 & ~n12475 ;
  assign n12477 = n910 & ~n12476 ;
  assign n12478 = n914 & ~n12477 ;
  assign n12479 = n918 & ~n12478 ;
  assign n12480 = n922 & ~n12479 ;
  assign n12481 = n926 & ~n12480 ;
  assign n12482 = n930 & ~n12481 ;
  assign n12483 = n2472 & ~n12482 ;
  assign n12484 = n2474 & ~n12483 ;
  assign n12485 = n3014 & ~n12484 ;
  assign n12486 = n1284 & ~n12485 ;
  assign n12487 = n1288 & ~n12486 ;
  assign n12488 = n1292 & ~n12487 ;
  assign n12489 = n1296 & ~n12488 ;
  assign n12490 = n1300 & ~n12489 ;
  assign n12491 = n1304 & ~n12490 ;
  assign n12492 = n1308 & ~n12491 ;
  assign n12493 = n1312 & ~n12492 ;
  assign n12494 = n1316 & ~n12493 ;
  assign n12495 = n1320 & ~n12494 ;
  assign n12496 = n1324 & ~n12495 ;
  assign n12497 = n1328 & ~n12496 ;
  assign n12498 = n1332 & ~n12497 ;
  assign n12499 = n1336 & ~n12498 ;
  assign n12500 = n1340 & ~n12499 ;
  assign n12501 = n1344 & ~n12500 ;
  assign n12502 = n1348 & ~n12501 ;
  assign n12503 = n1352 & ~n12502 ;
  assign n12504 = n1356 & ~n12503 ;
  assign n12505 = n1360 & ~n12504 ;
  assign n12506 = n1364 & ~n12505 ;
  assign n12507 = n1368 & ~n12506 ;
  assign n12508 = n1372 & ~n12507 ;
  assign n12509 = n1376 & ~n12508 ;
  assign n12510 = n1380 & ~n12509 ;
  assign n12511 = n1384 & ~n12510 ;
  assign n12512 = n1388 & ~n12511 ;
  assign n12513 = n1392 & ~n12512 ;
  assign n12514 = n1396 & ~n12513 ;
  assign n12515 = n1400 & ~n12514 ;
  assign n12516 = n1404 & ~n12515 ;
  assign n12517 = n1408 & ~n12516 ;
  assign n12518 = n1412 & ~n12517 ;
  assign n12519 = n1416 & ~n12518 ;
  assign n12520 = n1420 & ~n12519 ;
  assign n12521 = n1424 & ~n12520 ;
  assign n12522 = n1428 & ~n12521 ;
  assign n12523 = ~x188 & ~n1430 ;
  assign n12524 = ~n12522 & n12523 ;
  assign n12527 = ~n12524 & ~x316 ;
  assign n12528 = ~n12526 & ~n12527 ;
  assign n12529 = n1100 & ~n1776 ;
  assign n12530 = n1105 & ~n12529 ;
  assign n12531 = n1109 & ~n12530 ;
  assign n12532 = n1113 & ~n12531 ;
  assign n12533 = n1117 & ~n12532 ;
  assign n12534 = n1121 & ~n12533 ;
  assign n12535 = n1125 & ~n12534 ;
  assign n12536 = n1129 & ~n12535 ;
  assign n12537 = n1133 & ~n12536 ;
  assign n12538 = n1137 & ~n12537 ;
  assign n12539 = n1141 & ~n12538 ;
  assign n12540 = n1145 & ~n12539 ;
  assign n12541 = n1149 & ~n12540 ;
  assign n12542 = n1153 & ~n12541 ;
  assign n12543 = n1157 & ~n12542 ;
  assign n12544 = n1161 & ~n12543 ;
  assign n12545 = n1165 & ~n12544 ;
  assign n12546 = n1169 & ~n12545 ;
  assign n12547 = n1173 & ~n12546 ;
  assign n12548 = n1177 & ~n12547 ;
  assign n12549 = n1181 & ~n12548 ;
  assign n12550 = n1185 & ~n12549 ;
  assign n12551 = n1189 & ~n12550 ;
  assign n12552 = n1193 & ~n12551 ;
  assign n12553 = n1197 & ~n12552 ;
  assign n12554 = n1201 & ~n12553 ;
  assign n12555 = n1205 & ~n12554 ;
  assign n12556 = n1209 & ~n12555 ;
  assign n12557 = n1213 & ~n12556 ;
  assign n12558 = n1217 & ~n12557 ;
  assign n12559 = n1221 & ~n12558 ;
  assign n12560 = n1225 & ~n12559 ;
  assign n12561 = n1229 & ~n12560 ;
  assign n12562 = n1233 & ~n12561 ;
  assign n12563 = n1237 & ~n12562 ;
  assign n12564 = n1241 & ~n12563 ;
  assign n12565 = n1245 & ~n12564 ;
  assign n12566 = n1249 & ~n12565 ;
  assign n12567 = n1253 & ~n12566 ;
  assign n12568 = n1257 & ~n12567 ;
  assign n12569 = n1261 & ~n12568 ;
  assign n12570 = n1265 & ~n12569 ;
  assign n12571 = n1269 & ~n12570 ;
  assign n12572 = n1273 & ~n12571 ;
  assign n12573 = n2566 & ~n12572 ;
  assign n12574 = n2568 & ~n12573 ;
  assign n12575 = n3105 & ~n12574 ;
  assign n12576 = n1625 & ~n12575 ;
  assign n12577 = n1629 & ~n12576 ;
  assign n12578 = n1633 & ~n12577 ;
  assign n12579 = n1637 & ~n12578 ;
  assign n12580 = n1641 & ~n12579 ;
  assign n12581 = n1645 & ~n12580 ;
  assign n12582 = n1649 & ~n12581 ;
  assign n12583 = n1653 & ~n12582 ;
  assign n12584 = n1657 & ~n12583 ;
  assign n12585 = n1661 & ~n12584 ;
  assign n12586 = n1665 & ~n12585 ;
  assign n12587 = n1669 & ~n12586 ;
  assign n12588 = n1673 & ~n12587 ;
  assign n12589 = n1677 & ~n12588 ;
  assign n12590 = n1681 & ~n12589 ;
  assign n12591 = n1685 & ~n12590 ;
  assign n12592 = n1689 & ~n12591 ;
  assign n12593 = n1693 & ~n12592 ;
  assign n12594 = n1697 & ~n12593 ;
  assign n12595 = n1701 & ~n12594 ;
  assign n12596 = n1705 & ~n12595 ;
  assign n12597 = n1709 & ~n12596 ;
  assign n12598 = n1713 & ~n12597 ;
  assign n12599 = n1717 & ~n12598 ;
  assign n12600 = n1721 & ~n12599 ;
  assign n12601 = n1725 & ~n12600 ;
  assign n12602 = n1729 & ~n12601 ;
  assign n12603 = n1733 & ~n12602 ;
  assign n12604 = n1737 & ~n12603 ;
  assign n12605 = n1741 & ~n12604 ;
  assign n12606 = n1745 & ~n12605 ;
  assign n12607 = n1749 & ~n12606 ;
  assign n12608 = n1753 & ~n12607 ;
  assign n12609 = n1757 & ~n12608 ;
  assign n12610 = n1761 & ~n12609 ;
  assign n12611 = n1765 & ~n12610 ;
  assign n12612 = n1769 & ~n12611 ;
  assign n12613 = x189 & ~n1771 ;
  assign n12614 = ~n12612 & n12613 ;
  assign n12702 = n12614 & x317 ;
  assign n12615 = n1439 & ~n2113 ;
  assign n12616 = n1444 & ~n12615 ;
  assign n12617 = n1448 & ~n12616 ;
  assign n12618 = n1452 & ~n12617 ;
  assign n12619 = n1456 & ~n12618 ;
  assign n12620 = n1460 & ~n12619 ;
  assign n12621 = n1464 & ~n12620 ;
  assign n12622 = n1468 & ~n12621 ;
  assign n12623 = n1472 & ~n12622 ;
  assign n12624 = n1476 & ~n12623 ;
  assign n12625 = n1480 & ~n12624 ;
  assign n12626 = n1484 & ~n12625 ;
  assign n12627 = n1488 & ~n12626 ;
  assign n12628 = n1492 & ~n12627 ;
  assign n12629 = n1496 & ~n12628 ;
  assign n12630 = n1500 & ~n12629 ;
  assign n12631 = n1504 & ~n12630 ;
  assign n12632 = n1508 & ~n12631 ;
  assign n12633 = n1512 & ~n12632 ;
  assign n12634 = n1516 & ~n12633 ;
  assign n12635 = n1520 & ~n12634 ;
  assign n12636 = n1524 & ~n12635 ;
  assign n12637 = n1528 & ~n12636 ;
  assign n12638 = n1532 & ~n12637 ;
  assign n12639 = n1536 & ~n12638 ;
  assign n12640 = n1540 & ~n12639 ;
  assign n12641 = n1544 & ~n12640 ;
  assign n12642 = n1548 & ~n12641 ;
  assign n12643 = n1552 & ~n12642 ;
  assign n12644 = n1556 & ~n12643 ;
  assign n12645 = n1560 & ~n12644 ;
  assign n12646 = n1564 & ~n12645 ;
  assign n12647 = n1568 & ~n12646 ;
  assign n12648 = n1572 & ~n12647 ;
  assign n12649 = n1576 & ~n12648 ;
  assign n12650 = n1580 & ~n12649 ;
  assign n12651 = n1584 & ~n12650 ;
  assign n12652 = n1588 & ~n12651 ;
  assign n12653 = n1592 & ~n12652 ;
  assign n12654 = n1596 & ~n12653 ;
  assign n12655 = n1600 & ~n12654 ;
  assign n12656 = n1604 & ~n12655 ;
  assign n12657 = n1608 & ~n12656 ;
  assign n12658 = n1612 & ~n12657 ;
  assign n12659 = n2656 & ~n12658 ;
  assign n12660 = n2658 & ~n12659 ;
  assign n12661 = n3192 & ~n12660 ;
  assign n12662 = n1962 & ~n12661 ;
  assign n12663 = n1966 & ~n12662 ;
  assign n12664 = n1970 & ~n12663 ;
  assign n12665 = n1974 & ~n12664 ;
  assign n12666 = n1978 & ~n12665 ;
  assign n12667 = n1982 & ~n12666 ;
  assign n12668 = n1986 & ~n12667 ;
  assign n12669 = n1990 & ~n12668 ;
  assign n12670 = n1994 & ~n12669 ;
  assign n12671 = n1998 & ~n12670 ;
  assign n12672 = n2002 & ~n12671 ;
  assign n12673 = n2006 & ~n12672 ;
  assign n12674 = n2010 & ~n12673 ;
  assign n12675 = n2014 & ~n12674 ;
  assign n12676 = n2018 & ~n12675 ;
  assign n12677 = n2022 & ~n12676 ;
  assign n12678 = n2026 & ~n12677 ;
  assign n12679 = n2030 & ~n12678 ;
  assign n12680 = n2034 & ~n12679 ;
  assign n12681 = n2038 & ~n12680 ;
  assign n12682 = n2042 & ~n12681 ;
  assign n12683 = n2046 & ~n12682 ;
  assign n12684 = n2050 & ~n12683 ;
  assign n12685 = n2054 & ~n12684 ;
  assign n12686 = n2058 & ~n12685 ;
  assign n12687 = n2062 & ~n12686 ;
  assign n12688 = n2066 & ~n12687 ;
  assign n12689 = n2070 & ~n12688 ;
  assign n12690 = n2074 & ~n12689 ;
  assign n12691 = n2078 & ~n12690 ;
  assign n12692 = n2082 & ~n12691 ;
  assign n12693 = n2086 & ~n12692 ;
  assign n12694 = n2090 & ~n12693 ;
  assign n12695 = n2094 & ~n12694 ;
  assign n12696 = n2098 & ~n12695 ;
  assign n12697 = n2102 & ~n12696 ;
  assign n12698 = n2106 & ~n12697 ;
  assign n12699 = ~x189 & ~n2108 ;
  assign n12700 = ~n12698 & n12699 ;
  assign n12703 = ~n12700 & ~x317 ;
  assign n12704 = ~n12702 & ~n12703 ;
  assign n12705 = ~n422 & n1780 ;
  assign n12706 = n1785 & ~n12705 ;
  assign n12707 = n1789 & ~n12706 ;
  assign n12708 = n1793 & ~n12707 ;
  assign n12709 = n1797 & ~n12708 ;
  assign n12710 = n1801 & ~n12709 ;
  assign n12711 = n1805 & ~n12710 ;
  assign n12712 = n1809 & ~n12711 ;
  assign n12713 = n1813 & ~n12712 ;
  assign n12714 = n1817 & ~n12713 ;
  assign n12715 = n1821 & ~n12714 ;
  assign n12716 = n1825 & ~n12715 ;
  assign n12717 = n1829 & ~n12716 ;
  assign n12718 = n1833 & ~n12717 ;
  assign n12719 = n1837 & ~n12718 ;
  assign n12720 = n1841 & ~n12719 ;
  assign n12721 = n1845 & ~n12720 ;
  assign n12722 = n1849 & ~n12721 ;
  assign n12723 = n1853 & ~n12722 ;
  assign n12724 = n1857 & ~n12723 ;
  assign n12725 = n1861 & ~n12724 ;
  assign n12726 = n1865 & ~n12725 ;
  assign n12727 = n1869 & ~n12726 ;
  assign n12728 = n1873 & ~n12727 ;
  assign n12729 = n1877 & ~n12728 ;
  assign n12730 = n1881 & ~n12729 ;
  assign n12731 = n1885 & ~n12730 ;
  assign n12732 = n1889 & ~n12731 ;
  assign n12733 = n1893 & ~n12732 ;
  assign n12734 = n1897 & ~n12733 ;
  assign n12735 = n1901 & ~n12734 ;
  assign n12736 = n1905 & ~n12735 ;
  assign n12737 = n1909 & ~n12736 ;
  assign n12738 = n1913 & ~n12737 ;
  assign n12739 = n1917 & ~n12738 ;
  assign n12740 = n1921 & ~n12739 ;
  assign n12741 = n1925 & ~n12740 ;
  assign n12742 = n1929 & ~n12741 ;
  assign n12743 = n1933 & ~n12742 ;
  assign n12744 = n1937 & ~n12743 ;
  assign n12745 = n1941 & ~n12744 ;
  assign n12746 = n1945 & ~n12745 ;
  assign n12747 = n1949 & ~n12746 ;
  assign n12748 = n1953 & ~n12747 ;
  assign n12749 = n2749 & ~n12748 ;
  assign n12750 = n263 & ~n12749 ;
  assign n12751 = n267 & ~n12750 ;
  assign n12752 = n271 & ~n12751 ;
  assign n12753 = n275 & ~n12752 ;
  assign n12754 = n279 & ~n12753 ;
  assign n12755 = n283 & ~n12754 ;
  assign n12756 = n287 & ~n12755 ;
  assign n12757 = n291 & ~n12756 ;
  assign n12758 = n295 & ~n12757 ;
  assign n12759 = n299 & ~n12758 ;
  assign n12760 = n303 & ~n12759 ;
  assign n12761 = n307 & ~n12760 ;
  assign n12762 = n311 & ~n12761 ;
  assign n12763 = n315 & ~n12762 ;
  assign n12764 = n319 & ~n12763 ;
  assign n12765 = n323 & ~n12764 ;
  assign n12766 = n327 & ~n12765 ;
  assign n12767 = n331 & ~n12766 ;
  assign n12768 = n335 & ~n12767 ;
  assign n12769 = n339 & ~n12768 ;
  assign n12770 = n343 & ~n12769 ;
  assign n12771 = n347 & ~n12770 ;
  assign n12772 = n351 & ~n12771 ;
  assign n12773 = n355 & ~n12772 ;
  assign n12774 = n359 & ~n12773 ;
  assign n12775 = n363 & ~n12774 ;
  assign n12776 = n367 & ~n12775 ;
  assign n12777 = n371 & ~n12776 ;
  assign n12778 = n375 & ~n12777 ;
  assign n12779 = n379 & ~n12778 ;
  assign n12780 = n383 & ~n12779 ;
  assign n12781 = n387 & ~n12780 ;
  assign n12782 = n391 & ~n12781 ;
  assign n12783 = n395 & ~n12782 ;
  assign n12784 = n399 & ~n12783 ;
  assign n12785 = n403 & ~n12784 ;
  assign n12786 = n407 & ~n12785 ;
  assign n12787 = n411 & ~n12786 ;
  assign n12788 = n415 & ~n12787 ;
  assign n12789 = x190 & ~n417 ;
  assign n12790 = ~n12788 & n12789 ;
  assign n12878 = n12790 & x318 ;
  assign n12791 = ~n761 & n2117 ;
  assign n12792 = n2122 & ~n12791 ;
  assign n12793 = n2126 & ~n12792 ;
  assign n12794 = n2130 & ~n12793 ;
  assign n12795 = n2134 & ~n12794 ;
  assign n12796 = n2138 & ~n12795 ;
  assign n12797 = n2142 & ~n12796 ;
  assign n12798 = n2146 & ~n12797 ;
  assign n12799 = n2150 & ~n12798 ;
  assign n12800 = n2154 & ~n12799 ;
  assign n12801 = n2158 & ~n12800 ;
  assign n12802 = n2162 & ~n12801 ;
  assign n12803 = n2166 & ~n12802 ;
  assign n12804 = n2170 & ~n12803 ;
  assign n12805 = n2174 & ~n12804 ;
  assign n12806 = n2178 & ~n12805 ;
  assign n12807 = n2182 & ~n12806 ;
  assign n12808 = n2186 & ~n12807 ;
  assign n12809 = n2190 & ~n12808 ;
  assign n12810 = n2194 & ~n12809 ;
  assign n12811 = n2198 & ~n12810 ;
  assign n12812 = n2202 & ~n12811 ;
  assign n12813 = n2206 & ~n12812 ;
  assign n12814 = n2210 & ~n12813 ;
  assign n12815 = n2214 & ~n12814 ;
  assign n12816 = n2218 & ~n12815 ;
  assign n12817 = n2222 & ~n12816 ;
  assign n12818 = n2226 & ~n12817 ;
  assign n12819 = n2230 & ~n12818 ;
  assign n12820 = n2234 & ~n12819 ;
  assign n12821 = n2238 & ~n12820 ;
  assign n12822 = n2242 & ~n12821 ;
  assign n12823 = n2246 & ~n12822 ;
  assign n12824 = n2250 & ~n12823 ;
  assign n12825 = n2254 & ~n12824 ;
  assign n12826 = n2258 & ~n12825 ;
  assign n12827 = n2262 & ~n12826 ;
  assign n12828 = n2266 & ~n12827 ;
  assign n12829 = n2270 & ~n12828 ;
  assign n12830 = n2274 & ~n12829 ;
  assign n12831 = n2278 & ~n12830 ;
  assign n12832 = n2282 & ~n12831 ;
  assign n12833 = n2286 & ~n12832 ;
  assign n12834 = n2290 & ~n12833 ;
  assign n12835 = n2836 & ~n12834 ;
  assign n12836 = n602 & ~n12835 ;
  assign n12837 = n606 & ~n12836 ;
  assign n12838 = n610 & ~n12837 ;
  assign n12839 = n614 & ~n12838 ;
  assign n12840 = n618 & ~n12839 ;
  assign n12841 = n622 & ~n12840 ;
  assign n12842 = n626 & ~n12841 ;
  assign n12843 = n630 & ~n12842 ;
  assign n12844 = n634 & ~n12843 ;
  assign n12845 = n638 & ~n12844 ;
  assign n12846 = n642 & ~n12845 ;
  assign n12847 = n646 & ~n12846 ;
  assign n12848 = n650 & ~n12847 ;
  assign n12849 = n654 & ~n12848 ;
  assign n12850 = n658 & ~n12849 ;
  assign n12851 = n662 & ~n12850 ;
  assign n12852 = n666 & ~n12851 ;
  assign n12853 = n670 & ~n12852 ;
  assign n12854 = n674 & ~n12853 ;
  assign n12855 = n678 & ~n12854 ;
  assign n12856 = n682 & ~n12855 ;
  assign n12857 = n686 & ~n12856 ;
  assign n12858 = n690 & ~n12857 ;
  assign n12859 = n694 & ~n12858 ;
  assign n12860 = n698 & ~n12859 ;
  assign n12861 = n702 & ~n12860 ;
  assign n12862 = n706 & ~n12861 ;
  assign n12863 = n710 & ~n12862 ;
  assign n12864 = n714 & ~n12863 ;
  assign n12865 = n718 & ~n12864 ;
  assign n12866 = n722 & ~n12865 ;
  assign n12867 = n726 & ~n12866 ;
  assign n12868 = n730 & ~n12867 ;
  assign n12869 = n734 & ~n12868 ;
  assign n12870 = n738 & ~n12869 ;
  assign n12871 = n742 & ~n12870 ;
  assign n12872 = n746 & ~n12871 ;
  assign n12873 = n750 & ~n12872 ;
  assign n12874 = n754 & ~n12873 ;
  assign n12875 = ~x190 & ~n756 ;
  assign n12876 = ~n12874 & n12875 ;
  assign n12879 = ~n12876 & ~x318 ;
  assign n12880 = ~n12878 & ~n12879 ;
  assign n12881 = n426 & ~n1104 ;
  assign n12882 = n431 & ~n12881 ;
  assign n12883 = n435 & ~n12882 ;
  assign n12884 = n439 & ~n12883 ;
  assign n12885 = n443 & ~n12884 ;
  assign n12886 = n447 & ~n12885 ;
  assign n12887 = n451 & ~n12886 ;
  assign n12888 = n455 & ~n12887 ;
  assign n12889 = n459 & ~n12888 ;
  assign n12890 = n463 & ~n12889 ;
  assign n12891 = n467 & ~n12890 ;
  assign n12892 = n471 & ~n12891 ;
  assign n12893 = n475 & ~n12892 ;
  assign n12894 = n479 & ~n12893 ;
  assign n12895 = n483 & ~n12894 ;
  assign n12896 = n487 & ~n12895 ;
  assign n12897 = n491 & ~n12896 ;
  assign n12898 = n495 & ~n12897 ;
  assign n12899 = n499 & ~n12898 ;
  assign n12900 = n503 & ~n12899 ;
  assign n12901 = n507 & ~n12900 ;
  assign n12902 = n511 & ~n12901 ;
  assign n12903 = n515 & ~n12902 ;
  assign n12904 = n519 & ~n12903 ;
  assign n12905 = n523 & ~n12904 ;
  assign n12906 = n527 & ~n12905 ;
  assign n12907 = n531 & ~n12906 ;
  assign n12908 = n535 & ~n12907 ;
  assign n12909 = n539 & ~n12908 ;
  assign n12910 = n543 & ~n12909 ;
  assign n12911 = n547 & ~n12910 ;
  assign n12912 = n551 & ~n12911 ;
  assign n12913 = n555 & ~n12912 ;
  assign n12914 = n559 & ~n12913 ;
  assign n12915 = n563 & ~n12914 ;
  assign n12916 = n567 & ~n12915 ;
  assign n12917 = n571 & ~n12916 ;
  assign n12918 = n575 & ~n12917 ;
  assign n12919 = n579 & ~n12918 ;
  assign n12920 = n583 & ~n12919 ;
  assign n12921 = n587 & ~n12920 ;
  assign n12922 = n591 & ~n12921 ;
  assign n12923 = n2382 & ~n12922 ;
  assign n12924 = n2384 & ~n12923 ;
  assign n12925 = n2927 & ~n12924 ;
  assign n12926 = n945 & ~n12925 ;
  assign n12927 = n949 & ~n12926 ;
  assign n12928 = n953 & ~n12927 ;
  assign n12929 = n957 & ~n12928 ;
  assign n12930 = n961 & ~n12929 ;
  assign n12931 = n965 & ~n12930 ;
  assign n12932 = n969 & ~n12931 ;
  assign n12933 = n973 & ~n12932 ;
  assign n12934 = n977 & ~n12933 ;
  assign n12935 = n981 & ~n12934 ;
  assign n12936 = n985 & ~n12935 ;
  assign n12937 = n989 & ~n12936 ;
  assign n12938 = n993 & ~n12937 ;
  assign n12939 = n997 & ~n12938 ;
  assign n12940 = n1001 & ~n12939 ;
  assign n12941 = n1005 & ~n12940 ;
  assign n12942 = n1009 & ~n12941 ;
  assign n12943 = n1013 & ~n12942 ;
  assign n12944 = n1017 & ~n12943 ;
  assign n12945 = n1021 & ~n12944 ;
  assign n12946 = n1025 & ~n12945 ;
  assign n12947 = n1029 & ~n12946 ;
  assign n12948 = n1033 & ~n12947 ;
  assign n12949 = n1037 & ~n12948 ;
  assign n12950 = n1041 & ~n12949 ;
  assign n12951 = n1045 & ~n12950 ;
  assign n12952 = n1049 & ~n12951 ;
  assign n12953 = n1053 & ~n12952 ;
  assign n12954 = n1057 & ~n12953 ;
  assign n12955 = n1061 & ~n12954 ;
  assign n12956 = n1065 & ~n12955 ;
  assign n12957 = n1069 & ~n12956 ;
  assign n12958 = n1073 & ~n12957 ;
  assign n12959 = n1077 & ~n12958 ;
  assign n12960 = n1081 & ~n12959 ;
  assign n12961 = n1085 & ~n12960 ;
  assign n12962 = n1089 & ~n12961 ;
  assign n12963 = n1093 & ~n12962 ;
  assign n12964 = n1097 & ~n12963 ;
  assign n12965 = x191 & ~n1099 ;
  assign n12966 = ~n12964 & n12965 ;
  assign n13054 = n12966 & x319 ;
  assign n12967 = n765 & ~n1443 ;
  assign n12968 = n770 & ~n12967 ;
  assign n12969 = n774 & ~n12968 ;
  assign n12970 = n778 & ~n12969 ;
  assign n12971 = n782 & ~n12970 ;
  assign n12972 = n786 & ~n12971 ;
  assign n12973 = n790 & ~n12972 ;
  assign n12974 = n794 & ~n12973 ;
  assign n12975 = n798 & ~n12974 ;
  assign n12976 = n802 & ~n12975 ;
  assign n12977 = n806 & ~n12976 ;
  assign n12978 = n810 & ~n12977 ;
  assign n12979 = n814 & ~n12978 ;
  assign n12980 = n818 & ~n12979 ;
  assign n12981 = n822 & ~n12980 ;
  assign n12982 = n826 & ~n12981 ;
  assign n12983 = n830 & ~n12982 ;
  assign n12984 = n834 & ~n12983 ;
  assign n12985 = n838 & ~n12984 ;
  assign n12986 = n842 & ~n12985 ;
  assign n12987 = n846 & ~n12986 ;
  assign n12988 = n850 & ~n12987 ;
  assign n12989 = n854 & ~n12988 ;
  assign n12990 = n858 & ~n12989 ;
  assign n12991 = n862 & ~n12990 ;
  assign n12992 = n866 & ~n12991 ;
  assign n12993 = n870 & ~n12992 ;
  assign n12994 = n874 & ~n12993 ;
  assign n12995 = n878 & ~n12994 ;
  assign n12996 = n882 & ~n12995 ;
  assign n12997 = n886 & ~n12996 ;
  assign n12998 = n890 & ~n12997 ;
  assign n12999 = n894 & ~n12998 ;
  assign n13000 = n898 & ~n12999 ;
  assign n13001 = n902 & ~n13000 ;
  assign n13002 = n906 & ~n13001 ;
  assign n13003 = n910 & ~n13002 ;
  assign n13004 = n914 & ~n13003 ;
  assign n13005 = n918 & ~n13004 ;
  assign n13006 = n922 & ~n13005 ;
  assign n13007 = n926 & ~n13006 ;
  assign n13008 = n930 & ~n13007 ;
  assign n13009 = n2472 & ~n13008 ;
  assign n13010 = n2474 & ~n13009 ;
  assign n13011 = n3014 & ~n13010 ;
  assign n13012 = n1284 & ~n13011 ;
  assign n13013 = n1288 & ~n13012 ;
  assign n13014 = n1292 & ~n13013 ;
  assign n13015 = n1296 & ~n13014 ;
  assign n13016 = n1300 & ~n13015 ;
  assign n13017 = n1304 & ~n13016 ;
  assign n13018 = n1308 & ~n13017 ;
  assign n13019 = n1312 & ~n13018 ;
  assign n13020 = n1316 & ~n13019 ;
  assign n13021 = n1320 & ~n13020 ;
  assign n13022 = n1324 & ~n13021 ;
  assign n13023 = n1328 & ~n13022 ;
  assign n13024 = n1332 & ~n13023 ;
  assign n13025 = n1336 & ~n13024 ;
  assign n13026 = n1340 & ~n13025 ;
  assign n13027 = n1344 & ~n13026 ;
  assign n13028 = n1348 & ~n13027 ;
  assign n13029 = n1352 & ~n13028 ;
  assign n13030 = n1356 & ~n13029 ;
  assign n13031 = n1360 & ~n13030 ;
  assign n13032 = n1364 & ~n13031 ;
  assign n13033 = n1368 & ~n13032 ;
  assign n13034 = n1372 & ~n13033 ;
  assign n13035 = n1376 & ~n13034 ;
  assign n13036 = n1380 & ~n13035 ;
  assign n13037 = n1384 & ~n13036 ;
  assign n13038 = n1388 & ~n13037 ;
  assign n13039 = n1392 & ~n13038 ;
  assign n13040 = n1396 & ~n13039 ;
  assign n13041 = n1400 & ~n13040 ;
  assign n13042 = n1404 & ~n13041 ;
  assign n13043 = n1408 & ~n13042 ;
  assign n13044 = n1412 & ~n13043 ;
  assign n13045 = n1416 & ~n13044 ;
  assign n13046 = n1420 & ~n13045 ;
  assign n13047 = n1424 & ~n13046 ;
  assign n13048 = n1428 & ~n13047 ;
  assign n13049 = n1432 & ~n13048 ;
  assign n13050 = n1436 & ~n13049 ;
  assign n13051 = ~x191 & ~n1438 ;
  assign n13052 = ~n13050 & n13051 ;
  assign n13055 = ~n13052 & ~x319 ;
  assign n13056 = ~n13054 & ~n13055 ;
  assign n13057 = n1108 & ~n1784 ;
  assign n13058 = n1113 & ~n13057 ;
  assign n13059 = n1117 & ~n13058 ;
  assign n13060 = n1121 & ~n13059 ;
  assign n13061 = n1125 & ~n13060 ;
  assign n13062 = n1129 & ~n13061 ;
  assign n13063 = n1133 & ~n13062 ;
  assign n13064 = n1137 & ~n13063 ;
  assign n13065 = n1141 & ~n13064 ;
  assign n13066 = n1145 & ~n13065 ;
  assign n13067 = n1149 & ~n13066 ;
  assign n13068 = n1153 & ~n13067 ;
  assign n13069 = n1157 & ~n13068 ;
  assign n13070 = n1161 & ~n13069 ;
  assign n13071 = n1165 & ~n13070 ;
  assign n13072 = n1169 & ~n13071 ;
  assign n13073 = n1173 & ~n13072 ;
  assign n13074 = n1177 & ~n13073 ;
  assign n13075 = n1181 & ~n13074 ;
  assign n13076 = n1185 & ~n13075 ;
  assign n13077 = n1189 & ~n13076 ;
  assign n13078 = n1193 & ~n13077 ;
  assign n13079 = n1197 & ~n13078 ;
  assign n13080 = n1201 & ~n13079 ;
  assign n13081 = n1205 & ~n13080 ;
  assign n13082 = n1209 & ~n13081 ;
  assign n13083 = n1213 & ~n13082 ;
  assign n13084 = n1217 & ~n13083 ;
  assign n13085 = n1221 & ~n13084 ;
  assign n13086 = n1225 & ~n13085 ;
  assign n13087 = n1229 & ~n13086 ;
  assign n13088 = n1233 & ~n13087 ;
  assign n13089 = n1237 & ~n13088 ;
  assign n13090 = n1241 & ~n13089 ;
  assign n13091 = n1245 & ~n13090 ;
  assign n13092 = n1249 & ~n13091 ;
  assign n13093 = n1253 & ~n13092 ;
  assign n13094 = n1257 & ~n13093 ;
  assign n13095 = n1261 & ~n13094 ;
  assign n13096 = n1265 & ~n13095 ;
  assign n13097 = n1269 & ~n13096 ;
  assign n13098 = n1273 & ~n13097 ;
  assign n13099 = n2566 & ~n13098 ;
  assign n13100 = n2568 & ~n13099 ;
  assign n13101 = n3105 & ~n13100 ;
  assign n13102 = n1625 & ~n13101 ;
  assign n13103 = n1629 & ~n13102 ;
  assign n13104 = n1633 & ~n13103 ;
  assign n13105 = n1637 & ~n13104 ;
  assign n13106 = n1641 & ~n13105 ;
  assign n13107 = n1645 & ~n13106 ;
  assign n13108 = n1649 & ~n13107 ;
  assign n13109 = n1653 & ~n13108 ;
  assign n13110 = n1657 & ~n13109 ;
  assign n13111 = n1661 & ~n13110 ;
  assign n13112 = n1665 & ~n13111 ;
  assign n13113 = n1669 & ~n13112 ;
  assign n13114 = n1673 & ~n13113 ;
  assign n13115 = n1677 & ~n13114 ;
  assign n13116 = n1681 & ~n13115 ;
  assign n13117 = n1685 & ~n13116 ;
  assign n13118 = n1689 & ~n13117 ;
  assign n13119 = n1693 & ~n13118 ;
  assign n13120 = n1697 & ~n13119 ;
  assign n13121 = n1701 & ~n13120 ;
  assign n13122 = n1705 & ~n13121 ;
  assign n13123 = n1709 & ~n13122 ;
  assign n13124 = n1713 & ~n13123 ;
  assign n13125 = n1717 & ~n13124 ;
  assign n13126 = n1721 & ~n13125 ;
  assign n13127 = n1725 & ~n13126 ;
  assign n13128 = n1729 & ~n13127 ;
  assign n13129 = n1733 & ~n13128 ;
  assign n13130 = n1737 & ~n13129 ;
  assign n13131 = n1741 & ~n13130 ;
  assign n13132 = n1745 & ~n13131 ;
  assign n13133 = n1749 & ~n13132 ;
  assign n13134 = n1753 & ~n13133 ;
  assign n13135 = n1757 & ~n13134 ;
  assign n13136 = n1761 & ~n13135 ;
  assign n13137 = n1765 & ~n13136 ;
  assign n13138 = n1769 & ~n13137 ;
  assign n13139 = n1773 & ~n13138 ;
  assign n13140 = n1777 & ~n13139 ;
  assign n13141 = x192 & ~n1779 ;
  assign n13142 = ~n13140 & n13141 ;
  assign n13230 = n13142 & x320 ;
  assign n13143 = n1447 & ~n2121 ;
  assign n13144 = n1452 & ~n13143 ;
  assign n13145 = n1456 & ~n13144 ;
  assign n13146 = n1460 & ~n13145 ;
  assign n13147 = n1464 & ~n13146 ;
  assign n13148 = n1468 & ~n13147 ;
  assign n13149 = n1472 & ~n13148 ;
  assign n13150 = n1476 & ~n13149 ;
  assign n13151 = n1480 & ~n13150 ;
  assign n13152 = n1484 & ~n13151 ;
  assign n13153 = n1488 & ~n13152 ;
  assign n13154 = n1492 & ~n13153 ;
  assign n13155 = n1496 & ~n13154 ;
  assign n13156 = n1500 & ~n13155 ;
  assign n13157 = n1504 & ~n13156 ;
  assign n13158 = n1508 & ~n13157 ;
  assign n13159 = n1512 & ~n13158 ;
  assign n13160 = n1516 & ~n13159 ;
  assign n13161 = n1520 & ~n13160 ;
  assign n13162 = n1524 & ~n13161 ;
  assign n13163 = n1528 & ~n13162 ;
  assign n13164 = n1532 & ~n13163 ;
  assign n13165 = n1536 & ~n13164 ;
  assign n13166 = n1540 & ~n13165 ;
  assign n13167 = n1544 & ~n13166 ;
  assign n13168 = n1548 & ~n13167 ;
  assign n13169 = n1552 & ~n13168 ;
  assign n13170 = n1556 & ~n13169 ;
  assign n13171 = n1560 & ~n13170 ;
  assign n13172 = n1564 & ~n13171 ;
  assign n13173 = n1568 & ~n13172 ;
  assign n13174 = n1572 & ~n13173 ;
  assign n13175 = n1576 & ~n13174 ;
  assign n13176 = n1580 & ~n13175 ;
  assign n13177 = n1584 & ~n13176 ;
  assign n13178 = n1588 & ~n13177 ;
  assign n13179 = n1592 & ~n13178 ;
  assign n13180 = n1596 & ~n13179 ;
  assign n13181 = n1600 & ~n13180 ;
  assign n13182 = n1604 & ~n13181 ;
  assign n13183 = n1608 & ~n13182 ;
  assign n13184 = n1612 & ~n13183 ;
  assign n13185 = n2656 & ~n13184 ;
  assign n13186 = n2658 & ~n13185 ;
  assign n13187 = n3192 & ~n13186 ;
  assign n13188 = n1962 & ~n13187 ;
  assign n13189 = n1966 & ~n13188 ;
  assign n13190 = n1970 & ~n13189 ;
  assign n13191 = n1974 & ~n13190 ;
  assign n13192 = n1978 & ~n13191 ;
  assign n13193 = n1982 & ~n13192 ;
  assign n13194 = n1986 & ~n13193 ;
  assign n13195 = n1990 & ~n13194 ;
  assign n13196 = n1994 & ~n13195 ;
  assign n13197 = n1998 & ~n13196 ;
  assign n13198 = n2002 & ~n13197 ;
  assign n13199 = n2006 & ~n13198 ;
  assign n13200 = n2010 & ~n13199 ;
  assign n13201 = n2014 & ~n13200 ;
  assign n13202 = n2018 & ~n13201 ;
  assign n13203 = n2022 & ~n13202 ;
  assign n13204 = n2026 & ~n13203 ;
  assign n13205 = n2030 & ~n13204 ;
  assign n13206 = n2034 & ~n13205 ;
  assign n13207 = n2038 & ~n13206 ;
  assign n13208 = n2042 & ~n13207 ;
  assign n13209 = n2046 & ~n13208 ;
  assign n13210 = n2050 & ~n13209 ;
  assign n13211 = n2054 & ~n13210 ;
  assign n13212 = n2058 & ~n13211 ;
  assign n13213 = n2062 & ~n13212 ;
  assign n13214 = n2066 & ~n13213 ;
  assign n13215 = n2070 & ~n13214 ;
  assign n13216 = n2074 & ~n13215 ;
  assign n13217 = n2078 & ~n13216 ;
  assign n13218 = n2082 & ~n13217 ;
  assign n13219 = n2086 & ~n13218 ;
  assign n13220 = n2090 & ~n13219 ;
  assign n13221 = n2094 & ~n13220 ;
  assign n13222 = n2098 & ~n13221 ;
  assign n13223 = n2102 & ~n13222 ;
  assign n13224 = n2106 & ~n13223 ;
  assign n13225 = n2110 & ~n13224 ;
  assign n13226 = n2114 & ~n13225 ;
  assign n13227 = ~x192 & ~n2116 ;
  assign n13228 = ~n13226 & n13227 ;
  assign n13231 = ~n13228 & ~x320 ;
  assign n13232 = ~n13230 & ~n13231 ;
  assign n13233 = ~n430 & n1788 ;
  assign n13234 = n1793 & ~n13233 ;
  assign n13235 = n1797 & ~n13234 ;
  assign n13236 = n1801 & ~n13235 ;
  assign n13237 = n1805 & ~n13236 ;
  assign n13238 = n1809 & ~n13237 ;
  assign n13239 = n1813 & ~n13238 ;
  assign n13240 = n1817 & ~n13239 ;
  assign n13241 = n1821 & ~n13240 ;
  assign n13242 = n1825 & ~n13241 ;
  assign n13243 = n1829 & ~n13242 ;
  assign n13244 = n1833 & ~n13243 ;
  assign n13245 = n1837 & ~n13244 ;
  assign n13246 = n1841 & ~n13245 ;
  assign n13247 = n1845 & ~n13246 ;
  assign n13248 = n1849 & ~n13247 ;
  assign n13249 = n1853 & ~n13248 ;
  assign n13250 = n1857 & ~n13249 ;
  assign n13251 = n1861 & ~n13250 ;
  assign n13252 = n1865 & ~n13251 ;
  assign n13253 = n1869 & ~n13252 ;
  assign n13254 = n1873 & ~n13253 ;
  assign n13255 = n1877 & ~n13254 ;
  assign n13256 = n1881 & ~n13255 ;
  assign n13257 = n1885 & ~n13256 ;
  assign n13258 = n1889 & ~n13257 ;
  assign n13259 = n1893 & ~n13258 ;
  assign n13260 = n1897 & ~n13259 ;
  assign n13261 = n1901 & ~n13260 ;
  assign n13262 = n1905 & ~n13261 ;
  assign n13263 = n1909 & ~n13262 ;
  assign n13264 = n1913 & ~n13263 ;
  assign n13265 = n1917 & ~n13264 ;
  assign n13266 = n1921 & ~n13265 ;
  assign n13267 = n1925 & ~n13266 ;
  assign n13268 = n1929 & ~n13267 ;
  assign n13269 = n1933 & ~n13268 ;
  assign n13270 = n1937 & ~n13269 ;
  assign n13271 = n1941 & ~n13270 ;
  assign n13272 = n1945 & ~n13271 ;
  assign n13273 = n1949 & ~n13272 ;
  assign n13274 = n1953 & ~n13273 ;
  assign n13275 = n2749 & ~n13274 ;
  assign n13276 = n263 & ~n13275 ;
  assign n13277 = n267 & ~n13276 ;
  assign n13278 = n271 & ~n13277 ;
  assign n13279 = n275 & ~n13278 ;
  assign n13280 = n279 & ~n13279 ;
  assign n13281 = n283 & ~n13280 ;
  assign n13282 = n287 & ~n13281 ;
  assign n13283 = n291 & ~n13282 ;
  assign n13284 = n295 & ~n13283 ;
  assign n13285 = n299 & ~n13284 ;
  assign n13286 = n303 & ~n13285 ;
  assign n13287 = n307 & ~n13286 ;
  assign n13288 = n311 & ~n13287 ;
  assign n13289 = n315 & ~n13288 ;
  assign n13290 = n319 & ~n13289 ;
  assign n13291 = n323 & ~n13290 ;
  assign n13292 = n327 & ~n13291 ;
  assign n13293 = n331 & ~n13292 ;
  assign n13294 = n335 & ~n13293 ;
  assign n13295 = n339 & ~n13294 ;
  assign n13296 = n343 & ~n13295 ;
  assign n13297 = n347 & ~n13296 ;
  assign n13298 = n351 & ~n13297 ;
  assign n13299 = n355 & ~n13298 ;
  assign n13300 = n359 & ~n13299 ;
  assign n13301 = n363 & ~n13300 ;
  assign n13302 = n367 & ~n13301 ;
  assign n13303 = n371 & ~n13302 ;
  assign n13304 = n375 & ~n13303 ;
  assign n13305 = n379 & ~n13304 ;
  assign n13306 = n383 & ~n13305 ;
  assign n13307 = n387 & ~n13306 ;
  assign n13308 = n391 & ~n13307 ;
  assign n13309 = n395 & ~n13308 ;
  assign n13310 = n399 & ~n13309 ;
  assign n13311 = n403 & ~n13310 ;
  assign n13312 = n407 & ~n13311 ;
  assign n13313 = n411 & ~n13312 ;
  assign n13314 = n415 & ~n13313 ;
  assign n13315 = n419 & ~n13314 ;
  assign n13316 = n423 & ~n13315 ;
  assign n13317 = x193 & ~n425 ;
  assign n13318 = ~n13316 & n13317 ;
  assign n13406 = n13318 & x321 ;
  assign n13319 = ~n769 & n2125 ;
  assign n13320 = n2130 & ~n13319 ;
  assign n13321 = n2134 & ~n13320 ;
  assign n13322 = n2138 & ~n13321 ;
  assign n13323 = n2142 & ~n13322 ;
  assign n13324 = n2146 & ~n13323 ;
  assign n13325 = n2150 & ~n13324 ;
  assign n13326 = n2154 & ~n13325 ;
  assign n13327 = n2158 & ~n13326 ;
  assign n13328 = n2162 & ~n13327 ;
  assign n13329 = n2166 & ~n13328 ;
  assign n13330 = n2170 & ~n13329 ;
  assign n13331 = n2174 & ~n13330 ;
  assign n13332 = n2178 & ~n13331 ;
  assign n13333 = n2182 & ~n13332 ;
  assign n13334 = n2186 & ~n13333 ;
  assign n13335 = n2190 & ~n13334 ;
  assign n13336 = n2194 & ~n13335 ;
  assign n13337 = n2198 & ~n13336 ;
  assign n13338 = n2202 & ~n13337 ;
  assign n13339 = n2206 & ~n13338 ;
  assign n13340 = n2210 & ~n13339 ;
  assign n13341 = n2214 & ~n13340 ;
  assign n13342 = n2218 & ~n13341 ;
  assign n13343 = n2222 & ~n13342 ;
  assign n13344 = n2226 & ~n13343 ;
  assign n13345 = n2230 & ~n13344 ;
  assign n13346 = n2234 & ~n13345 ;
  assign n13347 = n2238 & ~n13346 ;
  assign n13348 = n2242 & ~n13347 ;
  assign n13349 = n2246 & ~n13348 ;
  assign n13350 = n2250 & ~n13349 ;
  assign n13351 = n2254 & ~n13350 ;
  assign n13352 = n2258 & ~n13351 ;
  assign n13353 = n2262 & ~n13352 ;
  assign n13354 = n2266 & ~n13353 ;
  assign n13355 = n2270 & ~n13354 ;
  assign n13356 = n2274 & ~n13355 ;
  assign n13357 = n2278 & ~n13356 ;
  assign n13358 = n2282 & ~n13357 ;
  assign n13359 = n2286 & ~n13358 ;
  assign n13360 = n2290 & ~n13359 ;
  assign n13361 = n2836 & ~n13360 ;
  assign n13362 = n602 & ~n13361 ;
  assign n13363 = n606 & ~n13362 ;
  assign n13364 = n610 & ~n13363 ;
  assign n13365 = n614 & ~n13364 ;
  assign n13366 = n618 & ~n13365 ;
  assign n13367 = n622 & ~n13366 ;
  assign n13368 = n626 & ~n13367 ;
  assign n13369 = n630 & ~n13368 ;
  assign n13370 = n634 & ~n13369 ;
  assign n13371 = n638 & ~n13370 ;
  assign n13372 = n642 & ~n13371 ;
  assign n13373 = n646 & ~n13372 ;
  assign n13374 = n650 & ~n13373 ;
  assign n13375 = n654 & ~n13374 ;
  assign n13376 = n658 & ~n13375 ;
  assign n13377 = n662 & ~n13376 ;
  assign n13378 = n666 & ~n13377 ;
  assign n13379 = n670 & ~n13378 ;
  assign n13380 = n674 & ~n13379 ;
  assign n13381 = n678 & ~n13380 ;
  assign n13382 = n682 & ~n13381 ;
  assign n13383 = n686 & ~n13382 ;
  assign n13384 = n690 & ~n13383 ;
  assign n13385 = n694 & ~n13384 ;
  assign n13386 = n698 & ~n13385 ;
  assign n13387 = n702 & ~n13386 ;
  assign n13388 = n706 & ~n13387 ;
  assign n13389 = n710 & ~n13388 ;
  assign n13390 = n714 & ~n13389 ;
  assign n13391 = n718 & ~n13390 ;
  assign n13392 = n722 & ~n13391 ;
  assign n13393 = n726 & ~n13392 ;
  assign n13394 = n730 & ~n13393 ;
  assign n13395 = n734 & ~n13394 ;
  assign n13396 = n738 & ~n13395 ;
  assign n13397 = n742 & ~n13396 ;
  assign n13398 = n746 & ~n13397 ;
  assign n13399 = n750 & ~n13398 ;
  assign n13400 = n754 & ~n13399 ;
  assign n13401 = n758 & ~n13400 ;
  assign n13402 = n762 & ~n13401 ;
  assign n13403 = ~x193 & ~n764 ;
  assign n13404 = ~n13402 & n13403 ;
  assign n13407 = ~n13404 & ~x321 ;
  assign n13408 = ~n13406 & ~n13407 ;
  assign n13409 = n434 & ~n1112 ;
  assign n13410 = n439 & ~n13409 ;
  assign n13411 = n443 & ~n13410 ;
  assign n13412 = n447 & ~n13411 ;
  assign n13413 = n451 & ~n13412 ;
  assign n13414 = n455 & ~n13413 ;
  assign n13415 = n459 & ~n13414 ;
  assign n13416 = n463 & ~n13415 ;
  assign n13417 = n467 & ~n13416 ;
  assign n13418 = n471 & ~n13417 ;
  assign n13419 = n475 & ~n13418 ;
  assign n13420 = n479 & ~n13419 ;
  assign n13421 = n483 & ~n13420 ;
  assign n13422 = n487 & ~n13421 ;
  assign n13423 = n491 & ~n13422 ;
  assign n13424 = n495 & ~n13423 ;
  assign n13425 = n499 & ~n13424 ;
  assign n13426 = n503 & ~n13425 ;
  assign n13427 = n507 & ~n13426 ;
  assign n13428 = n511 & ~n13427 ;
  assign n13429 = n515 & ~n13428 ;
  assign n13430 = n519 & ~n13429 ;
  assign n13431 = n523 & ~n13430 ;
  assign n13432 = n527 & ~n13431 ;
  assign n13433 = n531 & ~n13432 ;
  assign n13434 = n535 & ~n13433 ;
  assign n13435 = n539 & ~n13434 ;
  assign n13436 = n543 & ~n13435 ;
  assign n13437 = n547 & ~n13436 ;
  assign n13438 = n551 & ~n13437 ;
  assign n13439 = n555 & ~n13438 ;
  assign n13440 = n559 & ~n13439 ;
  assign n13441 = n563 & ~n13440 ;
  assign n13442 = n567 & ~n13441 ;
  assign n13443 = n571 & ~n13442 ;
  assign n13444 = n575 & ~n13443 ;
  assign n13445 = n579 & ~n13444 ;
  assign n13446 = n583 & ~n13445 ;
  assign n13447 = n587 & ~n13446 ;
  assign n13448 = n591 & ~n13447 ;
  assign n13449 = n2382 & ~n13448 ;
  assign n13450 = n2384 & ~n13449 ;
  assign n13451 = n2927 & ~n13450 ;
  assign n13452 = n945 & ~n13451 ;
  assign n13453 = n949 & ~n13452 ;
  assign n13454 = n953 & ~n13453 ;
  assign n13455 = n957 & ~n13454 ;
  assign n13456 = n961 & ~n13455 ;
  assign n13457 = n965 & ~n13456 ;
  assign n13458 = n969 & ~n13457 ;
  assign n13459 = n973 & ~n13458 ;
  assign n13460 = n977 & ~n13459 ;
  assign n13461 = n981 & ~n13460 ;
  assign n13462 = n985 & ~n13461 ;
  assign n13463 = n989 & ~n13462 ;
  assign n13464 = n993 & ~n13463 ;
  assign n13465 = n997 & ~n13464 ;
  assign n13466 = n1001 & ~n13465 ;
  assign n13467 = n1005 & ~n13466 ;
  assign n13468 = n1009 & ~n13467 ;
  assign n13469 = n1013 & ~n13468 ;
  assign n13470 = n1017 & ~n13469 ;
  assign n13471 = n1021 & ~n13470 ;
  assign n13472 = n1025 & ~n13471 ;
  assign n13473 = n1029 & ~n13472 ;
  assign n13474 = n1033 & ~n13473 ;
  assign n13475 = n1037 & ~n13474 ;
  assign n13476 = n1041 & ~n13475 ;
  assign n13477 = n1045 & ~n13476 ;
  assign n13478 = n1049 & ~n13477 ;
  assign n13479 = n1053 & ~n13478 ;
  assign n13480 = n1057 & ~n13479 ;
  assign n13481 = n1061 & ~n13480 ;
  assign n13482 = n1065 & ~n13481 ;
  assign n13483 = n1069 & ~n13482 ;
  assign n13484 = n1073 & ~n13483 ;
  assign n13485 = n1077 & ~n13484 ;
  assign n13486 = n1081 & ~n13485 ;
  assign n13487 = n1085 & ~n13486 ;
  assign n13488 = n1089 & ~n13487 ;
  assign n13489 = n1093 & ~n13488 ;
  assign n13490 = n1097 & ~n13489 ;
  assign n13491 = n1101 & ~n13490 ;
  assign n13492 = n1105 & ~n13491 ;
  assign n13493 = x194 & ~n1107 ;
  assign n13494 = ~n13492 & n13493 ;
  assign n13582 = n13494 & x322 ;
  assign n13495 = n773 & ~n1451 ;
  assign n13496 = n778 & ~n13495 ;
  assign n13497 = n782 & ~n13496 ;
  assign n13498 = n786 & ~n13497 ;
  assign n13499 = n790 & ~n13498 ;
  assign n13500 = n794 & ~n13499 ;
  assign n13501 = n798 & ~n13500 ;
  assign n13502 = n802 & ~n13501 ;
  assign n13503 = n806 & ~n13502 ;
  assign n13504 = n810 & ~n13503 ;
  assign n13505 = n814 & ~n13504 ;
  assign n13506 = n818 & ~n13505 ;
  assign n13507 = n822 & ~n13506 ;
  assign n13508 = n826 & ~n13507 ;
  assign n13509 = n830 & ~n13508 ;
  assign n13510 = n834 & ~n13509 ;
  assign n13511 = n838 & ~n13510 ;
  assign n13512 = n842 & ~n13511 ;
  assign n13513 = n846 & ~n13512 ;
  assign n13514 = n850 & ~n13513 ;
  assign n13515 = n854 & ~n13514 ;
  assign n13516 = n858 & ~n13515 ;
  assign n13517 = n862 & ~n13516 ;
  assign n13518 = n866 & ~n13517 ;
  assign n13519 = n870 & ~n13518 ;
  assign n13520 = n874 & ~n13519 ;
  assign n13521 = n878 & ~n13520 ;
  assign n13522 = n882 & ~n13521 ;
  assign n13523 = n886 & ~n13522 ;
  assign n13524 = n890 & ~n13523 ;
  assign n13525 = n894 & ~n13524 ;
  assign n13526 = n898 & ~n13525 ;
  assign n13527 = n902 & ~n13526 ;
  assign n13528 = n906 & ~n13527 ;
  assign n13529 = n910 & ~n13528 ;
  assign n13530 = n914 & ~n13529 ;
  assign n13531 = n918 & ~n13530 ;
  assign n13532 = n922 & ~n13531 ;
  assign n13533 = n926 & ~n13532 ;
  assign n13534 = n930 & ~n13533 ;
  assign n13535 = n2472 & ~n13534 ;
  assign n13536 = n2474 & ~n13535 ;
  assign n13537 = n3014 & ~n13536 ;
  assign n13538 = n1284 & ~n13537 ;
  assign n13539 = n1288 & ~n13538 ;
  assign n13540 = n1292 & ~n13539 ;
  assign n13541 = n1296 & ~n13540 ;
  assign n13542 = n1300 & ~n13541 ;
  assign n13543 = n1304 & ~n13542 ;
  assign n13544 = n1308 & ~n13543 ;
  assign n13545 = n1312 & ~n13544 ;
  assign n13546 = n1316 & ~n13545 ;
  assign n13547 = n1320 & ~n13546 ;
  assign n13548 = n1324 & ~n13547 ;
  assign n13549 = n1328 & ~n13548 ;
  assign n13550 = n1332 & ~n13549 ;
  assign n13551 = n1336 & ~n13550 ;
  assign n13552 = n1340 & ~n13551 ;
  assign n13553 = n1344 & ~n13552 ;
  assign n13554 = n1348 & ~n13553 ;
  assign n13555 = n1352 & ~n13554 ;
  assign n13556 = n1356 & ~n13555 ;
  assign n13557 = n1360 & ~n13556 ;
  assign n13558 = n1364 & ~n13557 ;
  assign n13559 = n1368 & ~n13558 ;
  assign n13560 = n1372 & ~n13559 ;
  assign n13561 = n1376 & ~n13560 ;
  assign n13562 = n1380 & ~n13561 ;
  assign n13563 = n1384 & ~n13562 ;
  assign n13564 = n1388 & ~n13563 ;
  assign n13565 = n1392 & ~n13564 ;
  assign n13566 = n1396 & ~n13565 ;
  assign n13567 = n1400 & ~n13566 ;
  assign n13568 = n1404 & ~n13567 ;
  assign n13569 = n1408 & ~n13568 ;
  assign n13570 = n1412 & ~n13569 ;
  assign n13571 = n1416 & ~n13570 ;
  assign n13572 = n1420 & ~n13571 ;
  assign n13573 = n1424 & ~n13572 ;
  assign n13574 = n1428 & ~n13573 ;
  assign n13575 = n1432 & ~n13574 ;
  assign n13576 = n1436 & ~n13575 ;
  assign n13577 = n1440 & ~n13576 ;
  assign n13578 = n1444 & ~n13577 ;
  assign n13579 = ~x194 & ~n1446 ;
  assign n13580 = ~n13578 & n13579 ;
  assign n13583 = ~n13580 & ~x322 ;
  assign n13584 = ~n13582 & ~n13583 ;
  assign n13585 = n1116 & ~n1792 ;
  assign n13586 = n1121 & ~n13585 ;
  assign n13587 = n1125 & ~n13586 ;
  assign n13588 = n1129 & ~n13587 ;
  assign n13589 = n1133 & ~n13588 ;
  assign n13590 = n1137 & ~n13589 ;
  assign n13591 = n1141 & ~n13590 ;
  assign n13592 = n1145 & ~n13591 ;
  assign n13593 = n1149 & ~n13592 ;
  assign n13594 = n1153 & ~n13593 ;
  assign n13595 = n1157 & ~n13594 ;
  assign n13596 = n1161 & ~n13595 ;
  assign n13597 = n1165 & ~n13596 ;
  assign n13598 = n1169 & ~n13597 ;
  assign n13599 = n1173 & ~n13598 ;
  assign n13600 = n1177 & ~n13599 ;
  assign n13601 = n1181 & ~n13600 ;
  assign n13602 = n1185 & ~n13601 ;
  assign n13603 = n1189 & ~n13602 ;
  assign n13604 = n1193 & ~n13603 ;
  assign n13605 = n1197 & ~n13604 ;
  assign n13606 = n1201 & ~n13605 ;
  assign n13607 = n1205 & ~n13606 ;
  assign n13608 = n1209 & ~n13607 ;
  assign n13609 = n1213 & ~n13608 ;
  assign n13610 = n1217 & ~n13609 ;
  assign n13611 = n1221 & ~n13610 ;
  assign n13612 = n1225 & ~n13611 ;
  assign n13613 = n1229 & ~n13612 ;
  assign n13614 = n1233 & ~n13613 ;
  assign n13615 = n1237 & ~n13614 ;
  assign n13616 = n1241 & ~n13615 ;
  assign n13617 = n1245 & ~n13616 ;
  assign n13618 = n1249 & ~n13617 ;
  assign n13619 = n1253 & ~n13618 ;
  assign n13620 = n1257 & ~n13619 ;
  assign n13621 = n1261 & ~n13620 ;
  assign n13622 = n1265 & ~n13621 ;
  assign n13623 = n1269 & ~n13622 ;
  assign n13624 = n1273 & ~n13623 ;
  assign n13625 = n2566 & ~n13624 ;
  assign n13626 = n2568 & ~n13625 ;
  assign n13627 = n3105 & ~n13626 ;
  assign n13628 = n1625 & ~n13627 ;
  assign n13629 = n1629 & ~n13628 ;
  assign n13630 = n1633 & ~n13629 ;
  assign n13631 = n1637 & ~n13630 ;
  assign n13632 = n1641 & ~n13631 ;
  assign n13633 = n1645 & ~n13632 ;
  assign n13634 = n1649 & ~n13633 ;
  assign n13635 = n1653 & ~n13634 ;
  assign n13636 = n1657 & ~n13635 ;
  assign n13637 = n1661 & ~n13636 ;
  assign n13638 = n1665 & ~n13637 ;
  assign n13639 = n1669 & ~n13638 ;
  assign n13640 = n1673 & ~n13639 ;
  assign n13641 = n1677 & ~n13640 ;
  assign n13642 = n1681 & ~n13641 ;
  assign n13643 = n1685 & ~n13642 ;
  assign n13644 = n1689 & ~n13643 ;
  assign n13645 = n1693 & ~n13644 ;
  assign n13646 = n1697 & ~n13645 ;
  assign n13647 = n1701 & ~n13646 ;
  assign n13648 = n1705 & ~n13647 ;
  assign n13649 = n1709 & ~n13648 ;
  assign n13650 = n1713 & ~n13649 ;
  assign n13651 = n1717 & ~n13650 ;
  assign n13652 = n1721 & ~n13651 ;
  assign n13653 = n1725 & ~n13652 ;
  assign n13654 = n1729 & ~n13653 ;
  assign n13655 = n1733 & ~n13654 ;
  assign n13656 = n1737 & ~n13655 ;
  assign n13657 = n1741 & ~n13656 ;
  assign n13658 = n1745 & ~n13657 ;
  assign n13659 = n1749 & ~n13658 ;
  assign n13660 = n1753 & ~n13659 ;
  assign n13661 = n1757 & ~n13660 ;
  assign n13662 = n1761 & ~n13661 ;
  assign n13663 = n1765 & ~n13662 ;
  assign n13664 = n1769 & ~n13663 ;
  assign n13665 = n1773 & ~n13664 ;
  assign n13666 = n1777 & ~n13665 ;
  assign n13667 = n1781 & ~n13666 ;
  assign n13668 = n1785 & ~n13667 ;
  assign n13669 = x195 & ~n1787 ;
  assign n13670 = ~n13668 & n13669 ;
  assign n13758 = n13670 & x323 ;
  assign n13671 = n1455 & ~n2129 ;
  assign n13672 = n1460 & ~n13671 ;
  assign n13673 = n1464 & ~n13672 ;
  assign n13674 = n1468 & ~n13673 ;
  assign n13675 = n1472 & ~n13674 ;
  assign n13676 = n1476 & ~n13675 ;
  assign n13677 = n1480 & ~n13676 ;
  assign n13678 = n1484 & ~n13677 ;
  assign n13679 = n1488 & ~n13678 ;
  assign n13680 = n1492 & ~n13679 ;
  assign n13681 = n1496 & ~n13680 ;
  assign n13682 = n1500 & ~n13681 ;
  assign n13683 = n1504 & ~n13682 ;
  assign n13684 = n1508 & ~n13683 ;
  assign n13685 = n1512 & ~n13684 ;
  assign n13686 = n1516 & ~n13685 ;
  assign n13687 = n1520 & ~n13686 ;
  assign n13688 = n1524 & ~n13687 ;
  assign n13689 = n1528 & ~n13688 ;
  assign n13690 = n1532 & ~n13689 ;
  assign n13691 = n1536 & ~n13690 ;
  assign n13692 = n1540 & ~n13691 ;
  assign n13693 = n1544 & ~n13692 ;
  assign n13694 = n1548 & ~n13693 ;
  assign n13695 = n1552 & ~n13694 ;
  assign n13696 = n1556 & ~n13695 ;
  assign n13697 = n1560 & ~n13696 ;
  assign n13698 = n1564 & ~n13697 ;
  assign n13699 = n1568 & ~n13698 ;
  assign n13700 = n1572 & ~n13699 ;
  assign n13701 = n1576 & ~n13700 ;
  assign n13702 = n1580 & ~n13701 ;
  assign n13703 = n1584 & ~n13702 ;
  assign n13704 = n1588 & ~n13703 ;
  assign n13705 = n1592 & ~n13704 ;
  assign n13706 = n1596 & ~n13705 ;
  assign n13707 = n1600 & ~n13706 ;
  assign n13708 = n1604 & ~n13707 ;
  assign n13709 = n1608 & ~n13708 ;
  assign n13710 = n1612 & ~n13709 ;
  assign n13711 = n2656 & ~n13710 ;
  assign n13712 = n2658 & ~n13711 ;
  assign n13713 = n3192 & ~n13712 ;
  assign n13714 = n1962 & ~n13713 ;
  assign n13715 = n1966 & ~n13714 ;
  assign n13716 = n1970 & ~n13715 ;
  assign n13717 = n1974 & ~n13716 ;
  assign n13718 = n1978 & ~n13717 ;
  assign n13719 = n1982 & ~n13718 ;
  assign n13720 = n1986 & ~n13719 ;
  assign n13721 = n1990 & ~n13720 ;
  assign n13722 = n1994 & ~n13721 ;
  assign n13723 = n1998 & ~n13722 ;
  assign n13724 = n2002 & ~n13723 ;
  assign n13725 = n2006 & ~n13724 ;
  assign n13726 = n2010 & ~n13725 ;
  assign n13727 = n2014 & ~n13726 ;
  assign n13728 = n2018 & ~n13727 ;
  assign n13729 = n2022 & ~n13728 ;
  assign n13730 = n2026 & ~n13729 ;
  assign n13731 = n2030 & ~n13730 ;
  assign n13732 = n2034 & ~n13731 ;
  assign n13733 = n2038 & ~n13732 ;
  assign n13734 = n2042 & ~n13733 ;
  assign n13735 = n2046 & ~n13734 ;
  assign n13736 = n2050 & ~n13735 ;
  assign n13737 = n2054 & ~n13736 ;
  assign n13738 = n2058 & ~n13737 ;
  assign n13739 = n2062 & ~n13738 ;
  assign n13740 = n2066 & ~n13739 ;
  assign n13741 = n2070 & ~n13740 ;
  assign n13742 = n2074 & ~n13741 ;
  assign n13743 = n2078 & ~n13742 ;
  assign n13744 = n2082 & ~n13743 ;
  assign n13745 = n2086 & ~n13744 ;
  assign n13746 = n2090 & ~n13745 ;
  assign n13747 = n2094 & ~n13746 ;
  assign n13748 = n2098 & ~n13747 ;
  assign n13749 = n2102 & ~n13748 ;
  assign n13750 = n2106 & ~n13749 ;
  assign n13751 = n2110 & ~n13750 ;
  assign n13752 = n2114 & ~n13751 ;
  assign n13753 = n2118 & ~n13752 ;
  assign n13754 = n2122 & ~n13753 ;
  assign n13755 = ~x195 & ~n2124 ;
  assign n13756 = ~n13754 & n13755 ;
  assign n13759 = ~n13756 & ~x323 ;
  assign n13760 = ~n13758 & ~n13759 ;
  assign n13761 = ~n438 & n1796 ;
  assign n13762 = n1801 & ~n13761 ;
  assign n13763 = n1805 & ~n13762 ;
  assign n13764 = n1809 & ~n13763 ;
  assign n13765 = n1813 & ~n13764 ;
  assign n13766 = n1817 & ~n13765 ;
  assign n13767 = n1821 & ~n13766 ;
  assign n13768 = n1825 & ~n13767 ;
  assign n13769 = n1829 & ~n13768 ;
  assign n13770 = n1833 & ~n13769 ;
  assign n13771 = n1837 & ~n13770 ;
  assign n13772 = n1841 & ~n13771 ;
  assign n13773 = n1845 & ~n13772 ;
  assign n13774 = n1849 & ~n13773 ;
  assign n13775 = n1853 & ~n13774 ;
  assign n13776 = n1857 & ~n13775 ;
  assign n13777 = n1861 & ~n13776 ;
  assign n13778 = n1865 & ~n13777 ;
  assign n13779 = n1869 & ~n13778 ;
  assign n13780 = n1873 & ~n13779 ;
  assign n13781 = n1877 & ~n13780 ;
  assign n13782 = n1881 & ~n13781 ;
  assign n13783 = n1885 & ~n13782 ;
  assign n13784 = n1889 & ~n13783 ;
  assign n13785 = n1893 & ~n13784 ;
  assign n13786 = n1897 & ~n13785 ;
  assign n13787 = n1901 & ~n13786 ;
  assign n13788 = n1905 & ~n13787 ;
  assign n13789 = n1909 & ~n13788 ;
  assign n13790 = n1913 & ~n13789 ;
  assign n13791 = n1917 & ~n13790 ;
  assign n13792 = n1921 & ~n13791 ;
  assign n13793 = n1925 & ~n13792 ;
  assign n13794 = n1929 & ~n13793 ;
  assign n13795 = n1933 & ~n13794 ;
  assign n13796 = n1937 & ~n13795 ;
  assign n13797 = n1941 & ~n13796 ;
  assign n13798 = n1945 & ~n13797 ;
  assign n13799 = n1949 & ~n13798 ;
  assign n13800 = n1953 & ~n13799 ;
  assign n13801 = n2749 & ~n13800 ;
  assign n13802 = n263 & ~n13801 ;
  assign n13803 = n267 & ~n13802 ;
  assign n13804 = n271 & ~n13803 ;
  assign n13805 = n275 & ~n13804 ;
  assign n13806 = n279 & ~n13805 ;
  assign n13807 = n283 & ~n13806 ;
  assign n13808 = n287 & ~n13807 ;
  assign n13809 = n291 & ~n13808 ;
  assign n13810 = n295 & ~n13809 ;
  assign n13811 = n299 & ~n13810 ;
  assign n13812 = n303 & ~n13811 ;
  assign n13813 = n307 & ~n13812 ;
  assign n13814 = n311 & ~n13813 ;
  assign n13815 = n315 & ~n13814 ;
  assign n13816 = n319 & ~n13815 ;
  assign n13817 = n323 & ~n13816 ;
  assign n13818 = n327 & ~n13817 ;
  assign n13819 = n331 & ~n13818 ;
  assign n13820 = n335 & ~n13819 ;
  assign n13821 = n339 & ~n13820 ;
  assign n13822 = n343 & ~n13821 ;
  assign n13823 = n347 & ~n13822 ;
  assign n13824 = n351 & ~n13823 ;
  assign n13825 = n355 & ~n13824 ;
  assign n13826 = n359 & ~n13825 ;
  assign n13827 = n363 & ~n13826 ;
  assign n13828 = n367 & ~n13827 ;
  assign n13829 = n371 & ~n13828 ;
  assign n13830 = n375 & ~n13829 ;
  assign n13831 = n379 & ~n13830 ;
  assign n13832 = n383 & ~n13831 ;
  assign n13833 = n387 & ~n13832 ;
  assign n13834 = n391 & ~n13833 ;
  assign n13835 = n395 & ~n13834 ;
  assign n13836 = n399 & ~n13835 ;
  assign n13837 = n403 & ~n13836 ;
  assign n13838 = n407 & ~n13837 ;
  assign n13839 = n411 & ~n13838 ;
  assign n13840 = n415 & ~n13839 ;
  assign n13841 = n419 & ~n13840 ;
  assign n13842 = n423 & ~n13841 ;
  assign n13843 = n427 & ~n13842 ;
  assign n13844 = n431 & ~n13843 ;
  assign n13845 = x196 & ~n433 ;
  assign n13846 = ~n13844 & n13845 ;
  assign n13934 = n13846 & x324 ;
  assign n13847 = ~n777 & n2133 ;
  assign n13848 = n2138 & ~n13847 ;
  assign n13849 = n2142 & ~n13848 ;
  assign n13850 = n2146 & ~n13849 ;
  assign n13851 = n2150 & ~n13850 ;
  assign n13852 = n2154 & ~n13851 ;
  assign n13853 = n2158 & ~n13852 ;
  assign n13854 = n2162 & ~n13853 ;
  assign n13855 = n2166 & ~n13854 ;
  assign n13856 = n2170 & ~n13855 ;
  assign n13857 = n2174 & ~n13856 ;
  assign n13858 = n2178 & ~n13857 ;
  assign n13859 = n2182 & ~n13858 ;
  assign n13860 = n2186 & ~n13859 ;
  assign n13861 = n2190 & ~n13860 ;
  assign n13862 = n2194 & ~n13861 ;
  assign n13863 = n2198 & ~n13862 ;
  assign n13864 = n2202 & ~n13863 ;
  assign n13865 = n2206 & ~n13864 ;
  assign n13866 = n2210 & ~n13865 ;
  assign n13867 = n2214 & ~n13866 ;
  assign n13868 = n2218 & ~n13867 ;
  assign n13869 = n2222 & ~n13868 ;
  assign n13870 = n2226 & ~n13869 ;
  assign n13871 = n2230 & ~n13870 ;
  assign n13872 = n2234 & ~n13871 ;
  assign n13873 = n2238 & ~n13872 ;
  assign n13874 = n2242 & ~n13873 ;
  assign n13875 = n2246 & ~n13874 ;
  assign n13876 = n2250 & ~n13875 ;
  assign n13877 = n2254 & ~n13876 ;
  assign n13878 = n2258 & ~n13877 ;
  assign n13879 = n2262 & ~n13878 ;
  assign n13880 = n2266 & ~n13879 ;
  assign n13881 = n2270 & ~n13880 ;
  assign n13882 = n2274 & ~n13881 ;
  assign n13883 = n2278 & ~n13882 ;
  assign n13884 = n2282 & ~n13883 ;
  assign n13885 = n2286 & ~n13884 ;
  assign n13886 = n2290 & ~n13885 ;
  assign n13887 = n2836 & ~n13886 ;
  assign n13888 = n602 & ~n13887 ;
  assign n13889 = n606 & ~n13888 ;
  assign n13890 = n610 & ~n13889 ;
  assign n13891 = n614 & ~n13890 ;
  assign n13892 = n618 & ~n13891 ;
  assign n13893 = n622 & ~n13892 ;
  assign n13894 = n626 & ~n13893 ;
  assign n13895 = n630 & ~n13894 ;
  assign n13896 = n634 & ~n13895 ;
  assign n13897 = n638 & ~n13896 ;
  assign n13898 = n642 & ~n13897 ;
  assign n13899 = n646 & ~n13898 ;
  assign n13900 = n650 & ~n13899 ;
  assign n13901 = n654 & ~n13900 ;
  assign n13902 = n658 & ~n13901 ;
  assign n13903 = n662 & ~n13902 ;
  assign n13904 = n666 & ~n13903 ;
  assign n13905 = n670 & ~n13904 ;
  assign n13906 = n674 & ~n13905 ;
  assign n13907 = n678 & ~n13906 ;
  assign n13908 = n682 & ~n13907 ;
  assign n13909 = n686 & ~n13908 ;
  assign n13910 = n690 & ~n13909 ;
  assign n13911 = n694 & ~n13910 ;
  assign n13912 = n698 & ~n13911 ;
  assign n13913 = n702 & ~n13912 ;
  assign n13914 = n706 & ~n13913 ;
  assign n13915 = n710 & ~n13914 ;
  assign n13916 = n714 & ~n13915 ;
  assign n13917 = n718 & ~n13916 ;
  assign n13918 = n722 & ~n13917 ;
  assign n13919 = n726 & ~n13918 ;
  assign n13920 = n730 & ~n13919 ;
  assign n13921 = n734 & ~n13920 ;
  assign n13922 = n738 & ~n13921 ;
  assign n13923 = n742 & ~n13922 ;
  assign n13924 = n746 & ~n13923 ;
  assign n13925 = n750 & ~n13924 ;
  assign n13926 = n754 & ~n13925 ;
  assign n13927 = n758 & ~n13926 ;
  assign n13928 = n762 & ~n13927 ;
  assign n13929 = n766 & ~n13928 ;
  assign n13930 = n770 & ~n13929 ;
  assign n13931 = ~x196 & ~n772 ;
  assign n13932 = ~n13930 & n13931 ;
  assign n13935 = ~n13932 & ~x324 ;
  assign n13936 = ~n13934 & ~n13935 ;
  assign n13937 = n442 & ~n1120 ;
  assign n13938 = n447 & ~n13937 ;
  assign n13939 = n451 & ~n13938 ;
  assign n13940 = n455 & ~n13939 ;
  assign n13941 = n459 & ~n13940 ;
  assign n13942 = n463 & ~n13941 ;
  assign n13943 = n467 & ~n13942 ;
  assign n13944 = n471 & ~n13943 ;
  assign n13945 = n475 & ~n13944 ;
  assign n13946 = n479 & ~n13945 ;
  assign n13947 = n483 & ~n13946 ;
  assign n13948 = n487 & ~n13947 ;
  assign n13949 = n491 & ~n13948 ;
  assign n13950 = n495 & ~n13949 ;
  assign n13951 = n499 & ~n13950 ;
  assign n13952 = n503 & ~n13951 ;
  assign n13953 = n507 & ~n13952 ;
  assign n13954 = n511 & ~n13953 ;
  assign n13955 = n515 & ~n13954 ;
  assign n13956 = n519 & ~n13955 ;
  assign n13957 = n523 & ~n13956 ;
  assign n13958 = n527 & ~n13957 ;
  assign n13959 = n531 & ~n13958 ;
  assign n13960 = n535 & ~n13959 ;
  assign n13961 = n539 & ~n13960 ;
  assign n13962 = n543 & ~n13961 ;
  assign n13963 = n547 & ~n13962 ;
  assign n13964 = n551 & ~n13963 ;
  assign n13965 = n555 & ~n13964 ;
  assign n13966 = n559 & ~n13965 ;
  assign n13967 = n563 & ~n13966 ;
  assign n13968 = n567 & ~n13967 ;
  assign n13969 = n571 & ~n13968 ;
  assign n13970 = n575 & ~n13969 ;
  assign n13971 = n579 & ~n13970 ;
  assign n13972 = n583 & ~n13971 ;
  assign n13973 = n587 & ~n13972 ;
  assign n13974 = n591 & ~n13973 ;
  assign n13975 = n2382 & ~n13974 ;
  assign n13976 = n2384 & ~n13975 ;
  assign n13977 = n2927 & ~n13976 ;
  assign n13978 = n945 & ~n13977 ;
  assign n13979 = n949 & ~n13978 ;
  assign n13980 = n953 & ~n13979 ;
  assign n13981 = n957 & ~n13980 ;
  assign n13982 = n961 & ~n13981 ;
  assign n13983 = n965 & ~n13982 ;
  assign n13984 = n969 & ~n13983 ;
  assign n13985 = n973 & ~n13984 ;
  assign n13986 = n977 & ~n13985 ;
  assign n13987 = n981 & ~n13986 ;
  assign n13988 = n985 & ~n13987 ;
  assign n13989 = n989 & ~n13988 ;
  assign n13990 = n993 & ~n13989 ;
  assign n13991 = n997 & ~n13990 ;
  assign n13992 = n1001 & ~n13991 ;
  assign n13993 = n1005 & ~n13992 ;
  assign n13994 = n1009 & ~n13993 ;
  assign n13995 = n1013 & ~n13994 ;
  assign n13996 = n1017 & ~n13995 ;
  assign n13997 = n1021 & ~n13996 ;
  assign n13998 = n1025 & ~n13997 ;
  assign n13999 = n1029 & ~n13998 ;
  assign n14000 = n1033 & ~n13999 ;
  assign n14001 = n1037 & ~n14000 ;
  assign n14002 = n1041 & ~n14001 ;
  assign n14003 = n1045 & ~n14002 ;
  assign n14004 = n1049 & ~n14003 ;
  assign n14005 = n1053 & ~n14004 ;
  assign n14006 = n1057 & ~n14005 ;
  assign n14007 = n1061 & ~n14006 ;
  assign n14008 = n1065 & ~n14007 ;
  assign n14009 = n1069 & ~n14008 ;
  assign n14010 = n1073 & ~n14009 ;
  assign n14011 = n1077 & ~n14010 ;
  assign n14012 = n1081 & ~n14011 ;
  assign n14013 = n1085 & ~n14012 ;
  assign n14014 = n1089 & ~n14013 ;
  assign n14015 = n1093 & ~n14014 ;
  assign n14016 = n1097 & ~n14015 ;
  assign n14017 = n1101 & ~n14016 ;
  assign n14018 = n1105 & ~n14017 ;
  assign n14019 = n1109 & ~n14018 ;
  assign n14020 = n1113 & ~n14019 ;
  assign n14021 = x197 & ~n1115 ;
  assign n14022 = ~n14020 & n14021 ;
  assign n14110 = n14022 & x325 ;
  assign n14023 = n781 & ~n1459 ;
  assign n14024 = n786 & ~n14023 ;
  assign n14025 = n790 & ~n14024 ;
  assign n14026 = n794 & ~n14025 ;
  assign n14027 = n798 & ~n14026 ;
  assign n14028 = n802 & ~n14027 ;
  assign n14029 = n806 & ~n14028 ;
  assign n14030 = n810 & ~n14029 ;
  assign n14031 = n814 & ~n14030 ;
  assign n14032 = n818 & ~n14031 ;
  assign n14033 = n822 & ~n14032 ;
  assign n14034 = n826 & ~n14033 ;
  assign n14035 = n830 & ~n14034 ;
  assign n14036 = n834 & ~n14035 ;
  assign n14037 = n838 & ~n14036 ;
  assign n14038 = n842 & ~n14037 ;
  assign n14039 = n846 & ~n14038 ;
  assign n14040 = n850 & ~n14039 ;
  assign n14041 = n854 & ~n14040 ;
  assign n14042 = n858 & ~n14041 ;
  assign n14043 = n862 & ~n14042 ;
  assign n14044 = n866 & ~n14043 ;
  assign n14045 = n870 & ~n14044 ;
  assign n14046 = n874 & ~n14045 ;
  assign n14047 = n878 & ~n14046 ;
  assign n14048 = n882 & ~n14047 ;
  assign n14049 = n886 & ~n14048 ;
  assign n14050 = n890 & ~n14049 ;
  assign n14051 = n894 & ~n14050 ;
  assign n14052 = n898 & ~n14051 ;
  assign n14053 = n902 & ~n14052 ;
  assign n14054 = n906 & ~n14053 ;
  assign n14055 = n910 & ~n14054 ;
  assign n14056 = n914 & ~n14055 ;
  assign n14057 = n918 & ~n14056 ;
  assign n14058 = n922 & ~n14057 ;
  assign n14059 = n926 & ~n14058 ;
  assign n14060 = n930 & ~n14059 ;
  assign n14061 = n2472 & ~n14060 ;
  assign n14062 = n2474 & ~n14061 ;
  assign n14063 = n3014 & ~n14062 ;
  assign n14064 = n1284 & ~n14063 ;
  assign n14065 = n1288 & ~n14064 ;
  assign n14066 = n1292 & ~n14065 ;
  assign n14067 = n1296 & ~n14066 ;
  assign n14068 = n1300 & ~n14067 ;
  assign n14069 = n1304 & ~n14068 ;
  assign n14070 = n1308 & ~n14069 ;
  assign n14071 = n1312 & ~n14070 ;
  assign n14072 = n1316 & ~n14071 ;
  assign n14073 = n1320 & ~n14072 ;
  assign n14074 = n1324 & ~n14073 ;
  assign n14075 = n1328 & ~n14074 ;
  assign n14076 = n1332 & ~n14075 ;
  assign n14077 = n1336 & ~n14076 ;
  assign n14078 = n1340 & ~n14077 ;
  assign n14079 = n1344 & ~n14078 ;
  assign n14080 = n1348 & ~n14079 ;
  assign n14081 = n1352 & ~n14080 ;
  assign n14082 = n1356 & ~n14081 ;
  assign n14083 = n1360 & ~n14082 ;
  assign n14084 = n1364 & ~n14083 ;
  assign n14085 = n1368 & ~n14084 ;
  assign n14086 = n1372 & ~n14085 ;
  assign n14087 = n1376 & ~n14086 ;
  assign n14088 = n1380 & ~n14087 ;
  assign n14089 = n1384 & ~n14088 ;
  assign n14090 = n1388 & ~n14089 ;
  assign n14091 = n1392 & ~n14090 ;
  assign n14092 = n1396 & ~n14091 ;
  assign n14093 = n1400 & ~n14092 ;
  assign n14094 = n1404 & ~n14093 ;
  assign n14095 = n1408 & ~n14094 ;
  assign n14096 = n1412 & ~n14095 ;
  assign n14097 = n1416 & ~n14096 ;
  assign n14098 = n1420 & ~n14097 ;
  assign n14099 = n1424 & ~n14098 ;
  assign n14100 = n1428 & ~n14099 ;
  assign n14101 = n1432 & ~n14100 ;
  assign n14102 = n1436 & ~n14101 ;
  assign n14103 = n1440 & ~n14102 ;
  assign n14104 = n1444 & ~n14103 ;
  assign n14105 = n1448 & ~n14104 ;
  assign n14106 = n1452 & ~n14105 ;
  assign n14107 = ~x197 & ~n1454 ;
  assign n14108 = ~n14106 & n14107 ;
  assign n14111 = ~n14108 & ~x325 ;
  assign n14112 = ~n14110 & ~n14111 ;
  assign n14113 = n1124 & ~n1800 ;
  assign n14114 = n1129 & ~n14113 ;
  assign n14115 = n1133 & ~n14114 ;
  assign n14116 = n1137 & ~n14115 ;
  assign n14117 = n1141 & ~n14116 ;
  assign n14118 = n1145 & ~n14117 ;
  assign n14119 = n1149 & ~n14118 ;
  assign n14120 = n1153 & ~n14119 ;
  assign n14121 = n1157 & ~n14120 ;
  assign n14122 = n1161 & ~n14121 ;
  assign n14123 = n1165 & ~n14122 ;
  assign n14124 = n1169 & ~n14123 ;
  assign n14125 = n1173 & ~n14124 ;
  assign n14126 = n1177 & ~n14125 ;
  assign n14127 = n1181 & ~n14126 ;
  assign n14128 = n1185 & ~n14127 ;
  assign n14129 = n1189 & ~n14128 ;
  assign n14130 = n1193 & ~n14129 ;
  assign n14131 = n1197 & ~n14130 ;
  assign n14132 = n1201 & ~n14131 ;
  assign n14133 = n1205 & ~n14132 ;
  assign n14134 = n1209 & ~n14133 ;
  assign n14135 = n1213 & ~n14134 ;
  assign n14136 = n1217 & ~n14135 ;
  assign n14137 = n1221 & ~n14136 ;
  assign n14138 = n1225 & ~n14137 ;
  assign n14139 = n1229 & ~n14138 ;
  assign n14140 = n1233 & ~n14139 ;
  assign n14141 = n1237 & ~n14140 ;
  assign n14142 = n1241 & ~n14141 ;
  assign n14143 = n1245 & ~n14142 ;
  assign n14144 = n1249 & ~n14143 ;
  assign n14145 = n1253 & ~n14144 ;
  assign n14146 = n1257 & ~n14145 ;
  assign n14147 = n1261 & ~n14146 ;
  assign n14148 = n1265 & ~n14147 ;
  assign n14149 = n1269 & ~n14148 ;
  assign n14150 = n1273 & ~n14149 ;
  assign n14151 = n2566 & ~n14150 ;
  assign n14152 = n2568 & ~n14151 ;
  assign n14153 = n3105 & ~n14152 ;
  assign n14154 = n1625 & ~n14153 ;
  assign n14155 = n1629 & ~n14154 ;
  assign n14156 = n1633 & ~n14155 ;
  assign n14157 = n1637 & ~n14156 ;
  assign n14158 = n1641 & ~n14157 ;
  assign n14159 = n1645 & ~n14158 ;
  assign n14160 = n1649 & ~n14159 ;
  assign n14161 = n1653 & ~n14160 ;
  assign n14162 = n1657 & ~n14161 ;
  assign n14163 = n1661 & ~n14162 ;
  assign n14164 = n1665 & ~n14163 ;
  assign n14165 = n1669 & ~n14164 ;
  assign n14166 = n1673 & ~n14165 ;
  assign n14167 = n1677 & ~n14166 ;
  assign n14168 = n1681 & ~n14167 ;
  assign n14169 = n1685 & ~n14168 ;
  assign n14170 = n1689 & ~n14169 ;
  assign n14171 = n1693 & ~n14170 ;
  assign n14172 = n1697 & ~n14171 ;
  assign n14173 = n1701 & ~n14172 ;
  assign n14174 = n1705 & ~n14173 ;
  assign n14175 = n1709 & ~n14174 ;
  assign n14176 = n1713 & ~n14175 ;
  assign n14177 = n1717 & ~n14176 ;
  assign n14178 = n1721 & ~n14177 ;
  assign n14179 = n1725 & ~n14178 ;
  assign n14180 = n1729 & ~n14179 ;
  assign n14181 = n1733 & ~n14180 ;
  assign n14182 = n1737 & ~n14181 ;
  assign n14183 = n1741 & ~n14182 ;
  assign n14184 = n1745 & ~n14183 ;
  assign n14185 = n1749 & ~n14184 ;
  assign n14186 = n1753 & ~n14185 ;
  assign n14187 = n1757 & ~n14186 ;
  assign n14188 = n1761 & ~n14187 ;
  assign n14189 = n1765 & ~n14188 ;
  assign n14190 = n1769 & ~n14189 ;
  assign n14191 = n1773 & ~n14190 ;
  assign n14192 = n1777 & ~n14191 ;
  assign n14193 = n1781 & ~n14192 ;
  assign n14194 = n1785 & ~n14193 ;
  assign n14195 = n1789 & ~n14194 ;
  assign n14196 = n1793 & ~n14195 ;
  assign n14197 = x198 & ~n1795 ;
  assign n14198 = ~n14196 & n14197 ;
  assign n14286 = n14198 & x326 ;
  assign n14199 = n1463 & ~n2137 ;
  assign n14200 = n1468 & ~n14199 ;
  assign n14201 = n1472 & ~n14200 ;
  assign n14202 = n1476 & ~n14201 ;
  assign n14203 = n1480 & ~n14202 ;
  assign n14204 = n1484 & ~n14203 ;
  assign n14205 = n1488 & ~n14204 ;
  assign n14206 = n1492 & ~n14205 ;
  assign n14207 = n1496 & ~n14206 ;
  assign n14208 = n1500 & ~n14207 ;
  assign n14209 = n1504 & ~n14208 ;
  assign n14210 = n1508 & ~n14209 ;
  assign n14211 = n1512 & ~n14210 ;
  assign n14212 = n1516 & ~n14211 ;
  assign n14213 = n1520 & ~n14212 ;
  assign n14214 = n1524 & ~n14213 ;
  assign n14215 = n1528 & ~n14214 ;
  assign n14216 = n1532 & ~n14215 ;
  assign n14217 = n1536 & ~n14216 ;
  assign n14218 = n1540 & ~n14217 ;
  assign n14219 = n1544 & ~n14218 ;
  assign n14220 = n1548 & ~n14219 ;
  assign n14221 = n1552 & ~n14220 ;
  assign n14222 = n1556 & ~n14221 ;
  assign n14223 = n1560 & ~n14222 ;
  assign n14224 = n1564 & ~n14223 ;
  assign n14225 = n1568 & ~n14224 ;
  assign n14226 = n1572 & ~n14225 ;
  assign n14227 = n1576 & ~n14226 ;
  assign n14228 = n1580 & ~n14227 ;
  assign n14229 = n1584 & ~n14228 ;
  assign n14230 = n1588 & ~n14229 ;
  assign n14231 = n1592 & ~n14230 ;
  assign n14232 = n1596 & ~n14231 ;
  assign n14233 = n1600 & ~n14232 ;
  assign n14234 = n1604 & ~n14233 ;
  assign n14235 = n1608 & ~n14234 ;
  assign n14236 = n1612 & ~n14235 ;
  assign n14237 = n2656 & ~n14236 ;
  assign n14238 = n2658 & ~n14237 ;
  assign n14239 = n3192 & ~n14238 ;
  assign n14240 = n1962 & ~n14239 ;
  assign n14241 = n1966 & ~n14240 ;
  assign n14242 = n1970 & ~n14241 ;
  assign n14243 = n1974 & ~n14242 ;
  assign n14244 = n1978 & ~n14243 ;
  assign n14245 = n1982 & ~n14244 ;
  assign n14246 = n1986 & ~n14245 ;
  assign n14247 = n1990 & ~n14246 ;
  assign n14248 = n1994 & ~n14247 ;
  assign n14249 = n1998 & ~n14248 ;
  assign n14250 = n2002 & ~n14249 ;
  assign n14251 = n2006 & ~n14250 ;
  assign n14252 = n2010 & ~n14251 ;
  assign n14253 = n2014 & ~n14252 ;
  assign n14254 = n2018 & ~n14253 ;
  assign n14255 = n2022 & ~n14254 ;
  assign n14256 = n2026 & ~n14255 ;
  assign n14257 = n2030 & ~n14256 ;
  assign n14258 = n2034 & ~n14257 ;
  assign n14259 = n2038 & ~n14258 ;
  assign n14260 = n2042 & ~n14259 ;
  assign n14261 = n2046 & ~n14260 ;
  assign n14262 = n2050 & ~n14261 ;
  assign n14263 = n2054 & ~n14262 ;
  assign n14264 = n2058 & ~n14263 ;
  assign n14265 = n2062 & ~n14264 ;
  assign n14266 = n2066 & ~n14265 ;
  assign n14267 = n2070 & ~n14266 ;
  assign n14268 = n2074 & ~n14267 ;
  assign n14269 = n2078 & ~n14268 ;
  assign n14270 = n2082 & ~n14269 ;
  assign n14271 = n2086 & ~n14270 ;
  assign n14272 = n2090 & ~n14271 ;
  assign n14273 = n2094 & ~n14272 ;
  assign n14274 = n2098 & ~n14273 ;
  assign n14275 = n2102 & ~n14274 ;
  assign n14276 = n2106 & ~n14275 ;
  assign n14277 = n2110 & ~n14276 ;
  assign n14278 = n2114 & ~n14277 ;
  assign n14279 = n2118 & ~n14278 ;
  assign n14280 = n2122 & ~n14279 ;
  assign n14281 = n2126 & ~n14280 ;
  assign n14282 = n2130 & ~n14281 ;
  assign n14283 = ~x198 & ~n2132 ;
  assign n14284 = ~n14282 & n14283 ;
  assign n14287 = ~n14284 & ~x326 ;
  assign n14288 = ~n14286 & ~n14287 ;
  assign n14289 = ~n446 & n1804 ;
  assign n14290 = n1809 & ~n14289 ;
  assign n14291 = n1813 & ~n14290 ;
  assign n14292 = n1817 & ~n14291 ;
  assign n14293 = n1821 & ~n14292 ;
  assign n14294 = n1825 & ~n14293 ;
  assign n14295 = n1829 & ~n14294 ;
  assign n14296 = n1833 & ~n14295 ;
  assign n14297 = n1837 & ~n14296 ;
  assign n14298 = n1841 & ~n14297 ;
  assign n14299 = n1845 & ~n14298 ;
  assign n14300 = n1849 & ~n14299 ;
  assign n14301 = n1853 & ~n14300 ;
  assign n14302 = n1857 & ~n14301 ;
  assign n14303 = n1861 & ~n14302 ;
  assign n14304 = n1865 & ~n14303 ;
  assign n14305 = n1869 & ~n14304 ;
  assign n14306 = n1873 & ~n14305 ;
  assign n14307 = n1877 & ~n14306 ;
  assign n14308 = n1881 & ~n14307 ;
  assign n14309 = n1885 & ~n14308 ;
  assign n14310 = n1889 & ~n14309 ;
  assign n14311 = n1893 & ~n14310 ;
  assign n14312 = n1897 & ~n14311 ;
  assign n14313 = n1901 & ~n14312 ;
  assign n14314 = n1905 & ~n14313 ;
  assign n14315 = n1909 & ~n14314 ;
  assign n14316 = n1913 & ~n14315 ;
  assign n14317 = n1917 & ~n14316 ;
  assign n14318 = n1921 & ~n14317 ;
  assign n14319 = n1925 & ~n14318 ;
  assign n14320 = n1929 & ~n14319 ;
  assign n14321 = n1933 & ~n14320 ;
  assign n14322 = n1937 & ~n14321 ;
  assign n14323 = n1941 & ~n14322 ;
  assign n14324 = n1945 & ~n14323 ;
  assign n14325 = n1949 & ~n14324 ;
  assign n14326 = n1953 & ~n14325 ;
  assign n14327 = n2749 & ~n14326 ;
  assign n14328 = n263 & ~n14327 ;
  assign n14329 = n267 & ~n14328 ;
  assign n14330 = n271 & ~n14329 ;
  assign n14331 = n275 & ~n14330 ;
  assign n14332 = n279 & ~n14331 ;
  assign n14333 = n283 & ~n14332 ;
  assign n14334 = n287 & ~n14333 ;
  assign n14335 = n291 & ~n14334 ;
  assign n14336 = n295 & ~n14335 ;
  assign n14337 = n299 & ~n14336 ;
  assign n14338 = n303 & ~n14337 ;
  assign n14339 = n307 & ~n14338 ;
  assign n14340 = n311 & ~n14339 ;
  assign n14341 = n315 & ~n14340 ;
  assign n14342 = n319 & ~n14341 ;
  assign n14343 = n323 & ~n14342 ;
  assign n14344 = n327 & ~n14343 ;
  assign n14345 = n331 & ~n14344 ;
  assign n14346 = n335 & ~n14345 ;
  assign n14347 = n339 & ~n14346 ;
  assign n14348 = n343 & ~n14347 ;
  assign n14349 = n347 & ~n14348 ;
  assign n14350 = n351 & ~n14349 ;
  assign n14351 = n355 & ~n14350 ;
  assign n14352 = n359 & ~n14351 ;
  assign n14353 = n363 & ~n14352 ;
  assign n14354 = n367 & ~n14353 ;
  assign n14355 = n371 & ~n14354 ;
  assign n14356 = n375 & ~n14355 ;
  assign n14357 = n379 & ~n14356 ;
  assign n14358 = n383 & ~n14357 ;
  assign n14359 = n387 & ~n14358 ;
  assign n14360 = n391 & ~n14359 ;
  assign n14361 = n395 & ~n14360 ;
  assign n14362 = n399 & ~n14361 ;
  assign n14363 = n403 & ~n14362 ;
  assign n14364 = n407 & ~n14363 ;
  assign n14365 = n411 & ~n14364 ;
  assign n14366 = n415 & ~n14365 ;
  assign n14367 = n419 & ~n14366 ;
  assign n14368 = n423 & ~n14367 ;
  assign n14369 = n427 & ~n14368 ;
  assign n14370 = n431 & ~n14369 ;
  assign n14371 = n435 & ~n14370 ;
  assign n14372 = n439 & ~n14371 ;
  assign n14373 = x199 & ~n441 ;
  assign n14374 = ~n14372 & n14373 ;
  assign n14462 = n14374 & x327 ;
  assign n14375 = ~n785 & n2141 ;
  assign n14376 = n2146 & ~n14375 ;
  assign n14377 = n2150 & ~n14376 ;
  assign n14378 = n2154 & ~n14377 ;
  assign n14379 = n2158 & ~n14378 ;
  assign n14380 = n2162 & ~n14379 ;
  assign n14381 = n2166 & ~n14380 ;
  assign n14382 = n2170 & ~n14381 ;
  assign n14383 = n2174 & ~n14382 ;
  assign n14384 = n2178 & ~n14383 ;
  assign n14385 = n2182 & ~n14384 ;
  assign n14386 = n2186 & ~n14385 ;
  assign n14387 = n2190 & ~n14386 ;
  assign n14388 = n2194 & ~n14387 ;
  assign n14389 = n2198 & ~n14388 ;
  assign n14390 = n2202 & ~n14389 ;
  assign n14391 = n2206 & ~n14390 ;
  assign n14392 = n2210 & ~n14391 ;
  assign n14393 = n2214 & ~n14392 ;
  assign n14394 = n2218 & ~n14393 ;
  assign n14395 = n2222 & ~n14394 ;
  assign n14396 = n2226 & ~n14395 ;
  assign n14397 = n2230 & ~n14396 ;
  assign n14398 = n2234 & ~n14397 ;
  assign n14399 = n2238 & ~n14398 ;
  assign n14400 = n2242 & ~n14399 ;
  assign n14401 = n2246 & ~n14400 ;
  assign n14402 = n2250 & ~n14401 ;
  assign n14403 = n2254 & ~n14402 ;
  assign n14404 = n2258 & ~n14403 ;
  assign n14405 = n2262 & ~n14404 ;
  assign n14406 = n2266 & ~n14405 ;
  assign n14407 = n2270 & ~n14406 ;
  assign n14408 = n2274 & ~n14407 ;
  assign n14409 = n2278 & ~n14408 ;
  assign n14410 = n2282 & ~n14409 ;
  assign n14411 = n2286 & ~n14410 ;
  assign n14412 = n2290 & ~n14411 ;
  assign n14413 = n2836 & ~n14412 ;
  assign n14414 = n602 & ~n14413 ;
  assign n14415 = n606 & ~n14414 ;
  assign n14416 = n610 & ~n14415 ;
  assign n14417 = n614 & ~n14416 ;
  assign n14418 = n618 & ~n14417 ;
  assign n14419 = n622 & ~n14418 ;
  assign n14420 = n626 & ~n14419 ;
  assign n14421 = n630 & ~n14420 ;
  assign n14422 = n634 & ~n14421 ;
  assign n14423 = n638 & ~n14422 ;
  assign n14424 = n642 & ~n14423 ;
  assign n14425 = n646 & ~n14424 ;
  assign n14426 = n650 & ~n14425 ;
  assign n14427 = n654 & ~n14426 ;
  assign n14428 = n658 & ~n14427 ;
  assign n14429 = n662 & ~n14428 ;
  assign n14430 = n666 & ~n14429 ;
  assign n14431 = n670 & ~n14430 ;
  assign n14432 = n674 & ~n14431 ;
  assign n14433 = n678 & ~n14432 ;
  assign n14434 = n682 & ~n14433 ;
  assign n14435 = n686 & ~n14434 ;
  assign n14436 = n690 & ~n14435 ;
  assign n14437 = n694 & ~n14436 ;
  assign n14438 = n698 & ~n14437 ;
  assign n14439 = n702 & ~n14438 ;
  assign n14440 = n706 & ~n14439 ;
  assign n14441 = n710 & ~n14440 ;
  assign n14442 = n714 & ~n14441 ;
  assign n14443 = n718 & ~n14442 ;
  assign n14444 = n722 & ~n14443 ;
  assign n14445 = n726 & ~n14444 ;
  assign n14446 = n730 & ~n14445 ;
  assign n14447 = n734 & ~n14446 ;
  assign n14448 = n738 & ~n14447 ;
  assign n14449 = n742 & ~n14448 ;
  assign n14450 = n746 & ~n14449 ;
  assign n14451 = n750 & ~n14450 ;
  assign n14452 = n754 & ~n14451 ;
  assign n14453 = n758 & ~n14452 ;
  assign n14454 = n762 & ~n14453 ;
  assign n14455 = n766 & ~n14454 ;
  assign n14456 = n770 & ~n14455 ;
  assign n14457 = n774 & ~n14456 ;
  assign n14458 = n778 & ~n14457 ;
  assign n14459 = ~x199 & ~n780 ;
  assign n14460 = ~n14458 & n14459 ;
  assign n14463 = ~n14460 & ~x327 ;
  assign n14464 = ~n14462 & ~n14463 ;
  assign n14465 = n450 & ~n1128 ;
  assign n14466 = n455 & ~n14465 ;
  assign n14467 = n459 & ~n14466 ;
  assign n14468 = n463 & ~n14467 ;
  assign n14469 = n467 & ~n14468 ;
  assign n14470 = n471 & ~n14469 ;
  assign n14471 = n475 & ~n14470 ;
  assign n14472 = n479 & ~n14471 ;
  assign n14473 = n483 & ~n14472 ;
  assign n14474 = n487 & ~n14473 ;
  assign n14475 = n491 & ~n14474 ;
  assign n14476 = n495 & ~n14475 ;
  assign n14477 = n499 & ~n14476 ;
  assign n14478 = n503 & ~n14477 ;
  assign n14479 = n507 & ~n14478 ;
  assign n14480 = n511 & ~n14479 ;
  assign n14481 = n515 & ~n14480 ;
  assign n14482 = n519 & ~n14481 ;
  assign n14483 = n523 & ~n14482 ;
  assign n14484 = n527 & ~n14483 ;
  assign n14485 = n531 & ~n14484 ;
  assign n14486 = n535 & ~n14485 ;
  assign n14487 = n539 & ~n14486 ;
  assign n14488 = n543 & ~n14487 ;
  assign n14489 = n547 & ~n14488 ;
  assign n14490 = n551 & ~n14489 ;
  assign n14491 = n555 & ~n14490 ;
  assign n14492 = n559 & ~n14491 ;
  assign n14493 = n563 & ~n14492 ;
  assign n14494 = n567 & ~n14493 ;
  assign n14495 = n571 & ~n14494 ;
  assign n14496 = n575 & ~n14495 ;
  assign n14497 = n579 & ~n14496 ;
  assign n14498 = n583 & ~n14497 ;
  assign n14499 = n587 & ~n14498 ;
  assign n14500 = n591 & ~n14499 ;
  assign n14501 = n2382 & ~n14500 ;
  assign n14502 = n2384 & ~n14501 ;
  assign n14503 = n2927 & ~n14502 ;
  assign n14504 = n945 & ~n14503 ;
  assign n14505 = n949 & ~n14504 ;
  assign n14506 = n953 & ~n14505 ;
  assign n14507 = n957 & ~n14506 ;
  assign n14508 = n961 & ~n14507 ;
  assign n14509 = n965 & ~n14508 ;
  assign n14510 = n969 & ~n14509 ;
  assign n14511 = n973 & ~n14510 ;
  assign n14512 = n977 & ~n14511 ;
  assign n14513 = n981 & ~n14512 ;
  assign n14514 = n985 & ~n14513 ;
  assign n14515 = n989 & ~n14514 ;
  assign n14516 = n993 & ~n14515 ;
  assign n14517 = n997 & ~n14516 ;
  assign n14518 = n1001 & ~n14517 ;
  assign n14519 = n1005 & ~n14518 ;
  assign n14520 = n1009 & ~n14519 ;
  assign n14521 = n1013 & ~n14520 ;
  assign n14522 = n1017 & ~n14521 ;
  assign n14523 = n1021 & ~n14522 ;
  assign n14524 = n1025 & ~n14523 ;
  assign n14525 = n1029 & ~n14524 ;
  assign n14526 = n1033 & ~n14525 ;
  assign n14527 = n1037 & ~n14526 ;
  assign n14528 = n1041 & ~n14527 ;
  assign n14529 = n1045 & ~n14528 ;
  assign n14530 = n1049 & ~n14529 ;
  assign n14531 = n1053 & ~n14530 ;
  assign n14532 = n1057 & ~n14531 ;
  assign n14533 = n1061 & ~n14532 ;
  assign n14534 = n1065 & ~n14533 ;
  assign n14535 = n1069 & ~n14534 ;
  assign n14536 = n1073 & ~n14535 ;
  assign n14537 = n1077 & ~n14536 ;
  assign n14538 = n1081 & ~n14537 ;
  assign n14539 = n1085 & ~n14538 ;
  assign n14540 = n1089 & ~n14539 ;
  assign n14541 = n1093 & ~n14540 ;
  assign n14542 = n1097 & ~n14541 ;
  assign n14543 = n1101 & ~n14542 ;
  assign n14544 = n1105 & ~n14543 ;
  assign n14545 = n1109 & ~n14544 ;
  assign n14546 = n1113 & ~n14545 ;
  assign n14547 = n1117 & ~n14546 ;
  assign n14548 = n1121 & ~n14547 ;
  assign n14549 = x200 & ~n1123 ;
  assign n14550 = ~n14548 & n14549 ;
  assign n14638 = n14550 & x328 ;
  assign n14551 = n789 & ~n1467 ;
  assign n14552 = n794 & ~n14551 ;
  assign n14553 = n798 & ~n14552 ;
  assign n14554 = n802 & ~n14553 ;
  assign n14555 = n806 & ~n14554 ;
  assign n14556 = n810 & ~n14555 ;
  assign n14557 = n814 & ~n14556 ;
  assign n14558 = n818 & ~n14557 ;
  assign n14559 = n822 & ~n14558 ;
  assign n14560 = n826 & ~n14559 ;
  assign n14561 = n830 & ~n14560 ;
  assign n14562 = n834 & ~n14561 ;
  assign n14563 = n838 & ~n14562 ;
  assign n14564 = n842 & ~n14563 ;
  assign n14565 = n846 & ~n14564 ;
  assign n14566 = n850 & ~n14565 ;
  assign n14567 = n854 & ~n14566 ;
  assign n14568 = n858 & ~n14567 ;
  assign n14569 = n862 & ~n14568 ;
  assign n14570 = n866 & ~n14569 ;
  assign n14571 = n870 & ~n14570 ;
  assign n14572 = n874 & ~n14571 ;
  assign n14573 = n878 & ~n14572 ;
  assign n14574 = n882 & ~n14573 ;
  assign n14575 = n886 & ~n14574 ;
  assign n14576 = n890 & ~n14575 ;
  assign n14577 = n894 & ~n14576 ;
  assign n14578 = n898 & ~n14577 ;
  assign n14579 = n902 & ~n14578 ;
  assign n14580 = n906 & ~n14579 ;
  assign n14581 = n910 & ~n14580 ;
  assign n14582 = n914 & ~n14581 ;
  assign n14583 = n918 & ~n14582 ;
  assign n14584 = n922 & ~n14583 ;
  assign n14585 = n926 & ~n14584 ;
  assign n14586 = n930 & ~n14585 ;
  assign n14587 = n2472 & ~n14586 ;
  assign n14588 = n2474 & ~n14587 ;
  assign n14589 = n3014 & ~n14588 ;
  assign n14590 = n1284 & ~n14589 ;
  assign n14591 = n1288 & ~n14590 ;
  assign n14592 = n1292 & ~n14591 ;
  assign n14593 = n1296 & ~n14592 ;
  assign n14594 = n1300 & ~n14593 ;
  assign n14595 = n1304 & ~n14594 ;
  assign n14596 = n1308 & ~n14595 ;
  assign n14597 = n1312 & ~n14596 ;
  assign n14598 = n1316 & ~n14597 ;
  assign n14599 = n1320 & ~n14598 ;
  assign n14600 = n1324 & ~n14599 ;
  assign n14601 = n1328 & ~n14600 ;
  assign n14602 = n1332 & ~n14601 ;
  assign n14603 = n1336 & ~n14602 ;
  assign n14604 = n1340 & ~n14603 ;
  assign n14605 = n1344 & ~n14604 ;
  assign n14606 = n1348 & ~n14605 ;
  assign n14607 = n1352 & ~n14606 ;
  assign n14608 = n1356 & ~n14607 ;
  assign n14609 = n1360 & ~n14608 ;
  assign n14610 = n1364 & ~n14609 ;
  assign n14611 = n1368 & ~n14610 ;
  assign n14612 = n1372 & ~n14611 ;
  assign n14613 = n1376 & ~n14612 ;
  assign n14614 = n1380 & ~n14613 ;
  assign n14615 = n1384 & ~n14614 ;
  assign n14616 = n1388 & ~n14615 ;
  assign n14617 = n1392 & ~n14616 ;
  assign n14618 = n1396 & ~n14617 ;
  assign n14619 = n1400 & ~n14618 ;
  assign n14620 = n1404 & ~n14619 ;
  assign n14621 = n1408 & ~n14620 ;
  assign n14622 = n1412 & ~n14621 ;
  assign n14623 = n1416 & ~n14622 ;
  assign n14624 = n1420 & ~n14623 ;
  assign n14625 = n1424 & ~n14624 ;
  assign n14626 = n1428 & ~n14625 ;
  assign n14627 = n1432 & ~n14626 ;
  assign n14628 = n1436 & ~n14627 ;
  assign n14629 = n1440 & ~n14628 ;
  assign n14630 = n1444 & ~n14629 ;
  assign n14631 = n1448 & ~n14630 ;
  assign n14632 = n1452 & ~n14631 ;
  assign n14633 = n1456 & ~n14632 ;
  assign n14634 = n1460 & ~n14633 ;
  assign n14635 = ~x200 & ~n1462 ;
  assign n14636 = ~n14634 & n14635 ;
  assign n14639 = ~n14636 & ~x328 ;
  assign n14640 = ~n14638 & ~n14639 ;
  assign n14641 = n1132 & ~n1808 ;
  assign n14642 = n1137 & ~n14641 ;
  assign n14643 = n1141 & ~n14642 ;
  assign n14644 = n1145 & ~n14643 ;
  assign n14645 = n1149 & ~n14644 ;
  assign n14646 = n1153 & ~n14645 ;
  assign n14647 = n1157 & ~n14646 ;
  assign n14648 = n1161 & ~n14647 ;
  assign n14649 = n1165 & ~n14648 ;
  assign n14650 = n1169 & ~n14649 ;
  assign n14651 = n1173 & ~n14650 ;
  assign n14652 = n1177 & ~n14651 ;
  assign n14653 = n1181 & ~n14652 ;
  assign n14654 = n1185 & ~n14653 ;
  assign n14655 = n1189 & ~n14654 ;
  assign n14656 = n1193 & ~n14655 ;
  assign n14657 = n1197 & ~n14656 ;
  assign n14658 = n1201 & ~n14657 ;
  assign n14659 = n1205 & ~n14658 ;
  assign n14660 = n1209 & ~n14659 ;
  assign n14661 = n1213 & ~n14660 ;
  assign n14662 = n1217 & ~n14661 ;
  assign n14663 = n1221 & ~n14662 ;
  assign n14664 = n1225 & ~n14663 ;
  assign n14665 = n1229 & ~n14664 ;
  assign n14666 = n1233 & ~n14665 ;
  assign n14667 = n1237 & ~n14666 ;
  assign n14668 = n1241 & ~n14667 ;
  assign n14669 = n1245 & ~n14668 ;
  assign n14670 = n1249 & ~n14669 ;
  assign n14671 = n1253 & ~n14670 ;
  assign n14672 = n1257 & ~n14671 ;
  assign n14673 = n1261 & ~n14672 ;
  assign n14674 = n1265 & ~n14673 ;
  assign n14675 = n1269 & ~n14674 ;
  assign n14676 = n1273 & ~n14675 ;
  assign n14677 = n2566 & ~n14676 ;
  assign n14678 = n2568 & ~n14677 ;
  assign n14679 = n3105 & ~n14678 ;
  assign n14680 = n1625 & ~n14679 ;
  assign n14681 = n1629 & ~n14680 ;
  assign n14682 = n1633 & ~n14681 ;
  assign n14683 = n1637 & ~n14682 ;
  assign n14684 = n1641 & ~n14683 ;
  assign n14685 = n1645 & ~n14684 ;
  assign n14686 = n1649 & ~n14685 ;
  assign n14687 = n1653 & ~n14686 ;
  assign n14688 = n1657 & ~n14687 ;
  assign n14689 = n1661 & ~n14688 ;
  assign n14690 = n1665 & ~n14689 ;
  assign n14691 = n1669 & ~n14690 ;
  assign n14692 = n1673 & ~n14691 ;
  assign n14693 = n1677 & ~n14692 ;
  assign n14694 = n1681 & ~n14693 ;
  assign n14695 = n1685 & ~n14694 ;
  assign n14696 = n1689 & ~n14695 ;
  assign n14697 = n1693 & ~n14696 ;
  assign n14698 = n1697 & ~n14697 ;
  assign n14699 = n1701 & ~n14698 ;
  assign n14700 = n1705 & ~n14699 ;
  assign n14701 = n1709 & ~n14700 ;
  assign n14702 = n1713 & ~n14701 ;
  assign n14703 = n1717 & ~n14702 ;
  assign n14704 = n1721 & ~n14703 ;
  assign n14705 = n1725 & ~n14704 ;
  assign n14706 = n1729 & ~n14705 ;
  assign n14707 = n1733 & ~n14706 ;
  assign n14708 = n1737 & ~n14707 ;
  assign n14709 = n1741 & ~n14708 ;
  assign n14710 = n1745 & ~n14709 ;
  assign n14711 = n1749 & ~n14710 ;
  assign n14712 = n1753 & ~n14711 ;
  assign n14713 = n1757 & ~n14712 ;
  assign n14714 = n1761 & ~n14713 ;
  assign n14715 = n1765 & ~n14714 ;
  assign n14716 = n1769 & ~n14715 ;
  assign n14717 = n1773 & ~n14716 ;
  assign n14718 = n1777 & ~n14717 ;
  assign n14719 = n1781 & ~n14718 ;
  assign n14720 = n1785 & ~n14719 ;
  assign n14721 = n1789 & ~n14720 ;
  assign n14722 = n1793 & ~n14721 ;
  assign n14723 = n1797 & ~n14722 ;
  assign n14724 = n1801 & ~n14723 ;
  assign n14725 = x201 & ~n1803 ;
  assign n14726 = ~n14724 & n14725 ;
  assign n14814 = n14726 & x329 ;
  assign n14727 = n1471 & ~n2145 ;
  assign n14728 = n1476 & ~n14727 ;
  assign n14729 = n1480 & ~n14728 ;
  assign n14730 = n1484 & ~n14729 ;
  assign n14731 = n1488 & ~n14730 ;
  assign n14732 = n1492 & ~n14731 ;
  assign n14733 = n1496 & ~n14732 ;
  assign n14734 = n1500 & ~n14733 ;
  assign n14735 = n1504 & ~n14734 ;
  assign n14736 = n1508 & ~n14735 ;
  assign n14737 = n1512 & ~n14736 ;
  assign n14738 = n1516 & ~n14737 ;
  assign n14739 = n1520 & ~n14738 ;
  assign n14740 = n1524 & ~n14739 ;
  assign n14741 = n1528 & ~n14740 ;
  assign n14742 = n1532 & ~n14741 ;
  assign n14743 = n1536 & ~n14742 ;
  assign n14744 = n1540 & ~n14743 ;
  assign n14745 = n1544 & ~n14744 ;
  assign n14746 = n1548 & ~n14745 ;
  assign n14747 = n1552 & ~n14746 ;
  assign n14748 = n1556 & ~n14747 ;
  assign n14749 = n1560 & ~n14748 ;
  assign n14750 = n1564 & ~n14749 ;
  assign n14751 = n1568 & ~n14750 ;
  assign n14752 = n1572 & ~n14751 ;
  assign n14753 = n1576 & ~n14752 ;
  assign n14754 = n1580 & ~n14753 ;
  assign n14755 = n1584 & ~n14754 ;
  assign n14756 = n1588 & ~n14755 ;
  assign n14757 = n1592 & ~n14756 ;
  assign n14758 = n1596 & ~n14757 ;
  assign n14759 = n1600 & ~n14758 ;
  assign n14760 = n1604 & ~n14759 ;
  assign n14761 = n1608 & ~n14760 ;
  assign n14762 = n1612 & ~n14761 ;
  assign n14763 = n2656 & ~n14762 ;
  assign n14764 = n2658 & ~n14763 ;
  assign n14765 = n3192 & ~n14764 ;
  assign n14766 = n1962 & ~n14765 ;
  assign n14767 = n1966 & ~n14766 ;
  assign n14768 = n1970 & ~n14767 ;
  assign n14769 = n1974 & ~n14768 ;
  assign n14770 = n1978 & ~n14769 ;
  assign n14771 = n1982 & ~n14770 ;
  assign n14772 = n1986 & ~n14771 ;
  assign n14773 = n1990 & ~n14772 ;
  assign n14774 = n1994 & ~n14773 ;
  assign n14775 = n1998 & ~n14774 ;
  assign n14776 = n2002 & ~n14775 ;
  assign n14777 = n2006 & ~n14776 ;
  assign n14778 = n2010 & ~n14777 ;
  assign n14779 = n2014 & ~n14778 ;
  assign n14780 = n2018 & ~n14779 ;
  assign n14781 = n2022 & ~n14780 ;
  assign n14782 = n2026 & ~n14781 ;
  assign n14783 = n2030 & ~n14782 ;
  assign n14784 = n2034 & ~n14783 ;
  assign n14785 = n2038 & ~n14784 ;
  assign n14786 = n2042 & ~n14785 ;
  assign n14787 = n2046 & ~n14786 ;
  assign n14788 = n2050 & ~n14787 ;
  assign n14789 = n2054 & ~n14788 ;
  assign n14790 = n2058 & ~n14789 ;
  assign n14791 = n2062 & ~n14790 ;
  assign n14792 = n2066 & ~n14791 ;
  assign n14793 = n2070 & ~n14792 ;
  assign n14794 = n2074 & ~n14793 ;
  assign n14795 = n2078 & ~n14794 ;
  assign n14796 = n2082 & ~n14795 ;
  assign n14797 = n2086 & ~n14796 ;
  assign n14798 = n2090 & ~n14797 ;
  assign n14799 = n2094 & ~n14798 ;
  assign n14800 = n2098 & ~n14799 ;
  assign n14801 = n2102 & ~n14800 ;
  assign n14802 = n2106 & ~n14801 ;
  assign n14803 = n2110 & ~n14802 ;
  assign n14804 = n2114 & ~n14803 ;
  assign n14805 = n2118 & ~n14804 ;
  assign n14806 = n2122 & ~n14805 ;
  assign n14807 = n2126 & ~n14806 ;
  assign n14808 = n2130 & ~n14807 ;
  assign n14809 = n2134 & ~n14808 ;
  assign n14810 = n2138 & ~n14809 ;
  assign n14811 = ~x201 & ~n2140 ;
  assign n14812 = ~n14810 & n14811 ;
  assign n14815 = ~n14812 & ~x329 ;
  assign n14816 = ~n14814 & ~n14815 ;
  assign n14817 = ~n454 & n1812 ;
  assign n14818 = n1817 & ~n14817 ;
  assign n14819 = n1821 & ~n14818 ;
  assign n14820 = n1825 & ~n14819 ;
  assign n14821 = n1829 & ~n14820 ;
  assign n14822 = n1833 & ~n14821 ;
  assign n14823 = n1837 & ~n14822 ;
  assign n14824 = n1841 & ~n14823 ;
  assign n14825 = n1845 & ~n14824 ;
  assign n14826 = n1849 & ~n14825 ;
  assign n14827 = n1853 & ~n14826 ;
  assign n14828 = n1857 & ~n14827 ;
  assign n14829 = n1861 & ~n14828 ;
  assign n14830 = n1865 & ~n14829 ;
  assign n14831 = n1869 & ~n14830 ;
  assign n14832 = n1873 & ~n14831 ;
  assign n14833 = n1877 & ~n14832 ;
  assign n14834 = n1881 & ~n14833 ;
  assign n14835 = n1885 & ~n14834 ;
  assign n14836 = n1889 & ~n14835 ;
  assign n14837 = n1893 & ~n14836 ;
  assign n14838 = n1897 & ~n14837 ;
  assign n14839 = n1901 & ~n14838 ;
  assign n14840 = n1905 & ~n14839 ;
  assign n14841 = n1909 & ~n14840 ;
  assign n14842 = n1913 & ~n14841 ;
  assign n14843 = n1917 & ~n14842 ;
  assign n14844 = n1921 & ~n14843 ;
  assign n14845 = n1925 & ~n14844 ;
  assign n14846 = n1929 & ~n14845 ;
  assign n14847 = n1933 & ~n14846 ;
  assign n14848 = n1937 & ~n14847 ;
  assign n14849 = n1941 & ~n14848 ;
  assign n14850 = n1945 & ~n14849 ;
  assign n14851 = n1949 & ~n14850 ;
  assign n14852 = n1953 & ~n14851 ;
  assign n14853 = n2749 & ~n14852 ;
  assign n14854 = n263 & ~n14853 ;
  assign n14855 = n267 & ~n14854 ;
  assign n14856 = n271 & ~n14855 ;
  assign n14857 = n275 & ~n14856 ;
  assign n14858 = n279 & ~n14857 ;
  assign n14859 = n283 & ~n14858 ;
  assign n14860 = n287 & ~n14859 ;
  assign n14861 = n291 & ~n14860 ;
  assign n14862 = n295 & ~n14861 ;
  assign n14863 = n299 & ~n14862 ;
  assign n14864 = n303 & ~n14863 ;
  assign n14865 = n307 & ~n14864 ;
  assign n14866 = n311 & ~n14865 ;
  assign n14867 = n315 & ~n14866 ;
  assign n14868 = n319 & ~n14867 ;
  assign n14869 = n323 & ~n14868 ;
  assign n14870 = n327 & ~n14869 ;
  assign n14871 = n331 & ~n14870 ;
  assign n14872 = n335 & ~n14871 ;
  assign n14873 = n339 & ~n14872 ;
  assign n14874 = n343 & ~n14873 ;
  assign n14875 = n347 & ~n14874 ;
  assign n14876 = n351 & ~n14875 ;
  assign n14877 = n355 & ~n14876 ;
  assign n14878 = n359 & ~n14877 ;
  assign n14879 = n363 & ~n14878 ;
  assign n14880 = n367 & ~n14879 ;
  assign n14881 = n371 & ~n14880 ;
  assign n14882 = n375 & ~n14881 ;
  assign n14883 = n379 & ~n14882 ;
  assign n14884 = n383 & ~n14883 ;
  assign n14885 = n387 & ~n14884 ;
  assign n14886 = n391 & ~n14885 ;
  assign n14887 = n395 & ~n14886 ;
  assign n14888 = n399 & ~n14887 ;
  assign n14889 = n403 & ~n14888 ;
  assign n14890 = n407 & ~n14889 ;
  assign n14891 = n411 & ~n14890 ;
  assign n14892 = n415 & ~n14891 ;
  assign n14893 = n419 & ~n14892 ;
  assign n14894 = n423 & ~n14893 ;
  assign n14895 = n427 & ~n14894 ;
  assign n14896 = n431 & ~n14895 ;
  assign n14897 = n435 & ~n14896 ;
  assign n14898 = n439 & ~n14897 ;
  assign n14899 = n443 & ~n14898 ;
  assign n14900 = n447 & ~n14899 ;
  assign n14901 = x202 & ~n449 ;
  assign n14902 = ~n14900 & n14901 ;
  assign n14990 = n14902 & x330 ;
  assign n14903 = ~n793 & n2149 ;
  assign n14904 = n2154 & ~n14903 ;
  assign n14905 = n2158 & ~n14904 ;
  assign n14906 = n2162 & ~n14905 ;
  assign n14907 = n2166 & ~n14906 ;
  assign n14908 = n2170 & ~n14907 ;
  assign n14909 = n2174 & ~n14908 ;
  assign n14910 = n2178 & ~n14909 ;
  assign n14911 = n2182 & ~n14910 ;
  assign n14912 = n2186 & ~n14911 ;
  assign n14913 = n2190 & ~n14912 ;
  assign n14914 = n2194 & ~n14913 ;
  assign n14915 = n2198 & ~n14914 ;
  assign n14916 = n2202 & ~n14915 ;
  assign n14917 = n2206 & ~n14916 ;
  assign n14918 = n2210 & ~n14917 ;
  assign n14919 = n2214 & ~n14918 ;
  assign n14920 = n2218 & ~n14919 ;
  assign n14921 = n2222 & ~n14920 ;
  assign n14922 = n2226 & ~n14921 ;
  assign n14923 = n2230 & ~n14922 ;
  assign n14924 = n2234 & ~n14923 ;
  assign n14925 = n2238 & ~n14924 ;
  assign n14926 = n2242 & ~n14925 ;
  assign n14927 = n2246 & ~n14926 ;
  assign n14928 = n2250 & ~n14927 ;
  assign n14929 = n2254 & ~n14928 ;
  assign n14930 = n2258 & ~n14929 ;
  assign n14931 = n2262 & ~n14930 ;
  assign n14932 = n2266 & ~n14931 ;
  assign n14933 = n2270 & ~n14932 ;
  assign n14934 = n2274 & ~n14933 ;
  assign n14935 = n2278 & ~n14934 ;
  assign n14936 = n2282 & ~n14935 ;
  assign n14937 = n2286 & ~n14936 ;
  assign n14938 = n2290 & ~n14937 ;
  assign n14939 = n2836 & ~n14938 ;
  assign n14940 = n602 & ~n14939 ;
  assign n14941 = n606 & ~n14940 ;
  assign n14942 = n610 & ~n14941 ;
  assign n14943 = n614 & ~n14942 ;
  assign n14944 = n618 & ~n14943 ;
  assign n14945 = n622 & ~n14944 ;
  assign n14946 = n626 & ~n14945 ;
  assign n14947 = n630 & ~n14946 ;
  assign n14948 = n634 & ~n14947 ;
  assign n14949 = n638 & ~n14948 ;
  assign n14950 = n642 & ~n14949 ;
  assign n14951 = n646 & ~n14950 ;
  assign n14952 = n650 & ~n14951 ;
  assign n14953 = n654 & ~n14952 ;
  assign n14954 = n658 & ~n14953 ;
  assign n14955 = n662 & ~n14954 ;
  assign n14956 = n666 & ~n14955 ;
  assign n14957 = n670 & ~n14956 ;
  assign n14958 = n674 & ~n14957 ;
  assign n14959 = n678 & ~n14958 ;
  assign n14960 = n682 & ~n14959 ;
  assign n14961 = n686 & ~n14960 ;
  assign n14962 = n690 & ~n14961 ;
  assign n14963 = n694 & ~n14962 ;
  assign n14964 = n698 & ~n14963 ;
  assign n14965 = n702 & ~n14964 ;
  assign n14966 = n706 & ~n14965 ;
  assign n14967 = n710 & ~n14966 ;
  assign n14968 = n714 & ~n14967 ;
  assign n14969 = n718 & ~n14968 ;
  assign n14970 = n722 & ~n14969 ;
  assign n14971 = n726 & ~n14970 ;
  assign n14972 = n730 & ~n14971 ;
  assign n14973 = n734 & ~n14972 ;
  assign n14974 = n738 & ~n14973 ;
  assign n14975 = n742 & ~n14974 ;
  assign n14976 = n746 & ~n14975 ;
  assign n14977 = n750 & ~n14976 ;
  assign n14978 = n754 & ~n14977 ;
  assign n14979 = n758 & ~n14978 ;
  assign n14980 = n762 & ~n14979 ;
  assign n14981 = n766 & ~n14980 ;
  assign n14982 = n770 & ~n14981 ;
  assign n14983 = n774 & ~n14982 ;
  assign n14984 = n778 & ~n14983 ;
  assign n14985 = n782 & ~n14984 ;
  assign n14986 = n786 & ~n14985 ;
  assign n14987 = ~x202 & ~n788 ;
  assign n14988 = ~n14986 & n14987 ;
  assign n14991 = ~n14988 & ~x330 ;
  assign n14992 = ~n14990 & ~n14991 ;
  assign n14993 = n458 & ~n1136 ;
  assign n14994 = n463 & ~n14993 ;
  assign n14995 = n467 & ~n14994 ;
  assign n14996 = n471 & ~n14995 ;
  assign n14997 = n475 & ~n14996 ;
  assign n14998 = n479 & ~n14997 ;
  assign n14999 = n483 & ~n14998 ;
  assign n15000 = n487 & ~n14999 ;
  assign n15001 = n491 & ~n15000 ;
  assign n15002 = n495 & ~n15001 ;
  assign n15003 = n499 & ~n15002 ;
  assign n15004 = n503 & ~n15003 ;
  assign n15005 = n507 & ~n15004 ;
  assign n15006 = n511 & ~n15005 ;
  assign n15007 = n515 & ~n15006 ;
  assign n15008 = n519 & ~n15007 ;
  assign n15009 = n523 & ~n15008 ;
  assign n15010 = n527 & ~n15009 ;
  assign n15011 = n531 & ~n15010 ;
  assign n15012 = n535 & ~n15011 ;
  assign n15013 = n539 & ~n15012 ;
  assign n15014 = n543 & ~n15013 ;
  assign n15015 = n547 & ~n15014 ;
  assign n15016 = n551 & ~n15015 ;
  assign n15017 = n555 & ~n15016 ;
  assign n15018 = n559 & ~n15017 ;
  assign n15019 = n563 & ~n15018 ;
  assign n15020 = n567 & ~n15019 ;
  assign n15021 = n571 & ~n15020 ;
  assign n15022 = n575 & ~n15021 ;
  assign n15023 = n579 & ~n15022 ;
  assign n15024 = n583 & ~n15023 ;
  assign n15025 = n587 & ~n15024 ;
  assign n15026 = n591 & ~n15025 ;
  assign n15027 = n2382 & ~n15026 ;
  assign n15028 = n2384 & ~n15027 ;
  assign n15029 = n2927 & ~n15028 ;
  assign n15030 = n945 & ~n15029 ;
  assign n15031 = n949 & ~n15030 ;
  assign n15032 = n953 & ~n15031 ;
  assign n15033 = n957 & ~n15032 ;
  assign n15034 = n961 & ~n15033 ;
  assign n15035 = n965 & ~n15034 ;
  assign n15036 = n969 & ~n15035 ;
  assign n15037 = n973 & ~n15036 ;
  assign n15038 = n977 & ~n15037 ;
  assign n15039 = n981 & ~n15038 ;
  assign n15040 = n985 & ~n15039 ;
  assign n15041 = n989 & ~n15040 ;
  assign n15042 = n993 & ~n15041 ;
  assign n15043 = n997 & ~n15042 ;
  assign n15044 = n1001 & ~n15043 ;
  assign n15045 = n1005 & ~n15044 ;
  assign n15046 = n1009 & ~n15045 ;
  assign n15047 = n1013 & ~n15046 ;
  assign n15048 = n1017 & ~n15047 ;
  assign n15049 = n1021 & ~n15048 ;
  assign n15050 = n1025 & ~n15049 ;
  assign n15051 = n1029 & ~n15050 ;
  assign n15052 = n1033 & ~n15051 ;
  assign n15053 = n1037 & ~n15052 ;
  assign n15054 = n1041 & ~n15053 ;
  assign n15055 = n1045 & ~n15054 ;
  assign n15056 = n1049 & ~n15055 ;
  assign n15057 = n1053 & ~n15056 ;
  assign n15058 = n1057 & ~n15057 ;
  assign n15059 = n1061 & ~n15058 ;
  assign n15060 = n1065 & ~n15059 ;
  assign n15061 = n1069 & ~n15060 ;
  assign n15062 = n1073 & ~n15061 ;
  assign n15063 = n1077 & ~n15062 ;
  assign n15064 = n1081 & ~n15063 ;
  assign n15065 = n1085 & ~n15064 ;
  assign n15066 = n1089 & ~n15065 ;
  assign n15067 = n1093 & ~n15066 ;
  assign n15068 = n1097 & ~n15067 ;
  assign n15069 = n1101 & ~n15068 ;
  assign n15070 = n1105 & ~n15069 ;
  assign n15071 = n1109 & ~n15070 ;
  assign n15072 = n1113 & ~n15071 ;
  assign n15073 = n1117 & ~n15072 ;
  assign n15074 = n1121 & ~n15073 ;
  assign n15075 = n1125 & ~n15074 ;
  assign n15076 = n1129 & ~n15075 ;
  assign n15077 = x203 & ~n1131 ;
  assign n15078 = ~n15076 & n15077 ;
  assign n15166 = n15078 & x331 ;
  assign n15079 = n797 & ~n1475 ;
  assign n15080 = n802 & ~n15079 ;
  assign n15081 = n806 & ~n15080 ;
  assign n15082 = n810 & ~n15081 ;
  assign n15083 = n814 & ~n15082 ;
  assign n15084 = n818 & ~n15083 ;
  assign n15085 = n822 & ~n15084 ;
  assign n15086 = n826 & ~n15085 ;
  assign n15087 = n830 & ~n15086 ;
  assign n15088 = n834 & ~n15087 ;
  assign n15089 = n838 & ~n15088 ;
  assign n15090 = n842 & ~n15089 ;
  assign n15091 = n846 & ~n15090 ;
  assign n15092 = n850 & ~n15091 ;
  assign n15093 = n854 & ~n15092 ;
  assign n15094 = n858 & ~n15093 ;
  assign n15095 = n862 & ~n15094 ;
  assign n15096 = n866 & ~n15095 ;
  assign n15097 = n870 & ~n15096 ;
  assign n15098 = n874 & ~n15097 ;
  assign n15099 = n878 & ~n15098 ;
  assign n15100 = n882 & ~n15099 ;
  assign n15101 = n886 & ~n15100 ;
  assign n15102 = n890 & ~n15101 ;
  assign n15103 = n894 & ~n15102 ;
  assign n15104 = n898 & ~n15103 ;
  assign n15105 = n902 & ~n15104 ;
  assign n15106 = n906 & ~n15105 ;
  assign n15107 = n910 & ~n15106 ;
  assign n15108 = n914 & ~n15107 ;
  assign n15109 = n918 & ~n15108 ;
  assign n15110 = n922 & ~n15109 ;
  assign n15111 = n926 & ~n15110 ;
  assign n15112 = n930 & ~n15111 ;
  assign n15113 = n2472 & ~n15112 ;
  assign n15114 = n2474 & ~n15113 ;
  assign n15115 = n3014 & ~n15114 ;
  assign n15116 = n1284 & ~n15115 ;
  assign n15117 = n1288 & ~n15116 ;
  assign n15118 = n1292 & ~n15117 ;
  assign n15119 = n1296 & ~n15118 ;
  assign n15120 = n1300 & ~n15119 ;
  assign n15121 = n1304 & ~n15120 ;
  assign n15122 = n1308 & ~n15121 ;
  assign n15123 = n1312 & ~n15122 ;
  assign n15124 = n1316 & ~n15123 ;
  assign n15125 = n1320 & ~n15124 ;
  assign n15126 = n1324 & ~n15125 ;
  assign n15127 = n1328 & ~n15126 ;
  assign n15128 = n1332 & ~n15127 ;
  assign n15129 = n1336 & ~n15128 ;
  assign n15130 = n1340 & ~n15129 ;
  assign n15131 = n1344 & ~n15130 ;
  assign n15132 = n1348 & ~n15131 ;
  assign n15133 = n1352 & ~n15132 ;
  assign n15134 = n1356 & ~n15133 ;
  assign n15135 = n1360 & ~n15134 ;
  assign n15136 = n1364 & ~n15135 ;
  assign n15137 = n1368 & ~n15136 ;
  assign n15138 = n1372 & ~n15137 ;
  assign n15139 = n1376 & ~n15138 ;
  assign n15140 = n1380 & ~n15139 ;
  assign n15141 = n1384 & ~n15140 ;
  assign n15142 = n1388 & ~n15141 ;
  assign n15143 = n1392 & ~n15142 ;
  assign n15144 = n1396 & ~n15143 ;
  assign n15145 = n1400 & ~n15144 ;
  assign n15146 = n1404 & ~n15145 ;
  assign n15147 = n1408 & ~n15146 ;
  assign n15148 = n1412 & ~n15147 ;
  assign n15149 = n1416 & ~n15148 ;
  assign n15150 = n1420 & ~n15149 ;
  assign n15151 = n1424 & ~n15150 ;
  assign n15152 = n1428 & ~n15151 ;
  assign n15153 = n1432 & ~n15152 ;
  assign n15154 = n1436 & ~n15153 ;
  assign n15155 = n1440 & ~n15154 ;
  assign n15156 = n1444 & ~n15155 ;
  assign n15157 = n1448 & ~n15156 ;
  assign n15158 = n1452 & ~n15157 ;
  assign n15159 = n1456 & ~n15158 ;
  assign n15160 = n1460 & ~n15159 ;
  assign n15161 = n1464 & ~n15160 ;
  assign n15162 = n1468 & ~n15161 ;
  assign n15163 = ~x203 & ~n1470 ;
  assign n15164 = ~n15162 & n15163 ;
  assign n15167 = ~n15164 & ~x331 ;
  assign n15168 = ~n15166 & ~n15167 ;
  assign n15169 = n1140 & ~n1816 ;
  assign n15170 = n1145 & ~n15169 ;
  assign n15171 = n1149 & ~n15170 ;
  assign n15172 = n1153 & ~n15171 ;
  assign n15173 = n1157 & ~n15172 ;
  assign n15174 = n1161 & ~n15173 ;
  assign n15175 = n1165 & ~n15174 ;
  assign n15176 = n1169 & ~n15175 ;
  assign n15177 = n1173 & ~n15176 ;
  assign n15178 = n1177 & ~n15177 ;
  assign n15179 = n1181 & ~n15178 ;
  assign n15180 = n1185 & ~n15179 ;
  assign n15181 = n1189 & ~n15180 ;
  assign n15182 = n1193 & ~n15181 ;
  assign n15183 = n1197 & ~n15182 ;
  assign n15184 = n1201 & ~n15183 ;
  assign n15185 = n1205 & ~n15184 ;
  assign n15186 = n1209 & ~n15185 ;
  assign n15187 = n1213 & ~n15186 ;
  assign n15188 = n1217 & ~n15187 ;
  assign n15189 = n1221 & ~n15188 ;
  assign n15190 = n1225 & ~n15189 ;
  assign n15191 = n1229 & ~n15190 ;
  assign n15192 = n1233 & ~n15191 ;
  assign n15193 = n1237 & ~n15192 ;
  assign n15194 = n1241 & ~n15193 ;
  assign n15195 = n1245 & ~n15194 ;
  assign n15196 = n1249 & ~n15195 ;
  assign n15197 = n1253 & ~n15196 ;
  assign n15198 = n1257 & ~n15197 ;
  assign n15199 = n1261 & ~n15198 ;
  assign n15200 = n1265 & ~n15199 ;
  assign n15201 = n1269 & ~n15200 ;
  assign n15202 = n1273 & ~n15201 ;
  assign n15203 = n2566 & ~n15202 ;
  assign n15204 = n2568 & ~n15203 ;
  assign n15205 = n3105 & ~n15204 ;
  assign n15206 = n1625 & ~n15205 ;
  assign n15207 = n1629 & ~n15206 ;
  assign n15208 = n1633 & ~n15207 ;
  assign n15209 = n1637 & ~n15208 ;
  assign n15210 = n1641 & ~n15209 ;
  assign n15211 = n1645 & ~n15210 ;
  assign n15212 = n1649 & ~n15211 ;
  assign n15213 = n1653 & ~n15212 ;
  assign n15214 = n1657 & ~n15213 ;
  assign n15215 = n1661 & ~n15214 ;
  assign n15216 = n1665 & ~n15215 ;
  assign n15217 = n1669 & ~n15216 ;
  assign n15218 = n1673 & ~n15217 ;
  assign n15219 = n1677 & ~n15218 ;
  assign n15220 = n1681 & ~n15219 ;
  assign n15221 = n1685 & ~n15220 ;
  assign n15222 = n1689 & ~n15221 ;
  assign n15223 = n1693 & ~n15222 ;
  assign n15224 = n1697 & ~n15223 ;
  assign n15225 = n1701 & ~n15224 ;
  assign n15226 = n1705 & ~n15225 ;
  assign n15227 = n1709 & ~n15226 ;
  assign n15228 = n1713 & ~n15227 ;
  assign n15229 = n1717 & ~n15228 ;
  assign n15230 = n1721 & ~n15229 ;
  assign n15231 = n1725 & ~n15230 ;
  assign n15232 = n1729 & ~n15231 ;
  assign n15233 = n1733 & ~n15232 ;
  assign n15234 = n1737 & ~n15233 ;
  assign n15235 = n1741 & ~n15234 ;
  assign n15236 = n1745 & ~n15235 ;
  assign n15237 = n1749 & ~n15236 ;
  assign n15238 = n1753 & ~n15237 ;
  assign n15239 = n1757 & ~n15238 ;
  assign n15240 = n1761 & ~n15239 ;
  assign n15241 = n1765 & ~n15240 ;
  assign n15242 = n1769 & ~n15241 ;
  assign n15243 = n1773 & ~n15242 ;
  assign n15244 = n1777 & ~n15243 ;
  assign n15245 = n1781 & ~n15244 ;
  assign n15246 = n1785 & ~n15245 ;
  assign n15247 = n1789 & ~n15246 ;
  assign n15248 = n1793 & ~n15247 ;
  assign n15249 = n1797 & ~n15248 ;
  assign n15250 = n1801 & ~n15249 ;
  assign n15251 = n1805 & ~n15250 ;
  assign n15252 = n1809 & ~n15251 ;
  assign n15253 = x204 & ~n1811 ;
  assign n15254 = ~n15252 & n15253 ;
  assign n15342 = n15254 & x332 ;
  assign n15255 = n1479 & ~n2153 ;
  assign n15256 = n1484 & ~n15255 ;
  assign n15257 = n1488 & ~n15256 ;
  assign n15258 = n1492 & ~n15257 ;
  assign n15259 = n1496 & ~n15258 ;
  assign n15260 = n1500 & ~n15259 ;
  assign n15261 = n1504 & ~n15260 ;
  assign n15262 = n1508 & ~n15261 ;
  assign n15263 = n1512 & ~n15262 ;
  assign n15264 = n1516 & ~n15263 ;
  assign n15265 = n1520 & ~n15264 ;
  assign n15266 = n1524 & ~n15265 ;
  assign n15267 = n1528 & ~n15266 ;
  assign n15268 = n1532 & ~n15267 ;
  assign n15269 = n1536 & ~n15268 ;
  assign n15270 = n1540 & ~n15269 ;
  assign n15271 = n1544 & ~n15270 ;
  assign n15272 = n1548 & ~n15271 ;
  assign n15273 = n1552 & ~n15272 ;
  assign n15274 = n1556 & ~n15273 ;
  assign n15275 = n1560 & ~n15274 ;
  assign n15276 = n1564 & ~n15275 ;
  assign n15277 = n1568 & ~n15276 ;
  assign n15278 = n1572 & ~n15277 ;
  assign n15279 = n1576 & ~n15278 ;
  assign n15280 = n1580 & ~n15279 ;
  assign n15281 = n1584 & ~n15280 ;
  assign n15282 = n1588 & ~n15281 ;
  assign n15283 = n1592 & ~n15282 ;
  assign n15284 = n1596 & ~n15283 ;
  assign n15285 = n1600 & ~n15284 ;
  assign n15286 = n1604 & ~n15285 ;
  assign n15287 = n1608 & ~n15286 ;
  assign n15288 = n1612 & ~n15287 ;
  assign n15289 = n2656 & ~n15288 ;
  assign n15290 = n2658 & ~n15289 ;
  assign n15291 = n3192 & ~n15290 ;
  assign n15292 = n1962 & ~n15291 ;
  assign n15293 = n1966 & ~n15292 ;
  assign n15294 = n1970 & ~n15293 ;
  assign n15295 = n1974 & ~n15294 ;
  assign n15296 = n1978 & ~n15295 ;
  assign n15297 = n1982 & ~n15296 ;
  assign n15298 = n1986 & ~n15297 ;
  assign n15299 = n1990 & ~n15298 ;
  assign n15300 = n1994 & ~n15299 ;
  assign n15301 = n1998 & ~n15300 ;
  assign n15302 = n2002 & ~n15301 ;
  assign n15303 = n2006 & ~n15302 ;
  assign n15304 = n2010 & ~n15303 ;
  assign n15305 = n2014 & ~n15304 ;
  assign n15306 = n2018 & ~n15305 ;
  assign n15307 = n2022 & ~n15306 ;
  assign n15308 = n2026 & ~n15307 ;
  assign n15309 = n2030 & ~n15308 ;
  assign n15310 = n2034 & ~n15309 ;
  assign n15311 = n2038 & ~n15310 ;
  assign n15312 = n2042 & ~n15311 ;
  assign n15313 = n2046 & ~n15312 ;
  assign n15314 = n2050 & ~n15313 ;
  assign n15315 = n2054 & ~n15314 ;
  assign n15316 = n2058 & ~n15315 ;
  assign n15317 = n2062 & ~n15316 ;
  assign n15318 = n2066 & ~n15317 ;
  assign n15319 = n2070 & ~n15318 ;
  assign n15320 = n2074 & ~n15319 ;
  assign n15321 = n2078 & ~n15320 ;
  assign n15322 = n2082 & ~n15321 ;
  assign n15323 = n2086 & ~n15322 ;
  assign n15324 = n2090 & ~n15323 ;
  assign n15325 = n2094 & ~n15324 ;
  assign n15326 = n2098 & ~n15325 ;
  assign n15327 = n2102 & ~n15326 ;
  assign n15328 = n2106 & ~n15327 ;
  assign n15329 = n2110 & ~n15328 ;
  assign n15330 = n2114 & ~n15329 ;
  assign n15331 = n2118 & ~n15330 ;
  assign n15332 = n2122 & ~n15331 ;
  assign n15333 = n2126 & ~n15332 ;
  assign n15334 = n2130 & ~n15333 ;
  assign n15335 = n2134 & ~n15334 ;
  assign n15336 = n2138 & ~n15335 ;
  assign n15337 = n2142 & ~n15336 ;
  assign n15338 = n2146 & ~n15337 ;
  assign n15339 = ~x204 & ~n2148 ;
  assign n15340 = ~n15338 & n15339 ;
  assign n15343 = ~n15340 & ~x332 ;
  assign n15344 = ~n15342 & ~n15343 ;
  assign n15345 = ~n462 & n1820 ;
  assign n15346 = n1825 & ~n15345 ;
  assign n15347 = n1829 & ~n15346 ;
  assign n15348 = n1833 & ~n15347 ;
  assign n15349 = n1837 & ~n15348 ;
  assign n15350 = n1841 & ~n15349 ;
  assign n15351 = n1845 & ~n15350 ;
  assign n15352 = n1849 & ~n15351 ;
  assign n15353 = n1853 & ~n15352 ;
  assign n15354 = n1857 & ~n15353 ;
  assign n15355 = n1861 & ~n15354 ;
  assign n15356 = n1865 & ~n15355 ;
  assign n15357 = n1869 & ~n15356 ;
  assign n15358 = n1873 & ~n15357 ;
  assign n15359 = n1877 & ~n15358 ;
  assign n15360 = n1881 & ~n15359 ;
  assign n15361 = n1885 & ~n15360 ;
  assign n15362 = n1889 & ~n15361 ;
  assign n15363 = n1893 & ~n15362 ;
  assign n15364 = n1897 & ~n15363 ;
  assign n15365 = n1901 & ~n15364 ;
  assign n15366 = n1905 & ~n15365 ;
  assign n15367 = n1909 & ~n15366 ;
  assign n15368 = n1913 & ~n15367 ;
  assign n15369 = n1917 & ~n15368 ;
  assign n15370 = n1921 & ~n15369 ;
  assign n15371 = n1925 & ~n15370 ;
  assign n15372 = n1929 & ~n15371 ;
  assign n15373 = n1933 & ~n15372 ;
  assign n15374 = n1937 & ~n15373 ;
  assign n15375 = n1941 & ~n15374 ;
  assign n15376 = n1945 & ~n15375 ;
  assign n15377 = n1949 & ~n15376 ;
  assign n15378 = n1953 & ~n15377 ;
  assign n15379 = n2749 & ~n15378 ;
  assign n15380 = n263 & ~n15379 ;
  assign n15381 = n267 & ~n15380 ;
  assign n15382 = n271 & ~n15381 ;
  assign n15383 = n275 & ~n15382 ;
  assign n15384 = n279 & ~n15383 ;
  assign n15385 = n283 & ~n15384 ;
  assign n15386 = n287 & ~n15385 ;
  assign n15387 = n291 & ~n15386 ;
  assign n15388 = n295 & ~n15387 ;
  assign n15389 = n299 & ~n15388 ;
  assign n15390 = n303 & ~n15389 ;
  assign n15391 = n307 & ~n15390 ;
  assign n15392 = n311 & ~n15391 ;
  assign n15393 = n315 & ~n15392 ;
  assign n15394 = n319 & ~n15393 ;
  assign n15395 = n323 & ~n15394 ;
  assign n15396 = n327 & ~n15395 ;
  assign n15397 = n331 & ~n15396 ;
  assign n15398 = n335 & ~n15397 ;
  assign n15399 = n339 & ~n15398 ;
  assign n15400 = n343 & ~n15399 ;
  assign n15401 = n347 & ~n15400 ;
  assign n15402 = n351 & ~n15401 ;
  assign n15403 = n355 & ~n15402 ;
  assign n15404 = n359 & ~n15403 ;
  assign n15405 = n363 & ~n15404 ;
  assign n15406 = n367 & ~n15405 ;
  assign n15407 = n371 & ~n15406 ;
  assign n15408 = n375 & ~n15407 ;
  assign n15409 = n379 & ~n15408 ;
  assign n15410 = n383 & ~n15409 ;
  assign n15411 = n387 & ~n15410 ;
  assign n15412 = n391 & ~n15411 ;
  assign n15413 = n395 & ~n15412 ;
  assign n15414 = n399 & ~n15413 ;
  assign n15415 = n403 & ~n15414 ;
  assign n15416 = n407 & ~n15415 ;
  assign n15417 = n411 & ~n15416 ;
  assign n15418 = n415 & ~n15417 ;
  assign n15419 = n419 & ~n15418 ;
  assign n15420 = n423 & ~n15419 ;
  assign n15421 = n427 & ~n15420 ;
  assign n15422 = n431 & ~n15421 ;
  assign n15423 = n435 & ~n15422 ;
  assign n15424 = n439 & ~n15423 ;
  assign n15425 = n443 & ~n15424 ;
  assign n15426 = n447 & ~n15425 ;
  assign n15427 = n451 & ~n15426 ;
  assign n15428 = n455 & ~n15427 ;
  assign n15429 = x205 & ~n457 ;
  assign n15430 = ~n15428 & n15429 ;
  assign n15518 = n15430 & x333 ;
  assign n15431 = ~n801 & n2157 ;
  assign n15432 = n2162 & ~n15431 ;
  assign n15433 = n2166 & ~n15432 ;
  assign n15434 = n2170 & ~n15433 ;
  assign n15435 = n2174 & ~n15434 ;
  assign n15436 = n2178 & ~n15435 ;
  assign n15437 = n2182 & ~n15436 ;
  assign n15438 = n2186 & ~n15437 ;
  assign n15439 = n2190 & ~n15438 ;
  assign n15440 = n2194 & ~n15439 ;
  assign n15441 = n2198 & ~n15440 ;
  assign n15442 = n2202 & ~n15441 ;
  assign n15443 = n2206 & ~n15442 ;
  assign n15444 = n2210 & ~n15443 ;
  assign n15445 = n2214 & ~n15444 ;
  assign n15446 = n2218 & ~n15445 ;
  assign n15447 = n2222 & ~n15446 ;
  assign n15448 = n2226 & ~n15447 ;
  assign n15449 = n2230 & ~n15448 ;
  assign n15450 = n2234 & ~n15449 ;
  assign n15451 = n2238 & ~n15450 ;
  assign n15452 = n2242 & ~n15451 ;
  assign n15453 = n2246 & ~n15452 ;
  assign n15454 = n2250 & ~n15453 ;
  assign n15455 = n2254 & ~n15454 ;
  assign n15456 = n2258 & ~n15455 ;
  assign n15457 = n2262 & ~n15456 ;
  assign n15458 = n2266 & ~n15457 ;
  assign n15459 = n2270 & ~n15458 ;
  assign n15460 = n2274 & ~n15459 ;
  assign n15461 = n2278 & ~n15460 ;
  assign n15462 = n2282 & ~n15461 ;
  assign n15463 = n2286 & ~n15462 ;
  assign n15464 = n2290 & ~n15463 ;
  assign n15465 = n2836 & ~n15464 ;
  assign n15466 = n602 & ~n15465 ;
  assign n15467 = n606 & ~n15466 ;
  assign n15468 = n610 & ~n15467 ;
  assign n15469 = n614 & ~n15468 ;
  assign n15470 = n618 & ~n15469 ;
  assign n15471 = n622 & ~n15470 ;
  assign n15472 = n626 & ~n15471 ;
  assign n15473 = n630 & ~n15472 ;
  assign n15474 = n634 & ~n15473 ;
  assign n15475 = n638 & ~n15474 ;
  assign n15476 = n642 & ~n15475 ;
  assign n15477 = n646 & ~n15476 ;
  assign n15478 = n650 & ~n15477 ;
  assign n15479 = n654 & ~n15478 ;
  assign n15480 = n658 & ~n15479 ;
  assign n15481 = n662 & ~n15480 ;
  assign n15482 = n666 & ~n15481 ;
  assign n15483 = n670 & ~n15482 ;
  assign n15484 = n674 & ~n15483 ;
  assign n15485 = n678 & ~n15484 ;
  assign n15486 = n682 & ~n15485 ;
  assign n15487 = n686 & ~n15486 ;
  assign n15488 = n690 & ~n15487 ;
  assign n15489 = n694 & ~n15488 ;
  assign n15490 = n698 & ~n15489 ;
  assign n15491 = n702 & ~n15490 ;
  assign n15492 = n706 & ~n15491 ;
  assign n15493 = n710 & ~n15492 ;
  assign n15494 = n714 & ~n15493 ;
  assign n15495 = n718 & ~n15494 ;
  assign n15496 = n722 & ~n15495 ;
  assign n15497 = n726 & ~n15496 ;
  assign n15498 = n730 & ~n15497 ;
  assign n15499 = n734 & ~n15498 ;
  assign n15500 = n738 & ~n15499 ;
  assign n15501 = n742 & ~n15500 ;
  assign n15502 = n746 & ~n15501 ;
  assign n15503 = n750 & ~n15502 ;
  assign n15504 = n754 & ~n15503 ;
  assign n15505 = n758 & ~n15504 ;
  assign n15506 = n762 & ~n15505 ;
  assign n15507 = n766 & ~n15506 ;
  assign n15508 = n770 & ~n15507 ;
  assign n15509 = n774 & ~n15508 ;
  assign n15510 = n778 & ~n15509 ;
  assign n15511 = n782 & ~n15510 ;
  assign n15512 = n786 & ~n15511 ;
  assign n15513 = n790 & ~n15512 ;
  assign n15514 = n794 & ~n15513 ;
  assign n15515 = ~x205 & ~n796 ;
  assign n15516 = ~n15514 & n15515 ;
  assign n15519 = ~n15516 & ~x333 ;
  assign n15520 = ~n15518 & ~n15519 ;
  assign n15521 = n466 & ~n1144 ;
  assign n15522 = n471 & ~n15521 ;
  assign n15523 = n475 & ~n15522 ;
  assign n15524 = n479 & ~n15523 ;
  assign n15525 = n483 & ~n15524 ;
  assign n15526 = n487 & ~n15525 ;
  assign n15527 = n491 & ~n15526 ;
  assign n15528 = n495 & ~n15527 ;
  assign n15529 = n499 & ~n15528 ;
  assign n15530 = n503 & ~n15529 ;
  assign n15531 = n507 & ~n15530 ;
  assign n15532 = n511 & ~n15531 ;
  assign n15533 = n515 & ~n15532 ;
  assign n15534 = n519 & ~n15533 ;
  assign n15535 = n523 & ~n15534 ;
  assign n15536 = n527 & ~n15535 ;
  assign n15537 = n531 & ~n15536 ;
  assign n15538 = n535 & ~n15537 ;
  assign n15539 = n539 & ~n15538 ;
  assign n15540 = n543 & ~n15539 ;
  assign n15541 = n547 & ~n15540 ;
  assign n15542 = n551 & ~n15541 ;
  assign n15543 = n555 & ~n15542 ;
  assign n15544 = n559 & ~n15543 ;
  assign n15545 = n563 & ~n15544 ;
  assign n15546 = n567 & ~n15545 ;
  assign n15547 = n571 & ~n15546 ;
  assign n15548 = n575 & ~n15547 ;
  assign n15549 = n579 & ~n15548 ;
  assign n15550 = n583 & ~n15549 ;
  assign n15551 = n587 & ~n15550 ;
  assign n15552 = n591 & ~n15551 ;
  assign n15553 = n2382 & ~n15552 ;
  assign n15554 = n2384 & ~n15553 ;
  assign n15555 = n2927 & ~n15554 ;
  assign n15556 = n945 & ~n15555 ;
  assign n15557 = n949 & ~n15556 ;
  assign n15558 = n953 & ~n15557 ;
  assign n15559 = n957 & ~n15558 ;
  assign n15560 = n961 & ~n15559 ;
  assign n15561 = n965 & ~n15560 ;
  assign n15562 = n969 & ~n15561 ;
  assign n15563 = n973 & ~n15562 ;
  assign n15564 = n977 & ~n15563 ;
  assign n15565 = n981 & ~n15564 ;
  assign n15566 = n985 & ~n15565 ;
  assign n15567 = n989 & ~n15566 ;
  assign n15568 = n993 & ~n15567 ;
  assign n15569 = n997 & ~n15568 ;
  assign n15570 = n1001 & ~n15569 ;
  assign n15571 = n1005 & ~n15570 ;
  assign n15572 = n1009 & ~n15571 ;
  assign n15573 = n1013 & ~n15572 ;
  assign n15574 = n1017 & ~n15573 ;
  assign n15575 = n1021 & ~n15574 ;
  assign n15576 = n1025 & ~n15575 ;
  assign n15577 = n1029 & ~n15576 ;
  assign n15578 = n1033 & ~n15577 ;
  assign n15579 = n1037 & ~n15578 ;
  assign n15580 = n1041 & ~n15579 ;
  assign n15581 = n1045 & ~n15580 ;
  assign n15582 = n1049 & ~n15581 ;
  assign n15583 = n1053 & ~n15582 ;
  assign n15584 = n1057 & ~n15583 ;
  assign n15585 = n1061 & ~n15584 ;
  assign n15586 = n1065 & ~n15585 ;
  assign n15587 = n1069 & ~n15586 ;
  assign n15588 = n1073 & ~n15587 ;
  assign n15589 = n1077 & ~n15588 ;
  assign n15590 = n1081 & ~n15589 ;
  assign n15591 = n1085 & ~n15590 ;
  assign n15592 = n1089 & ~n15591 ;
  assign n15593 = n1093 & ~n15592 ;
  assign n15594 = n1097 & ~n15593 ;
  assign n15595 = n1101 & ~n15594 ;
  assign n15596 = n1105 & ~n15595 ;
  assign n15597 = n1109 & ~n15596 ;
  assign n15598 = n1113 & ~n15597 ;
  assign n15599 = n1117 & ~n15598 ;
  assign n15600 = n1121 & ~n15599 ;
  assign n15601 = n1125 & ~n15600 ;
  assign n15602 = n1129 & ~n15601 ;
  assign n15603 = n1133 & ~n15602 ;
  assign n15604 = n1137 & ~n15603 ;
  assign n15605 = x206 & ~n1139 ;
  assign n15606 = ~n15604 & n15605 ;
  assign n15694 = n15606 & x334 ;
  assign n15607 = n805 & ~n1483 ;
  assign n15608 = n810 & ~n15607 ;
  assign n15609 = n814 & ~n15608 ;
  assign n15610 = n818 & ~n15609 ;
  assign n15611 = n822 & ~n15610 ;
  assign n15612 = n826 & ~n15611 ;
  assign n15613 = n830 & ~n15612 ;
  assign n15614 = n834 & ~n15613 ;
  assign n15615 = n838 & ~n15614 ;
  assign n15616 = n842 & ~n15615 ;
  assign n15617 = n846 & ~n15616 ;
  assign n15618 = n850 & ~n15617 ;
  assign n15619 = n854 & ~n15618 ;
  assign n15620 = n858 & ~n15619 ;
  assign n15621 = n862 & ~n15620 ;
  assign n15622 = n866 & ~n15621 ;
  assign n15623 = n870 & ~n15622 ;
  assign n15624 = n874 & ~n15623 ;
  assign n15625 = n878 & ~n15624 ;
  assign n15626 = n882 & ~n15625 ;
  assign n15627 = n886 & ~n15626 ;
  assign n15628 = n890 & ~n15627 ;
  assign n15629 = n894 & ~n15628 ;
  assign n15630 = n898 & ~n15629 ;
  assign n15631 = n902 & ~n15630 ;
  assign n15632 = n906 & ~n15631 ;
  assign n15633 = n910 & ~n15632 ;
  assign n15634 = n914 & ~n15633 ;
  assign n15635 = n918 & ~n15634 ;
  assign n15636 = n922 & ~n15635 ;
  assign n15637 = n926 & ~n15636 ;
  assign n15638 = n930 & ~n15637 ;
  assign n15639 = n2472 & ~n15638 ;
  assign n15640 = n2474 & ~n15639 ;
  assign n15641 = n3014 & ~n15640 ;
  assign n15642 = n1284 & ~n15641 ;
  assign n15643 = n1288 & ~n15642 ;
  assign n15644 = n1292 & ~n15643 ;
  assign n15645 = n1296 & ~n15644 ;
  assign n15646 = n1300 & ~n15645 ;
  assign n15647 = n1304 & ~n15646 ;
  assign n15648 = n1308 & ~n15647 ;
  assign n15649 = n1312 & ~n15648 ;
  assign n15650 = n1316 & ~n15649 ;
  assign n15651 = n1320 & ~n15650 ;
  assign n15652 = n1324 & ~n15651 ;
  assign n15653 = n1328 & ~n15652 ;
  assign n15654 = n1332 & ~n15653 ;
  assign n15655 = n1336 & ~n15654 ;
  assign n15656 = n1340 & ~n15655 ;
  assign n15657 = n1344 & ~n15656 ;
  assign n15658 = n1348 & ~n15657 ;
  assign n15659 = n1352 & ~n15658 ;
  assign n15660 = n1356 & ~n15659 ;
  assign n15661 = n1360 & ~n15660 ;
  assign n15662 = n1364 & ~n15661 ;
  assign n15663 = n1368 & ~n15662 ;
  assign n15664 = n1372 & ~n15663 ;
  assign n15665 = n1376 & ~n15664 ;
  assign n15666 = n1380 & ~n15665 ;
  assign n15667 = n1384 & ~n15666 ;
  assign n15668 = n1388 & ~n15667 ;
  assign n15669 = n1392 & ~n15668 ;
  assign n15670 = n1396 & ~n15669 ;
  assign n15671 = n1400 & ~n15670 ;
  assign n15672 = n1404 & ~n15671 ;
  assign n15673 = n1408 & ~n15672 ;
  assign n15674 = n1412 & ~n15673 ;
  assign n15675 = n1416 & ~n15674 ;
  assign n15676 = n1420 & ~n15675 ;
  assign n15677 = n1424 & ~n15676 ;
  assign n15678 = n1428 & ~n15677 ;
  assign n15679 = n1432 & ~n15678 ;
  assign n15680 = n1436 & ~n15679 ;
  assign n15681 = n1440 & ~n15680 ;
  assign n15682 = n1444 & ~n15681 ;
  assign n15683 = n1448 & ~n15682 ;
  assign n15684 = n1452 & ~n15683 ;
  assign n15685 = n1456 & ~n15684 ;
  assign n15686 = n1460 & ~n15685 ;
  assign n15687 = n1464 & ~n15686 ;
  assign n15688 = n1468 & ~n15687 ;
  assign n15689 = n1472 & ~n15688 ;
  assign n15690 = n1476 & ~n15689 ;
  assign n15691 = ~x206 & ~n1478 ;
  assign n15692 = ~n15690 & n15691 ;
  assign n15695 = ~n15692 & ~x334 ;
  assign n15696 = ~n15694 & ~n15695 ;
  assign n15697 = n1148 & ~n1824 ;
  assign n15698 = n1153 & ~n15697 ;
  assign n15699 = n1157 & ~n15698 ;
  assign n15700 = n1161 & ~n15699 ;
  assign n15701 = n1165 & ~n15700 ;
  assign n15702 = n1169 & ~n15701 ;
  assign n15703 = n1173 & ~n15702 ;
  assign n15704 = n1177 & ~n15703 ;
  assign n15705 = n1181 & ~n15704 ;
  assign n15706 = n1185 & ~n15705 ;
  assign n15707 = n1189 & ~n15706 ;
  assign n15708 = n1193 & ~n15707 ;
  assign n15709 = n1197 & ~n15708 ;
  assign n15710 = n1201 & ~n15709 ;
  assign n15711 = n1205 & ~n15710 ;
  assign n15712 = n1209 & ~n15711 ;
  assign n15713 = n1213 & ~n15712 ;
  assign n15714 = n1217 & ~n15713 ;
  assign n15715 = n1221 & ~n15714 ;
  assign n15716 = n1225 & ~n15715 ;
  assign n15717 = n1229 & ~n15716 ;
  assign n15718 = n1233 & ~n15717 ;
  assign n15719 = n1237 & ~n15718 ;
  assign n15720 = n1241 & ~n15719 ;
  assign n15721 = n1245 & ~n15720 ;
  assign n15722 = n1249 & ~n15721 ;
  assign n15723 = n1253 & ~n15722 ;
  assign n15724 = n1257 & ~n15723 ;
  assign n15725 = n1261 & ~n15724 ;
  assign n15726 = n1265 & ~n15725 ;
  assign n15727 = n1269 & ~n15726 ;
  assign n15728 = n1273 & ~n15727 ;
  assign n15729 = n2566 & ~n15728 ;
  assign n15730 = n2568 & ~n15729 ;
  assign n15731 = n3105 & ~n15730 ;
  assign n15732 = n1625 & ~n15731 ;
  assign n15733 = n1629 & ~n15732 ;
  assign n15734 = n1633 & ~n15733 ;
  assign n15735 = n1637 & ~n15734 ;
  assign n15736 = n1641 & ~n15735 ;
  assign n15737 = n1645 & ~n15736 ;
  assign n15738 = n1649 & ~n15737 ;
  assign n15739 = n1653 & ~n15738 ;
  assign n15740 = n1657 & ~n15739 ;
  assign n15741 = n1661 & ~n15740 ;
  assign n15742 = n1665 & ~n15741 ;
  assign n15743 = n1669 & ~n15742 ;
  assign n15744 = n1673 & ~n15743 ;
  assign n15745 = n1677 & ~n15744 ;
  assign n15746 = n1681 & ~n15745 ;
  assign n15747 = n1685 & ~n15746 ;
  assign n15748 = n1689 & ~n15747 ;
  assign n15749 = n1693 & ~n15748 ;
  assign n15750 = n1697 & ~n15749 ;
  assign n15751 = n1701 & ~n15750 ;
  assign n15752 = n1705 & ~n15751 ;
  assign n15753 = n1709 & ~n15752 ;
  assign n15754 = n1713 & ~n15753 ;
  assign n15755 = n1717 & ~n15754 ;
  assign n15756 = n1721 & ~n15755 ;
  assign n15757 = n1725 & ~n15756 ;
  assign n15758 = n1729 & ~n15757 ;
  assign n15759 = n1733 & ~n15758 ;
  assign n15760 = n1737 & ~n15759 ;
  assign n15761 = n1741 & ~n15760 ;
  assign n15762 = n1745 & ~n15761 ;
  assign n15763 = n1749 & ~n15762 ;
  assign n15764 = n1753 & ~n15763 ;
  assign n15765 = n1757 & ~n15764 ;
  assign n15766 = n1761 & ~n15765 ;
  assign n15767 = n1765 & ~n15766 ;
  assign n15768 = n1769 & ~n15767 ;
  assign n15769 = n1773 & ~n15768 ;
  assign n15770 = n1777 & ~n15769 ;
  assign n15771 = n1781 & ~n15770 ;
  assign n15772 = n1785 & ~n15771 ;
  assign n15773 = n1789 & ~n15772 ;
  assign n15774 = n1793 & ~n15773 ;
  assign n15775 = n1797 & ~n15774 ;
  assign n15776 = n1801 & ~n15775 ;
  assign n15777 = n1805 & ~n15776 ;
  assign n15778 = n1809 & ~n15777 ;
  assign n15779 = n1813 & ~n15778 ;
  assign n15780 = n1817 & ~n15779 ;
  assign n15781 = x207 & ~n1819 ;
  assign n15782 = ~n15780 & n15781 ;
  assign n15870 = n15782 & x335 ;
  assign n15783 = n1487 & ~n2161 ;
  assign n15784 = n1492 & ~n15783 ;
  assign n15785 = n1496 & ~n15784 ;
  assign n15786 = n1500 & ~n15785 ;
  assign n15787 = n1504 & ~n15786 ;
  assign n15788 = n1508 & ~n15787 ;
  assign n15789 = n1512 & ~n15788 ;
  assign n15790 = n1516 & ~n15789 ;
  assign n15791 = n1520 & ~n15790 ;
  assign n15792 = n1524 & ~n15791 ;
  assign n15793 = n1528 & ~n15792 ;
  assign n15794 = n1532 & ~n15793 ;
  assign n15795 = n1536 & ~n15794 ;
  assign n15796 = n1540 & ~n15795 ;
  assign n15797 = n1544 & ~n15796 ;
  assign n15798 = n1548 & ~n15797 ;
  assign n15799 = n1552 & ~n15798 ;
  assign n15800 = n1556 & ~n15799 ;
  assign n15801 = n1560 & ~n15800 ;
  assign n15802 = n1564 & ~n15801 ;
  assign n15803 = n1568 & ~n15802 ;
  assign n15804 = n1572 & ~n15803 ;
  assign n15805 = n1576 & ~n15804 ;
  assign n15806 = n1580 & ~n15805 ;
  assign n15807 = n1584 & ~n15806 ;
  assign n15808 = n1588 & ~n15807 ;
  assign n15809 = n1592 & ~n15808 ;
  assign n15810 = n1596 & ~n15809 ;
  assign n15811 = n1600 & ~n15810 ;
  assign n15812 = n1604 & ~n15811 ;
  assign n15813 = n1608 & ~n15812 ;
  assign n15814 = n1612 & ~n15813 ;
  assign n15815 = n2656 & ~n15814 ;
  assign n15816 = n2658 & ~n15815 ;
  assign n15817 = n3192 & ~n15816 ;
  assign n15818 = n1962 & ~n15817 ;
  assign n15819 = n1966 & ~n15818 ;
  assign n15820 = n1970 & ~n15819 ;
  assign n15821 = n1974 & ~n15820 ;
  assign n15822 = n1978 & ~n15821 ;
  assign n15823 = n1982 & ~n15822 ;
  assign n15824 = n1986 & ~n15823 ;
  assign n15825 = n1990 & ~n15824 ;
  assign n15826 = n1994 & ~n15825 ;
  assign n15827 = n1998 & ~n15826 ;
  assign n15828 = n2002 & ~n15827 ;
  assign n15829 = n2006 & ~n15828 ;
  assign n15830 = n2010 & ~n15829 ;
  assign n15831 = n2014 & ~n15830 ;
  assign n15832 = n2018 & ~n15831 ;
  assign n15833 = n2022 & ~n15832 ;
  assign n15834 = n2026 & ~n15833 ;
  assign n15835 = n2030 & ~n15834 ;
  assign n15836 = n2034 & ~n15835 ;
  assign n15837 = n2038 & ~n15836 ;
  assign n15838 = n2042 & ~n15837 ;
  assign n15839 = n2046 & ~n15838 ;
  assign n15840 = n2050 & ~n15839 ;
  assign n15841 = n2054 & ~n15840 ;
  assign n15842 = n2058 & ~n15841 ;
  assign n15843 = n2062 & ~n15842 ;
  assign n15844 = n2066 & ~n15843 ;
  assign n15845 = n2070 & ~n15844 ;
  assign n15846 = n2074 & ~n15845 ;
  assign n15847 = n2078 & ~n15846 ;
  assign n15848 = n2082 & ~n15847 ;
  assign n15849 = n2086 & ~n15848 ;
  assign n15850 = n2090 & ~n15849 ;
  assign n15851 = n2094 & ~n15850 ;
  assign n15852 = n2098 & ~n15851 ;
  assign n15853 = n2102 & ~n15852 ;
  assign n15854 = n2106 & ~n15853 ;
  assign n15855 = n2110 & ~n15854 ;
  assign n15856 = n2114 & ~n15855 ;
  assign n15857 = n2118 & ~n15856 ;
  assign n15858 = n2122 & ~n15857 ;
  assign n15859 = n2126 & ~n15858 ;
  assign n15860 = n2130 & ~n15859 ;
  assign n15861 = n2134 & ~n15860 ;
  assign n15862 = n2138 & ~n15861 ;
  assign n15863 = n2142 & ~n15862 ;
  assign n15864 = n2146 & ~n15863 ;
  assign n15865 = n2150 & ~n15864 ;
  assign n15866 = n2154 & ~n15865 ;
  assign n15867 = ~x207 & ~n2156 ;
  assign n15868 = ~n15866 & n15867 ;
  assign n15871 = ~n15868 & ~x335 ;
  assign n15872 = ~n15870 & ~n15871 ;
  assign n15873 = ~n470 & n1828 ;
  assign n15874 = n1833 & ~n15873 ;
  assign n15875 = n1837 & ~n15874 ;
  assign n15876 = n1841 & ~n15875 ;
  assign n15877 = n1845 & ~n15876 ;
  assign n15878 = n1849 & ~n15877 ;
  assign n15879 = n1853 & ~n15878 ;
  assign n15880 = n1857 & ~n15879 ;
  assign n15881 = n1861 & ~n15880 ;
  assign n15882 = n1865 & ~n15881 ;
  assign n15883 = n1869 & ~n15882 ;
  assign n15884 = n1873 & ~n15883 ;
  assign n15885 = n1877 & ~n15884 ;
  assign n15886 = n1881 & ~n15885 ;
  assign n15887 = n1885 & ~n15886 ;
  assign n15888 = n1889 & ~n15887 ;
  assign n15889 = n1893 & ~n15888 ;
  assign n15890 = n1897 & ~n15889 ;
  assign n15891 = n1901 & ~n15890 ;
  assign n15892 = n1905 & ~n15891 ;
  assign n15893 = n1909 & ~n15892 ;
  assign n15894 = n1913 & ~n15893 ;
  assign n15895 = n1917 & ~n15894 ;
  assign n15896 = n1921 & ~n15895 ;
  assign n15897 = n1925 & ~n15896 ;
  assign n15898 = n1929 & ~n15897 ;
  assign n15899 = n1933 & ~n15898 ;
  assign n15900 = n1937 & ~n15899 ;
  assign n15901 = n1941 & ~n15900 ;
  assign n15902 = n1945 & ~n15901 ;
  assign n15903 = n1949 & ~n15902 ;
  assign n15904 = n1953 & ~n15903 ;
  assign n15905 = n2749 & ~n15904 ;
  assign n15906 = n263 & ~n15905 ;
  assign n15907 = n267 & ~n15906 ;
  assign n15908 = n271 & ~n15907 ;
  assign n15909 = n275 & ~n15908 ;
  assign n15910 = n279 & ~n15909 ;
  assign n15911 = n283 & ~n15910 ;
  assign n15912 = n287 & ~n15911 ;
  assign n15913 = n291 & ~n15912 ;
  assign n15914 = n295 & ~n15913 ;
  assign n15915 = n299 & ~n15914 ;
  assign n15916 = n303 & ~n15915 ;
  assign n15917 = n307 & ~n15916 ;
  assign n15918 = n311 & ~n15917 ;
  assign n15919 = n315 & ~n15918 ;
  assign n15920 = n319 & ~n15919 ;
  assign n15921 = n323 & ~n15920 ;
  assign n15922 = n327 & ~n15921 ;
  assign n15923 = n331 & ~n15922 ;
  assign n15924 = n335 & ~n15923 ;
  assign n15925 = n339 & ~n15924 ;
  assign n15926 = n343 & ~n15925 ;
  assign n15927 = n347 & ~n15926 ;
  assign n15928 = n351 & ~n15927 ;
  assign n15929 = n355 & ~n15928 ;
  assign n15930 = n359 & ~n15929 ;
  assign n15931 = n363 & ~n15930 ;
  assign n15932 = n367 & ~n15931 ;
  assign n15933 = n371 & ~n15932 ;
  assign n15934 = n375 & ~n15933 ;
  assign n15935 = n379 & ~n15934 ;
  assign n15936 = n383 & ~n15935 ;
  assign n15937 = n387 & ~n15936 ;
  assign n15938 = n391 & ~n15937 ;
  assign n15939 = n395 & ~n15938 ;
  assign n15940 = n399 & ~n15939 ;
  assign n15941 = n403 & ~n15940 ;
  assign n15942 = n407 & ~n15941 ;
  assign n15943 = n411 & ~n15942 ;
  assign n15944 = n415 & ~n15943 ;
  assign n15945 = n419 & ~n15944 ;
  assign n15946 = n423 & ~n15945 ;
  assign n15947 = n427 & ~n15946 ;
  assign n15948 = n431 & ~n15947 ;
  assign n15949 = n435 & ~n15948 ;
  assign n15950 = n439 & ~n15949 ;
  assign n15951 = n443 & ~n15950 ;
  assign n15952 = n447 & ~n15951 ;
  assign n15953 = n451 & ~n15952 ;
  assign n15954 = n455 & ~n15953 ;
  assign n15955 = n459 & ~n15954 ;
  assign n15956 = n463 & ~n15955 ;
  assign n15957 = x208 & ~n465 ;
  assign n15958 = ~n15956 & n15957 ;
  assign n16046 = n15958 & x336 ;
  assign n15959 = ~n809 & n2165 ;
  assign n15960 = n2170 & ~n15959 ;
  assign n15961 = n2174 & ~n15960 ;
  assign n15962 = n2178 & ~n15961 ;
  assign n15963 = n2182 & ~n15962 ;
  assign n15964 = n2186 & ~n15963 ;
  assign n15965 = n2190 & ~n15964 ;
  assign n15966 = n2194 & ~n15965 ;
  assign n15967 = n2198 & ~n15966 ;
  assign n15968 = n2202 & ~n15967 ;
  assign n15969 = n2206 & ~n15968 ;
  assign n15970 = n2210 & ~n15969 ;
  assign n15971 = n2214 & ~n15970 ;
  assign n15972 = n2218 & ~n15971 ;
  assign n15973 = n2222 & ~n15972 ;
  assign n15974 = n2226 & ~n15973 ;
  assign n15975 = n2230 & ~n15974 ;
  assign n15976 = n2234 & ~n15975 ;
  assign n15977 = n2238 & ~n15976 ;
  assign n15978 = n2242 & ~n15977 ;
  assign n15979 = n2246 & ~n15978 ;
  assign n15980 = n2250 & ~n15979 ;
  assign n15981 = n2254 & ~n15980 ;
  assign n15982 = n2258 & ~n15981 ;
  assign n15983 = n2262 & ~n15982 ;
  assign n15984 = n2266 & ~n15983 ;
  assign n15985 = n2270 & ~n15984 ;
  assign n15986 = n2274 & ~n15985 ;
  assign n15987 = n2278 & ~n15986 ;
  assign n15988 = n2282 & ~n15987 ;
  assign n15989 = n2286 & ~n15988 ;
  assign n15990 = n2290 & ~n15989 ;
  assign n15991 = n2836 & ~n15990 ;
  assign n15992 = n602 & ~n15991 ;
  assign n15993 = n606 & ~n15992 ;
  assign n15994 = n610 & ~n15993 ;
  assign n15995 = n614 & ~n15994 ;
  assign n15996 = n618 & ~n15995 ;
  assign n15997 = n622 & ~n15996 ;
  assign n15998 = n626 & ~n15997 ;
  assign n15999 = n630 & ~n15998 ;
  assign n16000 = n634 & ~n15999 ;
  assign n16001 = n638 & ~n16000 ;
  assign n16002 = n642 & ~n16001 ;
  assign n16003 = n646 & ~n16002 ;
  assign n16004 = n650 & ~n16003 ;
  assign n16005 = n654 & ~n16004 ;
  assign n16006 = n658 & ~n16005 ;
  assign n16007 = n662 & ~n16006 ;
  assign n16008 = n666 & ~n16007 ;
  assign n16009 = n670 & ~n16008 ;
  assign n16010 = n674 & ~n16009 ;
  assign n16011 = n678 & ~n16010 ;
  assign n16012 = n682 & ~n16011 ;
  assign n16013 = n686 & ~n16012 ;
  assign n16014 = n690 & ~n16013 ;
  assign n16015 = n694 & ~n16014 ;
  assign n16016 = n698 & ~n16015 ;
  assign n16017 = n702 & ~n16016 ;
  assign n16018 = n706 & ~n16017 ;
  assign n16019 = n710 & ~n16018 ;
  assign n16020 = n714 & ~n16019 ;
  assign n16021 = n718 & ~n16020 ;
  assign n16022 = n722 & ~n16021 ;
  assign n16023 = n726 & ~n16022 ;
  assign n16024 = n730 & ~n16023 ;
  assign n16025 = n734 & ~n16024 ;
  assign n16026 = n738 & ~n16025 ;
  assign n16027 = n742 & ~n16026 ;
  assign n16028 = n746 & ~n16027 ;
  assign n16029 = n750 & ~n16028 ;
  assign n16030 = n754 & ~n16029 ;
  assign n16031 = n758 & ~n16030 ;
  assign n16032 = n762 & ~n16031 ;
  assign n16033 = n766 & ~n16032 ;
  assign n16034 = n770 & ~n16033 ;
  assign n16035 = n774 & ~n16034 ;
  assign n16036 = n778 & ~n16035 ;
  assign n16037 = n782 & ~n16036 ;
  assign n16038 = n786 & ~n16037 ;
  assign n16039 = n790 & ~n16038 ;
  assign n16040 = n794 & ~n16039 ;
  assign n16041 = n798 & ~n16040 ;
  assign n16042 = n802 & ~n16041 ;
  assign n16043 = ~x208 & ~n804 ;
  assign n16044 = ~n16042 & n16043 ;
  assign n16047 = ~n16044 & ~x336 ;
  assign n16048 = ~n16046 & ~n16047 ;
  assign n16049 = n474 & ~n1152 ;
  assign n16050 = n479 & ~n16049 ;
  assign n16051 = n483 & ~n16050 ;
  assign n16052 = n487 & ~n16051 ;
  assign n16053 = n491 & ~n16052 ;
  assign n16054 = n495 & ~n16053 ;
  assign n16055 = n499 & ~n16054 ;
  assign n16056 = n503 & ~n16055 ;
  assign n16057 = n507 & ~n16056 ;
  assign n16058 = n511 & ~n16057 ;
  assign n16059 = n515 & ~n16058 ;
  assign n16060 = n519 & ~n16059 ;
  assign n16061 = n523 & ~n16060 ;
  assign n16062 = n527 & ~n16061 ;
  assign n16063 = n531 & ~n16062 ;
  assign n16064 = n535 & ~n16063 ;
  assign n16065 = n539 & ~n16064 ;
  assign n16066 = n543 & ~n16065 ;
  assign n16067 = n547 & ~n16066 ;
  assign n16068 = n551 & ~n16067 ;
  assign n16069 = n555 & ~n16068 ;
  assign n16070 = n559 & ~n16069 ;
  assign n16071 = n563 & ~n16070 ;
  assign n16072 = n567 & ~n16071 ;
  assign n16073 = n571 & ~n16072 ;
  assign n16074 = n575 & ~n16073 ;
  assign n16075 = n579 & ~n16074 ;
  assign n16076 = n583 & ~n16075 ;
  assign n16077 = n587 & ~n16076 ;
  assign n16078 = n591 & ~n16077 ;
  assign n16079 = n2382 & ~n16078 ;
  assign n16080 = n2384 & ~n16079 ;
  assign n16081 = n2927 & ~n16080 ;
  assign n16082 = n945 & ~n16081 ;
  assign n16083 = n949 & ~n16082 ;
  assign n16084 = n953 & ~n16083 ;
  assign n16085 = n957 & ~n16084 ;
  assign n16086 = n961 & ~n16085 ;
  assign n16087 = n965 & ~n16086 ;
  assign n16088 = n969 & ~n16087 ;
  assign n16089 = n973 & ~n16088 ;
  assign n16090 = n977 & ~n16089 ;
  assign n16091 = n981 & ~n16090 ;
  assign n16092 = n985 & ~n16091 ;
  assign n16093 = n989 & ~n16092 ;
  assign n16094 = n993 & ~n16093 ;
  assign n16095 = n997 & ~n16094 ;
  assign n16096 = n1001 & ~n16095 ;
  assign n16097 = n1005 & ~n16096 ;
  assign n16098 = n1009 & ~n16097 ;
  assign n16099 = n1013 & ~n16098 ;
  assign n16100 = n1017 & ~n16099 ;
  assign n16101 = n1021 & ~n16100 ;
  assign n16102 = n1025 & ~n16101 ;
  assign n16103 = n1029 & ~n16102 ;
  assign n16104 = n1033 & ~n16103 ;
  assign n16105 = n1037 & ~n16104 ;
  assign n16106 = n1041 & ~n16105 ;
  assign n16107 = n1045 & ~n16106 ;
  assign n16108 = n1049 & ~n16107 ;
  assign n16109 = n1053 & ~n16108 ;
  assign n16110 = n1057 & ~n16109 ;
  assign n16111 = n1061 & ~n16110 ;
  assign n16112 = n1065 & ~n16111 ;
  assign n16113 = n1069 & ~n16112 ;
  assign n16114 = n1073 & ~n16113 ;
  assign n16115 = n1077 & ~n16114 ;
  assign n16116 = n1081 & ~n16115 ;
  assign n16117 = n1085 & ~n16116 ;
  assign n16118 = n1089 & ~n16117 ;
  assign n16119 = n1093 & ~n16118 ;
  assign n16120 = n1097 & ~n16119 ;
  assign n16121 = n1101 & ~n16120 ;
  assign n16122 = n1105 & ~n16121 ;
  assign n16123 = n1109 & ~n16122 ;
  assign n16124 = n1113 & ~n16123 ;
  assign n16125 = n1117 & ~n16124 ;
  assign n16126 = n1121 & ~n16125 ;
  assign n16127 = n1125 & ~n16126 ;
  assign n16128 = n1129 & ~n16127 ;
  assign n16129 = n1133 & ~n16128 ;
  assign n16130 = n1137 & ~n16129 ;
  assign n16131 = n1141 & ~n16130 ;
  assign n16132 = n1145 & ~n16131 ;
  assign n16133 = x209 & ~n1147 ;
  assign n16134 = ~n16132 & n16133 ;
  assign n16222 = n16134 & x337 ;
  assign n16135 = n813 & ~n1491 ;
  assign n16136 = n818 & ~n16135 ;
  assign n16137 = n822 & ~n16136 ;
  assign n16138 = n826 & ~n16137 ;
  assign n16139 = n830 & ~n16138 ;
  assign n16140 = n834 & ~n16139 ;
  assign n16141 = n838 & ~n16140 ;
  assign n16142 = n842 & ~n16141 ;
  assign n16143 = n846 & ~n16142 ;
  assign n16144 = n850 & ~n16143 ;
  assign n16145 = n854 & ~n16144 ;
  assign n16146 = n858 & ~n16145 ;
  assign n16147 = n862 & ~n16146 ;
  assign n16148 = n866 & ~n16147 ;
  assign n16149 = n870 & ~n16148 ;
  assign n16150 = n874 & ~n16149 ;
  assign n16151 = n878 & ~n16150 ;
  assign n16152 = n882 & ~n16151 ;
  assign n16153 = n886 & ~n16152 ;
  assign n16154 = n890 & ~n16153 ;
  assign n16155 = n894 & ~n16154 ;
  assign n16156 = n898 & ~n16155 ;
  assign n16157 = n902 & ~n16156 ;
  assign n16158 = n906 & ~n16157 ;
  assign n16159 = n910 & ~n16158 ;
  assign n16160 = n914 & ~n16159 ;
  assign n16161 = n918 & ~n16160 ;
  assign n16162 = n922 & ~n16161 ;
  assign n16163 = n926 & ~n16162 ;
  assign n16164 = n930 & ~n16163 ;
  assign n16165 = n2472 & ~n16164 ;
  assign n16166 = n2474 & ~n16165 ;
  assign n16167 = n3014 & ~n16166 ;
  assign n16168 = n1284 & ~n16167 ;
  assign n16169 = n1288 & ~n16168 ;
  assign n16170 = n1292 & ~n16169 ;
  assign n16171 = n1296 & ~n16170 ;
  assign n16172 = n1300 & ~n16171 ;
  assign n16173 = n1304 & ~n16172 ;
  assign n16174 = n1308 & ~n16173 ;
  assign n16175 = n1312 & ~n16174 ;
  assign n16176 = n1316 & ~n16175 ;
  assign n16177 = n1320 & ~n16176 ;
  assign n16178 = n1324 & ~n16177 ;
  assign n16179 = n1328 & ~n16178 ;
  assign n16180 = n1332 & ~n16179 ;
  assign n16181 = n1336 & ~n16180 ;
  assign n16182 = n1340 & ~n16181 ;
  assign n16183 = n1344 & ~n16182 ;
  assign n16184 = n1348 & ~n16183 ;
  assign n16185 = n1352 & ~n16184 ;
  assign n16186 = n1356 & ~n16185 ;
  assign n16187 = n1360 & ~n16186 ;
  assign n16188 = n1364 & ~n16187 ;
  assign n16189 = n1368 & ~n16188 ;
  assign n16190 = n1372 & ~n16189 ;
  assign n16191 = n1376 & ~n16190 ;
  assign n16192 = n1380 & ~n16191 ;
  assign n16193 = n1384 & ~n16192 ;
  assign n16194 = n1388 & ~n16193 ;
  assign n16195 = n1392 & ~n16194 ;
  assign n16196 = n1396 & ~n16195 ;
  assign n16197 = n1400 & ~n16196 ;
  assign n16198 = n1404 & ~n16197 ;
  assign n16199 = n1408 & ~n16198 ;
  assign n16200 = n1412 & ~n16199 ;
  assign n16201 = n1416 & ~n16200 ;
  assign n16202 = n1420 & ~n16201 ;
  assign n16203 = n1424 & ~n16202 ;
  assign n16204 = n1428 & ~n16203 ;
  assign n16205 = n1432 & ~n16204 ;
  assign n16206 = n1436 & ~n16205 ;
  assign n16207 = n1440 & ~n16206 ;
  assign n16208 = n1444 & ~n16207 ;
  assign n16209 = n1448 & ~n16208 ;
  assign n16210 = n1452 & ~n16209 ;
  assign n16211 = n1456 & ~n16210 ;
  assign n16212 = n1460 & ~n16211 ;
  assign n16213 = n1464 & ~n16212 ;
  assign n16214 = n1468 & ~n16213 ;
  assign n16215 = n1472 & ~n16214 ;
  assign n16216 = n1476 & ~n16215 ;
  assign n16217 = n1480 & ~n16216 ;
  assign n16218 = n1484 & ~n16217 ;
  assign n16219 = ~x209 & ~n1486 ;
  assign n16220 = ~n16218 & n16219 ;
  assign n16223 = ~n16220 & ~x337 ;
  assign n16224 = ~n16222 & ~n16223 ;
  assign n16225 = n1156 & ~n1832 ;
  assign n16226 = n1161 & ~n16225 ;
  assign n16227 = n1165 & ~n16226 ;
  assign n16228 = n1169 & ~n16227 ;
  assign n16229 = n1173 & ~n16228 ;
  assign n16230 = n1177 & ~n16229 ;
  assign n16231 = n1181 & ~n16230 ;
  assign n16232 = n1185 & ~n16231 ;
  assign n16233 = n1189 & ~n16232 ;
  assign n16234 = n1193 & ~n16233 ;
  assign n16235 = n1197 & ~n16234 ;
  assign n16236 = n1201 & ~n16235 ;
  assign n16237 = n1205 & ~n16236 ;
  assign n16238 = n1209 & ~n16237 ;
  assign n16239 = n1213 & ~n16238 ;
  assign n16240 = n1217 & ~n16239 ;
  assign n16241 = n1221 & ~n16240 ;
  assign n16242 = n1225 & ~n16241 ;
  assign n16243 = n1229 & ~n16242 ;
  assign n16244 = n1233 & ~n16243 ;
  assign n16245 = n1237 & ~n16244 ;
  assign n16246 = n1241 & ~n16245 ;
  assign n16247 = n1245 & ~n16246 ;
  assign n16248 = n1249 & ~n16247 ;
  assign n16249 = n1253 & ~n16248 ;
  assign n16250 = n1257 & ~n16249 ;
  assign n16251 = n1261 & ~n16250 ;
  assign n16252 = n1265 & ~n16251 ;
  assign n16253 = n1269 & ~n16252 ;
  assign n16254 = n1273 & ~n16253 ;
  assign n16255 = n2566 & ~n16254 ;
  assign n16256 = n2568 & ~n16255 ;
  assign n16257 = n3105 & ~n16256 ;
  assign n16258 = n1625 & ~n16257 ;
  assign n16259 = n1629 & ~n16258 ;
  assign n16260 = n1633 & ~n16259 ;
  assign n16261 = n1637 & ~n16260 ;
  assign n16262 = n1641 & ~n16261 ;
  assign n16263 = n1645 & ~n16262 ;
  assign n16264 = n1649 & ~n16263 ;
  assign n16265 = n1653 & ~n16264 ;
  assign n16266 = n1657 & ~n16265 ;
  assign n16267 = n1661 & ~n16266 ;
  assign n16268 = n1665 & ~n16267 ;
  assign n16269 = n1669 & ~n16268 ;
  assign n16270 = n1673 & ~n16269 ;
  assign n16271 = n1677 & ~n16270 ;
  assign n16272 = n1681 & ~n16271 ;
  assign n16273 = n1685 & ~n16272 ;
  assign n16274 = n1689 & ~n16273 ;
  assign n16275 = n1693 & ~n16274 ;
  assign n16276 = n1697 & ~n16275 ;
  assign n16277 = n1701 & ~n16276 ;
  assign n16278 = n1705 & ~n16277 ;
  assign n16279 = n1709 & ~n16278 ;
  assign n16280 = n1713 & ~n16279 ;
  assign n16281 = n1717 & ~n16280 ;
  assign n16282 = n1721 & ~n16281 ;
  assign n16283 = n1725 & ~n16282 ;
  assign n16284 = n1729 & ~n16283 ;
  assign n16285 = n1733 & ~n16284 ;
  assign n16286 = n1737 & ~n16285 ;
  assign n16287 = n1741 & ~n16286 ;
  assign n16288 = n1745 & ~n16287 ;
  assign n16289 = n1749 & ~n16288 ;
  assign n16290 = n1753 & ~n16289 ;
  assign n16291 = n1757 & ~n16290 ;
  assign n16292 = n1761 & ~n16291 ;
  assign n16293 = n1765 & ~n16292 ;
  assign n16294 = n1769 & ~n16293 ;
  assign n16295 = n1773 & ~n16294 ;
  assign n16296 = n1777 & ~n16295 ;
  assign n16297 = n1781 & ~n16296 ;
  assign n16298 = n1785 & ~n16297 ;
  assign n16299 = n1789 & ~n16298 ;
  assign n16300 = n1793 & ~n16299 ;
  assign n16301 = n1797 & ~n16300 ;
  assign n16302 = n1801 & ~n16301 ;
  assign n16303 = n1805 & ~n16302 ;
  assign n16304 = n1809 & ~n16303 ;
  assign n16305 = n1813 & ~n16304 ;
  assign n16306 = n1817 & ~n16305 ;
  assign n16307 = n1821 & ~n16306 ;
  assign n16308 = n1825 & ~n16307 ;
  assign n16309 = x210 & ~n1827 ;
  assign n16310 = ~n16308 & n16309 ;
  assign n16398 = n16310 & x338 ;
  assign n16311 = n1495 & ~n2169 ;
  assign n16312 = n1500 & ~n16311 ;
  assign n16313 = n1504 & ~n16312 ;
  assign n16314 = n1508 & ~n16313 ;
  assign n16315 = n1512 & ~n16314 ;
  assign n16316 = n1516 & ~n16315 ;
  assign n16317 = n1520 & ~n16316 ;
  assign n16318 = n1524 & ~n16317 ;
  assign n16319 = n1528 & ~n16318 ;
  assign n16320 = n1532 & ~n16319 ;
  assign n16321 = n1536 & ~n16320 ;
  assign n16322 = n1540 & ~n16321 ;
  assign n16323 = n1544 & ~n16322 ;
  assign n16324 = n1548 & ~n16323 ;
  assign n16325 = n1552 & ~n16324 ;
  assign n16326 = n1556 & ~n16325 ;
  assign n16327 = n1560 & ~n16326 ;
  assign n16328 = n1564 & ~n16327 ;
  assign n16329 = n1568 & ~n16328 ;
  assign n16330 = n1572 & ~n16329 ;
  assign n16331 = n1576 & ~n16330 ;
  assign n16332 = n1580 & ~n16331 ;
  assign n16333 = n1584 & ~n16332 ;
  assign n16334 = n1588 & ~n16333 ;
  assign n16335 = n1592 & ~n16334 ;
  assign n16336 = n1596 & ~n16335 ;
  assign n16337 = n1600 & ~n16336 ;
  assign n16338 = n1604 & ~n16337 ;
  assign n16339 = n1608 & ~n16338 ;
  assign n16340 = n1612 & ~n16339 ;
  assign n16341 = n2656 & ~n16340 ;
  assign n16342 = n2658 & ~n16341 ;
  assign n16343 = n3192 & ~n16342 ;
  assign n16344 = n1962 & ~n16343 ;
  assign n16345 = n1966 & ~n16344 ;
  assign n16346 = n1970 & ~n16345 ;
  assign n16347 = n1974 & ~n16346 ;
  assign n16348 = n1978 & ~n16347 ;
  assign n16349 = n1982 & ~n16348 ;
  assign n16350 = n1986 & ~n16349 ;
  assign n16351 = n1990 & ~n16350 ;
  assign n16352 = n1994 & ~n16351 ;
  assign n16353 = n1998 & ~n16352 ;
  assign n16354 = n2002 & ~n16353 ;
  assign n16355 = n2006 & ~n16354 ;
  assign n16356 = n2010 & ~n16355 ;
  assign n16357 = n2014 & ~n16356 ;
  assign n16358 = n2018 & ~n16357 ;
  assign n16359 = n2022 & ~n16358 ;
  assign n16360 = n2026 & ~n16359 ;
  assign n16361 = n2030 & ~n16360 ;
  assign n16362 = n2034 & ~n16361 ;
  assign n16363 = n2038 & ~n16362 ;
  assign n16364 = n2042 & ~n16363 ;
  assign n16365 = n2046 & ~n16364 ;
  assign n16366 = n2050 & ~n16365 ;
  assign n16367 = n2054 & ~n16366 ;
  assign n16368 = n2058 & ~n16367 ;
  assign n16369 = n2062 & ~n16368 ;
  assign n16370 = n2066 & ~n16369 ;
  assign n16371 = n2070 & ~n16370 ;
  assign n16372 = n2074 & ~n16371 ;
  assign n16373 = n2078 & ~n16372 ;
  assign n16374 = n2082 & ~n16373 ;
  assign n16375 = n2086 & ~n16374 ;
  assign n16376 = n2090 & ~n16375 ;
  assign n16377 = n2094 & ~n16376 ;
  assign n16378 = n2098 & ~n16377 ;
  assign n16379 = n2102 & ~n16378 ;
  assign n16380 = n2106 & ~n16379 ;
  assign n16381 = n2110 & ~n16380 ;
  assign n16382 = n2114 & ~n16381 ;
  assign n16383 = n2118 & ~n16382 ;
  assign n16384 = n2122 & ~n16383 ;
  assign n16385 = n2126 & ~n16384 ;
  assign n16386 = n2130 & ~n16385 ;
  assign n16387 = n2134 & ~n16386 ;
  assign n16388 = n2138 & ~n16387 ;
  assign n16389 = n2142 & ~n16388 ;
  assign n16390 = n2146 & ~n16389 ;
  assign n16391 = n2150 & ~n16390 ;
  assign n16392 = n2154 & ~n16391 ;
  assign n16393 = n2158 & ~n16392 ;
  assign n16394 = n2162 & ~n16393 ;
  assign n16395 = ~x210 & ~n2164 ;
  assign n16396 = ~n16394 & n16395 ;
  assign n16399 = ~n16396 & ~x338 ;
  assign n16400 = ~n16398 & ~n16399 ;
  assign n16401 = ~n478 & n1836 ;
  assign n16402 = n1841 & ~n16401 ;
  assign n16403 = n1845 & ~n16402 ;
  assign n16404 = n1849 & ~n16403 ;
  assign n16405 = n1853 & ~n16404 ;
  assign n16406 = n1857 & ~n16405 ;
  assign n16407 = n1861 & ~n16406 ;
  assign n16408 = n1865 & ~n16407 ;
  assign n16409 = n1869 & ~n16408 ;
  assign n16410 = n1873 & ~n16409 ;
  assign n16411 = n1877 & ~n16410 ;
  assign n16412 = n1881 & ~n16411 ;
  assign n16413 = n1885 & ~n16412 ;
  assign n16414 = n1889 & ~n16413 ;
  assign n16415 = n1893 & ~n16414 ;
  assign n16416 = n1897 & ~n16415 ;
  assign n16417 = n1901 & ~n16416 ;
  assign n16418 = n1905 & ~n16417 ;
  assign n16419 = n1909 & ~n16418 ;
  assign n16420 = n1913 & ~n16419 ;
  assign n16421 = n1917 & ~n16420 ;
  assign n16422 = n1921 & ~n16421 ;
  assign n16423 = n1925 & ~n16422 ;
  assign n16424 = n1929 & ~n16423 ;
  assign n16425 = n1933 & ~n16424 ;
  assign n16426 = n1937 & ~n16425 ;
  assign n16427 = n1941 & ~n16426 ;
  assign n16428 = n1945 & ~n16427 ;
  assign n16429 = n1949 & ~n16428 ;
  assign n16430 = n1953 & ~n16429 ;
  assign n16431 = n2749 & ~n16430 ;
  assign n16432 = n263 & ~n16431 ;
  assign n16433 = n267 & ~n16432 ;
  assign n16434 = n271 & ~n16433 ;
  assign n16435 = n275 & ~n16434 ;
  assign n16436 = n279 & ~n16435 ;
  assign n16437 = n283 & ~n16436 ;
  assign n16438 = n287 & ~n16437 ;
  assign n16439 = n291 & ~n16438 ;
  assign n16440 = n295 & ~n16439 ;
  assign n16441 = n299 & ~n16440 ;
  assign n16442 = n303 & ~n16441 ;
  assign n16443 = n307 & ~n16442 ;
  assign n16444 = n311 & ~n16443 ;
  assign n16445 = n315 & ~n16444 ;
  assign n16446 = n319 & ~n16445 ;
  assign n16447 = n323 & ~n16446 ;
  assign n16448 = n327 & ~n16447 ;
  assign n16449 = n331 & ~n16448 ;
  assign n16450 = n335 & ~n16449 ;
  assign n16451 = n339 & ~n16450 ;
  assign n16452 = n343 & ~n16451 ;
  assign n16453 = n347 & ~n16452 ;
  assign n16454 = n351 & ~n16453 ;
  assign n16455 = n355 & ~n16454 ;
  assign n16456 = n359 & ~n16455 ;
  assign n16457 = n363 & ~n16456 ;
  assign n16458 = n367 & ~n16457 ;
  assign n16459 = n371 & ~n16458 ;
  assign n16460 = n375 & ~n16459 ;
  assign n16461 = n379 & ~n16460 ;
  assign n16462 = n383 & ~n16461 ;
  assign n16463 = n387 & ~n16462 ;
  assign n16464 = n391 & ~n16463 ;
  assign n16465 = n395 & ~n16464 ;
  assign n16466 = n399 & ~n16465 ;
  assign n16467 = n403 & ~n16466 ;
  assign n16468 = n407 & ~n16467 ;
  assign n16469 = n411 & ~n16468 ;
  assign n16470 = n415 & ~n16469 ;
  assign n16471 = n419 & ~n16470 ;
  assign n16472 = n423 & ~n16471 ;
  assign n16473 = n427 & ~n16472 ;
  assign n16474 = n431 & ~n16473 ;
  assign n16475 = n435 & ~n16474 ;
  assign n16476 = n439 & ~n16475 ;
  assign n16477 = n443 & ~n16476 ;
  assign n16478 = n447 & ~n16477 ;
  assign n16479 = n451 & ~n16478 ;
  assign n16480 = n455 & ~n16479 ;
  assign n16481 = n459 & ~n16480 ;
  assign n16482 = n463 & ~n16481 ;
  assign n16483 = n467 & ~n16482 ;
  assign n16484 = n471 & ~n16483 ;
  assign n16485 = x211 & ~n473 ;
  assign n16486 = ~n16484 & n16485 ;
  assign n16574 = n16486 & x339 ;
  assign n16487 = ~n817 & n2173 ;
  assign n16488 = n2178 & ~n16487 ;
  assign n16489 = n2182 & ~n16488 ;
  assign n16490 = n2186 & ~n16489 ;
  assign n16491 = n2190 & ~n16490 ;
  assign n16492 = n2194 & ~n16491 ;
  assign n16493 = n2198 & ~n16492 ;
  assign n16494 = n2202 & ~n16493 ;
  assign n16495 = n2206 & ~n16494 ;
  assign n16496 = n2210 & ~n16495 ;
  assign n16497 = n2214 & ~n16496 ;
  assign n16498 = n2218 & ~n16497 ;
  assign n16499 = n2222 & ~n16498 ;
  assign n16500 = n2226 & ~n16499 ;
  assign n16501 = n2230 & ~n16500 ;
  assign n16502 = n2234 & ~n16501 ;
  assign n16503 = n2238 & ~n16502 ;
  assign n16504 = n2242 & ~n16503 ;
  assign n16505 = n2246 & ~n16504 ;
  assign n16506 = n2250 & ~n16505 ;
  assign n16507 = n2254 & ~n16506 ;
  assign n16508 = n2258 & ~n16507 ;
  assign n16509 = n2262 & ~n16508 ;
  assign n16510 = n2266 & ~n16509 ;
  assign n16511 = n2270 & ~n16510 ;
  assign n16512 = n2274 & ~n16511 ;
  assign n16513 = n2278 & ~n16512 ;
  assign n16514 = n2282 & ~n16513 ;
  assign n16515 = n2286 & ~n16514 ;
  assign n16516 = n2290 & ~n16515 ;
  assign n16517 = n2836 & ~n16516 ;
  assign n16518 = n602 & ~n16517 ;
  assign n16519 = n606 & ~n16518 ;
  assign n16520 = n610 & ~n16519 ;
  assign n16521 = n614 & ~n16520 ;
  assign n16522 = n618 & ~n16521 ;
  assign n16523 = n622 & ~n16522 ;
  assign n16524 = n626 & ~n16523 ;
  assign n16525 = n630 & ~n16524 ;
  assign n16526 = n634 & ~n16525 ;
  assign n16527 = n638 & ~n16526 ;
  assign n16528 = n642 & ~n16527 ;
  assign n16529 = n646 & ~n16528 ;
  assign n16530 = n650 & ~n16529 ;
  assign n16531 = n654 & ~n16530 ;
  assign n16532 = n658 & ~n16531 ;
  assign n16533 = n662 & ~n16532 ;
  assign n16534 = n666 & ~n16533 ;
  assign n16535 = n670 & ~n16534 ;
  assign n16536 = n674 & ~n16535 ;
  assign n16537 = n678 & ~n16536 ;
  assign n16538 = n682 & ~n16537 ;
  assign n16539 = n686 & ~n16538 ;
  assign n16540 = n690 & ~n16539 ;
  assign n16541 = n694 & ~n16540 ;
  assign n16542 = n698 & ~n16541 ;
  assign n16543 = n702 & ~n16542 ;
  assign n16544 = n706 & ~n16543 ;
  assign n16545 = n710 & ~n16544 ;
  assign n16546 = n714 & ~n16545 ;
  assign n16547 = n718 & ~n16546 ;
  assign n16548 = n722 & ~n16547 ;
  assign n16549 = n726 & ~n16548 ;
  assign n16550 = n730 & ~n16549 ;
  assign n16551 = n734 & ~n16550 ;
  assign n16552 = n738 & ~n16551 ;
  assign n16553 = n742 & ~n16552 ;
  assign n16554 = n746 & ~n16553 ;
  assign n16555 = n750 & ~n16554 ;
  assign n16556 = n754 & ~n16555 ;
  assign n16557 = n758 & ~n16556 ;
  assign n16558 = n762 & ~n16557 ;
  assign n16559 = n766 & ~n16558 ;
  assign n16560 = n770 & ~n16559 ;
  assign n16561 = n774 & ~n16560 ;
  assign n16562 = n778 & ~n16561 ;
  assign n16563 = n782 & ~n16562 ;
  assign n16564 = n786 & ~n16563 ;
  assign n16565 = n790 & ~n16564 ;
  assign n16566 = n794 & ~n16565 ;
  assign n16567 = n798 & ~n16566 ;
  assign n16568 = n802 & ~n16567 ;
  assign n16569 = n806 & ~n16568 ;
  assign n16570 = n810 & ~n16569 ;
  assign n16571 = ~x211 & ~n812 ;
  assign n16572 = ~n16570 & n16571 ;
  assign n16575 = ~n16572 & ~x339 ;
  assign n16576 = ~n16574 & ~n16575 ;
  assign n16577 = n482 & ~n1160 ;
  assign n16578 = n487 & ~n16577 ;
  assign n16579 = n491 & ~n16578 ;
  assign n16580 = n495 & ~n16579 ;
  assign n16581 = n499 & ~n16580 ;
  assign n16582 = n503 & ~n16581 ;
  assign n16583 = n507 & ~n16582 ;
  assign n16584 = n511 & ~n16583 ;
  assign n16585 = n515 & ~n16584 ;
  assign n16586 = n519 & ~n16585 ;
  assign n16587 = n523 & ~n16586 ;
  assign n16588 = n527 & ~n16587 ;
  assign n16589 = n531 & ~n16588 ;
  assign n16590 = n535 & ~n16589 ;
  assign n16591 = n539 & ~n16590 ;
  assign n16592 = n543 & ~n16591 ;
  assign n16593 = n547 & ~n16592 ;
  assign n16594 = n551 & ~n16593 ;
  assign n16595 = n555 & ~n16594 ;
  assign n16596 = n559 & ~n16595 ;
  assign n16597 = n563 & ~n16596 ;
  assign n16598 = n567 & ~n16597 ;
  assign n16599 = n571 & ~n16598 ;
  assign n16600 = n575 & ~n16599 ;
  assign n16601 = n579 & ~n16600 ;
  assign n16602 = n583 & ~n16601 ;
  assign n16603 = n587 & ~n16602 ;
  assign n16604 = n591 & ~n16603 ;
  assign n16605 = n2382 & ~n16604 ;
  assign n16606 = n2384 & ~n16605 ;
  assign n16607 = n2927 & ~n16606 ;
  assign n16608 = n945 & ~n16607 ;
  assign n16609 = n949 & ~n16608 ;
  assign n16610 = n953 & ~n16609 ;
  assign n16611 = n957 & ~n16610 ;
  assign n16612 = n961 & ~n16611 ;
  assign n16613 = n965 & ~n16612 ;
  assign n16614 = n969 & ~n16613 ;
  assign n16615 = n973 & ~n16614 ;
  assign n16616 = n977 & ~n16615 ;
  assign n16617 = n981 & ~n16616 ;
  assign n16618 = n985 & ~n16617 ;
  assign n16619 = n989 & ~n16618 ;
  assign n16620 = n993 & ~n16619 ;
  assign n16621 = n997 & ~n16620 ;
  assign n16622 = n1001 & ~n16621 ;
  assign n16623 = n1005 & ~n16622 ;
  assign n16624 = n1009 & ~n16623 ;
  assign n16625 = n1013 & ~n16624 ;
  assign n16626 = n1017 & ~n16625 ;
  assign n16627 = n1021 & ~n16626 ;
  assign n16628 = n1025 & ~n16627 ;
  assign n16629 = n1029 & ~n16628 ;
  assign n16630 = n1033 & ~n16629 ;
  assign n16631 = n1037 & ~n16630 ;
  assign n16632 = n1041 & ~n16631 ;
  assign n16633 = n1045 & ~n16632 ;
  assign n16634 = n1049 & ~n16633 ;
  assign n16635 = n1053 & ~n16634 ;
  assign n16636 = n1057 & ~n16635 ;
  assign n16637 = n1061 & ~n16636 ;
  assign n16638 = n1065 & ~n16637 ;
  assign n16639 = n1069 & ~n16638 ;
  assign n16640 = n1073 & ~n16639 ;
  assign n16641 = n1077 & ~n16640 ;
  assign n16642 = n1081 & ~n16641 ;
  assign n16643 = n1085 & ~n16642 ;
  assign n16644 = n1089 & ~n16643 ;
  assign n16645 = n1093 & ~n16644 ;
  assign n16646 = n1097 & ~n16645 ;
  assign n16647 = n1101 & ~n16646 ;
  assign n16648 = n1105 & ~n16647 ;
  assign n16649 = n1109 & ~n16648 ;
  assign n16650 = n1113 & ~n16649 ;
  assign n16651 = n1117 & ~n16650 ;
  assign n16652 = n1121 & ~n16651 ;
  assign n16653 = n1125 & ~n16652 ;
  assign n16654 = n1129 & ~n16653 ;
  assign n16655 = n1133 & ~n16654 ;
  assign n16656 = n1137 & ~n16655 ;
  assign n16657 = n1141 & ~n16656 ;
  assign n16658 = n1145 & ~n16657 ;
  assign n16659 = n1149 & ~n16658 ;
  assign n16660 = n1153 & ~n16659 ;
  assign n16661 = x212 & ~n1155 ;
  assign n16662 = ~n16660 & n16661 ;
  assign n16750 = n16662 & x340 ;
  assign n16663 = n821 & ~n1499 ;
  assign n16664 = n826 & ~n16663 ;
  assign n16665 = n830 & ~n16664 ;
  assign n16666 = n834 & ~n16665 ;
  assign n16667 = n838 & ~n16666 ;
  assign n16668 = n842 & ~n16667 ;
  assign n16669 = n846 & ~n16668 ;
  assign n16670 = n850 & ~n16669 ;
  assign n16671 = n854 & ~n16670 ;
  assign n16672 = n858 & ~n16671 ;
  assign n16673 = n862 & ~n16672 ;
  assign n16674 = n866 & ~n16673 ;
  assign n16675 = n870 & ~n16674 ;
  assign n16676 = n874 & ~n16675 ;
  assign n16677 = n878 & ~n16676 ;
  assign n16678 = n882 & ~n16677 ;
  assign n16679 = n886 & ~n16678 ;
  assign n16680 = n890 & ~n16679 ;
  assign n16681 = n894 & ~n16680 ;
  assign n16682 = n898 & ~n16681 ;
  assign n16683 = n902 & ~n16682 ;
  assign n16684 = n906 & ~n16683 ;
  assign n16685 = n910 & ~n16684 ;
  assign n16686 = n914 & ~n16685 ;
  assign n16687 = n918 & ~n16686 ;
  assign n16688 = n922 & ~n16687 ;
  assign n16689 = n926 & ~n16688 ;
  assign n16690 = n930 & ~n16689 ;
  assign n16691 = n2472 & ~n16690 ;
  assign n16692 = n2474 & ~n16691 ;
  assign n16693 = n3014 & ~n16692 ;
  assign n16694 = n1284 & ~n16693 ;
  assign n16695 = n1288 & ~n16694 ;
  assign n16696 = n1292 & ~n16695 ;
  assign n16697 = n1296 & ~n16696 ;
  assign n16698 = n1300 & ~n16697 ;
  assign n16699 = n1304 & ~n16698 ;
  assign n16700 = n1308 & ~n16699 ;
  assign n16701 = n1312 & ~n16700 ;
  assign n16702 = n1316 & ~n16701 ;
  assign n16703 = n1320 & ~n16702 ;
  assign n16704 = n1324 & ~n16703 ;
  assign n16705 = n1328 & ~n16704 ;
  assign n16706 = n1332 & ~n16705 ;
  assign n16707 = n1336 & ~n16706 ;
  assign n16708 = n1340 & ~n16707 ;
  assign n16709 = n1344 & ~n16708 ;
  assign n16710 = n1348 & ~n16709 ;
  assign n16711 = n1352 & ~n16710 ;
  assign n16712 = n1356 & ~n16711 ;
  assign n16713 = n1360 & ~n16712 ;
  assign n16714 = n1364 & ~n16713 ;
  assign n16715 = n1368 & ~n16714 ;
  assign n16716 = n1372 & ~n16715 ;
  assign n16717 = n1376 & ~n16716 ;
  assign n16718 = n1380 & ~n16717 ;
  assign n16719 = n1384 & ~n16718 ;
  assign n16720 = n1388 & ~n16719 ;
  assign n16721 = n1392 & ~n16720 ;
  assign n16722 = n1396 & ~n16721 ;
  assign n16723 = n1400 & ~n16722 ;
  assign n16724 = n1404 & ~n16723 ;
  assign n16725 = n1408 & ~n16724 ;
  assign n16726 = n1412 & ~n16725 ;
  assign n16727 = n1416 & ~n16726 ;
  assign n16728 = n1420 & ~n16727 ;
  assign n16729 = n1424 & ~n16728 ;
  assign n16730 = n1428 & ~n16729 ;
  assign n16731 = n1432 & ~n16730 ;
  assign n16732 = n1436 & ~n16731 ;
  assign n16733 = n1440 & ~n16732 ;
  assign n16734 = n1444 & ~n16733 ;
  assign n16735 = n1448 & ~n16734 ;
  assign n16736 = n1452 & ~n16735 ;
  assign n16737 = n1456 & ~n16736 ;
  assign n16738 = n1460 & ~n16737 ;
  assign n16739 = n1464 & ~n16738 ;
  assign n16740 = n1468 & ~n16739 ;
  assign n16741 = n1472 & ~n16740 ;
  assign n16742 = n1476 & ~n16741 ;
  assign n16743 = n1480 & ~n16742 ;
  assign n16744 = n1484 & ~n16743 ;
  assign n16745 = n1488 & ~n16744 ;
  assign n16746 = n1492 & ~n16745 ;
  assign n16747 = ~x212 & ~n1494 ;
  assign n16748 = ~n16746 & n16747 ;
  assign n16751 = ~n16748 & ~x340 ;
  assign n16752 = ~n16750 & ~n16751 ;
  assign n16753 = n1164 & ~n1840 ;
  assign n16754 = n1169 & ~n16753 ;
  assign n16755 = n1173 & ~n16754 ;
  assign n16756 = n1177 & ~n16755 ;
  assign n16757 = n1181 & ~n16756 ;
  assign n16758 = n1185 & ~n16757 ;
  assign n16759 = n1189 & ~n16758 ;
  assign n16760 = n1193 & ~n16759 ;
  assign n16761 = n1197 & ~n16760 ;
  assign n16762 = n1201 & ~n16761 ;
  assign n16763 = n1205 & ~n16762 ;
  assign n16764 = n1209 & ~n16763 ;
  assign n16765 = n1213 & ~n16764 ;
  assign n16766 = n1217 & ~n16765 ;
  assign n16767 = n1221 & ~n16766 ;
  assign n16768 = n1225 & ~n16767 ;
  assign n16769 = n1229 & ~n16768 ;
  assign n16770 = n1233 & ~n16769 ;
  assign n16771 = n1237 & ~n16770 ;
  assign n16772 = n1241 & ~n16771 ;
  assign n16773 = n1245 & ~n16772 ;
  assign n16774 = n1249 & ~n16773 ;
  assign n16775 = n1253 & ~n16774 ;
  assign n16776 = n1257 & ~n16775 ;
  assign n16777 = n1261 & ~n16776 ;
  assign n16778 = n1265 & ~n16777 ;
  assign n16779 = n1269 & ~n16778 ;
  assign n16780 = n1273 & ~n16779 ;
  assign n16781 = n2566 & ~n16780 ;
  assign n16782 = n2568 & ~n16781 ;
  assign n16783 = n3105 & ~n16782 ;
  assign n16784 = n1625 & ~n16783 ;
  assign n16785 = n1629 & ~n16784 ;
  assign n16786 = n1633 & ~n16785 ;
  assign n16787 = n1637 & ~n16786 ;
  assign n16788 = n1641 & ~n16787 ;
  assign n16789 = n1645 & ~n16788 ;
  assign n16790 = n1649 & ~n16789 ;
  assign n16791 = n1653 & ~n16790 ;
  assign n16792 = n1657 & ~n16791 ;
  assign n16793 = n1661 & ~n16792 ;
  assign n16794 = n1665 & ~n16793 ;
  assign n16795 = n1669 & ~n16794 ;
  assign n16796 = n1673 & ~n16795 ;
  assign n16797 = n1677 & ~n16796 ;
  assign n16798 = n1681 & ~n16797 ;
  assign n16799 = n1685 & ~n16798 ;
  assign n16800 = n1689 & ~n16799 ;
  assign n16801 = n1693 & ~n16800 ;
  assign n16802 = n1697 & ~n16801 ;
  assign n16803 = n1701 & ~n16802 ;
  assign n16804 = n1705 & ~n16803 ;
  assign n16805 = n1709 & ~n16804 ;
  assign n16806 = n1713 & ~n16805 ;
  assign n16807 = n1717 & ~n16806 ;
  assign n16808 = n1721 & ~n16807 ;
  assign n16809 = n1725 & ~n16808 ;
  assign n16810 = n1729 & ~n16809 ;
  assign n16811 = n1733 & ~n16810 ;
  assign n16812 = n1737 & ~n16811 ;
  assign n16813 = n1741 & ~n16812 ;
  assign n16814 = n1745 & ~n16813 ;
  assign n16815 = n1749 & ~n16814 ;
  assign n16816 = n1753 & ~n16815 ;
  assign n16817 = n1757 & ~n16816 ;
  assign n16818 = n1761 & ~n16817 ;
  assign n16819 = n1765 & ~n16818 ;
  assign n16820 = n1769 & ~n16819 ;
  assign n16821 = n1773 & ~n16820 ;
  assign n16822 = n1777 & ~n16821 ;
  assign n16823 = n1781 & ~n16822 ;
  assign n16824 = n1785 & ~n16823 ;
  assign n16825 = n1789 & ~n16824 ;
  assign n16826 = n1793 & ~n16825 ;
  assign n16827 = n1797 & ~n16826 ;
  assign n16828 = n1801 & ~n16827 ;
  assign n16829 = n1805 & ~n16828 ;
  assign n16830 = n1809 & ~n16829 ;
  assign n16831 = n1813 & ~n16830 ;
  assign n16832 = n1817 & ~n16831 ;
  assign n16833 = n1821 & ~n16832 ;
  assign n16834 = n1825 & ~n16833 ;
  assign n16835 = n1829 & ~n16834 ;
  assign n16836 = n1833 & ~n16835 ;
  assign n16837 = x213 & ~n1835 ;
  assign n16838 = ~n16836 & n16837 ;
  assign n16926 = n16838 & x341 ;
  assign n16839 = n1503 & ~n2177 ;
  assign n16840 = n1508 & ~n16839 ;
  assign n16841 = n1512 & ~n16840 ;
  assign n16842 = n1516 & ~n16841 ;
  assign n16843 = n1520 & ~n16842 ;
  assign n16844 = n1524 & ~n16843 ;
  assign n16845 = n1528 & ~n16844 ;
  assign n16846 = n1532 & ~n16845 ;
  assign n16847 = n1536 & ~n16846 ;
  assign n16848 = n1540 & ~n16847 ;
  assign n16849 = n1544 & ~n16848 ;
  assign n16850 = n1548 & ~n16849 ;
  assign n16851 = n1552 & ~n16850 ;
  assign n16852 = n1556 & ~n16851 ;
  assign n16853 = n1560 & ~n16852 ;
  assign n16854 = n1564 & ~n16853 ;
  assign n16855 = n1568 & ~n16854 ;
  assign n16856 = n1572 & ~n16855 ;
  assign n16857 = n1576 & ~n16856 ;
  assign n16858 = n1580 & ~n16857 ;
  assign n16859 = n1584 & ~n16858 ;
  assign n16860 = n1588 & ~n16859 ;
  assign n16861 = n1592 & ~n16860 ;
  assign n16862 = n1596 & ~n16861 ;
  assign n16863 = n1600 & ~n16862 ;
  assign n16864 = n1604 & ~n16863 ;
  assign n16865 = n1608 & ~n16864 ;
  assign n16866 = n1612 & ~n16865 ;
  assign n16867 = n2656 & ~n16866 ;
  assign n16868 = n2658 & ~n16867 ;
  assign n16869 = n3192 & ~n16868 ;
  assign n16870 = n1962 & ~n16869 ;
  assign n16871 = n1966 & ~n16870 ;
  assign n16872 = n1970 & ~n16871 ;
  assign n16873 = n1974 & ~n16872 ;
  assign n16874 = n1978 & ~n16873 ;
  assign n16875 = n1982 & ~n16874 ;
  assign n16876 = n1986 & ~n16875 ;
  assign n16877 = n1990 & ~n16876 ;
  assign n16878 = n1994 & ~n16877 ;
  assign n16879 = n1998 & ~n16878 ;
  assign n16880 = n2002 & ~n16879 ;
  assign n16881 = n2006 & ~n16880 ;
  assign n16882 = n2010 & ~n16881 ;
  assign n16883 = n2014 & ~n16882 ;
  assign n16884 = n2018 & ~n16883 ;
  assign n16885 = n2022 & ~n16884 ;
  assign n16886 = n2026 & ~n16885 ;
  assign n16887 = n2030 & ~n16886 ;
  assign n16888 = n2034 & ~n16887 ;
  assign n16889 = n2038 & ~n16888 ;
  assign n16890 = n2042 & ~n16889 ;
  assign n16891 = n2046 & ~n16890 ;
  assign n16892 = n2050 & ~n16891 ;
  assign n16893 = n2054 & ~n16892 ;
  assign n16894 = n2058 & ~n16893 ;
  assign n16895 = n2062 & ~n16894 ;
  assign n16896 = n2066 & ~n16895 ;
  assign n16897 = n2070 & ~n16896 ;
  assign n16898 = n2074 & ~n16897 ;
  assign n16899 = n2078 & ~n16898 ;
  assign n16900 = n2082 & ~n16899 ;
  assign n16901 = n2086 & ~n16900 ;
  assign n16902 = n2090 & ~n16901 ;
  assign n16903 = n2094 & ~n16902 ;
  assign n16904 = n2098 & ~n16903 ;
  assign n16905 = n2102 & ~n16904 ;
  assign n16906 = n2106 & ~n16905 ;
  assign n16907 = n2110 & ~n16906 ;
  assign n16908 = n2114 & ~n16907 ;
  assign n16909 = n2118 & ~n16908 ;
  assign n16910 = n2122 & ~n16909 ;
  assign n16911 = n2126 & ~n16910 ;
  assign n16912 = n2130 & ~n16911 ;
  assign n16913 = n2134 & ~n16912 ;
  assign n16914 = n2138 & ~n16913 ;
  assign n16915 = n2142 & ~n16914 ;
  assign n16916 = n2146 & ~n16915 ;
  assign n16917 = n2150 & ~n16916 ;
  assign n16918 = n2154 & ~n16917 ;
  assign n16919 = n2158 & ~n16918 ;
  assign n16920 = n2162 & ~n16919 ;
  assign n16921 = n2166 & ~n16920 ;
  assign n16922 = n2170 & ~n16921 ;
  assign n16923 = ~x213 & ~n2172 ;
  assign n16924 = ~n16922 & n16923 ;
  assign n16927 = ~n16924 & ~x341 ;
  assign n16928 = ~n16926 & ~n16927 ;
  assign n16929 = ~n486 & n1844 ;
  assign n16930 = n1849 & ~n16929 ;
  assign n16931 = n1853 & ~n16930 ;
  assign n16932 = n1857 & ~n16931 ;
  assign n16933 = n1861 & ~n16932 ;
  assign n16934 = n1865 & ~n16933 ;
  assign n16935 = n1869 & ~n16934 ;
  assign n16936 = n1873 & ~n16935 ;
  assign n16937 = n1877 & ~n16936 ;
  assign n16938 = n1881 & ~n16937 ;
  assign n16939 = n1885 & ~n16938 ;
  assign n16940 = n1889 & ~n16939 ;
  assign n16941 = n1893 & ~n16940 ;
  assign n16942 = n1897 & ~n16941 ;
  assign n16943 = n1901 & ~n16942 ;
  assign n16944 = n1905 & ~n16943 ;
  assign n16945 = n1909 & ~n16944 ;
  assign n16946 = n1913 & ~n16945 ;
  assign n16947 = n1917 & ~n16946 ;
  assign n16948 = n1921 & ~n16947 ;
  assign n16949 = n1925 & ~n16948 ;
  assign n16950 = n1929 & ~n16949 ;
  assign n16951 = n1933 & ~n16950 ;
  assign n16952 = n1937 & ~n16951 ;
  assign n16953 = n1941 & ~n16952 ;
  assign n16954 = n1945 & ~n16953 ;
  assign n16955 = n1949 & ~n16954 ;
  assign n16956 = n1953 & ~n16955 ;
  assign n16957 = n2749 & ~n16956 ;
  assign n16958 = n263 & ~n16957 ;
  assign n16959 = n267 & ~n16958 ;
  assign n16960 = n271 & ~n16959 ;
  assign n16961 = n275 & ~n16960 ;
  assign n16962 = n279 & ~n16961 ;
  assign n16963 = n283 & ~n16962 ;
  assign n16964 = n287 & ~n16963 ;
  assign n16965 = n291 & ~n16964 ;
  assign n16966 = n295 & ~n16965 ;
  assign n16967 = n299 & ~n16966 ;
  assign n16968 = n303 & ~n16967 ;
  assign n16969 = n307 & ~n16968 ;
  assign n16970 = n311 & ~n16969 ;
  assign n16971 = n315 & ~n16970 ;
  assign n16972 = n319 & ~n16971 ;
  assign n16973 = n323 & ~n16972 ;
  assign n16974 = n327 & ~n16973 ;
  assign n16975 = n331 & ~n16974 ;
  assign n16976 = n335 & ~n16975 ;
  assign n16977 = n339 & ~n16976 ;
  assign n16978 = n343 & ~n16977 ;
  assign n16979 = n347 & ~n16978 ;
  assign n16980 = n351 & ~n16979 ;
  assign n16981 = n355 & ~n16980 ;
  assign n16982 = n359 & ~n16981 ;
  assign n16983 = n363 & ~n16982 ;
  assign n16984 = n367 & ~n16983 ;
  assign n16985 = n371 & ~n16984 ;
  assign n16986 = n375 & ~n16985 ;
  assign n16987 = n379 & ~n16986 ;
  assign n16988 = n383 & ~n16987 ;
  assign n16989 = n387 & ~n16988 ;
  assign n16990 = n391 & ~n16989 ;
  assign n16991 = n395 & ~n16990 ;
  assign n16992 = n399 & ~n16991 ;
  assign n16993 = n403 & ~n16992 ;
  assign n16994 = n407 & ~n16993 ;
  assign n16995 = n411 & ~n16994 ;
  assign n16996 = n415 & ~n16995 ;
  assign n16997 = n419 & ~n16996 ;
  assign n16998 = n423 & ~n16997 ;
  assign n16999 = n427 & ~n16998 ;
  assign n17000 = n431 & ~n16999 ;
  assign n17001 = n435 & ~n17000 ;
  assign n17002 = n439 & ~n17001 ;
  assign n17003 = n443 & ~n17002 ;
  assign n17004 = n447 & ~n17003 ;
  assign n17005 = n451 & ~n17004 ;
  assign n17006 = n455 & ~n17005 ;
  assign n17007 = n459 & ~n17006 ;
  assign n17008 = n463 & ~n17007 ;
  assign n17009 = n467 & ~n17008 ;
  assign n17010 = n471 & ~n17009 ;
  assign n17011 = n475 & ~n17010 ;
  assign n17012 = n479 & ~n17011 ;
  assign n17013 = x214 & ~n481 ;
  assign n17014 = ~n17012 & n17013 ;
  assign n17102 = n17014 & x342 ;
  assign n17015 = ~n825 & n2181 ;
  assign n17016 = n2186 & ~n17015 ;
  assign n17017 = n2190 & ~n17016 ;
  assign n17018 = n2194 & ~n17017 ;
  assign n17019 = n2198 & ~n17018 ;
  assign n17020 = n2202 & ~n17019 ;
  assign n17021 = n2206 & ~n17020 ;
  assign n17022 = n2210 & ~n17021 ;
  assign n17023 = n2214 & ~n17022 ;
  assign n17024 = n2218 & ~n17023 ;
  assign n17025 = n2222 & ~n17024 ;
  assign n17026 = n2226 & ~n17025 ;
  assign n17027 = n2230 & ~n17026 ;
  assign n17028 = n2234 & ~n17027 ;
  assign n17029 = n2238 & ~n17028 ;
  assign n17030 = n2242 & ~n17029 ;
  assign n17031 = n2246 & ~n17030 ;
  assign n17032 = n2250 & ~n17031 ;
  assign n17033 = n2254 & ~n17032 ;
  assign n17034 = n2258 & ~n17033 ;
  assign n17035 = n2262 & ~n17034 ;
  assign n17036 = n2266 & ~n17035 ;
  assign n17037 = n2270 & ~n17036 ;
  assign n17038 = n2274 & ~n17037 ;
  assign n17039 = n2278 & ~n17038 ;
  assign n17040 = n2282 & ~n17039 ;
  assign n17041 = n2286 & ~n17040 ;
  assign n17042 = n2290 & ~n17041 ;
  assign n17043 = n2836 & ~n17042 ;
  assign n17044 = n602 & ~n17043 ;
  assign n17045 = n606 & ~n17044 ;
  assign n17046 = n610 & ~n17045 ;
  assign n17047 = n614 & ~n17046 ;
  assign n17048 = n618 & ~n17047 ;
  assign n17049 = n622 & ~n17048 ;
  assign n17050 = n626 & ~n17049 ;
  assign n17051 = n630 & ~n17050 ;
  assign n17052 = n634 & ~n17051 ;
  assign n17053 = n638 & ~n17052 ;
  assign n17054 = n642 & ~n17053 ;
  assign n17055 = n646 & ~n17054 ;
  assign n17056 = n650 & ~n17055 ;
  assign n17057 = n654 & ~n17056 ;
  assign n17058 = n658 & ~n17057 ;
  assign n17059 = n662 & ~n17058 ;
  assign n17060 = n666 & ~n17059 ;
  assign n17061 = n670 & ~n17060 ;
  assign n17062 = n674 & ~n17061 ;
  assign n17063 = n678 & ~n17062 ;
  assign n17064 = n682 & ~n17063 ;
  assign n17065 = n686 & ~n17064 ;
  assign n17066 = n690 & ~n17065 ;
  assign n17067 = n694 & ~n17066 ;
  assign n17068 = n698 & ~n17067 ;
  assign n17069 = n702 & ~n17068 ;
  assign n17070 = n706 & ~n17069 ;
  assign n17071 = n710 & ~n17070 ;
  assign n17072 = n714 & ~n17071 ;
  assign n17073 = n718 & ~n17072 ;
  assign n17074 = n722 & ~n17073 ;
  assign n17075 = n726 & ~n17074 ;
  assign n17076 = n730 & ~n17075 ;
  assign n17077 = n734 & ~n17076 ;
  assign n17078 = n738 & ~n17077 ;
  assign n17079 = n742 & ~n17078 ;
  assign n17080 = n746 & ~n17079 ;
  assign n17081 = n750 & ~n17080 ;
  assign n17082 = n754 & ~n17081 ;
  assign n17083 = n758 & ~n17082 ;
  assign n17084 = n762 & ~n17083 ;
  assign n17085 = n766 & ~n17084 ;
  assign n17086 = n770 & ~n17085 ;
  assign n17087 = n774 & ~n17086 ;
  assign n17088 = n778 & ~n17087 ;
  assign n17089 = n782 & ~n17088 ;
  assign n17090 = n786 & ~n17089 ;
  assign n17091 = n790 & ~n17090 ;
  assign n17092 = n794 & ~n17091 ;
  assign n17093 = n798 & ~n17092 ;
  assign n17094 = n802 & ~n17093 ;
  assign n17095 = n806 & ~n17094 ;
  assign n17096 = n810 & ~n17095 ;
  assign n17097 = n814 & ~n17096 ;
  assign n17098 = n818 & ~n17097 ;
  assign n17099 = ~x214 & ~n820 ;
  assign n17100 = ~n17098 & n17099 ;
  assign n17103 = ~n17100 & ~x342 ;
  assign n17104 = ~n17102 & ~n17103 ;
  assign n17105 = n490 & ~n1168 ;
  assign n17106 = n495 & ~n17105 ;
  assign n17107 = n499 & ~n17106 ;
  assign n17108 = n503 & ~n17107 ;
  assign n17109 = n507 & ~n17108 ;
  assign n17110 = n511 & ~n17109 ;
  assign n17111 = n515 & ~n17110 ;
  assign n17112 = n519 & ~n17111 ;
  assign n17113 = n523 & ~n17112 ;
  assign n17114 = n527 & ~n17113 ;
  assign n17115 = n531 & ~n17114 ;
  assign n17116 = n535 & ~n17115 ;
  assign n17117 = n539 & ~n17116 ;
  assign n17118 = n543 & ~n17117 ;
  assign n17119 = n547 & ~n17118 ;
  assign n17120 = n551 & ~n17119 ;
  assign n17121 = n555 & ~n17120 ;
  assign n17122 = n559 & ~n17121 ;
  assign n17123 = n563 & ~n17122 ;
  assign n17124 = n567 & ~n17123 ;
  assign n17125 = n571 & ~n17124 ;
  assign n17126 = n575 & ~n17125 ;
  assign n17127 = n579 & ~n17126 ;
  assign n17128 = n583 & ~n17127 ;
  assign n17129 = n587 & ~n17128 ;
  assign n17130 = n591 & ~n17129 ;
  assign n17131 = n2382 & ~n17130 ;
  assign n17132 = n2384 & ~n17131 ;
  assign n17133 = n2927 & ~n17132 ;
  assign n17134 = n945 & ~n17133 ;
  assign n17135 = n949 & ~n17134 ;
  assign n17136 = n953 & ~n17135 ;
  assign n17137 = n957 & ~n17136 ;
  assign n17138 = n961 & ~n17137 ;
  assign n17139 = n965 & ~n17138 ;
  assign n17140 = n969 & ~n17139 ;
  assign n17141 = n973 & ~n17140 ;
  assign n17142 = n977 & ~n17141 ;
  assign n17143 = n981 & ~n17142 ;
  assign n17144 = n985 & ~n17143 ;
  assign n17145 = n989 & ~n17144 ;
  assign n17146 = n993 & ~n17145 ;
  assign n17147 = n997 & ~n17146 ;
  assign n17148 = n1001 & ~n17147 ;
  assign n17149 = n1005 & ~n17148 ;
  assign n17150 = n1009 & ~n17149 ;
  assign n17151 = n1013 & ~n17150 ;
  assign n17152 = n1017 & ~n17151 ;
  assign n17153 = n1021 & ~n17152 ;
  assign n17154 = n1025 & ~n17153 ;
  assign n17155 = n1029 & ~n17154 ;
  assign n17156 = n1033 & ~n17155 ;
  assign n17157 = n1037 & ~n17156 ;
  assign n17158 = n1041 & ~n17157 ;
  assign n17159 = n1045 & ~n17158 ;
  assign n17160 = n1049 & ~n17159 ;
  assign n17161 = n1053 & ~n17160 ;
  assign n17162 = n1057 & ~n17161 ;
  assign n17163 = n1061 & ~n17162 ;
  assign n17164 = n1065 & ~n17163 ;
  assign n17165 = n1069 & ~n17164 ;
  assign n17166 = n1073 & ~n17165 ;
  assign n17167 = n1077 & ~n17166 ;
  assign n17168 = n1081 & ~n17167 ;
  assign n17169 = n1085 & ~n17168 ;
  assign n17170 = n1089 & ~n17169 ;
  assign n17171 = n1093 & ~n17170 ;
  assign n17172 = n1097 & ~n17171 ;
  assign n17173 = n1101 & ~n17172 ;
  assign n17174 = n1105 & ~n17173 ;
  assign n17175 = n1109 & ~n17174 ;
  assign n17176 = n1113 & ~n17175 ;
  assign n17177 = n1117 & ~n17176 ;
  assign n17178 = n1121 & ~n17177 ;
  assign n17179 = n1125 & ~n17178 ;
  assign n17180 = n1129 & ~n17179 ;
  assign n17181 = n1133 & ~n17180 ;
  assign n17182 = n1137 & ~n17181 ;
  assign n17183 = n1141 & ~n17182 ;
  assign n17184 = n1145 & ~n17183 ;
  assign n17185 = n1149 & ~n17184 ;
  assign n17186 = n1153 & ~n17185 ;
  assign n17187 = n1157 & ~n17186 ;
  assign n17188 = n1161 & ~n17187 ;
  assign n17189 = x215 & ~n1163 ;
  assign n17190 = ~n17188 & n17189 ;
  assign n17278 = n17190 & x343 ;
  assign n17191 = n829 & ~n1507 ;
  assign n17192 = n834 & ~n17191 ;
  assign n17193 = n838 & ~n17192 ;
  assign n17194 = n842 & ~n17193 ;
  assign n17195 = n846 & ~n17194 ;
  assign n17196 = n850 & ~n17195 ;
  assign n17197 = n854 & ~n17196 ;
  assign n17198 = n858 & ~n17197 ;
  assign n17199 = n862 & ~n17198 ;
  assign n17200 = n866 & ~n17199 ;
  assign n17201 = n870 & ~n17200 ;
  assign n17202 = n874 & ~n17201 ;
  assign n17203 = n878 & ~n17202 ;
  assign n17204 = n882 & ~n17203 ;
  assign n17205 = n886 & ~n17204 ;
  assign n17206 = n890 & ~n17205 ;
  assign n17207 = n894 & ~n17206 ;
  assign n17208 = n898 & ~n17207 ;
  assign n17209 = n902 & ~n17208 ;
  assign n17210 = n906 & ~n17209 ;
  assign n17211 = n910 & ~n17210 ;
  assign n17212 = n914 & ~n17211 ;
  assign n17213 = n918 & ~n17212 ;
  assign n17214 = n922 & ~n17213 ;
  assign n17215 = n926 & ~n17214 ;
  assign n17216 = n930 & ~n17215 ;
  assign n17217 = n2472 & ~n17216 ;
  assign n17218 = n2474 & ~n17217 ;
  assign n17219 = n3014 & ~n17218 ;
  assign n17220 = n1284 & ~n17219 ;
  assign n17221 = n1288 & ~n17220 ;
  assign n17222 = n1292 & ~n17221 ;
  assign n17223 = n1296 & ~n17222 ;
  assign n17224 = n1300 & ~n17223 ;
  assign n17225 = n1304 & ~n17224 ;
  assign n17226 = n1308 & ~n17225 ;
  assign n17227 = n1312 & ~n17226 ;
  assign n17228 = n1316 & ~n17227 ;
  assign n17229 = n1320 & ~n17228 ;
  assign n17230 = n1324 & ~n17229 ;
  assign n17231 = n1328 & ~n17230 ;
  assign n17232 = n1332 & ~n17231 ;
  assign n17233 = n1336 & ~n17232 ;
  assign n17234 = n1340 & ~n17233 ;
  assign n17235 = n1344 & ~n17234 ;
  assign n17236 = n1348 & ~n17235 ;
  assign n17237 = n1352 & ~n17236 ;
  assign n17238 = n1356 & ~n17237 ;
  assign n17239 = n1360 & ~n17238 ;
  assign n17240 = n1364 & ~n17239 ;
  assign n17241 = n1368 & ~n17240 ;
  assign n17242 = n1372 & ~n17241 ;
  assign n17243 = n1376 & ~n17242 ;
  assign n17244 = n1380 & ~n17243 ;
  assign n17245 = n1384 & ~n17244 ;
  assign n17246 = n1388 & ~n17245 ;
  assign n17247 = n1392 & ~n17246 ;
  assign n17248 = n1396 & ~n17247 ;
  assign n17249 = n1400 & ~n17248 ;
  assign n17250 = n1404 & ~n17249 ;
  assign n17251 = n1408 & ~n17250 ;
  assign n17252 = n1412 & ~n17251 ;
  assign n17253 = n1416 & ~n17252 ;
  assign n17254 = n1420 & ~n17253 ;
  assign n17255 = n1424 & ~n17254 ;
  assign n17256 = n1428 & ~n17255 ;
  assign n17257 = n1432 & ~n17256 ;
  assign n17258 = n1436 & ~n17257 ;
  assign n17259 = n1440 & ~n17258 ;
  assign n17260 = n1444 & ~n17259 ;
  assign n17261 = n1448 & ~n17260 ;
  assign n17262 = n1452 & ~n17261 ;
  assign n17263 = n1456 & ~n17262 ;
  assign n17264 = n1460 & ~n17263 ;
  assign n17265 = n1464 & ~n17264 ;
  assign n17266 = n1468 & ~n17265 ;
  assign n17267 = n1472 & ~n17266 ;
  assign n17268 = n1476 & ~n17267 ;
  assign n17269 = n1480 & ~n17268 ;
  assign n17270 = n1484 & ~n17269 ;
  assign n17271 = n1488 & ~n17270 ;
  assign n17272 = n1492 & ~n17271 ;
  assign n17273 = n1496 & ~n17272 ;
  assign n17274 = n1500 & ~n17273 ;
  assign n17275 = ~x215 & ~n1502 ;
  assign n17276 = ~n17274 & n17275 ;
  assign n17279 = ~n17276 & ~x343 ;
  assign n17280 = ~n17278 & ~n17279 ;
  assign n17281 = n1172 & ~n1848 ;
  assign n17282 = n1177 & ~n17281 ;
  assign n17283 = n1181 & ~n17282 ;
  assign n17284 = n1185 & ~n17283 ;
  assign n17285 = n1189 & ~n17284 ;
  assign n17286 = n1193 & ~n17285 ;
  assign n17287 = n1197 & ~n17286 ;
  assign n17288 = n1201 & ~n17287 ;
  assign n17289 = n1205 & ~n17288 ;
  assign n17290 = n1209 & ~n17289 ;
  assign n17291 = n1213 & ~n17290 ;
  assign n17292 = n1217 & ~n17291 ;
  assign n17293 = n1221 & ~n17292 ;
  assign n17294 = n1225 & ~n17293 ;
  assign n17295 = n1229 & ~n17294 ;
  assign n17296 = n1233 & ~n17295 ;
  assign n17297 = n1237 & ~n17296 ;
  assign n17298 = n1241 & ~n17297 ;
  assign n17299 = n1245 & ~n17298 ;
  assign n17300 = n1249 & ~n17299 ;
  assign n17301 = n1253 & ~n17300 ;
  assign n17302 = n1257 & ~n17301 ;
  assign n17303 = n1261 & ~n17302 ;
  assign n17304 = n1265 & ~n17303 ;
  assign n17305 = n1269 & ~n17304 ;
  assign n17306 = n1273 & ~n17305 ;
  assign n17307 = n2566 & ~n17306 ;
  assign n17308 = n2568 & ~n17307 ;
  assign n17309 = n3105 & ~n17308 ;
  assign n17310 = n1625 & ~n17309 ;
  assign n17311 = n1629 & ~n17310 ;
  assign n17312 = n1633 & ~n17311 ;
  assign n17313 = n1637 & ~n17312 ;
  assign n17314 = n1641 & ~n17313 ;
  assign n17315 = n1645 & ~n17314 ;
  assign n17316 = n1649 & ~n17315 ;
  assign n17317 = n1653 & ~n17316 ;
  assign n17318 = n1657 & ~n17317 ;
  assign n17319 = n1661 & ~n17318 ;
  assign n17320 = n1665 & ~n17319 ;
  assign n17321 = n1669 & ~n17320 ;
  assign n17322 = n1673 & ~n17321 ;
  assign n17323 = n1677 & ~n17322 ;
  assign n17324 = n1681 & ~n17323 ;
  assign n17325 = n1685 & ~n17324 ;
  assign n17326 = n1689 & ~n17325 ;
  assign n17327 = n1693 & ~n17326 ;
  assign n17328 = n1697 & ~n17327 ;
  assign n17329 = n1701 & ~n17328 ;
  assign n17330 = n1705 & ~n17329 ;
  assign n17331 = n1709 & ~n17330 ;
  assign n17332 = n1713 & ~n17331 ;
  assign n17333 = n1717 & ~n17332 ;
  assign n17334 = n1721 & ~n17333 ;
  assign n17335 = n1725 & ~n17334 ;
  assign n17336 = n1729 & ~n17335 ;
  assign n17337 = n1733 & ~n17336 ;
  assign n17338 = n1737 & ~n17337 ;
  assign n17339 = n1741 & ~n17338 ;
  assign n17340 = n1745 & ~n17339 ;
  assign n17341 = n1749 & ~n17340 ;
  assign n17342 = n1753 & ~n17341 ;
  assign n17343 = n1757 & ~n17342 ;
  assign n17344 = n1761 & ~n17343 ;
  assign n17345 = n1765 & ~n17344 ;
  assign n17346 = n1769 & ~n17345 ;
  assign n17347 = n1773 & ~n17346 ;
  assign n17348 = n1777 & ~n17347 ;
  assign n17349 = n1781 & ~n17348 ;
  assign n17350 = n1785 & ~n17349 ;
  assign n17351 = n1789 & ~n17350 ;
  assign n17352 = n1793 & ~n17351 ;
  assign n17353 = n1797 & ~n17352 ;
  assign n17354 = n1801 & ~n17353 ;
  assign n17355 = n1805 & ~n17354 ;
  assign n17356 = n1809 & ~n17355 ;
  assign n17357 = n1813 & ~n17356 ;
  assign n17358 = n1817 & ~n17357 ;
  assign n17359 = n1821 & ~n17358 ;
  assign n17360 = n1825 & ~n17359 ;
  assign n17361 = n1829 & ~n17360 ;
  assign n17362 = n1833 & ~n17361 ;
  assign n17363 = n1837 & ~n17362 ;
  assign n17364 = n1841 & ~n17363 ;
  assign n17365 = x216 & ~n1843 ;
  assign n17366 = ~n17364 & n17365 ;
  assign n17454 = n17366 & x344 ;
  assign n17367 = n1511 & ~n2185 ;
  assign n17368 = n1516 & ~n17367 ;
  assign n17369 = n1520 & ~n17368 ;
  assign n17370 = n1524 & ~n17369 ;
  assign n17371 = n1528 & ~n17370 ;
  assign n17372 = n1532 & ~n17371 ;
  assign n17373 = n1536 & ~n17372 ;
  assign n17374 = n1540 & ~n17373 ;
  assign n17375 = n1544 & ~n17374 ;
  assign n17376 = n1548 & ~n17375 ;
  assign n17377 = n1552 & ~n17376 ;
  assign n17378 = n1556 & ~n17377 ;
  assign n17379 = n1560 & ~n17378 ;
  assign n17380 = n1564 & ~n17379 ;
  assign n17381 = n1568 & ~n17380 ;
  assign n17382 = n1572 & ~n17381 ;
  assign n17383 = n1576 & ~n17382 ;
  assign n17384 = n1580 & ~n17383 ;
  assign n17385 = n1584 & ~n17384 ;
  assign n17386 = n1588 & ~n17385 ;
  assign n17387 = n1592 & ~n17386 ;
  assign n17388 = n1596 & ~n17387 ;
  assign n17389 = n1600 & ~n17388 ;
  assign n17390 = n1604 & ~n17389 ;
  assign n17391 = n1608 & ~n17390 ;
  assign n17392 = n1612 & ~n17391 ;
  assign n17393 = n2656 & ~n17392 ;
  assign n17394 = n2658 & ~n17393 ;
  assign n17395 = n3192 & ~n17394 ;
  assign n17396 = n1962 & ~n17395 ;
  assign n17397 = n1966 & ~n17396 ;
  assign n17398 = n1970 & ~n17397 ;
  assign n17399 = n1974 & ~n17398 ;
  assign n17400 = n1978 & ~n17399 ;
  assign n17401 = n1982 & ~n17400 ;
  assign n17402 = n1986 & ~n17401 ;
  assign n17403 = n1990 & ~n17402 ;
  assign n17404 = n1994 & ~n17403 ;
  assign n17405 = n1998 & ~n17404 ;
  assign n17406 = n2002 & ~n17405 ;
  assign n17407 = n2006 & ~n17406 ;
  assign n17408 = n2010 & ~n17407 ;
  assign n17409 = n2014 & ~n17408 ;
  assign n17410 = n2018 & ~n17409 ;
  assign n17411 = n2022 & ~n17410 ;
  assign n17412 = n2026 & ~n17411 ;
  assign n17413 = n2030 & ~n17412 ;
  assign n17414 = n2034 & ~n17413 ;
  assign n17415 = n2038 & ~n17414 ;
  assign n17416 = n2042 & ~n17415 ;
  assign n17417 = n2046 & ~n17416 ;
  assign n17418 = n2050 & ~n17417 ;
  assign n17419 = n2054 & ~n17418 ;
  assign n17420 = n2058 & ~n17419 ;
  assign n17421 = n2062 & ~n17420 ;
  assign n17422 = n2066 & ~n17421 ;
  assign n17423 = n2070 & ~n17422 ;
  assign n17424 = n2074 & ~n17423 ;
  assign n17425 = n2078 & ~n17424 ;
  assign n17426 = n2082 & ~n17425 ;
  assign n17427 = n2086 & ~n17426 ;
  assign n17428 = n2090 & ~n17427 ;
  assign n17429 = n2094 & ~n17428 ;
  assign n17430 = n2098 & ~n17429 ;
  assign n17431 = n2102 & ~n17430 ;
  assign n17432 = n2106 & ~n17431 ;
  assign n17433 = n2110 & ~n17432 ;
  assign n17434 = n2114 & ~n17433 ;
  assign n17435 = n2118 & ~n17434 ;
  assign n17436 = n2122 & ~n17435 ;
  assign n17437 = n2126 & ~n17436 ;
  assign n17438 = n2130 & ~n17437 ;
  assign n17439 = n2134 & ~n17438 ;
  assign n17440 = n2138 & ~n17439 ;
  assign n17441 = n2142 & ~n17440 ;
  assign n17442 = n2146 & ~n17441 ;
  assign n17443 = n2150 & ~n17442 ;
  assign n17444 = n2154 & ~n17443 ;
  assign n17445 = n2158 & ~n17444 ;
  assign n17446 = n2162 & ~n17445 ;
  assign n17447 = n2166 & ~n17446 ;
  assign n17448 = n2170 & ~n17447 ;
  assign n17449 = n2174 & ~n17448 ;
  assign n17450 = n2178 & ~n17449 ;
  assign n17451 = ~x216 & ~n2180 ;
  assign n17452 = ~n17450 & n17451 ;
  assign n17455 = ~n17452 & ~x344 ;
  assign n17456 = ~n17454 & ~n17455 ;
  assign n17457 = ~n494 & n1852 ;
  assign n17458 = n1857 & ~n17457 ;
  assign n17459 = n1861 & ~n17458 ;
  assign n17460 = n1865 & ~n17459 ;
  assign n17461 = n1869 & ~n17460 ;
  assign n17462 = n1873 & ~n17461 ;
  assign n17463 = n1877 & ~n17462 ;
  assign n17464 = n1881 & ~n17463 ;
  assign n17465 = n1885 & ~n17464 ;
  assign n17466 = n1889 & ~n17465 ;
  assign n17467 = n1893 & ~n17466 ;
  assign n17468 = n1897 & ~n17467 ;
  assign n17469 = n1901 & ~n17468 ;
  assign n17470 = n1905 & ~n17469 ;
  assign n17471 = n1909 & ~n17470 ;
  assign n17472 = n1913 & ~n17471 ;
  assign n17473 = n1917 & ~n17472 ;
  assign n17474 = n1921 & ~n17473 ;
  assign n17475 = n1925 & ~n17474 ;
  assign n17476 = n1929 & ~n17475 ;
  assign n17477 = n1933 & ~n17476 ;
  assign n17478 = n1937 & ~n17477 ;
  assign n17479 = n1941 & ~n17478 ;
  assign n17480 = n1945 & ~n17479 ;
  assign n17481 = n1949 & ~n17480 ;
  assign n17482 = n1953 & ~n17481 ;
  assign n17483 = n2749 & ~n17482 ;
  assign n17484 = n263 & ~n17483 ;
  assign n17485 = n267 & ~n17484 ;
  assign n17486 = n271 & ~n17485 ;
  assign n17487 = n275 & ~n17486 ;
  assign n17488 = n279 & ~n17487 ;
  assign n17489 = n283 & ~n17488 ;
  assign n17490 = n287 & ~n17489 ;
  assign n17491 = n291 & ~n17490 ;
  assign n17492 = n295 & ~n17491 ;
  assign n17493 = n299 & ~n17492 ;
  assign n17494 = n303 & ~n17493 ;
  assign n17495 = n307 & ~n17494 ;
  assign n17496 = n311 & ~n17495 ;
  assign n17497 = n315 & ~n17496 ;
  assign n17498 = n319 & ~n17497 ;
  assign n17499 = n323 & ~n17498 ;
  assign n17500 = n327 & ~n17499 ;
  assign n17501 = n331 & ~n17500 ;
  assign n17502 = n335 & ~n17501 ;
  assign n17503 = n339 & ~n17502 ;
  assign n17504 = n343 & ~n17503 ;
  assign n17505 = n347 & ~n17504 ;
  assign n17506 = n351 & ~n17505 ;
  assign n17507 = n355 & ~n17506 ;
  assign n17508 = n359 & ~n17507 ;
  assign n17509 = n363 & ~n17508 ;
  assign n17510 = n367 & ~n17509 ;
  assign n17511 = n371 & ~n17510 ;
  assign n17512 = n375 & ~n17511 ;
  assign n17513 = n379 & ~n17512 ;
  assign n17514 = n383 & ~n17513 ;
  assign n17515 = n387 & ~n17514 ;
  assign n17516 = n391 & ~n17515 ;
  assign n17517 = n395 & ~n17516 ;
  assign n17518 = n399 & ~n17517 ;
  assign n17519 = n403 & ~n17518 ;
  assign n17520 = n407 & ~n17519 ;
  assign n17521 = n411 & ~n17520 ;
  assign n17522 = n415 & ~n17521 ;
  assign n17523 = n419 & ~n17522 ;
  assign n17524 = n423 & ~n17523 ;
  assign n17525 = n427 & ~n17524 ;
  assign n17526 = n431 & ~n17525 ;
  assign n17527 = n435 & ~n17526 ;
  assign n17528 = n439 & ~n17527 ;
  assign n17529 = n443 & ~n17528 ;
  assign n17530 = n447 & ~n17529 ;
  assign n17531 = n451 & ~n17530 ;
  assign n17532 = n455 & ~n17531 ;
  assign n17533 = n459 & ~n17532 ;
  assign n17534 = n463 & ~n17533 ;
  assign n17535 = n467 & ~n17534 ;
  assign n17536 = n471 & ~n17535 ;
  assign n17537 = n475 & ~n17536 ;
  assign n17538 = n479 & ~n17537 ;
  assign n17539 = n483 & ~n17538 ;
  assign n17540 = n487 & ~n17539 ;
  assign n17541 = x217 & ~n489 ;
  assign n17542 = ~n17540 & n17541 ;
  assign n17630 = n17542 & x345 ;
  assign n17543 = ~n833 & n2189 ;
  assign n17544 = n2194 & ~n17543 ;
  assign n17545 = n2198 & ~n17544 ;
  assign n17546 = n2202 & ~n17545 ;
  assign n17547 = n2206 & ~n17546 ;
  assign n17548 = n2210 & ~n17547 ;
  assign n17549 = n2214 & ~n17548 ;
  assign n17550 = n2218 & ~n17549 ;
  assign n17551 = n2222 & ~n17550 ;
  assign n17552 = n2226 & ~n17551 ;
  assign n17553 = n2230 & ~n17552 ;
  assign n17554 = n2234 & ~n17553 ;
  assign n17555 = n2238 & ~n17554 ;
  assign n17556 = n2242 & ~n17555 ;
  assign n17557 = n2246 & ~n17556 ;
  assign n17558 = n2250 & ~n17557 ;
  assign n17559 = n2254 & ~n17558 ;
  assign n17560 = n2258 & ~n17559 ;
  assign n17561 = n2262 & ~n17560 ;
  assign n17562 = n2266 & ~n17561 ;
  assign n17563 = n2270 & ~n17562 ;
  assign n17564 = n2274 & ~n17563 ;
  assign n17565 = n2278 & ~n17564 ;
  assign n17566 = n2282 & ~n17565 ;
  assign n17567 = n2286 & ~n17566 ;
  assign n17568 = n2290 & ~n17567 ;
  assign n17569 = n2836 & ~n17568 ;
  assign n17570 = n602 & ~n17569 ;
  assign n17571 = n606 & ~n17570 ;
  assign n17572 = n610 & ~n17571 ;
  assign n17573 = n614 & ~n17572 ;
  assign n17574 = n618 & ~n17573 ;
  assign n17575 = n622 & ~n17574 ;
  assign n17576 = n626 & ~n17575 ;
  assign n17577 = n630 & ~n17576 ;
  assign n17578 = n634 & ~n17577 ;
  assign n17579 = n638 & ~n17578 ;
  assign n17580 = n642 & ~n17579 ;
  assign n17581 = n646 & ~n17580 ;
  assign n17582 = n650 & ~n17581 ;
  assign n17583 = n654 & ~n17582 ;
  assign n17584 = n658 & ~n17583 ;
  assign n17585 = n662 & ~n17584 ;
  assign n17586 = n666 & ~n17585 ;
  assign n17587 = n670 & ~n17586 ;
  assign n17588 = n674 & ~n17587 ;
  assign n17589 = n678 & ~n17588 ;
  assign n17590 = n682 & ~n17589 ;
  assign n17591 = n686 & ~n17590 ;
  assign n17592 = n690 & ~n17591 ;
  assign n17593 = n694 & ~n17592 ;
  assign n17594 = n698 & ~n17593 ;
  assign n17595 = n702 & ~n17594 ;
  assign n17596 = n706 & ~n17595 ;
  assign n17597 = n710 & ~n17596 ;
  assign n17598 = n714 & ~n17597 ;
  assign n17599 = n718 & ~n17598 ;
  assign n17600 = n722 & ~n17599 ;
  assign n17601 = n726 & ~n17600 ;
  assign n17602 = n730 & ~n17601 ;
  assign n17603 = n734 & ~n17602 ;
  assign n17604 = n738 & ~n17603 ;
  assign n17605 = n742 & ~n17604 ;
  assign n17606 = n746 & ~n17605 ;
  assign n17607 = n750 & ~n17606 ;
  assign n17608 = n754 & ~n17607 ;
  assign n17609 = n758 & ~n17608 ;
  assign n17610 = n762 & ~n17609 ;
  assign n17611 = n766 & ~n17610 ;
  assign n17612 = n770 & ~n17611 ;
  assign n17613 = n774 & ~n17612 ;
  assign n17614 = n778 & ~n17613 ;
  assign n17615 = n782 & ~n17614 ;
  assign n17616 = n786 & ~n17615 ;
  assign n17617 = n790 & ~n17616 ;
  assign n17618 = n794 & ~n17617 ;
  assign n17619 = n798 & ~n17618 ;
  assign n17620 = n802 & ~n17619 ;
  assign n17621 = n806 & ~n17620 ;
  assign n17622 = n810 & ~n17621 ;
  assign n17623 = n814 & ~n17622 ;
  assign n17624 = n818 & ~n17623 ;
  assign n17625 = n822 & ~n17624 ;
  assign n17626 = n826 & ~n17625 ;
  assign n17627 = ~x217 & ~n828 ;
  assign n17628 = ~n17626 & n17627 ;
  assign n17631 = ~n17628 & ~x345 ;
  assign n17632 = ~n17630 & ~n17631 ;
  assign n17633 = n498 & ~n1176 ;
  assign n17634 = n503 & ~n17633 ;
  assign n17635 = n507 & ~n17634 ;
  assign n17636 = n511 & ~n17635 ;
  assign n17637 = n515 & ~n17636 ;
  assign n17638 = n519 & ~n17637 ;
  assign n17639 = n523 & ~n17638 ;
  assign n17640 = n527 & ~n17639 ;
  assign n17641 = n531 & ~n17640 ;
  assign n17642 = n535 & ~n17641 ;
  assign n17643 = n539 & ~n17642 ;
  assign n17644 = n543 & ~n17643 ;
  assign n17645 = n547 & ~n17644 ;
  assign n17646 = n551 & ~n17645 ;
  assign n17647 = n555 & ~n17646 ;
  assign n17648 = n559 & ~n17647 ;
  assign n17649 = n563 & ~n17648 ;
  assign n17650 = n567 & ~n17649 ;
  assign n17651 = n571 & ~n17650 ;
  assign n17652 = n575 & ~n17651 ;
  assign n17653 = n579 & ~n17652 ;
  assign n17654 = n583 & ~n17653 ;
  assign n17655 = n587 & ~n17654 ;
  assign n17656 = n591 & ~n17655 ;
  assign n17657 = n2382 & ~n17656 ;
  assign n17658 = n2384 & ~n17657 ;
  assign n17659 = n2927 & ~n17658 ;
  assign n17660 = n945 & ~n17659 ;
  assign n17661 = n949 & ~n17660 ;
  assign n17662 = n953 & ~n17661 ;
  assign n17663 = n957 & ~n17662 ;
  assign n17664 = n961 & ~n17663 ;
  assign n17665 = n965 & ~n17664 ;
  assign n17666 = n969 & ~n17665 ;
  assign n17667 = n973 & ~n17666 ;
  assign n17668 = n977 & ~n17667 ;
  assign n17669 = n981 & ~n17668 ;
  assign n17670 = n985 & ~n17669 ;
  assign n17671 = n989 & ~n17670 ;
  assign n17672 = n993 & ~n17671 ;
  assign n17673 = n997 & ~n17672 ;
  assign n17674 = n1001 & ~n17673 ;
  assign n17675 = n1005 & ~n17674 ;
  assign n17676 = n1009 & ~n17675 ;
  assign n17677 = n1013 & ~n17676 ;
  assign n17678 = n1017 & ~n17677 ;
  assign n17679 = n1021 & ~n17678 ;
  assign n17680 = n1025 & ~n17679 ;
  assign n17681 = n1029 & ~n17680 ;
  assign n17682 = n1033 & ~n17681 ;
  assign n17683 = n1037 & ~n17682 ;
  assign n17684 = n1041 & ~n17683 ;
  assign n17685 = n1045 & ~n17684 ;
  assign n17686 = n1049 & ~n17685 ;
  assign n17687 = n1053 & ~n17686 ;
  assign n17688 = n1057 & ~n17687 ;
  assign n17689 = n1061 & ~n17688 ;
  assign n17690 = n1065 & ~n17689 ;
  assign n17691 = n1069 & ~n17690 ;
  assign n17692 = n1073 & ~n17691 ;
  assign n17693 = n1077 & ~n17692 ;
  assign n17694 = n1081 & ~n17693 ;
  assign n17695 = n1085 & ~n17694 ;
  assign n17696 = n1089 & ~n17695 ;
  assign n17697 = n1093 & ~n17696 ;
  assign n17698 = n1097 & ~n17697 ;
  assign n17699 = n1101 & ~n17698 ;
  assign n17700 = n1105 & ~n17699 ;
  assign n17701 = n1109 & ~n17700 ;
  assign n17702 = n1113 & ~n17701 ;
  assign n17703 = n1117 & ~n17702 ;
  assign n17704 = n1121 & ~n17703 ;
  assign n17705 = n1125 & ~n17704 ;
  assign n17706 = n1129 & ~n17705 ;
  assign n17707 = n1133 & ~n17706 ;
  assign n17708 = n1137 & ~n17707 ;
  assign n17709 = n1141 & ~n17708 ;
  assign n17710 = n1145 & ~n17709 ;
  assign n17711 = n1149 & ~n17710 ;
  assign n17712 = n1153 & ~n17711 ;
  assign n17713 = n1157 & ~n17712 ;
  assign n17714 = n1161 & ~n17713 ;
  assign n17715 = n1165 & ~n17714 ;
  assign n17716 = n1169 & ~n17715 ;
  assign n17717 = x218 & ~n1171 ;
  assign n17718 = ~n17716 & n17717 ;
  assign n17806 = n17718 & x346 ;
  assign n17719 = n837 & ~n1515 ;
  assign n17720 = n842 & ~n17719 ;
  assign n17721 = n846 & ~n17720 ;
  assign n17722 = n850 & ~n17721 ;
  assign n17723 = n854 & ~n17722 ;
  assign n17724 = n858 & ~n17723 ;
  assign n17725 = n862 & ~n17724 ;
  assign n17726 = n866 & ~n17725 ;
  assign n17727 = n870 & ~n17726 ;
  assign n17728 = n874 & ~n17727 ;
  assign n17729 = n878 & ~n17728 ;
  assign n17730 = n882 & ~n17729 ;
  assign n17731 = n886 & ~n17730 ;
  assign n17732 = n890 & ~n17731 ;
  assign n17733 = n894 & ~n17732 ;
  assign n17734 = n898 & ~n17733 ;
  assign n17735 = n902 & ~n17734 ;
  assign n17736 = n906 & ~n17735 ;
  assign n17737 = n910 & ~n17736 ;
  assign n17738 = n914 & ~n17737 ;
  assign n17739 = n918 & ~n17738 ;
  assign n17740 = n922 & ~n17739 ;
  assign n17741 = n926 & ~n17740 ;
  assign n17742 = n930 & ~n17741 ;
  assign n17743 = n2472 & ~n17742 ;
  assign n17744 = n2474 & ~n17743 ;
  assign n17745 = n3014 & ~n17744 ;
  assign n17746 = n1284 & ~n17745 ;
  assign n17747 = n1288 & ~n17746 ;
  assign n17748 = n1292 & ~n17747 ;
  assign n17749 = n1296 & ~n17748 ;
  assign n17750 = n1300 & ~n17749 ;
  assign n17751 = n1304 & ~n17750 ;
  assign n17752 = n1308 & ~n17751 ;
  assign n17753 = n1312 & ~n17752 ;
  assign n17754 = n1316 & ~n17753 ;
  assign n17755 = n1320 & ~n17754 ;
  assign n17756 = n1324 & ~n17755 ;
  assign n17757 = n1328 & ~n17756 ;
  assign n17758 = n1332 & ~n17757 ;
  assign n17759 = n1336 & ~n17758 ;
  assign n17760 = n1340 & ~n17759 ;
  assign n17761 = n1344 & ~n17760 ;
  assign n17762 = n1348 & ~n17761 ;
  assign n17763 = n1352 & ~n17762 ;
  assign n17764 = n1356 & ~n17763 ;
  assign n17765 = n1360 & ~n17764 ;
  assign n17766 = n1364 & ~n17765 ;
  assign n17767 = n1368 & ~n17766 ;
  assign n17768 = n1372 & ~n17767 ;
  assign n17769 = n1376 & ~n17768 ;
  assign n17770 = n1380 & ~n17769 ;
  assign n17771 = n1384 & ~n17770 ;
  assign n17772 = n1388 & ~n17771 ;
  assign n17773 = n1392 & ~n17772 ;
  assign n17774 = n1396 & ~n17773 ;
  assign n17775 = n1400 & ~n17774 ;
  assign n17776 = n1404 & ~n17775 ;
  assign n17777 = n1408 & ~n17776 ;
  assign n17778 = n1412 & ~n17777 ;
  assign n17779 = n1416 & ~n17778 ;
  assign n17780 = n1420 & ~n17779 ;
  assign n17781 = n1424 & ~n17780 ;
  assign n17782 = n1428 & ~n17781 ;
  assign n17783 = n1432 & ~n17782 ;
  assign n17784 = n1436 & ~n17783 ;
  assign n17785 = n1440 & ~n17784 ;
  assign n17786 = n1444 & ~n17785 ;
  assign n17787 = n1448 & ~n17786 ;
  assign n17788 = n1452 & ~n17787 ;
  assign n17789 = n1456 & ~n17788 ;
  assign n17790 = n1460 & ~n17789 ;
  assign n17791 = n1464 & ~n17790 ;
  assign n17792 = n1468 & ~n17791 ;
  assign n17793 = n1472 & ~n17792 ;
  assign n17794 = n1476 & ~n17793 ;
  assign n17795 = n1480 & ~n17794 ;
  assign n17796 = n1484 & ~n17795 ;
  assign n17797 = n1488 & ~n17796 ;
  assign n17798 = n1492 & ~n17797 ;
  assign n17799 = n1496 & ~n17798 ;
  assign n17800 = n1500 & ~n17799 ;
  assign n17801 = n1504 & ~n17800 ;
  assign n17802 = n1508 & ~n17801 ;
  assign n17803 = ~x218 & ~n1510 ;
  assign n17804 = ~n17802 & n17803 ;
  assign n17807 = ~n17804 & ~x346 ;
  assign n17808 = ~n17806 & ~n17807 ;
  assign n17809 = n1180 & ~n1856 ;
  assign n17810 = n1185 & ~n17809 ;
  assign n17811 = n1189 & ~n17810 ;
  assign n17812 = n1193 & ~n17811 ;
  assign n17813 = n1197 & ~n17812 ;
  assign n17814 = n1201 & ~n17813 ;
  assign n17815 = n1205 & ~n17814 ;
  assign n17816 = n1209 & ~n17815 ;
  assign n17817 = n1213 & ~n17816 ;
  assign n17818 = n1217 & ~n17817 ;
  assign n17819 = n1221 & ~n17818 ;
  assign n17820 = n1225 & ~n17819 ;
  assign n17821 = n1229 & ~n17820 ;
  assign n17822 = n1233 & ~n17821 ;
  assign n17823 = n1237 & ~n17822 ;
  assign n17824 = n1241 & ~n17823 ;
  assign n17825 = n1245 & ~n17824 ;
  assign n17826 = n1249 & ~n17825 ;
  assign n17827 = n1253 & ~n17826 ;
  assign n17828 = n1257 & ~n17827 ;
  assign n17829 = n1261 & ~n17828 ;
  assign n17830 = n1265 & ~n17829 ;
  assign n17831 = n1269 & ~n17830 ;
  assign n17832 = n1273 & ~n17831 ;
  assign n17833 = n2566 & ~n17832 ;
  assign n17834 = n2568 & ~n17833 ;
  assign n17835 = n3105 & ~n17834 ;
  assign n17836 = n1625 & ~n17835 ;
  assign n17837 = n1629 & ~n17836 ;
  assign n17838 = n1633 & ~n17837 ;
  assign n17839 = n1637 & ~n17838 ;
  assign n17840 = n1641 & ~n17839 ;
  assign n17841 = n1645 & ~n17840 ;
  assign n17842 = n1649 & ~n17841 ;
  assign n17843 = n1653 & ~n17842 ;
  assign n17844 = n1657 & ~n17843 ;
  assign n17845 = n1661 & ~n17844 ;
  assign n17846 = n1665 & ~n17845 ;
  assign n17847 = n1669 & ~n17846 ;
  assign n17848 = n1673 & ~n17847 ;
  assign n17849 = n1677 & ~n17848 ;
  assign n17850 = n1681 & ~n17849 ;
  assign n17851 = n1685 & ~n17850 ;
  assign n17852 = n1689 & ~n17851 ;
  assign n17853 = n1693 & ~n17852 ;
  assign n17854 = n1697 & ~n17853 ;
  assign n17855 = n1701 & ~n17854 ;
  assign n17856 = n1705 & ~n17855 ;
  assign n17857 = n1709 & ~n17856 ;
  assign n17858 = n1713 & ~n17857 ;
  assign n17859 = n1717 & ~n17858 ;
  assign n17860 = n1721 & ~n17859 ;
  assign n17861 = n1725 & ~n17860 ;
  assign n17862 = n1729 & ~n17861 ;
  assign n17863 = n1733 & ~n17862 ;
  assign n17864 = n1737 & ~n17863 ;
  assign n17865 = n1741 & ~n17864 ;
  assign n17866 = n1745 & ~n17865 ;
  assign n17867 = n1749 & ~n17866 ;
  assign n17868 = n1753 & ~n17867 ;
  assign n17869 = n1757 & ~n17868 ;
  assign n17870 = n1761 & ~n17869 ;
  assign n17871 = n1765 & ~n17870 ;
  assign n17872 = n1769 & ~n17871 ;
  assign n17873 = n1773 & ~n17872 ;
  assign n17874 = n1777 & ~n17873 ;
  assign n17875 = n1781 & ~n17874 ;
  assign n17876 = n1785 & ~n17875 ;
  assign n17877 = n1789 & ~n17876 ;
  assign n17878 = n1793 & ~n17877 ;
  assign n17879 = n1797 & ~n17878 ;
  assign n17880 = n1801 & ~n17879 ;
  assign n17881 = n1805 & ~n17880 ;
  assign n17882 = n1809 & ~n17881 ;
  assign n17883 = n1813 & ~n17882 ;
  assign n17884 = n1817 & ~n17883 ;
  assign n17885 = n1821 & ~n17884 ;
  assign n17886 = n1825 & ~n17885 ;
  assign n17887 = n1829 & ~n17886 ;
  assign n17888 = n1833 & ~n17887 ;
  assign n17889 = n1837 & ~n17888 ;
  assign n17890 = n1841 & ~n17889 ;
  assign n17891 = n1845 & ~n17890 ;
  assign n17892 = n1849 & ~n17891 ;
  assign n17893 = x219 & ~n1851 ;
  assign n17894 = ~n17892 & n17893 ;
  assign n17982 = n17894 & x347 ;
  assign n17895 = n1519 & ~n2193 ;
  assign n17896 = n1524 & ~n17895 ;
  assign n17897 = n1528 & ~n17896 ;
  assign n17898 = n1532 & ~n17897 ;
  assign n17899 = n1536 & ~n17898 ;
  assign n17900 = n1540 & ~n17899 ;
  assign n17901 = n1544 & ~n17900 ;
  assign n17902 = n1548 & ~n17901 ;
  assign n17903 = n1552 & ~n17902 ;
  assign n17904 = n1556 & ~n17903 ;
  assign n17905 = n1560 & ~n17904 ;
  assign n17906 = n1564 & ~n17905 ;
  assign n17907 = n1568 & ~n17906 ;
  assign n17908 = n1572 & ~n17907 ;
  assign n17909 = n1576 & ~n17908 ;
  assign n17910 = n1580 & ~n17909 ;
  assign n17911 = n1584 & ~n17910 ;
  assign n17912 = n1588 & ~n17911 ;
  assign n17913 = n1592 & ~n17912 ;
  assign n17914 = n1596 & ~n17913 ;
  assign n17915 = n1600 & ~n17914 ;
  assign n17916 = n1604 & ~n17915 ;
  assign n17917 = n1608 & ~n17916 ;
  assign n17918 = n1612 & ~n17917 ;
  assign n17919 = n2656 & ~n17918 ;
  assign n17920 = n2658 & ~n17919 ;
  assign n17921 = n3192 & ~n17920 ;
  assign n17922 = n1962 & ~n17921 ;
  assign n17923 = n1966 & ~n17922 ;
  assign n17924 = n1970 & ~n17923 ;
  assign n17925 = n1974 & ~n17924 ;
  assign n17926 = n1978 & ~n17925 ;
  assign n17927 = n1982 & ~n17926 ;
  assign n17928 = n1986 & ~n17927 ;
  assign n17929 = n1990 & ~n17928 ;
  assign n17930 = n1994 & ~n17929 ;
  assign n17931 = n1998 & ~n17930 ;
  assign n17932 = n2002 & ~n17931 ;
  assign n17933 = n2006 & ~n17932 ;
  assign n17934 = n2010 & ~n17933 ;
  assign n17935 = n2014 & ~n17934 ;
  assign n17936 = n2018 & ~n17935 ;
  assign n17937 = n2022 & ~n17936 ;
  assign n17938 = n2026 & ~n17937 ;
  assign n17939 = n2030 & ~n17938 ;
  assign n17940 = n2034 & ~n17939 ;
  assign n17941 = n2038 & ~n17940 ;
  assign n17942 = n2042 & ~n17941 ;
  assign n17943 = n2046 & ~n17942 ;
  assign n17944 = n2050 & ~n17943 ;
  assign n17945 = n2054 & ~n17944 ;
  assign n17946 = n2058 & ~n17945 ;
  assign n17947 = n2062 & ~n17946 ;
  assign n17948 = n2066 & ~n17947 ;
  assign n17949 = n2070 & ~n17948 ;
  assign n17950 = n2074 & ~n17949 ;
  assign n17951 = n2078 & ~n17950 ;
  assign n17952 = n2082 & ~n17951 ;
  assign n17953 = n2086 & ~n17952 ;
  assign n17954 = n2090 & ~n17953 ;
  assign n17955 = n2094 & ~n17954 ;
  assign n17956 = n2098 & ~n17955 ;
  assign n17957 = n2102 & ~n17956 ;
  assign n17958 = n2106 & ~n17957 ;
  assign n17959 = n2110 & ~n17958 ;
  assign n17960 = n2114 & ~n17959 ;
  assign n17961 = n2118 & ~n17960 ;
  assign n17962 = n2122 & ~n17961 ;
  assign n17963 = n2126 & ~n17962 ;
  assign n17964 = n2130 & ~n17963 ;
  assign n17965 = n2134 & ~n17964 ;
  assign n17966 = n2138 & ~n17965 ;
  assign n17967 = n2142 & ~n17966 ;
  assign n17968 = n2146 & ~n17967 ;
  assign n17969 = n2150 & ~n17968 ;
  assign n17970 = n2154 & ~n17969 ;
  assign n17971 = n2158 & ~n17970 ;
  assign n17972 = n2162 & ~n17971 ;
  assign n17973 = n2166 & ~n17972 ;
  assign n17974 = n2170 & ~n17973 ;
  assign n17975 = n2174 & ~n17974 ;
  assign n17976 = n2178 & ~n17975 ;
  assign n17977 = n2182 & ~n17976 ;
  assign n17978 = n2186 & ~n17977 ;
  assign n17979 = ~x219 & ~n2188 ;
  assign n17980 = ~n17978 & n17979 ;
  assign n17983 = ~n17980 & ~x347 ;
  assign n17984 = ~n17982 & ~n17983 ;
  assign n17985 = ~n502 & n1860 ;
  assign n17986 = n1865 & ~n17985 ;
  assign n17987 = n1869 & ~n17986 ;
  assign n17988 = n1873 & ~n17987 ;
  assign n17989 = n1877 & ~n17988 ;
  assign n17990 = n1881 & ~n17989 ;
  assign n17991 = n1885 & ~n17990 ;
  assign n17992 = n1889 & ~n17991 ;
  assign n17993 = n1893 & ~n17992 ;
  assign n17994 = n1897 & ~n17993 ;
  assign n17995 = n1901 & ~n17994 ;
  assign n17996 = n1905 & ~n17995 ;
  assign n17997 = n1909 & ~n17996 ;
  assign n17998 = n1913 & ~n17997 ;
  assign n17999 = n1917 & ~n17998 ;
  assign n18000 = n1921 & ~n17999 ;
  assign n18001 = n1925 & ~n18000 ;
  assign n18002 = n1929 & ~n18001 ;
  assign n18003 = n1933 & ~n18002 ;
  assign n18004 = n1937 & ~n18003 ;
  assign n18005 = n1941 & ~n18004 ;
  assign n18006 = n1945 & ~n18005 ;
  assign n18007 = n1949 & ~n18006 ;
  assign n18008 = n1953 & ~n18007 ;
  assign n18009 = n2749 & ~n18008 ;
  assign n18010 = n263 & ~n18009 ;
  assign n18011 = n267 & ~n18010 ;
  assign n18012 = n271 & ~n18011 ;
  assign n18013 = n275 & ~n18012 ;
  assign n18014 = n279 & ~n18013 ;
  assign n18015 = n283 & ~n18014 ;
  assign n18016 = n287 & ~n18015 ;
  assign n18017 = n291 & ~n18016 ;
  assign n18018 = n295 & ~n18017 ;
  assign n18019 = n299 & ~n18018 ;
  assign n18020 = n303 & ~n18019 ;
  assign n18021 = n307 & ~n18020 ;
  assign n18022 = n311 & ~n18021 ;
  assign n18023 = n315 & ~n18022 ;
  assign n18024 = n319 & ~n18023 ;
  assign n18025 = n323 & ~n18024 ;
  assign n18026 = n327 & ~n18025 ;
  assign n18027 = n331 & ~n18026 ;
  assign n18028 = n335 & ~n18027 ;
  assign n18029 = n339 & ~n18028 ;
  assign n18030 = n343 & ~n18029 ;
  assign n18031 = n347 & ~n18030 ;
  assign n18032 = n351 & ~n18031 ;
  assign n18033 = n355 & ~n18032 ;
  assign n18034 = n359 & ~n18033 ;
  assign n18035 = n363 & ~n18034 ;
  assign n18036 = n367 & ~n18035 ;
  assign n18037 = n371 & ~n18036 ;
  assign n18038 = n375 & ~n18037 ;
  assign n18039 = n379 & ~n18038 ;
  assign n18040 = n383 & ~n18039 ;
  assign n18041 = n387 & ~n18040 ;
  assign n18042 = n391 & ~n18041 ;
  assign n18043 = n395 & ~n18042 ;
  assign n18044 = n399 & ~n18043 ;
  assign n18045 = n403 & ~n18044 ;
  assign n18046 = n407 & ~n18045 ;
  assign n18047 = n411 & ~n18046 ;
  assign n18048 = n415 & ~n18047 ;
  assign n18049 = n419 & ~n18048 ;
  assign n18050 = n423 & ~n18049 ;
  assign n18051 = n427 & ~n18050 ;
  assign n18052 = n431 & ~n18051 ;
  assign n18053 = n435 & ~n18052 ;
  assign n18054 = n439 & ~n18053 ;
  assign n18055 = n443 & ~n18054 ;
  assign n18056 = n447 & ~n18055 ;
  assign n18057 = n451 & ~n18056 ;
  assign n18058 = n455 & ~n18057 ;
  assign n18059 = n459 & ~n18058 ;
  assign n18060 = n463 & ~n18059 ;
  assign n18061 = n467 & ~n18060 ;
  assign n18062 = n471 & ~n18061 ;
  assign n18063 = n475 & ~n18062 ;
  assign n18064 = n479 & ~n18063 ;
  assign n18065 = n483 & ~n18064 ;
  assign n18066 = n487 & ~n18065 ;
  assign n18067 = n491 & ~n18066 ;
  assign n18068 = n495 & ~n18067 ;
  assign n18069 = x220 & ~n497 ;
  assign n18070 = ~n18068 & n18069 ;
  assign n18158 = n18070 & x348 ;
  assign n18071 = ~n841 & n2197 ;
  assign n18072 = n2202 & ~n18071 ;
  assign n18073 = n2206 & ~n18072 ;
  assign n18074 = n2210 & ~n18073 ;
  assign n18075 = n2214 & ~n18074 ;
  assign n18076 = n2218 & ~n18075 ;
  assign n18077 = n2222 & ~n18076 ;
  assign n18078 = n2226 & ~n18077 ;
  assign n18079 = n2230 & ~n18078 ;
  assign n18080 = n2234 & ~n18079 ;
  assign n18081 = n2238 & ~n18080 ;
  assign n18082 = n2242 & ~n18081 ;
  assign n18083 = n2246 & ~n18082 ;
  assign n18084 = n2250 & ~n18083 ;
  assign n18085 = n2254 & ~n18084 ;
  assign n18086 = n2258 & ~n18085 ;
  assign n18087 = n2262 & ~n18086 ;
  assign n18088 = n2266 & ~n18087 ;
  assign n18089 = n2270 & ~n18088 ;
  assign n18090 = n2274 & ~n18089 ;
  assign n18091 = n2278 & ~n18090 ;
  assign n18092 = n2282 & ~n18091 ;
  assign n18093 = n2286 & ~n18092 ;
  assign n18094 = n2290 & ~n18093 ;
  assign n18095 = n2836 & ~n18094 ;
  assign n18096 = n602 & ~n18095 ;
  assign n18097 = n606 & ~n18096 ;
  assign n18098 = n610 & ~n18097 ;
  assign n18099 = n614 & ~n18098 ;
  assign n18100 = n618 & ~n18099 ;
  assign n18101 = n622 & ~n18100 ;
  assign n18102 = n626 & ~n18101 ;
  assign n18103 = n630 & ~n18102 ;
  assign n18104 = n634 & ~n18103 ;
  assign n18105 = n638 & ~n18104 ;
  assign n18106 = n642 & ~n18105 ;
  assign n18107 = n646 & ~n18106 ;
  assign n18108 = n650 & ~n18107 ;
  assign n18109 = n654 & ~n18108 ;
  assign n18110 = n658 & ~n18109 ;
  assign n18111 = n662 & ~n18110 ;
  assign n18112 = n666 & ~n18111 ;
  assign n18113 = n670 & ~n18112 ;
  assign n18114 = n674 & ~n18113 ;
  assign n18115 = n678 & ~n18114 ;
  assign n18116 = n682 & ~n18115 ;
  assign n18117 = n686 & ~n18116 ;
  assign n18118 = n690 & ~n18117 ;
  assign n18119 = n694 & ~n18118 ;
  assign n18120 = n698 & ~n18119 ;
  assign n18121 = n702 & ~n18120 ;
  assign n18122 = n706 & ~n18121 ;
  assign n18123 = n710 & ~n18122 ;
  assign n18124 = n714 & ~n18123 ;
  assign n18125 = n718 & ~n18124 ;
  assign n18126 = n722 & ~n18125 ;
  assign n18127 = n726 & ~n18126 ;
  assign n18128 = n730 & ~n18127 ;
  assign n18129 = n734 & ~n18128 ;
  assign n18130 = n738 & ~n18129 ;
  assign n18131 = n742 & ~n18130 ;
  assign n18132 = n746 & ~n18131 ;
  assign n18133 = n750 & ~n18132 ;
  assign n18134 = n754 & ~n18133 ;
  assign n18135 = n758 & ~n18134 ;
  assign n18136 = n762 & ~n18135 ;
  assign n18137 = n766 & ~n18136 ;
  assign n18138 = n770 & ~n18137 ;
  assign n18139 = n774 & ~n18138 ;
  assign n18140 = n778 & ~n18139 ;
  assign n18141 = n782 & ~n18140 ;
  assign n18142 = n786 & ~n18141 ;
  assign n18143 = n790 & ~n18142 ;
  assign n18144 = n794 & ~n18143 ;
  assign n18145 = n798 & ~n18144 ;
  assign n18146 = n802 & ~n18145 ;
  assign n18147 = n806 & ~n18146 ;
  assign n18148 = n810 & ~n18147 ;
  assign n18149 = n814 & ~n18148 ;
  assign n18150 = n818 & ~n18149 ;
  assign n18151 = n822 & ~n18150 ;
  assign n18152 = n826 & ~n18151 ;
  assign n18153 = n830 & ~n18152 ;
  assign n18154 = n834 & ~n18153 ;
  assign n18155 = ~x220 & ~n836 ;
  assign n18156 = ~n18154 & n18155 ;
  assign n18159 = ~n18156 & ~x348 ;
  assign n18160 = ~n18158 & ~n18159 ;
  assign n18161 = n506 & ~n1184 ;
  assign n18162 = n511 & ~n18161 ;
  assign n18163 = n515 & ~n18162 ;
  assign n18164 = n519 & ~n18163 ;
  assign n18165 = n523 & ~n18164 ;
  assign n18166 = n527 & ~n18165 ;
  assign n18167 = n531 & ~n18166 ;
  assign n18168 = n535 & ~n18167 ;
  assign n18169 = n539 & ~n18168 ;
  assign n18170 = n543 & ~n18169 ;
  assign n18171 = n547 & ~n18170 ;
  assign n18172 = n551 & ~n18171 ;
  assign n18173 = n555 & ~n18172 ;
  assign n18174 = n559 & ~n18173 ;
  assign n18175 = n563 & ~n18174 ;
  assign n18176 = n567 & ~n18175 ;
  assign n18177 = n571 & ~n18176 ;
  assign n18178 = n575 & ~n18177 ;
  assign n18179 = n579 & ~n18178 ;
  assign n18180 = n583 & ~n18179 ;
  assign n18181 = n587 & ~n18180 ;
  assign n18182 = n591 & ~n18181 ;
  assign n18183 = n2382 & ~n18182 ;
  assign n18184 = n2384 & ~n18183 ;
  assign n18185 = n2927 & ~n18184 ;
  assign n18186 = n945 & ~n18185 ;
  assign n18187 = n949 & ~n18186 ;
  assign n18188 = n953 & ~n18187 ;
  assign n18189 = n957 & ~n18188 ;
  assign n18190 = n961 & ~n18189 ;
  assign n18191 = n965 & ~n18190 ;
  assign n18192 = n969 & ~n18191 ;
  assign n18193 = n973 & ~n18192 ;
  assign n18194 = n977 & ~n18193 ;
  assign n18195 = n981 & ~n18194 ;
  assign n18196 = n985 & ~n18195 ;
  assign n18197 = n989 & ~n18196 ;
  assign n18198 = n993 & ~n18197 ;
  assign n18199 = n997 & ~n18198 ;
  assign n18200 = n1001 & ~n18199 ;
  assign n18201 = n1005 & ~n18200 ;
  assign n18202 = n1009 & ~n18201 ;
  assign n18203 = n1013 & ~n18202 ;
  assign n18204 = n1017 & ~n18203 ;
  assign n18205 = n1021 & ~n18204 ;
  assign n18206 = n1025 & ~n18205 ;
  assign n18207 = n1029 & ~n18206 ;
  assign n18208 = n1033 & ~n18207 ;
  assign n18209 = n1037 & ~n18208 ;
  assign n18210 = n1041 & ~n18209 ;
  assign n18211 = n1045 & ~n18210 ;
  assign n18212 = n1049 & ~n18211 ;
  assign n18213 = n1053 & ~n18212 ;
  assign n18214 = n1057 & ~n18213 ;
  assign n18215 = n1061 & ~n18214 ;
  assign n18216 = n1065 & ~n18215 ;
  assign n18217 = n1069 & ~n18216 ;
  assign n18218 = n1073 & ~n18217 ;
  assign n18219 = n1077 & ~n18218 ;
  assign n18220 = n1081 & ~n18219 ;
  assign n18221 = n1085 & ~n18220 ;
  assign n18222 = n1089 & ~n18221 ;
  assign n18223 = n1093 & ~n18222 ;
  assign n18224 = n1097 & ~n18223 ;
  assign n18225 = n1101 & ~n18224 ;
  assign n18226 = n1105 & ~n18225 ;
  assign n18227 = n1109 & ~n18226 ;
  assign n18228 = n1113 & ~n18227 ;
  assign n18229 = n1117 & ~n18228 ;
  assign n18230 = n1121 & ~n18229 ;
  assign n18231 = n1125 & ~n18230 ;
  assign n18232 = n1129 & ~n18231 ;
  assign n18233 = n1133 & ~n18232 ;
  assign n18234 = n1137 & ~n18233 ;
  assign n18235 = n1141 & ~n18234 ;
  assign n18236 = n1145 & ~n18235 ;
  assign n18237 = n1149 & ~n18236 ;
  assign n18238 = n1153 & ~n18237 ;
  assign n18239 = n1157 & ~n18238 ;
  assign n18240 = n1161 & ~n18239 ;
  assign n18241 = n1165 & ~n18240 ;
  assign n18242 = n1169 & ~n18241 ;
  assign n18243 = n1173 & ~n18242 ;
  assign n18244 = n1177 & ~n18243 ;
  assign n18245 = x221 & ~n1179 ;
  assign n18246 = ~n18244 & n18245 ;
  assign n18334 = n18246 & x349 ;
  assign n18247 = n845 & ~n1523 ;
  assign n18248 = n850 & ~n18247 ;
  assign n18249 = n854 & ~n18248 ;
  assign n18250 = n858 & ~n18249 ;
  assign n18251 = n862 & ~n18250 ;
  assign n18252 = n866 & ~n18251 ;
  assign n18253 = n870 & ~n18252 ;
  assign n18254 = n874 & ~n18253 ;
  assign n18255 = n878 & ~n18254 ;
  assign n18256 = n882 & ~n18255 ;
  assign n18257 = n886 & ~n18256 ;
  assign n18258 = n890 & ~n18257 ;
  assign n18259 = n894 & ~n18258 ;
  assign n18260 = n898 & ~n18259 ;
  assign n18261 = n902 & ~n18260 ;
  assign n18262 = n906 & ~n18261 ;
  assign n18263 = n910 & ~n18262 ;
  assign n18264 = n914 & ~n18263 ;
  assign n18265 = n918 & ~n18264 ;
  assign n18266 = n922 & ~n18265 ;
  assign n18267 = n926 & ~n18266 ;
  assign n18268 = n930 & ~n18267 ;
  assign n18269 = n2472 & ~n18268 ;
  assign n18270 = n2474 & ~n18269 ;
  assign n18271 = n3014 & ~n18270 ;
  assign n18272 = n1284 & ~n18271 ;
  assign n18273 = n1288 & ~n18272 ;
  assign n18274 = n1292 & ~n18273 ;
  assign n18275 = n1296 & ~n18274 ;
  assign n18276 = n1300 & ~n18275 ;
  assign n18277 = n1304 & ~n18276 ;
  assign n18278 = n1308 & ~n18277 ;
  assign n18279 = n1312 & ~n18278 ;
  assign n18280 = n1316 & ~n18279 ;
  assign n18281 = n1320 & ~n18280 ;
  assign n18282 = n1324 & ~n18281 ;
  assign n18283 = n1328 & ~n18282 ;
  assign n18284 = n1332 & ~n18283 ;
  assign n18285 = n1336 & ~n18284 ;
  assign n18286 = n1340 & ~n18285 ;
  assign n18287 = n1344 & ~n18286 ;
  assign n18288 = n1348 & ~n18287 ;
  assign n18289 = n1352 & ~n18288 ;
  assign n18290 = n1356 & ~n18289 ;
  assign n18291 = n1360 & ~n18290 ;
  assign n18292 = n1364 & ~n18291 ;
  assign n18293 = n1368 & ~n18292 ;
  assign n18294 = n1372 & ~n18293 ;
  assign n18295 = n1376 & ~n18294 ;
  assign n18296 = n1380 & ~n18295 ;
  assign n18297 = n1384 & ~n18296 ;
  assign n18298 = n1388 & ~n18297 ;
  assign n18299 = n1392 & ~n18298 ;
  assign n18300 = n1396 & ~n18299 ;
  assign n18301 = n1400 & ~n18300 ;
  assign n18302 = n1404 & ~n18301 ;
  assign n18303 = n1408 & ~n18302 ;
  assign n18304 = n1412 & ~n18303 ;
  assign n18305 = n1416 & ~n18304 ;
  assign n18306 = n1420 & ~n18305 ;
  assign n18307 = n1424 & ~n18306 ;
  assign n18308 = n1428 & ~n18307 ;
  assign n18309 = n1432 & ~n18308 ;
  assign n18310 = n1436 & ~n18309 ;
  assign n18311 = n1440 & ~n18310 ;
  assign n18312 = n1444 & ~n18311 ;
  assign n18313 = n1448 & ~n18312 ;
  assign n18314 = n1452 & ~n18313 ;
  assign n18315 = n1456 & ~n18314 ;
  assign n18316 = n1460 & ~n18315 ;
  assign n18317 = n1464 & ~n18316 ;
  assign n18318 = n1468 & ~n18317 ;
  assign n18319 = n1472 & ~n18318 ;
  assign n18320 = n1476 & ~n18319 ;
  assign n18321 = n1480 & ~n18320 ;
  assign n18322 = n1484 & ~n18321 ;
  assign n18323 = n1488 & ~n18322 ;
  assign n18324 = n1492 & ~n18323 ;
  assign n18325 = n1496 & ~n18324 ;
  assign n18326 = n1500 & ~n18325 ;
  assign n18327 = n1504 & ~n18326 ;
  assign n18328 = n1508 & ~n18327 ;
  assign n18329 = n1512 & ~n18328 ;
  assign n18330 = n1516 & ~n18329 ;
  assign n18331 = ~x221 & ~n1518 ;
  assign n18332 = ~n18330 & n18331 ;
  assign n18335 = ~n18332 & ~x349 ;
  assign n18336 = ~n18334 & ~n18335 ;
  assign n18337 = n1188 & ~n1864 ;
  assign n18338 = n1193 & ~n18337 ;
  assign n18339 = n1197 & ~n18338 ;
  assign n18340 = n1201 & ~n18339 ;
  assign n18341 = n1205 & ~n18340 ;
  assign n18342 = n1209 & ~n18341 ;
  assign n18343 = n1213 & ~n18342 ;
  assign n18344 = n1217 & ~n18343 ;
  assign n18345 = n1221 & ~n18344 ;
  assign n18346 = n1225 & ~n18345 ;
  assign n18347 = n1229 & ~n18346 ;
  assign n18348 = n1233 & ~n18347 ;
  assign n18349 = n1237 & ~n18348 ;
  assign n18350 = n1241 & ~n18349 ;
  assign n18351 = n1245 & ~n18350 ;
  assign n18352 = n1249 & ~n18351 ;
  assign n18353 = n1253 & ~n18352 ;
  assign n18354 = n1257 & ~n18353 ;
  assign n18355 = n1261 & ~n18354 ;
  assign n18356 = n1265 & ~n18355 ;
  assign n18357 = n1269 & ~n18356 ;
  assign n18358 = n1273 & ~n18357 ;
  assign n18359 = n2566 & ~n18358 ;
  assign n18360 = n2568 & ~n18359 ;
  assign n18361 = n3105 & ~n18360 ;
  assign n18362 = n1625 & ~n18361 ;
  assign n18363 = n1629 & ~n18362 ;
  assign n18364 = n1633 & ~n18363 ;
  assign n18365 = n1637 & ~n18364 ;
  assign n18366 = n1641 & ~n18365 ;
  assign n18367 = n1645 & ~n18366 ;
  assign n18368 = n1649 & ~n18367 ;
  assign n18369 = n1653 & ~n18368 ;
  assign n18370 = n1657 & ~n18369 ;
  assign n18371 = n1661 & ~n18370 ;
  assign n18372 = n1665 & ~n18371 ;
  assign n18373 = n1669 & ~n18372 ;
  assign n18374 = n1673 & ~n18373 ;
  assign n18375 = n1677 & ~n18374 ;
  assign n18376 = n1681 & ~n18375 ;
  assign n18377 = n1685 & ~n18376 ;
  assign n18378 = n1689 & ~n18377 ;
  assign n18379 = n1693 & ~n18378 ;
  assign n18380 = n1697 & ~n18379 ;
  assign n18381 = n1701 & ~n18380 ;
  assign n18382 = n1705 & ~n18381 ;
  assign n18383 = n1709 & ~n18382 ;
  assign n18384 = n1713 & ~n18383 ;
  assign n18385 = n1717 & ~n18384 ;
  assign n18386 = n1721 & ~n18385 ;
  assign n18387 = n1725 & ~n18386 ;
  assign n18388 = n1729 & ~n18387 ;
  assign n18389 = n1733 & ~n18388 ;
  assign n18390 = n1737 & ~n18389 ;
  assign n18391 = n1741 & ~n18390 ;
  assign n18392 = n1745 & ~n18391 ;
  assign n18393 = n1749 & ~n18392 ;
  assign n18394 = n1753 & ~n18393 ;
  assign n18395 = n1757 & ~n18394 ;
  assign n18396 = n1761 & ~n18395 ;
  assign n18397 = n1765 & ~n18396 ;
  assign n18398 = n1769 & ~n18397 ;
  assign n18399 = n1773 & ~n18398 ;
  assign n18400 = n1777 & ~n18399 ;
  assign n18401 = n1781 & ~n18400 ;
  assign n18402 = n1785 & ~n18401 ;
  assign n18403 = n1789 & ~n18402 ;
  assign n18404 = n1793 & ~n18403 ;
  assign n18405 = n1797 & ~n18404 ;
  assign n18406 = n1801 & ~n18405 ;
  assign n18407 = n1805 & ~n18406 ;
  assign n18408 = n1809 & ~n18407 ;
  assign n18409 = n1813 & ~n18408 ;
  assign n18410 = n1817 & ~n18409 ;
  assign n18411 = n1821 & ~n18410 ;
  assign n18412 = n1825 & ~n18411 ;
  assign n18413 = n1829 & ~n18412 ;
  assign n18414 = n1833 & ~n18413 ;
  assign n18415 = n1837 & ~n18414 ;
  assign n18416 = n1841 & ~n18415 ;
  assign n18417 = n1845 & ~n18416 ;
  assign n18418 = n1849 & ~n18417 ;
  assign n18419 = n1853 & ~n18418 ;
  assign n18420 = n1857 & ~n18419 ;
  assign n18421 = x222 & ~n1859 ;
  assign n18422 = ~n18420 & n18421 ;
  assign n18510 = n18422 & x350 ;
  assign n18423 = n1527 & ~n2201 ;
  assign n18424 = n1532 & ~n18423 ;
  assign n18425 = n1536 & ~n18424 ;
  assign n18426 = n1540 & ~n18425 ;
  assign n18427 = n1544 & ~n18426 ;
  assign n18428 = n1548 & ~n18427 ;
  assign n18429 = n1552 & ~n18428 ;
  assign n18430 = n1556 & ~n18429 ;
  assign n18431 = n1560 & ~n18430 ;
  assign n18432 = n1564 & ~n18431 ;
  assign n18433 = n1568 & ~n18432 ;
  assign n18434 = n1572 & ~n18433 ;
  assign n18435 = n1576 & ~n18434 ;
  assign n18436 = n1580 & ~n18435 ;
  assign n18437 = n1584 & ~n18436 ;
  assign n18438 = n1588 & ~n18437 ;
  assign n18439 = n1592 & ~n18438 ;
  assign n18440 = n1596 & ~n18439 ;
  assign n18441 = n1600 & ~n18440 ;
  assign n18442 = n1604 & ~n18441 ;
  assign n18443 = n1608 & ~n18442 ;
  assign n18444 = n1612 & ~n18443 ;
  assign n18445 = n2656 & ~n18444 ;
  assign n18446 = n2658 & ~n18445 ;
  assign n18447 = n3192 & ~n18446 ;
  assign n18448 = n1962 & ~n18447 ;
  assign n18449 = n1966 & ~n18448 ;
  assign n18450 = n1970 & ~n18449 ;
  assign n18451 = n1974 & ~n18450 ;
  assign n18452 = n1978 & ~n18451 ;
  assign n18453 = n1982 & ~n18452 ;
  assign n18454 = n1986 & ~n18453 ;
  assign n18455 = n1990 & ~n18454 ;
  assign n18456 = n1994 & ~n18455 ;
  assign n18457 = n1998 & ~n18456 ;
  assign n18458 = n2002 & ~n18457 ;
  assign n18459 = n2006 & ~n18458 ;
  assign n18460 = n2010 & ~n18459 ;
  assign n18461 = n2014 & ~n18460 ;
  assign n18462 = n2018 & ~n18461 ;
  assign n18463 = n2022 & ~n18462 ;
  assign n18464 = n2026 & ~n18463 ;
  assign n18465 = n2030 & ~n18464 ;
  assign n18466 = n2034 & ~n18465 ;
  assign n18467 = n2038 & ~n18466 ;
  assign n18468 = n2042 & ~n18467 ;
  assign n18469 = n2046 & ~n18468 ;
  assign n18470 = n2050 & ~n18469 ;
  assign n18471 = n2054 & ~n18470 ;
  assign n18472 = n2058 & ~n18471 ;
  assign n18473 = n2062 & ~n18472 ;
  assign n18474 = n2066 & ~n18473 ;
  assign n18475 = n2070 & ~n18474 ;
  assign n18476 = n2074 & ~n18475 ;
  assign n18477 = n2078 & ~n18476 ;
  assign n18478 = n2082 & ~n18477 ;
  assign n18479 = n2086 & ~n18478 ;
  assign n18480 = n2090 & ~n18479 ;
  assign n18481 = n2094 & ~n18480 ;
  assign n18482 = n2098 & ~n18481 ;
  assign n18483 = n2102 & ~n18482 ;
  assign n18484 = n2106 & ~n18483 ;
  assign n18485 = n2110 & ~n18484 ;
  assign n18486 = n2114 & ~n18485 ;
  assign n18487 = n2118 & ~n18486 ;
  assign n18488 = n2122 & ~n18487 ;
  assign n18489 = n2126 & ~n18488 ;
  assign n18490 = n2130 & ~n18489 ;
  assign n18491 = n2134 & ~n18490 ;
  assign n18492 = n2138 & ~n18491 ;
  assign n18493 = n2142 & ~n18492 ;
  assign n18494 = n2146 & ~n18493 ;
  assign n18495 = n2150 & ~n18494 ;
  assign n18496 = n2154 & ~n18495 ;
  assign n18497 = n2158 & ~n18496 ;
  assign n18498 = n2162 & ~n18497 ;
  assign n18499 = n2166 & ~n18498 ;
  assign n18500 = n2170 & ~n18499 ;
  assign n18501 = n2174 & ~n18500 ;
  assign n18502 = n2178 & ~n18501 ;
  assign n18503 = n2182 & ~n18502 ;
  assign n18504 = n2186 & ~n18503 ;
  assign n18505 = n2190 & ~n18504 ;
  assign n18506 = n2194 & ~n18505 ;
  assign n18507 = ~x222 & ~n2196 ;
  assign n18508 = ~n18506 & n18507 ;
  assign n18511 = ~n18508 & ~x350 ;
  assign n18512 = ~n18510 & ~n18511 ;
  assign n18513 = ~n510 & n1868 ;
  assign n18514 = n1873 & ~n18513 ;
  assign n18515 = n1877 & ~n18514 ;
  assign n18516 = n1881 & ~n18515 ;
  assign n18517 = n1885 & ~n18516 ;
  assign n18518 = n1889 & ~n18517 ;
  assign n18519 = n1893 & ~n18518 ;
  assign n18520 = n1897 & ~n18519 ;
  assign n18521 = n1901 & ~n18520 ;
  assign n18522 = n1905 & ~n18521 ;
  assign n18523 = n1909 & ~n18522 ;
  assign n18524 = n1913 & ~n18523 ;
  assign n18525 = n1917 & ~n18524 ;
  assign n18526 = n1921 & ~n18525 ;
  assign n18527 = n1925 & ~n18526 ;
  assign n18528 = n1929 & ~n18527 ;
  assign n18529 = n1933 & ~n18528 ;
  assign n18530 = n1937 & ~n18529 ;
  assign n18531 = n1941 & ~n18530 ;
  assign n18532 = n1945 & ~n18531 ;
  assign n18533 = n1949 & ~n18532 ;
  assign n18534 = n1953 & ~n18533 ;
  assign n18535 = n2749 & ~n18534 ;
  assign n18536 = n263 & ~n18535 ;
  assign n18537 = n267 & ~n18536 ;
  assign n18538 = n271 & ~n18537 ;
  assign n18539 = n275 & ~n18538 ;
  assign n18540 = n279 & ~n18539 ;
  assign n18541 = n283 & ~n18540 ;
  assign n18542 = n287 & ~n18541 ;
  assign n18543 = n291 & ~n18542 ;
  assign n18544 = n295 & ~n18543 ;
  assign n18545 = n299 & ~n18544 ;
  assign n18546 = n303 & ~n18545 ;
  assign n18547 = n307 & ~n18546 ;
  assign n18548 = n311 & ~n18547 ;
  assign n18549 = n315 & ~n18548 ;
  assign n18550 = n319 & ~n18549 ;
  assign n18551 = n323 & ~n18550 ;
  assign n18552 = n327 & ~n18551 ;
  assign n18553 = n331 & ~n18552 ;
  assign n18554 = n335 & ~n18553 ;
  assign n18555 = n339 & ~n18554 ;
  assign n18556 = n343 & ~n18555 ;
  assign n18557 = n347 & ~n18556 ;
  assign n18558 = n351 & ~n18557 ;
  assign n18559 = n355 & ~n18558 ;
  assign n18560 = n359 & ~n18559 ;
  assign n18561 = n363 & ~n18560 ;
  assign n18562 = n367 & ~n18561 ;
  assign n18563 = n371 & ~n18562 ;
  assign n18564 = n375 & ~n18563 ;
  assign n18565 = n379 & ~n18564 ;
  assign n18566 = n383 & ~n18565 ;
  assign n18567 = n387 & ~n18566 ;
  assign n18568 = n391 & ~n18567 ;
  assign n18569 = n395 & ~n18568 ;
  assign n18570 = n399 & ~n18569 ;
  assign n18571 = n403 & ~n18570 ;
  assign n18572 = n407 & ~n18571 ;
  assign n18573 = n411 & ~n18572 ;
  assign n18574 = n415 & ~n18573 ;
  assign n18575 = n419 & ~n18574 ;
  assign n18576 = n423 & ~n18575 ;
  assign n18577 = n427 & ~n18576 ;
  assign n18578 = n431 & ~n18577 ;
  assign n18579 = n435 & ~n18578 ;
  assign n18580 = n439 & ~n18579 ;
  assign n18581 = n443 & ~n18580 ;
  assign n18582 = n447 & ~n18581 ;
  assign n18583 = n451 & ~n18582 ;
  assign n18584 = n455 & ~n18583 ;
  assign n18585 = n459 & ~n18584 ;
  assign n18586 = n463 & ~n18585 ;
  assign n18587 = n467 & ~n18586 ;
  assign n18588 = n471 & ~n18587 ;
  assign n18589 = n475 & ~n18588 ;
  assign n18590 = n479 & ~n18589 ;
  assign n18591 = n483 & ~n18590 ;
  assign n18592 = n487 & ~n18591 ;
  assign n18593 = n491 & ~n18592 ;
  assign n18594 = n495 & ~n18593 ;
  assign n18595 = n499 & ~n18594 ;
  assign n18596 = n503 & ~n18595 ;
  assign n18597 = x223 & ~n505 ;
  assign n18598 = ~n18596 & n18597 ;
  assign n18686 = n18598 & x351 ;
  assign n18599 = ~n849 & n2205 ;
  assign n18600 = n2210 & ~n18599 ;
  assign n18601 = n2214 & ~n18600 ;
  assign n18602 = n2218 & ~n18601 ;
  assign n18603 = n2222 & ~n18602 ;
  assign n18604 = n2226 & ~n18603 ;
  assign n18605 = n2230 & ~n18604 ;
  assign n18606 = n2234 & ~n18605 ;
  assign n18607 = n2238 & ~n18606 ;
  assign n18608 = n2242 & ~n18607 ;
  assign n18609 = n2246 & ~n18608 ;
  assign n18610 = n2250 & ~n18609 ;
  assign n18611 = n2254 & ~n18610 ;
  assign n18612 = n2258 & ~n18611 ;
  assign n18613 = n2262 & ~n18612 ;
  assign n18614 = n2266 & ~n18613 ;
  assign n18615 = n2270 & ~n18614 ;
  assign n18616 = n2274 & ~n18615 ;
  assign n18617 = n2278 & ~n18616 ;
  assign n18618 = n2282 & ~n18617 ;
  assign n18619 = n2286 & ~n18618 ;
  assign n18620 = n2290 & ~n18619 ;
  assign n18621 = n2836 & ~n18620 ;
  assign n18622 = n602 & ~n18621 ;
  assign n18623 = n606 & ~n18622 ;
  assign n18624 = n610 & ~n18623 ;
  assign n18625 = n614 & ~n18624 ;
  assign n18626 = n618 & ~n18625 ;
  assign n18627 = n622 & ~n18626 ;
  assign n18628 = n626 & ~n18627 ;
  assign n18629 = n630 & ~n18628 ;
  assign n18630 = n634 & ~n18629 ;
  assign n18631 = n638 & ~n18630 ;
  assign n18632 = n642 & ~n18631 ;
  assign n18633 = n646 & ~n18632 ;
  assign n18634 = n650 & ~n18633 ;
  assign n18635 = n654 & ~n18634 ;
  assign n18636 = n658 & ~n18635 ;
  assign n18637 = n662 & ~n18636 ;
  assign n18638 = n666 & ~n18637 ;
  assign n18639 = n670 & ~n18638 ;
  assign n18640 = n674 & ~n18639 ;
  assign n18641 = n678 & ~n18640 ;
  assign n18642 = n682 & ~n18641 ;
  assign n18643 = n686 & ~n18642 ;
  assign n18644 = n690 & ~n18643 ;
  assign n18645 = n694 & ~n18644 ;
  assign n18646 = n698 & ~n18645 ;
  assign n18647 = n702 & ~n18646 ;
  assign n18648 = n706 & ~n18647 ;
  assign n18649 = n710 & ~n18648 ;
  assign n18650 = n714 & ~n18649 ;
  assign n18651 = n718 & ~n18650 ;
  assign n18652 = n722 & ~n18651 ;
  assign n18653 = n726 & ~n18652 ;
  assign n18654 = n730 & ~n18653 ;
  assign n18655 = n734 & ~n18654 ;
  assign n18656 = n738 & ~n18655 ;
  assign n18657 = n742 & ~n18656 ;
  assign n18658 = n746 & ~n18657 ;
  assign n18659 = n750 & ~n18658 ;
  assign n18660 = n754 & ~n18659 ;
  assign n18661 = n758 & ~n18660 ;
  assign n18662 = n762 & ~n18661 ;
  assign n18663 = n766 & ~n18662 ;
  assign n18664 = n770 & ~n18663 ;
  assign n18665 = n774 & ~n18664 ;
  assign n18666 = n778 & ~n18665 ;
  assign n18667 = n782 & ~n18666 ;
  assign n18668 = n786 & ~n18667 ;
  assign n18669 = n790 & ~n18668 ;
  assign n18670 = n794 & ~n18669 ;
  assign n18671 = n798 & ~n18670 ;
  assign n18672 = n802 & ~n18671 ;
  assign n18673 = n806 & ~n18672 ;
  assign n18674 = n810 & ~n18673 ;
  assign n18675 = n814 & ~n18674 ;
  assign n18676 = n818 & ~n18675 ;
  assign n18677 = n822 & ~n18676 ;
  assign n18678 = n826 & ~n18677 ;
  assign n18679 = n830 & ~n18678 ;
  assign n18680 = n834 & ~n18679 ;
  assign n18681 = n838 & ~n18680 ;
  assign n18682 = n842 & ~n18681 ;
  assign n18683 = ~x223 & ~n844 ;
  assign n18684 = ~n18682 & n18683 ;
  assign n18687 = ~n18684 & ~x351 ;
  assign n18688 = ~n18686 & ~n18687 ;
  assign n18689 = n514 & ~n1192 ;
  assign n18690 = n519 & ~n18689 ;
  assign n18691 = n523 & ~n18690 ;
  assign n18692 = n527 & ~n18691 ;
  assign n18693 = n531 & ~n18692 ;
  assign n18694 = n535 & ~n18693 ;
  assign n18695 = n539 & ~n18694 ;
  assign n18696 = n543 & ~n18695 ;
  assign n18697 = n547 & ~n18696 ;
  assign n18698 = n551 & ~n18697 ;
  assign n18699 = n555 & ~n18698 ;
  assign n18700 = n559 & ~n18699 ;
  assign n18701 = n563 & ~n18700 ;
  assign n18702 = n567 & ~n18701 ;
  assign n18703 = n571 & ~n18702 ;
  assign n18704 = n575 & ~n18703 ;
  assign n18705 = n579 & ~n18704 ;
  assign n18706 = n583 & ~n18705 ;
  assign n18707 = n587 & ~n18706 ;
  assign n18708 = n591 & ~n18707 ;
  assign n18709 = n2382 & ~n18708 ;
  assign n18710 = n2384 & ~n18709 ;
  assign n18711 = n2927 & ~n18710 ;
  assign n18712 = n945 & ~n18711 ;
  assign n18713 = n949 & ~n18712 ;
  assign n18714 = n953 & ~n18713 ;
  assign n18715 = n957 & ~n18714 ;
  assign n18716 = n961 & ~n18715 ;
  assign n18717 = n965 & ~n18716 ;
  assign n18718 = n969 & ~n18717 ;
  assign n18719 = n973 & ~n18718 ;
  assign n18720 = n977 & ~n18719 ;
  assign n18721 = n981 & ~n18720 ;
  assign n18722 = n985 & ~n18721 ;
  assign n18723 = n989 & ~n18722 ;
  assign n18724 = n993 & ~n18723 ;
  assign n18725 = n997 & ~n18724 ;
  assign n18726 = n1001 & ~n18725 ;
  assign n18727 = n1005 & ~n18726 ;
  assign n18728 = n1009 & ~n18727 ;
  assign n18729 = n1013 & ~n18728 ;
  assign n18730 = n1017 & ~n18729 ;
  assign n18731 = n1021 & ~n18730 ;
  assign n18732 = n1025 & ~n18731 ;
  assign n18733 = n1029 & ~n18732 ;
  assign n18734 = n1033 & ~n18733 ;
  assign n18735 = n1037 & ~n18734 ;
  assign n18736 = n1041 & ~n18735 ;
  assign n18737 = n1045 & ~n18736 ;
  assign n18738 = n1049 & ~n18737 ;
  assign n18739 = n1053 & ~n18738 ;
  assign n18740 = n1057 & ~n18739 ;
  assign n18741 = n1061 & ~n18740 ;
  assign n18742 = n1065 & ~n18741 ;
  assign n18743 = n1069 & ~n18742 ;
  assign n18744 = n1073 & ~n18743 ;
  assign n18745 = n1077 & ~n18744 ;
  assign n18746 = n1081 & ~n18745 ;
  assign n18747 = n1085 & ~n18746 ;
  assign n18748 = n1089 & ~n18747 ;
  assign n18749 = n1093 & ~n18748 ;
  assign n18750 = n1097 & ~n18749 ;
  assign n18751 = n1101 & ~n18750 ;
  assign n18752 = n1105 & ~n18751 ;
  assign n18753 = n1109 & ~n18752 ;
  assign n18754 = n1113 & ~n18753 ;
  assign n18755 = n1117 & ~n18754 ;
  assign n18756 = n1121 & ~n18755 ;
  assign n18757 = n1125 & ~n18756 ;
  assign n18758 = n1129 & ~n18757 ;
  assign n18759 = n1133 & ~n18758 ;
  assign n18760 = n1137 & ~n18759 ;
  assign n18761 = n1141 & ~n18760 ;
  assign n18762 = n1145 & ~n18761 ;
  assign n18763 = n1149 & ~n18762 ;
  assign n18764 = n1153 & ~n18763 ;
  assign n18765 = n1157 & ~n18764 ;
  assign n18766 = n1161 & ~n18765 ;
  assign n18767 = n1165 & ~n18766 ;
  assign n18768 = n1169 & ~n18767 ;
  assign n18769 = n1173 & ~n18768 ;
  assign n18770 = n1177 & ~n18769 ;
  assign n18771 = n1181 & ~n18770 ;
  assign n18772 = n1185 & ~n18771 ;
  assign n18773 = x224 & ~n1187 ;
  assign n18774 = ~n18772 & n18773 ;
  assign n18862 = n18774 & x352 ;
  assign n18775 = n853 & ~n1531 ;
  assign n18776 = n858 & ~n18775 ;
  assign n18777 = n862 & ~n18776 ;
  assign n18778 = n866 & ~n18777 ;
  assign n18779 = n870 & ~n18778 ;
  assign n18780 = n874 & ~n18779 ;
  assign n18781 = n878 & ~n18780 ;
  assign n18782 = n882 & ~n18781 ;
  assign n18783 = n886 & ~n18782 ;
  assign n18784 = n890 & ~n18783 ;
  assign n18785 = n894 & ~n18784 ;
  assign n18786 = n898 & ~n18785 ;
  assign n18787 = n902 & ~n18786 ;
  assign n18788 = n906 & ~n18787 ;
  assign n18789 = n910 & ~n18788 ;
  assign n18790 = n914 & ~n18789 ;
  assign n18791 = n918 & ~n18790 ;
  assign n18792 = n922 & ~n18791 ;
  assign n18793 = n926 & ~n18792 ;
  assign n18794 = n930 & ~n18793 ;
  assign n18795 = n2472 & ~n18794 ;
  assign n18796 = n2474 & ~n18795 ;
  assign n18797 = n3014 & ~n18796 ;
  assign n18798 = n1284 & ~n18797 ;
  assign n18799 = n1288 & ~n18798 ;
  assign n18800 = n1292 & ~n18799 ;
  assign n18801 = n1296 & ~n18800 ;
  assign n18802 = n1300 & ~n18801 ;
  assign n18803 = n1304 & ~n18802 ;
  assign n18804 = n1308 & ~n18803 ;
  assign n18805 = n1312 & ~n18804 ;
  assign n18806 = n1316 & ~n18805 ;
  assign n18807 = n1320 & ~n18806 ;
  assign n18808 = n1324 & ~n18807 ;
  assign n18809 = n1328 & ~n18808 ;
  assign n18810 = n1332 & ~n18809 ;
  assign n18811 = n1336 & ~n18810 ;
  assign n18812 = n1340 & ~n18811 ;
  assign n18813 = n1344 & ~n18812 ;
  assign n18814 = n1348 & ~n18813 ;
  assign n18815 = n1352 & ~n18814 ;
  assign n18816 = n1356 & ~n18815 ;
  assign n18817 = n1360 & ~n18816 ;
  assign n18818 = n1364 & ~n18817 ;
  assign n18819 = n1368 & ~n18818 ;
  assign n18820 = n1372 & ~n18819 ;
  assign n18821 = n1376 & ~n18820 ;
  assign n18822 = n1380 & ~n18821 ;
  assign n18823 = n1384 & ~n18822 ;
  assign n18824 = n1388 & ~n18823 ;
  assign n18825 = n1392 & ~n18824 ;
  assign n18826 = n1396 & ~n18825 ;
  assign n18827 = n1400 & ~n18826 ;
  assign n18828 = n1404 & ~n18827 ;
  assign n18829 = n1408 & ~n18828 ;
  assign n18830 = n1412 & ~n18829 ;
  assign n18831 = n1416 & ~n18830 ;
  assign n18832 = n1420 & ~n18831 ;
  assign n18833 = n1424 & ~n18832 ;
  assign n18834 = n1428 & ~n18833 ;
  assign n18835 = n1432 & ~n18834 ;
  assign n18836 = n1436 & ~n18835 ;
  assign n18837 = n1440 & ~n18836 ;
  assign n18838 = n1444 & ~n18837 ;
  assign n18839 = n1448 & ~n18838 ;
  assign n18840 = n1452 & ~n18839 ;
  assign n18841 = n1456 & ~n18840 ;
  assign n18842 = n1460 & ~n18841 ;
  assign n18843 = n1464 & ~n18842 ;
  assign n18844 = n1468 & ~n18843 ;
  assign n18845 = n1472 & ~n18844 ;
  assign n18846 = n1476 & ~n18845 ;
  assign n18847 = n1480 & ~n18846 ;
  assign n18848 = n1484 & ~n18847 ;
  assign n18849 = n1488 & ~n18848 ;
  assign n18850 = n1492 & ~n18849 ;
  assign n18851 = n1496 & ~n18850 ;
  assign n18852 = n1500 & ~n18851 ;
  assign n18853 = n1504 & ~n18852 ;
  assign n18854 = n1508 & ~n18853 ;
  assign n18855 = n1512 & ~n18854 ;
  assign n18856 = n1516 & ~n18855 ;
  assign n18857 = n1520 & ~n18856 ;
  assign n18858 = n1524 & ~n18857 ;
  assign n18859 = ~x224 & ~n1526 ;
  assign n18860 = ~n18858 & n18859 ;
  assign n18863 = ~n18860 & ~x352 ;
  assign n18864 = ~n18862 & ~n18863 ;
  assign n18865 = n1196 & ~n1872 ;
  assign n18866 = n1201 & ~n18865 ;
  assign n18867 = n1205 & ~n18866 ;
  assign n18868 = n1209 & ~n18867 ;
  assign n18869 = n1213 & ~n18868 ;
  assign n18870 = n1217 & ~n18869 ;
  assign n18871 = n1221 & ~n18870 ;
  assign n18872 = n1225 & ~n18871 ;
  assign n18873 = n1229 & ~n18872 ;
  assign n18874 = n1233 & ~n18873 ;
  assign n18875 = n1237 & ~n18874 ;
  assign n18876 = n1241 & ~n18875 ;
  assign n18877 = n1245 & ~n18876 ;
  assign n18878 = n1249 & ~n18877 ;
  assign n18879 = n1253 & ~n18878 ;
  assign n18880 = n1257 & ~n18879 ;
  assign n18881 = n1261 & ~n18880 ;
  assign n18882 = n1265 & ~n18881 ;
  assign n18883 = n1269 & ~n18882 ;
  assign n18884 = n1273 & ~n18883 ;
  assign n18885 = n2566 & ~n18884 ;
  assign n18886 = n2568 & ~n18885 ;
  assign n18887 = n3105 & ~n18886 ;
  assign n18888 = n1625 & ~n18887 ;
  assign n18889 = n1629 & ~n18888 ;
  assign n18890 = n1633 & ~n18889 ;
  assign n18891 = n1637 & ~n18890 ;
  assign n18892 = n1641 & ~n18891 ;
  assign n18893 = n1645 & ~n18892 ;
  assign n18894 = n1649 & ~n18893 ;
  assign n18895 = n1653 & ~n18894 ;
  assign n18896 = n1657 & ~n18895 ;
  assign n18897 = n1661 & ~n18896 ;
  assign n18898 = n1665 & ~n18897 ;
  assign n18899 = n1669 & ~n18898 ;
  assign n18900 = n1673 & ~n18899 ;
  assign n18901 = n1677 & ~n18900 ;
  assign n18902 = n1681 & ~n18901 ;
  assign n18903 = n1685 & ~n18902 ;
  assign n18904 = n1689 & ~n18903 ;
  assign n18905 = n1693 & ~n18904 ;
  assign n18906 = n1697 & ~n18905 ;
  assign n18907 = n1701 & ~n18906 ;
  assign n18908 = n1705 & ~n18907 ;
  assign n18909 = n1709 & ~n18908 ;
  assign n18910 = n1713 & ~n18909 ;
  assign n18911 = n1717 & ~n18910 ;
  assign n18912 = n1721 & ~n18911 ;
  assign n18913 = n1725 & ~n18912 ;
  assign n18914 = n1729 & ~n18913 ;
  assign n18915 = n1733 & ~n18914 ;
  assign n18916 = n1737 & ~n18915 ;
  assign n18917 = n1741 & ~n18916 ;
  assign n18918 = n1745 & ~n18917 ;
  assign n18919 = n1749 & ~n18918 ;
  assign n18920 = n1753 & ~n18919 ;
  assign n18921 = n1757 & ~n18920 ;
  assign n18922 = n1761 & ~n18921 ;
  assign n18923 = n1765 & ~n18922 ;
  assign n18924 = n1769 & ~n18923 ;
  assign n18925 = n1773 & ~n18924 ;
  assign n18926 = n1777 & ~n18925 ;
  assign n18927 = n1781 & ~n18926 ;
  assign n18928 = n1785 & ~n18927 ;
  assign n18929 = n1789 & ~n18928 ;
  assign n18930 = n1793 & ~n18929 ;
  assign n18931 = n1797 & ~n18930 ;
  assign n18932 = n1801 & ~n18931 ;
  assign n18933 = n1805 & ~n18932 ;
  assign n18934 = n1809 & ~n18933 ;
  assign n18935 = n1813 & ~n18934 ;
  assign n18936 = n1817 & ~n18935 ;
  assign n18937 = n1821 & ~n18936 ;
  assign n18938 = n1825 & ~n18937 ;
  assign n18939 = n1829 & ~n18938 ;
  assign n18940 = n1833 & ~n18939 ;
  assign n18941 = n1837 & ~n18940 ;
  assign n18942 = n1841 & ~n18941 ;
  assign n18943 = n1845 & ~n18942 ;
  assign n18944 = n1849 & ~n18943 ;
  assign n18945 = n1853 & ~n18944 ;
  assign n18946 = n1857 & ~n18945 ;
  assign n18947 = n1861 & ~n18946 ;
  assign n18948 = n1865 & ~n18947 ;
  assign n18949 = x225 & ~n1867 ;
  assign n18950 = ~n18948 & n18949 ;
  assign n19038 = n18950 & x353 ;
  assign n18951 = n1535 & ~n2209 ;
  assign n18952 = n1540 & ~n18951 ;
  assign n18953 = n1544 & ~n18952 ;
  assign n18954 = n1548 & ~n18953 ;
  assign n18955 = n1552 & ~n18954 ;
  assign n18956 = n1556 & ~n18955 ;
  assign n18957 = n1560 & ~n18956 ;
  assign n18958 = n1564 & ~n18957 ;
  assign n18959 = n1568 & ~n18958 ;
  assign n18960 = n1572 & ~n18959 ;
  assign n18961 = n1576 & ~n18960 ;
  assign n18962 = n1580 & ~n18961 ;
  assign n18963 = n1584 & ~n18962 ;
  assign n18964 = n1588 & ~n18963 ;
  assign n18965 = n1592 & ~n18964 ;
  assign n18966 = n1596 & ~n18965 ;
  assign n18967 = n1600 & ~n18966 ;
  assign n18968 = n1604 & ~n18967 ;
  assign n18969 = n1608 & ~n18968 ;
  assign n18970 = n1612 & ~n18969 ;
  assign n18971 = n2656 & ~n18970 ;
  assign n18972 = n2658 & ~n18971 ;
  assign n18973 = n3192 & ~n18972 ;
  assign n18974 = n1962 & ~n18973 ;
  assign n18975 = n1966 & ~n18974 ;
  assign n18976 = n1970 & ~n18975 ;
  assign n18977 = n1974 & ~n18976 ;
  assign n18978 = n1978 & ~n18977 ;
  assign n18979 = n1982 & ~n18978 ;
  assign n18980 = n1986 & ~n18979 ;
  assign n18981 = n1990 & ~n18980 ;
  assign n18982 = n1994 & ~n18981 ;
  assign n18983 = n1998 & ~n18982 ;
  assign n18984 = n2002 & ~n18983 ;
  assign n18985 = n2006 & ~n18984 ;
  assign n18986 = n2010 & ~n18985 ;
  assign n18987 = n2014 & ~n18986 ;
  assign n18988 = n2018 & ~n18987 ;
  assign n18989 = n2022 & ~n18988 ;
  assign n18990 = n2026 & ~n18989 ;
  assign n18991 = n2030 & ~n18990 ;
  assign n18992 = n2034 & ~n18991 ;
  assign n18993 = n2038 & ~n18992 ;
  assign n18994 = n2042 & ~n18993 ;
  assign n18995 = n2046 & ~n18994 ;
  assign n18996 = n2050 & ~n18995 ;
  assign n18997 = n2054 & ~n18996 ;
  assign n18998 = n2058 & ~n18997 ;
  assign n18999 = n2062 & ~n18998 ;
  assign n19000 = n2066 & ~n18999 ;
  assign n19001 = n2070 & ~n19000 ;
  assign n19002 = n2074 & ~n19001 ;
  assign n19003 = n2078 & ~n19002 ;
  assign n19004 = n2082 & ~n19003 ;
  assign n19005 = n2086 & ~n19004 ;
  assign n19006 = n2090 & ~n19005 ;
  assign n19007 = n2094 & ~n19006 ;
  assign n19008 = n2098 & ~n19007 ;
  assign n19009 = n2102 & ~n19008 ;
  assign n19010 = n2106 & ~n19009 ;
  assign n19011 = n2110 & ~n19010 ;
  assign n19012 = n2114 & ~n19011 ;
  assign n19013 = n2118 & ~n19012 ;
  assign n19014 = n2122 & ~n19013 ;
  assign n19015 = n2126 & ~n19014 ;
  assign n19016 = n2130 & ~n19015 ;
  assign n19017 = n2134 & ~n19016 ;
  assign n19018 = n2138 & ~n19017 ;
  assign n19019 = n2142 & ~n19018 ;
  assign n19020 = n2146 & ~n19019 ;
  assign n19021 = n2150 & ~n19020 ;
  assign n19022 = n2154 & ~n19021 ;
  assign n19023 = n2158 & ~n19022 ;
  assign n19024 = n2162 & ~n19023 ;
  assign n19025 = n2166 & ~n19024 ;
  assign n19026 = n2170 & ~n19025 ;
  assign n19027 = n2174 & ~n19026 ;
  assign n19028 = n2178 & ~n19027 ;
  assign n19029 = n2182 & ~n19028 ;
  assign n19030 = n2186 & ~n19029 ;
  assign n19031 = n2190 & ~n19030 ;
  assign n19032 = n2194 & ~n19031 ;
  assign n19033 = n2198 & ~n19032 ;
  assign n19034 = n2202 & ~n19033 ;
  assign n19035 = ~x225 & ~n2204 ;
  assign n19036 = ~n19034 & n19035 ;
  assign n19039 = ~n19036 & ~x353 ;
  assign n19040 = ~n19038 & ~n19039 ;
  assign n19041 = ~n518 & n1876 ;
  assign n19042 = n1881 & ~n19041 ;
  assign n19043 = n1885 & ~n19042 ;
  assign n19044 = n1889 & ~n19043 ;
  assign n19045 = n1893 & ~n19044 ;
  assign n19046 = n1897 & ~n19045 ;
  assign n19047 = n1901 & ~n19046 ;
  assign n19048 = n1905 & ~n19047 ;
  assign n19049 = n1909 & ~n19048 ;
  assign n19050 = n1913 & ~n19049 ;
  assign n19051 = n1917 & ~n19050 ;
  assign n19052 = n1921 & ~n19051 ;
  assign n19053 = n1925 & ~n19052 ;
  assign n19054 = n1929 & ~n19053 ;
  assign n19055 = n1933 & ~n19054 ;
  assign n19056 = n1937 & ~n19055 ;
  assign n19057 = n1941 & ~n19056 ;
  assign n19058 = n1945 & ~n19057 ;
  assign n19059 = n1949 & ~n19058 ;
  assign n19060 = n1953 & ~n19059 ;
  assign n19061 = n2749 & ~n19060 ;
  assign n19062 = n263 & ~n19061 ;
  assign n19063 = n267 & ~n19062 ;
  assign n19064 = n271 & ~n19063 ;
  assign n19065 = n275 & ~n19064 ;
  assign n19066 = n279 & ~n19065 ;
  assign n19067 = n283 & ~n19066 ;
  assign n19068 = n287 & ~n19067 ;
  assign n19069 = n291 & ~n19068 ;
  assign n19070 = n295 & ~n19069 ;
  assign n19071 = n299 & ~n19070 ;
  assign n19072 = n303 & ~n19071 ;
  assign n19073 = n307 & ~n19072 ;
  assign n19074 = n311 & ~n19073 ;
  assign n19075 = n315 & ~n19074 ;
  assign n19076 = n319 & ~n19075 ;
  assign n19077 = n323 & ~n19076 ;
  assign n19078 = n327 & ~n19077 ;
  assign n19079 = n331 & ~n19078 ;
  assign n19080 = n335 & ~n19079 ;
  assign n19081 = n339 & ~n19080 ;
  assign n19082 = n343 & ~n19081 ;
  assign n19083 = n347 & ~n19082 ;
  assign n19084 = n351 & ~n19083 ;
  assign n19085 = n355 & ~n19084 ;
  assign n19086 = n359 & ~n19085 ;
  assign n19087 = n363 & ~n19086 ;
  assign n19088 = n367 & ~n19087 ;
  assign n19089 = n371 & ~n19088 ;
  assign n19090 = n375 & ~n19089 ;
  assign n19091 = n379 & ~n19090 ;
  assign n19092 = n383 & ~n19091 ;
  assign n19093 = n387 & ~n19092 ;
  assign n19094 = n391 & ~n19093 ;
  assign n19095 = n395 & ~n19094 ;
  assign n19096 = n399 & ~n19095 ;
  assign n19097 = n403 & ~n19096 ;
  assign n19098 = n407 & ~n19097 ;
  assign n19099 = n411 & ~n19098 ;
  assign n19100 = n415 & ~n19099 ;
  assign n19101 = n419 & ~n19100 ;
  assign n19102 = n423 & ~n19101 ;
  assign n19103 = n427 & ~n19102 ;
  assign n19104 = n431 & ~n19103 ;
  assign n19105 = n435 & ~n19104 ;
  assign n19106 = n439 & ~n19105 ;
  assign n19107 = n443 & ~n19106 ;
  assign n19108 = n447 & ~n19107 ;
  assign n19109 = n451 & ~n19108 ;
  assign n19110 = n455 & ~n19109 ;
  assign n19111 = n459 & ~n19110 ;
  assign n19112 = n463 & ~n19111 ;
  assign n19113 = n467 & ~n19112 ;
  assign n19114 = n471 & ~n19113 ;
  assign n19115 = n475 & ~n19114 ;
  assign n19116 = n479 & ~n19115 ;
  assign n19117 = n483 & ~n19116 ;
  assign n19118 = n487 & ~n19117 ;
  assign n19119 = n491 & ~n19118 ;
  assign n19120 = n495 & ~n19119 ;
  assign n19121 = n499 & ~n19120 ;
  assign n19122 = n503 & ~n19121 ;
  assign n19123 = n507 & ~n19122 ;
  assign n19124 = n511 & ~n19123 ;
  assign n19125 = x226 & ~n513 ;
  assign n19126 = ~n19124 & n19125 ;
  assign n19214 = n19126 & x354 ;
  assign n19127 = ~n857 & n2213 ;
  assign n19128 = n2218 & ~n19127 ;
  assign n19129 = n2222 & ~n19128 ;
  assign n19130 = n2226 & ~n19129 ;
  assign n19131 = n2230 & ~n19130 ;
  assign n19132 = n2234 & ~n19131 ;
  assign n19133 = n2238 & ~n19132 ;
  assign n19134 = n2242 & ~n19133 ;
  assign n19135 = n2246 & ~n19134 ;
  assign n19136 = n2250 & ~n19135 ;
  assign n19137 = n2254 & ~n19136 ;
  assign n19138 = n2258 & ~n19137 ;
  assign n19139 = n2262 & ~n19138 ;
  assign n19140 = n2266 & ~n19139 ;
  assign n19141 = n2270 & ~n19140 ;
  assign n19142 = n2274 & ~n19141 ;
  assign n19143 = n2278 & ~n19142 ;
  assign n19144 = n2282 & ~n19143 ;
  assign n19145 = n2286 & ~n19144 ;
  assign n19146 = n2290 & ~n19145 ;
  assign n19147 = n2836 & ~n19146 ;
  assign n19148 = n602 & ~n19147 ;
  assign n19149 = n606 & ~n19148 ;
  assign n19150 = n610 & ~n19149 ;
  assign n19151 = n614 & ~n19150 ;
  assign n19152 = n618 & ~n19151 ;
  assign n19153 = n622 & ~n19152 ;
  assign n19154 = n626 & ~n19153 ;
  assign n19155 = n630 & ~n19154 ;
  assign n19156 = n634 & ~n19155 ;
  assign n19157 = n638 & ~n19156 ;
  assign n19158 = n642 & ~n19157 ;
  assign n19159 = n646 & ~n19158 ;
  assign n19160 = n650 & ~n19159 ;
  assign n19161 = n654 & ~n19160 ;
  assign n19162 = n658 & ~n19161 ;
  assign n19163 = n662 & ~n19162 ;
  assign n19164 = n666 & ~n19163 ;
  assign n19165 = n670 & ~n19164 ;
  assign n19166 = n674 & ~n19165 ;
  assign n19167 = n678 & ~n19166 ;
  assign n19168 = n682 & ~n19167 ;
  assign n19169 = n686 & ~n19168 ;
  assign n19170 = n690 & ~n19169 ;
  assign n19171 = n694 & ~n19170 ;
  assign n19172 = n698 & ~n19171 ;
  assign n19173 = n702 & ~n19172 ;
  assign n19174 = n706 & ~n19173 ;
  assign n19175 = n710 & ~n19174 ;
  assign n19176 = n714 & ~n19175 ;
  assign n19177 = n718 & ~n19176 ;
  assign n19178 = n722 & ~n19177 ;
  assign n19179 = n726 & ~n19178 ;
  assign n19180 = n730 & ~n19179 ;
  assign n19181 = n734 & ~n19180 ;
  assign n19182 = n738 & ~n19181 ;
  assign n19183 = n742 & ~n19182 ;
  assign n19184 = n746 & ~n19183 ;
  assign n19185 = n750 & ~n19184 ;
  assign n19186 = n754 & ~n19185 ;
  assign n19187 = n758 & ~n19186 ;
  assign n19188 = n762 & ~n19187 ;
  assign n19189 = n766 & ~n19188 ;
  assign n19190 = n770 & ~n19189 ;
  assign n19191 = n774 & ~n19190 ;
  assign n19192 = n778 & ~n19191 ;
  assign n19193 = n782 & ~n19192 ;
  assign n19194 = n786 & ~n19193 ;
  assign n19195 = n790 & ~n19194 ;
  assign n19196 = n794 & ~n19195 ;
  assign n19197 = n798 & ~n19196 ;
  assign n19198 = n802 & ~n19197 ;
  assign n19199 = n806 & ~n19198 ;
  assign n19200 = n810 & ~n19199 ;
  assign n19201 = n814 & ~n19200 ;
  assign n19202 = n818 & ~n19201 ;
  assign n19203 = n822 & ~n19202 ;
  assign n19204 = n826 & ~n19203 ;
  assign n19205 = n830 & ~n19204 ;
  assign n19206 = n834 & ~n19205 ;
  assign n19207 = n838 & ~n19206 ;
  assign n19208 = n842 & ~n19207 ;
  assign n19209 = n846 & ~n19208 ;
  assign n19210 = n850 & ~n19209 ;
  assign n19211 = ~x226 & ~n852 ;
  assign n19212 = ~n19210 & n19211 ;
  assign n19215 = ~n19212 & ~x354 ;
  assign n19216 = ~n19214 & ~n19215 ;
  assign n19217 = n522 & ~n1200 ;
  assign n19218 = n527 & ~n19217 ;
  assign n19219 = n531 & ~n19218 ;
  assign n19220 = n535 & ~n19219 ;
  assign n19221 = n539 & ~n19220 ;
  assign n19222 = n543 & ~n19221 ;
  assign n19223 = n547 & ~n19222 ;
  assign n19224 = n551 & ~n19223 ;
  assign n19225 = n555 & ~n19224 ;
  assign n19226 = n559 & ~n19225 ;
  assign n19227 = n563 & ~n19226 ;
  assign n19228 = n567 & ~n19227 ;
  assign n19229 = n571 & ~n19228 ;
  assign n19230 = n575 & ~n19229 ;
  assign n19231 = n579 & ~n19230 ;
  assign n19232 = n583 & ~n19231 ;
  assign n19233 = n587 & ~n19232 ;
  assign n19234 = n591 & ~n19233 ;
  assign n19235 = n2382 & ~n19234 ;
  assign n19236 = n2384 & ~n19235 ;
  assign n19237 = n2927 & ~n19236 ;
  assign n19238 = n945 & ~n19237 ;
  assign n19239 = n949 & ~n19238 ;
  assign n19240 = n953 & ~n19239 ;
  assign n19241 = n957 & ~n19240 ;
  assign n19242 = n961 & ~n19241 ;
  assign n19243 = n965 & ~n19242 ;
  assign n19244 = n969 & ~n19243 ;
  assign n19245 = n973 & ~n19244 ;
  assign n19246 = n977 & ~n19245 ;
  assign n19247 = n981 & ~n19246 ;
  assign n19248 = n985 & ~n19247 ;
  assign n19249 = n989 & ~n19248 ;
  assign n19250 = n993 & ~n19249 ;
  assign n19251 = n997 & ~n19250 ;
  assign n19252 = n1001 & ~n19251 ;
  assign n19253 = n1005 & ~n19252 ;
  assign n19254 = n1009 & ~n19253 ;
  assign n19255 = n1013 & ~n19254 ;
  assign n19256 = n1017 & ~n19255 ;
  assign n19257 = n1021 & ~n19256 ;
  assign n19258 = n1025 & ~n19257 ;
  assign n19259 = n1029 & ~n19258 ;
  assign n19260 = n1033 & ~n19259 ;
  assign n19261 = n1037 & ~n19260 ;
  assign n19262 = n1041 & ~n19261 ;
  assign n19263 = n1045 & ~n19262 ;
  assign n19264 = n1049 & ~n19263 ;
  assign n19265 = n1053 & ~n19264 ;
  assign n19266 = n1057 & ~n19265 ;
  assign n19267 = n1061 & ~n19266 ;
  assign n19268 = n1065 & ~n19267 ;
  assign n19269 = n1069 & ~n19268 ;
  assign n19270 = n1073 & ~n19269 ;
  assign n19271 = n1077 & ~n19270 ;
  assign n19272 = n1081 & ~n19271 ;
  assign n19273 = n1085 & ~n19272 ;
  assign n19274 = n1089 & ~n19273 ;
  assign n19275 = n1093 & ~n19274 ;
  assign n19276 = n1097 & ~n19275 ;
  assign n19277 = n1101 & ~n19276 ;
  assign n19278 = n1105 & ~n19277 ;
  assign n19279 = n1109 & ~n19278 ;
  assign n19280 = n1113 & ~n19279 ;
  assign n19281 = n1117 & ~n19280 ;
  assign n19282 = n1121 & ~n19281 ;
  assign n19283 = n1125 & ~n19282 ;
  assign n19284 = n1129 & ~n19283 ;
  assign n19285 = n1133 & ~n19284 ;
  assign n19286 = n1137 & ~n19285 ;
  assign n19287 = n1141 & ~n19286 ;
  assign n19288 = n1145 & ~n19287 ;
  assign n19289 = n1149 & ~n19288 ;
  assign n19290 = n1153 & ~n19289 ;
  assign n19291 = n1157 & ~n19290 ;
  assign n19292 = n1161 & ~n19291 ;
  assign n19293 = n1165 & ~n19292 ;
  assign n19294 = n1169 & ~n19293 ;
  assign n19295 = n1173 & ~n19294 ;
  assign n19296 = n1177 & ~n19295 ;
  assign n19297 = n1181 & ~n19296 ;
  assign n19298 = n1185 & ~n19297 ;
  assign n19299 = n1189 & ~n19298 ;
  assign n19300 = n1193 & ~n19299 ;
  assign n19301 = x227 & ~n1195 ;
  assign n19302 = ~n19300 & n19301 ;
  assign n19390 = n19302 & x355 ;
  assign n19303 = n861 & ~n1539 ;
  assign n19304 = n866 & ~n19303 ;
  assign n19305 = n870 & ~n19304 ;
  assign n19306 = n874 & ~n19305 ;
  assign n19307 = n878 & ~n19306 ;
  assign n19308 = n882 & ~n19307 ;
  assign n19309 = n886 & ~n19308 ;
  assign n19310 = n890 & ~n19309 ;
  assign n19311 = n894 & ~n19310 ;
  assign n19312 = n898 & ~n19311 ;
  assign n19313 = n902 & ~n19312 ;
  assign n19314 = n906 & ~n19313 ;
  assign n19315 = n910 & ~n19314 ;
  assign n19316 = n914 & ~n19315 ;
  assign n19317 = n918 & ~n19316 ;
  assign n19318 = n922 & ~n19317 ;
  assign n19319 = n926 & ~n19318 ;
  assign n19320 = n930 & ~n19319 ;
  assign n19321 = n2472 & ~n19320 ;
  assign n19322 = n2474 & ~n19321 ;
  assign n19323 = n3014 & ~n19322 ;
  assign n19324 = n1284 & ~n19323 ;
  assign n19325 = n1288 & ~n19324 ;
  assign n19326 = n1292 & ~n19325 ;
  assign n19327 = n1296 & ~n19326 ;
  assign n19328 = n1300 & ~n19327 ;
  assign n19329 = n1304 & ~n19328 ;
  assign n19330 = n1308 & ~n19329 ;
  assign n19331 = n1312 & ~n19330 ;
  assign n19332 = n1316 & ~n19331 ;
  assign n19333 = n1320 & ~n19332 ;
  assign n19334 = n1324 & ~n19333 ;
  assign n19335 = n1328 & ~n19334 ;
  assign n19336 = n1332 & ~n19335 ;
  assign n19337 = n1336 & ~n19336 ;
  assign n19338 = n1340 & ~n19337 ;
  assign n19339 = n1344 & ~n19338 ;
  assign n19340 = n1348 & ~n19339 ;
  assign n19341 = n1352 & ~n19340 ;
  assign n19342 = n1356 & ~n19341 ;
  assign n19343 = n1360 & ~n19342 ;
  assign n19344 = n1364 & ~n19343 ;
  assign n19345 = n1368 & ~n19344 ;
  assign n19346 = n1372 & ~n19345 ;
  assign n19347 = n1376 & ~n19346 ;
  assign n19348 = n1380 & ~n19347 ;
  assign n19349 = n1384 & ~n19348 ;
  assign n19350 = n1388 & ~n19349 ;
  assign n19351 = n1392 & ~n19350 ;
  assign n19352 = n1396 & ~n19351 ;
  assign n19353 = n1400 & ~n19352 ;
  assign n19354 = n1404 & ~n19353 ;
  assign n19355 = n1408 & ~n19354 ;
  assign n19356 = n1412 & ~n19355 ;
  assign n19357 = n1416 & ~n19356 ;
  assign n19358 = n1420 & ~n19357 ;
  assign n19359 = n1424 & ~n19358 ;
  assign n19360 = n1428 & ~n19359 ;
  assign n19361 = n1432 & ~n19360 ;
  assign n19362 = n1436 & ~n19361 ;
  assign n19363 = n1440 & ~n19362 ;
  assign n19364 = n1444 & ~n19363 ;
  assign n19365 = n1448 & ~n19364 ;
  assign n19366 = n1452 & ~n19365 ;
  assign n19367 = n1456 & ~n19366 ;
  assign n19368 = n1460 & ~n19367 ;
  assign n19369 = n1464 & ~n19368 ;
  assign n19370 = n1468 & ~n19369 ;
  assign n19371 = n1472 & ~n19370 ;
  assign n19372 = n1476 & ~n19371 ;
  assign n19373 = n1480 & ~n19372 ;
  assign n19374 = n1484 & ~n19373 ;
  assign n19375 = n1488 & ~n19374 ;
  assign n19376 = n1492 & ~n19375 ;
  assign n19377 = n1496 & ~n19376 ;
  assign n19378 = n1500 & ~n19377 ;
  assign n19379 = n1504 & ~n19378 ;
  assign n19380 = n1508 & ~n19379 ;
  assign n19381 = n1512 & ~n19380 ;
  assign n19382 = n1516 & ~n19381 ;
  assign n19383 = n1520 & ~n19382 ;
  assign n19384 = n1524 & ~n19383 ;
  assign n19385 = n1528 & ~n19384 ;
  assign n19386 = n1532 & ~n19385 ;
  assign n19387 = ~x227 & ~n1534 ;
  assign n19388 = ~n19386 & n19387 ;
  assign n19391 = ~n19388 & ~x355 ;
  assign n19392 = ~n19390 & ~n19391 ;
  assign n19393 = n1204 & ~n1880 ;
  assign n19394 = n1209 & ~n19393 ;
  assign n19395 = n1213 & ~n19394 ;
  assign n19396 = n1217 & ~n19395 ;
  assign n19397 = n1221 & ~n19396 ;
  assign n19398 = n1225 & ~n19397 ;
  assign n19399 = n1229 & ~n19398 ;
  assign n19400 = n1233 & ~n19399 ;
  assign n19401 = n1237 & ~n19400 ;
  assign n19402 = n1241 & ~n19401 ;
  assign n19403 = n1245 & ~n19402 ;
  assign n19404 = n1249 & ~n19403 ;
  assign n19405 = n1253 & ~n19404 ;
  assign n19406 = n1257 & ~n19405 ;
  assign n19407 = n1261 & ~n19406 ;
  assign n19408 = n1265 & ~n19407 ;
  assign n19409 = n1269 & ~n19408 ;
  assign n19410 = n1273 & ~n19409 ;
  assign n19411 = n2566 & ~n19410 ;
  assign n19412 = n2568 & ~n19411 ;
  assign n19413 = n3105 & ~n19412 ;
  assign n19414 = n1625 & ~n19413 ;
  assign n19415 = n1629 & ~n19414 ;
  assign n19416 = n1633 & ~n19415 ;
  assign n19417 = n1637 & ~n19416 ;
  assign n19418 = n1641 & ~n19417 ;
  assign n19419 = n1645 & ~n19418 ;
  assign n19420 = n1649 & ~n19419 ;
  assign n19421 = n1653 & ~n19420 ;
  assign n19422 = n1657 & ~n19421 ;
  assign n19423 = n1661 & ~n19422 ;
  assign n19424 = n1665 & ~n19423 ;
  assign n19425 = n1669 & ~n19424 ;
  assign n19426 = n1673 & ~n19425 ;
  assign n19427 = n1677 & ~n19426 ;
  assign n19428 = n1681 & ~n19427 ;
  assign n19429 = n1685 & ~n19428 ;
  assign n19430 = n1689 & ~n19429 ;
  assign n19431 = n1693 & ~n19430 ;
  assign n19432 = n1697 & ~n19431 ;
  assign n19433 = n1701 & ~n19432 ;
  assign n19434 = n1705 & ~n19433 ;
  assign n19435 = n1709 & ~n19434 ;
  assign n19436 = n1713 & ~n19435 ;
  assign n19437 = n1717 & ~n19436 ;
  assign n19438 = n1721 & ~n19437 ;
  assign n19439 = n1725 & ~n19438 ;
  assign n19440 = n1729 & ~n19439 ;
  assign n19441 = n1733 & ~n19440 ;
  assign n19442 = n1737 & ~n19441 ;
  assign n19443 = n1741 & ~n19442 ;
  assign n19444 = n1745 & ~n19443 ;
  assign n19445 = n1749 & ~n19444 ;
  assign n19446 = n1753 & ~n19445 ;
  assign n19447 = n1757 & ~n19446 ;
  assign n19448 = n1761 & ~n19447 ;
  assign n19449 = n1765 & ~n19448 ;
  assign n19450 = n1769 & ~n19449 ;
  assign n19451 = n1773 & ~n19450 ;
  assign n19452 = n1777 & ~n19451 ;
  assign n19453 = n1781 & ~n19452 ;
  assign n19454 = n1785 & ~n19453 ;
  assign n19455 = n1789 & ~n19454 ;
  assign n19456 = n1793 & ~n19455 ;
  assign n19457 = n1797 & ~n19456 ;
  assign n19458 = n1801 & ~n19457 ;
  assign n19459 = n1805 & ~n19458 ;
  assign n19460 = n1809 & ~n19459 ;
  assign n19461 = n1813 & ~n19460 ;
  assign n19462 = n1817 & ~n19461 ;
  assign n19463 = n1821 & ~n19462 ;
  assign n19464 = n1825 & ~n19463 ;
  assign n19465 = n1829 & ~n19464 ;
  assign n19466 = n1833 & ~n19465 ;
  assign n19467 = n1837 & ~n19466 ;
  assign n19468 = n1841 & ~n19467 ;
  assign n19469 = n1845 & ~n19468 ;
  assign n19470 = n1849 & ~n19469 ;
  assign n19471 = n1853 & ~n19470 ;
  assign n19472 = n1857 & ~n19471 ;
  assign n19473 = n1861 & ~n19472 ;
  assign n19474 = n1865 & ~n19473 ;
  assign n19475 = n1869 & ~n19474 ;
  assign n19476 = n1873 & ~n19475 ;
  assign n19477 = x228 & ~n1875 ;
  assign n19478 = ~n19476 & n19477 ;
  assign n19566 = n19478 & x356 ;
  assign n19479 = n1543 & ~n2217 ;
  assign n19480 = n1548 & ~n19479 ;
  assign n19481 = n1552 & ~n19480 ;
  assign n19482 = n1556 & ~n19481 ;
  assign n19483 = n1560 & ~n19482 ;
  assign n19484 = n1564 & ~n19483 ;
  assign n19485 = n1568 & ~n19484 ;
  assign n19486 = n1572 & ~n19485 ;
  assign n19487 = n1576 & ~n19486 ;
  assign n19488 = n1580 & ~n19487 ;
  assign n19489 = n1584 & ~n19488 ;
  assign n19490 = n1588 & ~n19489 ;
  assign n19491 = n1592 & ~n19490 ;
  assign n19492 = n1596 & ~n19491 ;
  assign n19493 = n1600 & ~n19492 ;
  assign n19494 = n1604 & ~n19493 ;
  assign n19495 = n1608 & ~n19494 ;
  assign n19496 = n1612 & ~n19495 ;
  assign n19497 = n2656 & ~n19496 ;
  assign n19498 = n2658 & ~n19497 ;
  assign n19499 = n3192 & ~n19498 ;
  assign n19500 = n1962 & ~n19499 ;
  assign n19501 = n1966 & ~n19500 ;
  assign n19502 = n1970 & ~n19501 ;
  assign n19503 = n1974 & ~n19502 ;
  assign n19504 = n1978 & ~n19503 ;
  assign n19505 = n1982 & ~n19504 ;
  assign n19506 = n1986 & ~n19505 ;
  assign n19507 = n1990 & ~n19506 ;
  assign n19508 = n1994 & ~n19507 ;
  assign n19509 = n1998 & ~n19508 ;
  assign n19510 = n2002 & ~n19509 ;
  assign n19511 = n2006 & ~n19510 ;
  assign n19512 = n2010 & ~n19511 ;
  assign n19513 = n2014 & ~n19512 ;
  assign n19514 = n2018 & ~n19513 ;
  assign n19515 = n2022 & ~n19514 ;
  assign n19516 = n2026 & ~n19515 ;
  assign n19517 = n2030 & ~n19516 ;
  assign n19518 = n2034 & ~n19517 ;
  assign n19519 = n2038 & ~n19518 ;
  assign n19520 = n2042 & ~n19519 ;
  assign n19521 = n2046 & ~n19520 ;
  assign n19522 = n2050 & ~n19521 ;
  assign n19523 = n2054 & ~n19522 ;
  assign n19524 = n2058 & ~n19523 ;
  assign n19525 = n2062 & ~n19524 ;
  assign n19526 = n2066 & ~n19525 ;
  assign n19527 = n2070 & ~n19526 ;
  assign n19528 = n2074 & ~n19527 ;
  assign n19529 = n2078 & ~n19528 ;
  assign n19530 = n2082 & ~n19529 ;
  assign n19531 = n2086 & ~n19530 ;
  assign n19532 = n2090 & ~n19531 ;
  assign n19533 = n2094 & ~n19532 ;
  assign n19534 = n2098 & ~n19533 ;
  assign n19535 = n2102 & ~n19534 ;
  assign n19536 = n2106 & ~n19535 ;
  assign n19537 = n2110 & ~n19536 ;
  assign n19538 = n2114 & ~n19537 ;
  assign n19539 = n2118 & ~n19538 ;
  assign n19540 = n2122 & ~n19539 ;
  assign n19541 = n2126 & ~n19540 ;
  assign n19542 = n2130 & ~n19541 ;
  assign n19543 = n2134 & ~n19542 ;
  assign n19544 = n2138 & ~n19543 ;
  assign n19545 = n2142 & ~n19544 ;
  assign n19546 = n2146 & ~n19545 ;
  assign n19547 = n2150 & ~n19546 ;
  assign n19548 = n2154 & ~n19547 ;
  assign n19549 = n2158 & ~n19548 ;
  assign n19550 = n2162 & ~n19549 ;
  assign n19551 = n2166 & ~n19550 ;
  assign n19552 = n2170 & ~n19551 ;
  assign n19553 = n2174 & ~n19552 ;
  assign n19554 = n2178 & ~n19553 ;
  assign n19555 = n2182 & ~n19554 ;
  assign n19556 = n2186 & ~n19555 ;
  assign n19557 = n2190 & ~n19556 ;
  assign n19558 = n2194 & ~n19557 ;
  assign n19559 = n2198 & ~n19558 ;
  assign n19560 = n2202 & ~n19559 ;
  assign n19561 = n2206 & ~n19560 ;
  assign n19562 = n2210 & ~n19561 ;
  assign n19563 = ~x228 & ~n2212 ;
  assign n19564 = ~n19562 & n19563 ;
  assign n19567 = ~n19564 & ~x356 ;
  assign n19568 = ~n19566 & ~n19567 ;
  assign n19569 = ~n526 & n1884 ;
  assign n19570 = n1889 & ~n19569 ;
  assign n19571 = n1893 & ~n19570 ;
  assign n19572 = n1897 & ~n19571 ;
  assign n19573 = n1901 & ~n19572 ;
  assign n19574 = n1905 & ~n19573 ;
  assign n19575 = n1909 & ~n19574 ;
  assign n19576 = n1913 & ~n19575 ;
  assign n19577 = n1917 & ~n19576 ;
  assign n19578 = n1921 & ~n19577 ;
  assign n19579 = n1925 & ~n19578 ;
  assign n19580 = n1929 & ~n19579 ;
  assign n19581 = n1933 & ~n19580 ;
  assign n19582 = n1937 & ~n19581 ;
  assign n19583 = n1941 & ~n19582 ;
  assign n19584 = n1945 & ~n19583 ;
  assign n19585 = n1949 & ~n19584 ;
  assign n19586 = n1953 & ~n19585 ;
  assign n19587 = n2749 & ~n19586 ;
  assign n19588 = n263 & ~n19587 ;
  assign n19589 = n267 & ~n19588 ;
  assign n19590 = n271 & ~n19589 ;
  assign n19591 = n275 & ~n19590 ;
  assign n19592 = n279 & ~n19591 ;
  assign n19593 = n283 & ~n19592 ;
  assign n19594 = n287 & ~n19593 ;
  assign n19595 = n291 & ~n19594 ;
  assign n19596 = n295 & ~n19595 ;
  assign n19597 = n299 & ~n19596 ;
  assign n19598 = n303 & ~n19597 ;
  assign n19599 = n307 & ~n19598 ;
  assign n19600 = n311 & ~n19599 ;
  assign n19601 = n315 & ~n19600 ;
  assign n19602 = n319 & ~n19601 ;
  assign n19603 = n323 & ~n19602 ;
  assign n19604 = n327 & ~n19603 ;
  assign n19605 = n331 & ~n19604 ;
  assign n19606 = n335 & ~n19605 ;
  assign n19607 = n339 & ~n19606 ;
  assign n19608 = n343 & ~n19607 ;
  assign n19609 = n347 & ~n19608 ;
  assign n19610 = n351 & ~n19609 ;
  assign n19611 = n355 & ~n19610 ;
  assign n19612 = n359 & ~n19611 ;
  assign n19613 = n363 & ~n19612 ;
  assign n19614 = n367 & ~n19613 ;
  assign n19615 = n371 & ~n19614 ;
  assign n19616 = n375 & ~n19615 ;
  assign n19617 = n379 & ~n19616 ;
  assign n19618 = n383 & ~n19617 ;
  assign n19619 = n387 & ~n19618 ;
  assign n19620 = n391 & ~n19619 ;
  assign n19621 = n395 & ~n19620 ;
  assign n19622 = n399 & ~n19621 ;
  assign n19623 = n403 & ~n19622 ;
  assign n19624 = n407 & ~n19623 ;
  assign n19625 = n411 & ~n19624 ;
  assign n19626 = n415 & ~n19625 ;
  assign n19627 = n419 & ~n19626 ;
  assign n19628 = n423 & ~n19627 ;
  assign n19629 = n427 & ~n19628 ;
  assign n19630 = n431 & ~n19629 ;
  assign n19631 = n435 & ~n19630 ;
  assign n19632 = n439 & ~n19631 ;
  assign n19633 = n443 & ~n19632 ;
  assign n19634 = n447 & ~n19633 ;
  assign n19635 = n451 & ~n19634 ;
  assign n19636 = n455 & ~n19635 ;
  assign n19637 = n459 & ~n19636 ;
  assign n19638 = n463 & ~n19637 ;
  assign n19639 = n467 & ~n19638 ;
  assign n19640 = n471 & ~n19639 ;
  assign n19641 = n475 & ~n19640 ;
  assign n19642 = n479 & ~n19641 ;
  assign n19643 = n483 & ~n19642 ;
  assign n19644 = n487 & ~n19643 ;
  assign n19645 = n491 & ~n19644 ;
  assign n19646 = n495 & ~n19645 ;
  assign n19647 = n499 & ~n19646 ;
  assign n19648 = n503 & ~n19647 ;
  assign n19649 = n507 & ~n19648 ;
  assign n19650 = n511 & ~n19649 ;
  assign n19651 = n515 & ~n19650 ;
  assign n19652 = n519 & ~n19651 ;
  assign n19653 = x229 & ~n521 ;
  assign n19654 = ~n19652 & n19653 ;
  assign n19742 = n19654 & x357 ;
  assign n19655 = ~n865 & n2221 ;
  assign n19656 = n2226 & ~n19655 ;
  assign n19657 = n2230 & ~n19656 ;
  assign n19658 = n2234 & ~n19657 ;
  assign n19659 = n2238 & ~n19658 ;
  assign n19660 = n2242 & ~n19659 ;
  assign n19661 = n2246 & ~n19660 ;
  assign n19662 = n2250 & ~n19661 ;
  assign n19663 = n2254 & ~n19662 ;
  assign n19664 = n2258 & ~n19663 ;
  assign n19665 = n2262 & ~n19664 ;
  assign n19666 = n2266 & ~n19665 ;
  assign n19667 = n2270 & ~n19666 ;
  assign n19668 = n2274 & ~n19667 ;
  assign n19669 = n2278 & ~n19668 ;
  assign n19670 = n2282 & ~n19669 ;
  assign n19671 = n2286 & ~n19670 ;
  assign n19672 = n2290 & ~n19671 ;
  assign n19673 = n2836 & ~n19672 ;
  assign n19674 = n602 & ~n19673 ;
  assign n19675 = n606 & ~n19674 ;
  assign n19676 = n610 & ~n19675 ;
  assign n19677 = n614 & ~n19676 ;
  assign n19678 = n618 & ~n19677 ;
  assign n19679 = n622 & ~n19678 ;
  assign n19680 = n626 & ~n19679 ;
  assign n19681 = n630 & ~n19680 ;
  assign n19682 = n634 & ~n19681 ;
  assign n19683 = n638 & ~n19682 ;
  assign n19684 = n642 & ~n19683 ;
  assign n19685 = n646 & ~n19684 ;
  assign n19686 = n650 & ~n19685 ;
  assign n19687 = n654 & ~n19686 ;
  assign n19688 = n658 & ~n19687 ;
  assign n19689 = n662 & ~n19688 ;
  assign n19690 = n666 & ~n19689 ;
  assign n19691 = n670 & ~n19690 ;
  assign n19692 = n674 & ~n19691 ;
  assign n19693 = n678 & ~n19692 ;
  assign n19694 = n682 & ~n19693 ;
  assign n19695 = n686 & ~n19694 ;
  assign n19696 = n690 & ~n19695 ;
  assign n19697 = n694 & ~n19696 ;
  assign n19698 = n698 & ~n19697 ;
  assign n19699 = n702 & ~n19698 ;
  assign n19700 = n706 & ~n19699 ;
  assign n19701 = n710 & ~n19700 ;
  assign n19702 = n714 & ~n19701 ;
  assign n19703 = n718 & ~n19702 ;
  assign n19704 = n722 & ~n19703 ;
  assign n19705 = n726 & ~n19704 ;
  assign n19706 = n730 & ~n19705 ;
  assign n19707 = n734 & ~n19706 ;
  assign n19708 = n738 & ~n19707 ;
  assign n19709 = n742 & ~n19708 ;
  assign n19710 = n746 & ~n19709 ;
  assign n19711 = n750 & ~n19710 ;
  assign n19712 = n754 & ~n19711 ;
  assign n19713 = n758 & ~n19712 ;
  assign n19714 = n762 & ~n19713 ;
  assign n19715 = n766 & ~n19714 ;
  assign n19716 = n770 & ~n19715 ;
  assign n19717 = n774 & ~n19716 ;
  assign n19718 = n778 & ~n19717 ;
  assign n19719 = n782 & ~n19718 ;
  assign n19720 = n786 & ~n19719 ;
  assign n19721 = n790 & ~n19720 ;
  assign n19722 = n794 & ~n19721 ;
  assign n19723 = n798 & ~n19722 ;
  assign n19724 = n802 & ~n19723 ;
  assign n19725 = n806 & ~n19724 ;
  assign n19726 = n810 & ~n19725 ;
  assign n19727 = n814 & ~n19726 ;
  assign n19728 = n818 & ~n19727 ;
  assign n19729 = n822 & ~n19728 ;
  assign n19730 = n826 & ~n19729 ;
  assign n19731 = n830 & ~n19730 ;
  assign n19732 = n834 & ~n19731 ;
  assign n19733 = n838 & ~n19732 ;
  assign n19734 = n842 & ~n19733 ;
  assign n19735 = n846 & ~n19734 ;
  assign n19736 = n850 & ~n19735 ;
  assign n19737 = n854 & ~n19736 ;
  assign n19738 = n858 & ~n19737 ;
  assign n19739 = ~x229 & ~n860 ;
  assign n19740 = ~n19738 & n19739 ;
  assign n19743 = ~n19740 & ~x357 ;
  assign n19744 = ~n19742 & ~n19743 ;
  assign n19745 = n530 & ~n1208 ;
  assign n19746 = n535 & ~n19745 ;
  assign n19747 = n539 & ~n19746 ;
  assign n19748 = n543 & ~n19747 ;
  assign n19749 = n547 & ~n19748 ;
  assign n19750 = n551 & ~n19749 ;
  assign n19751 = n555 & ~n19750 ;
  assign n19752 = n559 & ~n19751 ;
  assign n19753 = n563 & ~n19752 ;
  assign n19754 = n567 & ~n19753 ;
  assign n19755 = n571 & ~n19754 ;
  assign n19756 = n575 & ~n19755 ;
  assign n19757 = n579 & ~n19756 ;
  assign n19758 = n583 & ~n19757 ;
  assign n19759 = n587 & ~n19758 ;
  assign n19760 = n591 & ~n19759 ;
  assign n19761 = n2382 & ~n19760 ;
  assign n19762 = n2384 & ~n19761 ;
  assign n19763 = n2927 & ~n19762 ;
  assign n19764 = n945 & ~n19763 ;
  assign n19765 = n949 & ~n19764 ;
  assign n19766 = n953 & ~n19765 ;
  assign n19767 = n957 & ~n19766 ;
  assign n19768 = n961 & ~n19767 ;
  assign n19769 = n965 & ~n19768 ;
  assign n19770 = n969 & ~n19769 ;
  assign n19771 = n973 & ~n19770 ;
  assign n19772 = n977 & ~n19771 ;
  assign n19773 = n981 & ~n19772 ;
  assign n19774 = n985 & ~n19773 ;
  assign n19775 = n989 & ~n19774 ;
  assign n19776 = n993 & ~n19775 ;
  assign n19777 = n997 & ~n19776 ;
  assign n19778 = n1001 & ~n19777 ;
  assign n19779 = n1005 & ~n19778 ;
  assign n19780 = n1009 & ~n19779 ;
  assign n19781 = n1013 & ~n19780 ;
  assign n19782 = n1017 & ~n19781 ;
  assign n19783 = n1021 & ~n19782 ;
  assign n19784 = n1025 & ~n19783 ;
  assign n19785 = n1029 & ~n19784 ;
  assign n19786 = n1033 & ~n19785 ;
  assign n19787 = n1037 & ~n19786 ;
  assign n19788 = n1041 & ~n19787 ;
  assign n19789 = n1045 & ~n19788 ;
  assign n19790 = n1049 & ~n19789 ;
  assign n19791 = n1053 & ~n19790 ;
  assign n19792 = n1057 & ~n19791 ;
  assign n19793 = n1061 & ~n19792 ;
  assign n19794 = n1065 & ~n19793 ;
  assign n19795 = n1069 & ~n19794 ;
  assign n19796 = n1073 & ~n19795 ;
  assign n19797 = n1077 & ~n19796 ;
  assign n19798 = n1081 & ~n19797 ;
  assign n19799 = n1085 & ~n19798 ;
  assign n19800 = n1089 & ~n19799 ;
  assign n19801 = n1093 & ~n19800 ;
  assign n19802 = n1097 & ~n19801 ;
  assign n19803 = n1101 & ~n19802 ;
  assign n19804 = n1105 & ~n19803 ;
  assign n19805 = n1109 & ~n19804 ;
  assign n19806 = n1113 & ~n19805 ;
  assign n19807 = n1117 & ~n19806 ;
  assign n19808 = n1121 & ~n19807 ;
  assign n19809 = n1125 & ~n19808 ;
  assign n19810 = n1129 & ~n19809 ;
  assign n19811 = n1133 & ~n19810 ;
  assign n19812 = n1137 & ~n19811 ;
  assign n19813 = n1141 & ~n19812 ;
  assign n19814 = n1145 & ~n19813 ;
  assign n19815 = n1149 & ~n19814 ;
  assign n19816 = n1153 & ~n19815 ;
  assign n19817 = n1157 & ~n19816 ;
  assign n19818 = n1161 & ~n19817 ;
  assign n19819 = n1165 & ~n19818 ;
  assign n19820 = n1169 & ~n19819 ;
  assign n19821 = n1173 & ~n19820 ;
  assign n19822 = n1177 & ~n19821 ;
  assign n19823 = n1181 & ~n19822 ;
  assign n19824 = n1185 & ~n19823 ;
  assign n19825 = n1189 & ~n19824 ;
  assign n19826 = n1193 & ~n19825 ;
  assign n19827 = n1197 & ~n19826 ;
  assign n19828 = n1201 & ~n19827 ;
  assign n19829 = x230 & ~n1203 ;
  assign n19830 = ~n19828 & n19829 ;
  assign n19918 = n19830 & x358 ;
  assign n19831 = n869 & ~n1547 ;
  assign n19832 = n874 & ~n19831 ;
  assign n19833 = n878 & ~n19832 ;
  assign n19834 = n882 & ~n19833 ;
  assign n19835 = n886 & ~n19834 ;
  assign n19836 = n890 & ~n19835 ;
  assign n19837 = n894 & ~n19836 ;
  assign n19838 = n898 & ~n19837 ;
  assign n19839 = n902 & ~n19838 ;
  assign n19840 = n906 & ~n19839 ;
  assign n19841 = n910 & ~n19840 ;
  assign n19842 = n914 & ~n19841 ;
  assign n19843 = n918 & ~n19842 ;
  assign n19844 = n922 & ~n19843 ;
  assign n19845 = n926 & ~n19844 ;
  assign n19846 = n930 & ~n19845 ;
  assign n19847 = n2472 & ~n19846 ;
  assign n19848 = n2474 & ~n19847 ;
  assign n19849 = n3014 & ~n19848 ;
  assign n19850 = n1284 & ~n19849 ;
  assign n19851 = n1288 & ~n19850 ;
  assign n19852 = n1292 & ~n19851 ;
  assign n19853 = n1296 & ~n19852 ;
  assign n19854 = n1300 & ~n19853 ;
  assign n19855 = n1304 & ~n19854 ;
  assign n19856 = n1308 & ~n19855 ;
  assign n19857 = n1312 & ~n19856 ;
  assign n19858 = n1316 & ~n19857 ;
  assign n19859 = n1320 & ~n19858 ;
  assign n19860 = n1324 & ~n19859 ;
  assign n19861 = n1328 & ~n19860 ;
  assign n19862 = n1332 & ~n19861 ;
  assign n19863 = n1336 & ~n19862 ;
  assign n19864 = n1340 & ~n19863 ;
  assign n19865 = n1344 & ~n19864 ;
  assign n19866 = n1348 & ~n19865 ;
  assign n19867 = n1352 & ~n19866 ;
  assign n19868 = n1356 & ~n19867 ;
  assign n19869 = n1360 & ~n19868 ;
  assign n19870 = n1364 & ~n19869 ;
  assign n19871 = n1368 & ~n19870 ;
  assign n19872 = n1372 & ~n19871 ;
  assign n19873 = n1376 & ~n19872 ;
  assign n19874 = n1380 & ~n19873 ;
  assign n19875 = n1384 & ~n19874 ;
  assign n19876 = n1388 & ~n19875 ;
  assign n19877 = n1392 & ~n19876 ;
  assign n19878 = n1396 & ~n19877 ;
  assign n19879 = n1400 & ~n19878 ;
  assign n19880 = n1404 & ~n19879 ;
  assign n19881 = n1408 & ~n19880 ;
  assign n19882 = n1412 & ~n19881 ;
  assign n19883 = n1416 & ~n19882 ;
  assign n19884 = n1420 & ~n19883 ;
  assign n19885 = n1424 & ~n19884 ;
  assign n19886 = n1428 & ~n19885 ;
  assign n19887 = n1432 & ~n19886 ;
  assign n19888 = n1436 & ~n19887 ;
  assign n19889 = n1440 & ~n19888 ;
  assign n19890 = n1444 & ~n19889 ;
  assign n19891 = n1448 & ~n19890 ;
  assign n19892 = n1452 & ~n19891 ;
  assign n19893 = n1456 & ~n19892 ;
  assign n19894 = n1460 & ~n19893 ;
  assign n19895 = n1464 & ~n19894 ;
  assign n19896 = n1468 & ~n19895 ;
  assign n19897 = n1472 & ~n19896 ;
  assign n19898 = n1476 & ~n19897 ;
  assign n19899 = n1480 & ~n19898 ;
  assign n19900 = n1484 & ~n19899 ;
  assign n19901 = n1488 & ~n19900 ;
  assign n19902 = n1492 & ~n19901 ;
  assign n19903 = n1496 & ~n19902 ;
  assign n19904 = n1500 & ~n19903 ;
  assign n19905 = n1504 & ~n19904 ;
  assign n19906 = n1508 & ~n19905 ;
  assign n19907 = n1512 & ~n19906 ;
  assign n19908 = n1516 & ~n19907 ;
  assign n19909 = n1520 & ~n19908 ;
  assign n19910 = n1524 & ~n19909 ;
  assign n19911 = n1528 & ~n19910 ;
  assign n19912 = n1532 & ~n19911 ;
  assign n19913 = n1536 & ~n19912 ;
  assign n19914 = n1540 & ~n19913 ;
  assign n19915 = ~x230 & ~n1542 ;
  assign n19916 = ~n19914 & n19915 ;
  assign n19919 = ~n19916 & ~x358 ;
  assign n19920 = ~n19918 & ~n19919 ;
  assign n19921 = n1212 & ~n1888 ;
  assign n19922 = n1217 & ~n19921 ;
  assign n19923 = n1221 & ~n19922 ;
  assign n19924 = n1225 & ~n19923 ;
  assign n19925 = n1229 & ~n19924 ;
  assign n19926 = n1233 & ~n19925 ;
  assign n19927 = n1237 & ~n19926 ;
  assign n19928 = n1241 & ~n19927 ;
  assign n19929 = n1245 & ~n19928 ;
  assign n19930 = n1249 & ~n19929 ;
  assign n19931 = n1253 & ~n19930 ;
  assign n19932 = n1257 & ~n19931 ;
  assign n19933 = n1261 & ~n19932 ;
  assign n19934 = n1265 & ~n19933 ;
  assign n19935 = n1269 & ~n19934 ;
  assign n19936 = n1273 & ~n19935 ;
  assign n19937 = n2566 & ~n19936 ;
  assign n19938 = n2568 & ~n19937 ;
  assign n19939 = n3105 & ~n19938 ;
  assign n19940 = n1625 & ~n19939 ;
  assign n19941 = n1629 & ~n19940 ;
  assign n19942 = n1633 & ~n19941 ;
  assign n19943 = n1637 & ~n19942 ;
  assign n19944 = n1641 & ~n19943 ;
  assign n19945 = n1645 & ~n19944 ;
  assign n19946 = n1649 & ~n19945 ;
  assign n19947 = n1653 & ~n19946 ;
  assign n19948 = n1657 & ~n19947 ;
  assign n19949 = n1661 & ~n19948 ;
  assign n19950 = n1665 & ~n19949 ;
  assign n19951 = n1669 & ~n19950 ;
  assign n19952 = n1673 & ~n19951 ;
  assign n19953 = n1677 & ~n19952 ;
  assign n19954 = n1681 & ~n19953 ;
  assign n19955 = n1685 & ~n19954 ;
  assign n19956 = n1689 & ~n19955 ;
  assign n19957 = n1693 & ~n19956 ;
  assign n19958 = n1697 & ~n19957 ;
  assign n19959 = n1701 & ~n19958 ;
  assign n19960 = n1705 & ~n19959 ;
  assign n19961 = n1709 & ~n19960 ;
  assign n19962 = n1713 & ~n19961 ;
  assign n19963 = n1717 & ~n19962 ;
  assign n19964 = n1721 & ~n19963 ;
  assign n19965 = n1725 & ~n19964 ;
  assign n19966 = n1729 & ~n19965 ;
  assign n19967 = n1733 & ~n19966 ;
  assign n19968 = n1737 & ~n19967 ;
  assign n19969 = n1741 & ~n19968 ;
  assign n19970 = n1745 & ~n19969 ;
  assign n19971 = n1749 & ~n19970 ;
  assign n19972 = n1753 & ~n19971 ;
  assign n19973 = n1757 & ~n19972 ;
  assign n19974 = n1761 & ~n19973 ;
  assign n19975 = n1765 & ~n19974 ;
  assign n19976 = n1769 & ~n19975 ;
  assign n19977 = n1773 & ~n19976 ;
  assign n19978 = n1777 & ~n19977 ;
  assign n19979 = n1781 & ~n19978 ;
  assign n19980 = n1785 & ~n19979 ;
  assign n19981 = n1789 & ~n19980 ;
  assign n19982 = n1793 & ~n19981 ;
  assign n19983 = n1797 & ~n19982 ;
  assign n19984 = n1801 & ~n19983 ;
  assign n19985 = n1805 & ~n19984 ;
  assign n19986 = n1809 & ~n19985 ;
  assign n19987 = n1813 & ~n19986 ;
  assign n19988 = n1817 & ~n19987 ;
  assign n19989 = n1821 & ~n19988 ;
  assign n19990 = n1825 & ~n19989 ;
  assign n19991 = n1829 & ~n19990 ;
  assign n19992 = n1833 & ~n19991 ;
  assign n19993 = n1837 & ~n19992 ;
  assign n19994 = n1841 & ~n19993 ;
  assign n19995 = n1845 & ~n19994 ;
  assign n19996 = n1849 & ~n19995 ;
  assign n19997 = n1853 & ~n19996 ;
  assign n19998 = n1857 & ~n19997 ;
  assign n19999 = n1861 & ~n19998 ;
  assign n20000 = n1865 & ~n19999 ;
  assign n20001 = n1869 & ~n20000 ;
  assign n20002 = n1873 & ~n20001 ;
  assign n20003 = n1877 & ~n20002 ;
  assign n20004 = n1881 & ~n20003 ;
  assign n20005 = x231 & ~n1883 ;
  assign n20006 = ~n20004 & n20005 ;
  assign n20094 = n20006 & x359 ;
  assign n20007 = n1551 & ~n2225 ;
  assign n20008 = n1556 & ~n20007 ;
  assign n20009 = n1560 & ~n20008 ;
  assign n20010 = n1564 & ~n20009 ;
  assign n20011 = n1568 & ~n20010 ;
  assign n20012 = n1572 & ~n20011 ;
  assign n20013 = n1576 & ~n20012 ;
  assign n20014 = n1580 & ~n20013 ;
  assign n20015 = n1584 & ~n20014 ;
  assign n20016 = n1588 & ~n20015 ;
  assign n20017 = n1592 & ~n20016 ;
  assign n20018 = n1596 & ~n20017 ;
  assign n20019 = n1600 & ~n20018 ;
  assign n20020 = n1604 & ~n20019 ;
  assign n20021 = n1608 & ~n20020 ;
  assign n20022 = n1612 & ~n20021 ;
  assign n20023 = n2656 & ~n20022 ;
  assign n20024 = n2658 & ~n20023 ;
  assign n20025 = n3192 & ~n20024 ;
  assign n20026 = n1962 & ~n20025 ;
  assign n20027 = n1966 & ~n20026 ;
  assign n20028 = n1970 & ~n20027 ;
  assign n20029 = n1974 & ~n20028 ;
  assign n20030 = n1978 & ~n20029 ;
  assign n20031 = n1982 & ~n20030 ;
  assign n20032 = n1986 & ~n20031 ;
  assign n20033 = n1990 & ~n20032 ;
  assign n20034 = n1994 & ~n20033 ;
  assign n20035 = n1998 & ~n20034 ;
  assign n20036 = n2002 & ~n20035 ;
  assign n20037 = n2006 & ~n20036 ;
  assign n20038 = n2010 & ~n20037 ;
  assign n20039 = n2014 & ~n20038 ;
  assign n20040 = n2018 & ~n20039 ;
  assign n20041 = n2022 & ~n20040 ;
  assign n20042 = n2026 & ~n20041 ;
  assign n20043 = n2030 & ~n20042 ;
  assign n20044 = n2034 & ~n20043 ;
  assign n20045 = n2038 & ~n20044 ;
  assign n20046 = n2042 & ~n20045 ;
  assign n20047 = n2046 & ~n20046 ;
  assign n20048 = n2050 & ~n20047 ;
  assign n20049 = n2054 & ~n20048 ;
  assign n20050 = n2058 & ~n20049 ;
  assign n20051 = n2062 & ~n20050 ;
  assign n20052 = n2066 & ~n20051 ;
  assign n20053 = n2070 & ~n20052 ;
  assign n20054 = n2074 & ~n20053 ;
  assign n20055 = n2078 & ~n20054 ;
  assign n20056 = n2082 & ~n20055 ;
  assign n20057 = n2086 & ~n20056 ;
  assign n20058 = n2090 & ~n20057 ;
  assign n20059 = n2094 & ~n20058 ;
  assign n20060 = n2098 & ~n20059 ;
  assign n20061 = n2102 & ~n20060 ;
  assign n20062 = n2106 & ~n20061 ;
  assign n20063 = n2110 & ~n20062 ;
  assign n20064 = n2114 & ~n20063 ;
  assign n20065 = n2118 & ~n20064 ;
  assign n20066 = n2122 & ~n20065 ;
  assign n20067 = n2126 & ~n20066 ;
  assign n20068 = n2130 & ~n20067 ;
  assign n20069 = n2134 & ~n20068 ;
  assign n20070 = n2138 & ~n20069 ;
  assign n20071 = n2142 & ~n20070 ;
  assign n20072 = n2146 & ~n20071 ;
  assign n20073 = n2150 & ~n20072 ;
  assign n20074 = n2154 & ~n20073 ;
  assign n20075 = n2158 & ~n20074 ;
  assign n20076 = n2162 & ~n20075 ;
  assign n20077 = n2166 & ~n20076 ;
  assign n20078 = n2170 & ~n20077 ;
  assign n20079 = n2174 & ~n20078 ;
  assign n20080 = n2178 & ~n20079 ;
  assign n20081 = n2182 & ~n20080 ;
  assign n20082 = n2186 & ~n20081 ;
  assign n20083 = n2190 & ~n20082 ;
  assign n20084 = n2194 & ~n20083 ;
  assign n20085 = n2198 & ~n20084 ;
  assign n20086 = n2202 & ~n20085 ;
  assign n20087 = n2206 & ~n20086 ;
  assign n20088 = n2210 & ~n20087 ;
  assign n20089 = n2214 & ~n20088 ;
  assign n20090 = n2218 & ~n20089 ;
  assign n20091 = ~x231 & ~n2220 ;
  assign n20092 = ~n20090 & n20091 ;
  assign n20095 = ~n20092 & ~x359 ;
  assign n20096 = ~n20094 & ~n20095 ;
  assign n20097 = ~n534 & n1892 ;
  assign n20098 = n1897 & ~n20097 ;
  assign n20099 = n1901 & ~n20098 ;
  assign n20100 = n1905 & ~n20099 ;
  assign n20101 = n1909 & ~n20100 ;
  assign n20102 = n1913 & ~n20101 ;
  assign n20103 = n1917 & ~n20102 ;
  assign n20104 = n1921 & ~n20103 ;
  assign n20105 = n1925 & ~n20104 ;
  assign n20106 = n1929 & ~n20105 ;
  assign n20107 = n1933 & ~n20106 ;
  assign n20108 = n1937 & ~n20107 ;
  assign n20109 = n1941 & ~n20108 ;
  assign n20110 = n1945 & ~n20109 ;
  assign n20111 = n1949 & ~n20110 ;
  assign n20112 = n1953 & ~n20111 ;
  assign n20113 = n2749 & ~n20112 ;
  assign n20114 = n263 & ~n20113 ;
  assign n20115 = n267 & ~n20114 ;
  assign n20116 = n271 & ~n20115 ;
  assign n20117 = n275 & ~n20116 ;
  assign n20118 = n279 & ~n20117 ;
  assign n20119 = n283 & ~n20118 ;
  assign n20120 = n287 & ~n20119 ;
  assign n20121 = n291 & ~n20120 ;
  assign n20122 = n295 & ~n20121 ;
  assign n20123 = n299 & ~n20122 ;
  assign n20124 = n303 & ~n20123 ;
  assign n20125 = n307 & ~n20124 ;
  assign n20126 = n311 & ~n20125 ;
  assign n20127 = n315 & ~n20126 ;
  assign n20128 = n319 & ~n20127 ;
  assign n20129 = n323 & ~n20128 ;
  assign n20130 = n327 & ~n20129 ;
  assign n20131 = n331 & ~n20130 ;
  assign n20132 = n335 & ~n20131 ;
  assign n20133 = n339 & ~n20132 ;
  assign n20134 = n343 & ~n20133 ;
  assign n20135 = n347 & ~n20134 ;
  assign n20136 = n351 & ~n20135 ;
  assign n20137 = n355 & ~n20136 ;
  assign n20138 = n359 & ~n20137 ;
  assign n20139 = n363 & ~n20138 ;
  assign n20140 = n367 & ~n20139 ;
  assign n20141 = n371 & ~n20140 ;
  assign n20142 = n375 & ~n20141 ;
  assign n20143 = n379 & ~n20142 ;
  assign n20144 = n383 & ~n20143 ;
  assign n20145 = n387 & ~n20144 ;
  assign n20146 = n391 & ~n20145 ;
  assign n20147 = n395 & ~n20146 ;
  assign n20148 = n399 & ~n20147 ;
  assign n20149 = n403 & ~n20148 ;
  assign n20150 = n407 & ~n20149 ;
  assign n20151 = n411 & ~n20150 ;
  assign n20152 = n415 & ~n20151 ;
  assign n20153 = n419 & ~n20152 ;
  assign n20154 = n423 & ~n20153 ;
  assign n20155 = n427 & ~n20154 ;
  assign n20156 = n431 & ~n20155 ;
  assign n20157 = n435 & ~n20156 ;
  assign n20158 = n439 & ~n20157 ;
  assign n20159 = n443 & ~n20158 ;
  assign n20160 = n447 & ~n20159 ;
  assign n20161 = n451 & ~n20160 ;
  assign n20162 = n455 & ~n20161 ;
  assign n20163 = n459 & ~n20162 ;
  assign n20164 = n463 & ~n20163 ;
  assign n20165 = n467 & ~n20164 ;
  assign n20166 = n471 & ~n20165 ;
  assign n20167 = n475 & ~n20166 ;
  assign n20168 = n479 & ~n20167 ;
  assign n20169 = n483 & ~n20168 ;
  assign n20170 = n487 & ~n20169 ;
  assign n20171 = n491 & ~n20170 ;
  assign n20172 = n495 & ~n20171 ;
  assign n20173 = n499 & ~n20172 ;
  assign n20174 = n503 & ~n20173 ;
  assign n20175 = n507 & ~n20174 ;
  assign n20176 = n511 & ~n20175 ;
  assign n20177 = n515 & ~n20176 ;
  assign n20178 = n519 & ~n20177 ;
  assign n20179 = n523 & ~n20178 ;
  assign n20180 = n527 & ~n20179 ;
  assign n20181 = x232 & ~n529 ;
  assign n20182 = ~n20180 & n20181 ;
  assign n20270 = n20182 & x360 ;
  assign n20183 = ~n873 & n2229 ;
  assign n20184 = n2234 & ~n20183 ;
  assign n20185 = n2238 & ~n20184 ;
  assign n20186 = n2242 & ~n20185 ;
  assign n20187 = n2246 & ~n20186 ;
  assign n20188 = n2250 & ~n20187 ;
  assign n20189 = n2254 & ~n20188 ;
  assign n20190 = n2258 & ~n20189 ;
  assign n20191 = n2262 & ~n20190 ;
  assign n20192 = n2266 & ~n20191 ;
  assign n20193 = n2270 & ~n20192 ;
  assign n20194 = n2274 & ~n20193 ;
  assign n20195 = n2278 & ~n20194 ;
  assign n20196 = n2282 & ~n20195 ;
  assign n20197 = n2286 & ~n20196 ;
  assign n20198 = n2290 & ~n20197 ;
  assign n20199 = n2836 & ~n20198 ;
  assign n20200 = n602 & ~n20199 ;
  assign n20201 = n606 & ~n20200 ;
  assign n20202 = n610 & ~n20201 ;
  assign n20203 = n614 & ~n20202 ;
  assign n20204 = n618 & ~n20203 ;
  assign n20205 = n622 & ~n20204 ;
  assign n20206 = n626 & ~n20205 ;
  assign n20207 = n630 & ~n20206 ;
  assign n20208 = n634 & ~n20207 ;
  assign n20209 = n638 & ~n20208 ;
  assign n20210 = n642 & ~n20209 ;
  assign n20211 = n646 & ~n20210 ;
  assign n20212 = n650 & ~n20211 ;
  assign n20213 = n654 & ~n20212 ;
  assign n20214 = n658 & ~n20213 ;
  assign n20215 = n662 & ~n20214 ;
  assign n20216 = n666 & ~n20215 ;
  assign n20217 = n670 & ~n20216 ;
  assign n20218 = n674 & ~n20217 ;
  assign n20219 = n678 & ~n20218 ;
  assign n20220 = n682 & ~n20219 ;
  assign n20221 = n686 & ~n20220 ;
  assign n20222 = n690 & ~n20221 ;
  assign n20223 = n694 & ~n20222 ;
  assign n20224 = n698 & ~n20223 ;
  assign n20225 = n702 & ~n20224 ;
  assign n20226 = n706 & ~n20225 ;
  assign n20227 = n710 & ~n20226 ;
  assign n20228 = n714 & ~n20227 ;
  assign n20229 = n718 & ~n20228 ;
  assign n20230 = n722 & ~n20229 ;
  assign n20231 = n726 & ~n20230 ;
  assign n20232 = n730 & ~n20231 ;
  assign n20233 = n734 & ~n20232 ;
  assign n20234 = n738 & ~n20233 ;
  assign n20235 = n742 & ~n20234 ;
  assign n20236 = n746 & ~n20235 ;
  assign n20237 = n750 & ~n20236 ;
  assign n20238 = n754 & ~n20237 ;
  assign n20239 = n758 & ~n20238 ;
  assign n20240 = n762 & ~n20239 ;
  assign n20241 = n766 & ~n20240 ;
  assign n20242 = n770 & ~n20241 ;
  assign n20243 = n774 & ~n20242 ;
  assign n20244 = n778 & ~n20243 ;
  assign n20245 = n782 & ~n20244 ;
  assign n20246 = n786 & ~n20245 ;
  assign n20247 = n790 & ~n20246 ;
  assign n20248 = n794 & ~n20247 ;
  assign n20249 = n798 & ~n20248 ;
  assign n20250 = n802 & ~n20249 ;
  assign n20251 = n806 & ~n20250 ;
  assign n20252 = n810 & ~n20251 ;
  assign n20253 = n814 & ~n20252 ;
  assign n20254 = n818 & ~n20253 ;
  assign n20255 = n822 & ~n20254 ;
  assign n20256 = n826 & ~n20255 ;
  assign n20257 = n830 & ~n20256 ;
  assign n20258 = n834 & ~n20257 ;
  assign n20259 = n838 & ~n20258 ;
  assign n20260 = n842 & ~n20259 ;
  assign n20261 = n846 & ~n20260 ;
  assign n20262 = n850 & ~n20261 ;
  assign n20263 = n854 & ~n20262 ;
  assign n20264 = n858 & ~n20263 ;
  assign n20265 = n862 & ~n20264 ;
  assign n20266 = n866 & ~n20265 ;
  assign n20267 = ~x232 & ~n868 ;
  assign n20268 = ~n20266 & n20267 ;
  assign n20271 = ~n20268 & ~x360 ;
  assign n20272 = ~n20270 & ~n20271 ;
  assign n20273 = n538 & ~n1216 ;
  assign n20274 = n543 & ~n20273 ;
  assign n20275 = n547 & ~n20274 ;
  assign n20276 = n551 & ~n20275 ;
  assign n20277 = n555 & ~n20276 ;
  assign n20278 = n559 & ~n20277 ;
  assign n20279 = n563 & ~n20278 ;
  assign n20280 = n567 & ~n20279 ;
  assign n20281 = n571 & ~n20280 ;
  assign n20282 = n575 & ~n20281 ;
  assign n20283 = n579 & ~n20282 ;
  assign n20284 = n583 & ~n20283 ;
  assign n20285 = n587 & ~n20284 ;
  assign n20286 = n591 & ~n20285 ;
  assign n20287 = n2382 & ~n20286 ;
  assign n20288 = n2384 & ~n20287 ;
  assign n20289 = n2927 & ~n20288 ;
  assign n20290 = n945 & ~n20289 ;
  assign n20291 = n949 & ~n20290 ;
  assign n20292 = n953 & ~n20291 ;
  assign n20293 = n957 & ~n20292 ;
  assign n20294 = n961 & ~n20293 ;
  assign n20295 = n965 & ~n20294 ;
  assign n20296 = n969 & ~n20295 ;
  assign n20297 = n973 & ~n20296 ;
  assign n20298 = n977 & ~n20297 ;
  assign n20299 = n981 & ~n20298 ;
  assign n20300 = n985 & ~n20299 ;
  assign n20301 = n989 & ~n20300 ;
  assign n20302 = n993 & ~n20301 ;
  assign n20303 = n997 & ~n20302 ;
  assign n20304 = n1001 & ~n20303 ;
  assign n20305 = n1005 & ~n20304 ;
  assign n20306 = n1009 & ~n20305 ;
  assign n20307 = n1013 & ~n20306 ;
  assign n20308 = n1017 & ~n20307 ;
  assign n20309 = n1021 & ~n20308 ;
  assign n20310 = n1025 & ~n20309 ;
  assign n20311 = n1029 & ~n20310 ;
  assign n20312 = n1033 & ~n20311 ;
  assign n20313 = n1037 & ~n20312 ;
  assign n20314 = n1041 & ~n20313 ;
  assign n20315 = n1045 & ~n20314 ;
  assign n20316 = n1049 & ~n20315 ;
  assign n20317 = n1053 & ~n20316 ;
  assign n20318 = n1057 & ~n20317 ;
  assign n20319 = n1061 & ~n20318 ;
  assign n20320 = n1065 & ~n20319 ;
  assign n20321 = n1069 & ~n20320 ;
  assign n20322 = n1073 & ~n20321 ;
  assign n20323 = n1077 & ~n20322 ;
  assign n20324 = n1081 & ~n20323 ;
  assign n20325 = n1085 & ~n20324 ;
  assign n20326 = n1089 & ~n20325 ;
  assign n20327 = n1093 & ~n20326 ;
  assign n20328 = n1097 & ~n20327 ;
  assign n20329 = n1101 & ~n20328 ;
  assign n20330 = n1105 & ~n20329 ;
  assign n20331 = n1109 & ~n20330 ;
  assign n20332 = n1113 & ~n20331 ;
  assign n20333 = n1117 & ~n20332 ;
  assign n20334 = n1121 & ~n20333 ;
  assign n20335 = n1125 & ~n20334 ;
  assign n20336 = n1129 & ~n20335 ;
  assign n20337 = n1133 & ~n20336 ;
  assign n20338 = n1137 & ~n20337 ;
  assign n20339 = n1141 & ~n20338 ;
  assign n20340 = n1145 & ~n20339 ;
  assign n20341 = n1149 & ~n20340 ;
  assign n20342 = n1153 & ~n20341 ;
  assign n20343 = n1157 & ~n20342 ;
  assign n20344 = n1161 & ~n20343 ;
  assign n20345 = n1165 & ~n20344 ;
  assign n20346 = n1169 & ~n20345 ;
  assign n20347 = n1173 & ~n20346 ;
  assign n20348 = n1177 & ~n20347 ;
  assign n20349 = n1181 & ~n20348 ;
  assign n20350 = n1185 & ~n20349 ;
  assign n20351 = n1189 & ~n20350 ;
  assign n20352 = n1193 & ~n20351 ;
  assign n20353 = n1197 & ~n20352 ;
  assign n20354 = n1201 & ~n20353 ;
  assign n20355 = n1205 & ~n20354 ;
  assign n20356 = n1209 & ~n20355 ;
  assign n20357 = x233 & ~n1211 ;
  assign n20358 = ~n20356 & n20357 ;
  assign n20446 = n20358 & x361 ;
  assign n20359 = n877 & ~n1555 ;
  assign n20360 = n882 & ~n20359 ;
  assign n20361 = n886 & ~n20360 ;
  assign n20362 = n890 & ~n20361 ;
  assign n20363 = n894 & ~n20362 ;
  assign n20364 = n898 & ~n20363 ;
  assign n20365 = n902 & ~n20364 ;
  assign n20366 = n906 & ~n20365 ;
  assign n20367 = n910 & ~n20366 ;
  assign n20368 = n914 & ~n20367 ;
  assign n20369 = n918 & ~n20368 ;
  assign n20370 = n922 & ~n20369 ;
  assign n20371 = n926 & ~n20370 ;
  assign n20372 = n930 & ~n20371 ;
  assign n20373 = n2472 & ~n20372 ;
  assign n20374 = n2474 & ~n20373 ;
  assign n20375 = n3014 & ~n20374 ;
  assign n20376 = n1284 & ~n20375 ;
  assign n20377 = n1288 & ~n20376 ;
  assign n20378 = n1292 & ~n20377 ;
  assign n20379 = n1296 & ~n20378 ;
  assign n20380 = n1300 & ~n20379 ;
  assign n20381 = n1304 & ~n20380 ;
  assign n20382 = n1308 & ~n20381 ;
  assign n20383 = n1312 & ~n20382 ;
  assign n20384 = n1316 & ~n20383 ;
  assign n20385 = n1320 & ~n20384 ;
  assign n20386 = n1324 & ~n20385 ;
  assign n20387 = n1328 & ~n20386 ;
  assign n20388 = n1332 & ~n20387 ;
  assign n20389 = n1336 & ~n20388 ;
  assign n20390 = n1340 & ~n20389 ;
  assign n20391 = n1344 & ~n20390 ;
  assign n20392 = n1348 & ~n20391 ;
  assign n20393 = n1352 & ~n20392 ;
  assign n20394 = n1356 & ~n20393 ;
  assign n20395 = n1360 & ~n20394 ;
  assign n20396 = n1364 & ~n20395 ;
  assign n20397 = n1368 & ~n20396 ;
  assign n20398 = n1372 & ~n20397 ;
  assign n20399 = n1376 & ~n20398 ;
  assign n20400 = n1380 & ~n20399 ;
  assign n20401 = n1384 & ~n20400 ;
  assign n20402 = n1388 & ~n20401 ;
  assign n20403 = n1392 & ~n20402 ;
  assign n20404 = n1396 & ~n20403 ;
  assign n20405 = n1400 & ~n20404 ;
  assign n20406 = n1404 & ~n20405 ;
  assign n20407 = n1408 & ~n20406 ;
  assign n20408 = n1412 & ~n20407 ;
  assign n20409 = n1416 & ~n20408 ;
  assign n20410 = n1420 & ~n20409 ;
  assign n20411 = n1424 & ~n20410 ;
  assign n20412 = n1428 & ~n20411 ;
  assign n20413 = n1432 & ~n20412 ;
  assign n20414 = n1436 & ~n20413 ;
  assign n20415 = n1440 & ~n20414 ;
  assign n20416 = n1444 & ~n20415 ;
  assign n20417 = n1448 & ~n20416 ;
  assign n20418 = n1452 & ~n20417 ;
  assign n20419 = n1456 & ~n20418 ;
  assign n20420 = n1460 & ~n20419 ;
  assign n20421 = n1464 & ~n20420 ;
  assign n20422 = n1468 & ~n20421 ;
  assign n20423 = n1472 & ~n20422 ;
  assign n20424 = n1476 & ~n20423 ;
  assign n20425 = n1480 & ~n20424 ;
  assign n20426 = n1484 & ~n20425 ;
  assign n20427 = n1488 & ~n20426 ;
  assign n20428 = n1492 & ~n20427 ;
  assign n20429 = n1496 & ~n20428 ;
  assign n20430 = n1500 & ~n20429 ;
  assign n20431 = n1504 & ~n20430 ;
  assign n20432 = n1508 & ~n20431 ;
  assign n20433 = n1512 & ~n20432 ;
  assign n20434 = n1516 & ~n20433 ;
  assign n20435 = n1520 & ~n20434 ;
  assign n20436 = n1524 & ~n20435 ;
  assign n20437 = n1528 & ~n20436 ;
  assign n20438 = n1532 & ~n20437 ;
  assign n20439 = n1536 & ~n20438 ;
  assign n20440 = n1540 & ~n20439 ;
  assign n20441 = n1544 & ~n20440 ;
  assign n20442 = n1548 & ~n20441 ;
  assign n20443 = ~x233 & ~n1550 ;
  assign n20444 = ~n20442 & n20443 ;
  assign n20447 = ~n20444 & ~x361 ;
  assign n20448 = ~n20446 & ~n20447 ;
  assign n20449 = n1220 & ~n1896 ;
  assign n20450 = n1225 & ~n20449 ;
  assign n20451 = n1229 & ~n20450 ;
  assign n20452 = n1233 & ~n20451 ;
  assign n20453 = n1237 & ~n20452 ;
  assign n20454 = n1241 & ~n20453 ;
  assign n20455 = n1245 & ~n20454 ;
  assign n20456 = n1249 & ~n20455 ;
  assign n20457 = n1253 & ~n20456 ;
  assign n20458 = n1257 & ~n20457 ;
  assign n20459 = n1261 & ~n20458 ;
  assign n20460 = n1265 & ~n20459 ;
  assign n20461 = n1269 & ~n20460 ;
  assign n20462 = n1273 & ~n20461 ;
  assign n20463 = n2566 & ~n20462 ;
  assign n20464 = n2568 & ~n20463 ;
  assign n20465 = n3105 & ~n20464 ;
  assign n20466 = n1625 & ~n20465 ;
  assign n20467 = n1629 & ~n20466 ;
  assign n20468 = n1633 & ~n20467 ;
  assign n20469 = n1637 & ~n20468 ;
  assign n20470 = n1641 & ~n20469 ;
  assign n20471 = n1645 & ~n20470 ;
  assign n20472 = n1649 & ~n20471 ;
  assign n20473 = n1653 & ~n20472 ;
  assign n20474 = n1657 & ~n20473 ;
  assign n20475 = n1661 & ~n20474 ;
  assign n20476 = n1665 & ~n20475 ;
  assign n20477 = n1669 & ~n20476 ;
  assign n20478 = n1673 & ~n20477 ;
  assign n20479 = n1677 & ~n20478 ;
  assign n20480 = n1681 & ~n20479 ;
  assign n20481 = n1685 & ~n20480 ;
  assign n20482 = n1689 & ~n20481 ;
  assign n20483 = n1693 & ~n20482 ;
  assign n20484 = n1697 & ~n20483 ;
  assign n20485 = n1701 & ~n20484 ;
  assign n20486 = n1705 & ~n20485 ;
  assign n20487 = n1709 & ~n20486 ;
  assign n20488 = n1713 & ~n20487 ;
  assign n20489 = n1717 & ~n20488 ;
  assign n20490 = n1721 & ~n20489 ;
  assign n20491 = n1725 & ~n20490 ;
  assign n20492 = n1729 & ~n20491 ;
  assign n20493 = n1733 & ~n20492 ;
  assign n20494 = n1737 & ~n20493 ;
  assign n20495 = n1741 & ~n20494 ;
  assign n20496 = n1745 & ~n20495 ;
  assign n20497 = n1749 & ~n20496 ;
  assign n20498 = n1753 & ~n20497 ;
  assign n20499 = n1757 & ~n20498 ;
  assign n20500 = n1761 & ~n20499 ;
  assign n20501 = n1765 & ~n20500 ;
  assign n20502 = n1769 & ~n20501 ;
  assign n20503 = n1773 & ~n20502 ;
  assign n20504 = n1777 & ~n20503 ;
  assign n20505 = n1781 & ~n20504 ;
  assign n20506 = n1785 & ~n20505 ;
  assign n20507 = n1789 & ~n20506 ;
  assign n20508 = n1793 & ~n20507 ;
  assign n20509 = n1797 & ~n20508 ;
  assign n20510 = n1801 & ~n20509 ;
  assign n20511 = n1805 & ~n20510 ;
  assign n20512 = n1809 & ~n20511 ;
  assign n20513 = n1813 & ~n20512 ;
  assign n20514 = n1817 & ~n20513 ;
  assign n20515 = n1821 & ~n20514 ;
  assign n20516 = n1825 & ~n20515 ;
  assign n20517 = n1829 & ~n20516 ;
  assign n20518 = n1833 & ~n20517 ;
  assign n20519 = n1837 & ~n20518 ;
  assign n20520 = n1841 & ~n20519 ;
  assign n20521 = n1845 & ~n20520 ;
  assign n20522 = n1849 & ~n20521 ;
  assign n20523 = n1853 & ~n20522 ;
  assign n20524 = n1857 & ~n20523 ;
  assign n20525 = n1861 & ~n20524 ;
  assign n20526 = n1865 & ~n20525 ;
  assign n20527 = n1869 & ~n20526 ;
  assign n20528 = n1873 & ~n20527 ;
  assign n20529 = n1877 & ~n20528 ;
  assign n20530 = n1881 & ~n20529 ;
  assign n20531 = n1885 & ~n20530 ;
  assign n20532 = n1889 & ~n20531 ;
  assign n20533 = x234 & ~n1891 ;
  assign n20534 = ~n20532 & n20533 ;
  assign n20622 = n20534 & x362 ;
  assign n20535 = n1559 & ~n2233 ;
  assign n20536 = n1564 & ~n20535 ;
  assign n20537 = n1568 & ~n20536 ;
  assign n20538 = n1572 & ~n20537 ;
  assign n20539 = n1576 & ~n20538 ;
  assign n20540 = n1580 & ~n20539 ;
  assign n20541 = n1584 & ~n20540 ;
  assign n20542 = n1588 & ~n20541 ;
  assign n20543 = n1592 & ~n20542 ;
  assign n20544 = n1596 & ~n20543 ;
  assign n20545 = n1600 & ~n20544 ;
  assign n20546 = n1604 & ~n20545 ;
  assign n20547 = n1608 & ~n20546 ;
  assign n20548 = n1612 & ~n20547 ;
  assign n20549 = n2656 & ~n20548 ;
  assign n20550 = n2658 & ~n20549 ;
  assign n20551 = n3192 & ~n20550 ;
  assign n20552 = n1962 & ~n20551 ;
  assign n20553 = n1966 & ~n20552 ;
  assign n20554 = n1970 & ~n20553 ;
  assign n20555 = n1974 & ~n20554 ;
  assign n20556 = n1978 & ~n20555 ;
  assign n20557 = n1982 & ~n20556 ;
  assign n20558 = n1986 & ~n20557 ;
  assign n20559 = n1990 & ~n20558 ;
  assign n20560 = n1994 & ~n20559 ;
  assign n20561 = n1998 & ~n20560 ;
  assign n20562 = n2002 & ~n20561 ;
  assign n20563 = n2006 & ~n20562 ;
  assign n20564 = n2010 & ~n20563 ;
  assign n20565 = n2014 & ~n20564 ;
  assign n20566 = n2018 & ~n20565 ;
  assign n20567 = n2022 & ~n20566 ;
  assign n20568 = n2026 & ~n20567 ;
  assign n20569 = n2030 & ~n20568 ;
  assign n20570 = n2034 & ~n20569 ;
  assign n20571 = n2038 & ~n20570 ;
  assign n20572 = n2042 & ~n20571 ;
  assign n20573 = n2046 & ~n20572 ;
  assign n20574 = n2050 & ~n20573 ;
  assign n20575 = n2054 & ~n20574 ;
  assign n20576 = n2058 & ~n20575 ;
  assign n20577 = n2062 & ~n20576 ;
  assign n20578 = n2066 & ~n20577 ;
  assign n20579 = n2070 & ~n20578 ;
  assign n20580 = n2074 & ~n20579 ;
  assign n20581 = n2078 & ~n20580 ;
  assign n20582 = n2082 & ~n20581 ;
  assign n20583 = n2086 & ~n20582 ;
  assign n20584 = n2090 & ~n20583 ;
  assign n20585 = n2094 & ~n20584 ;
  assign n20586 = n2098 & ~n20585 ;
  assign n20587 = n2102 & ~n20586 ;
  assign n20588 = n2106 & ~n20587 ;
  assign n20589 = n2110 & ~n20588 ;
  assign n20590 = n2114 & ~n20589 ;
  assign n20591 = n2118 & ~n20590 ;
  assign n20592 = n2122 & ~n20591 ;
  assign n20593 = n2126 & ~n20592 ;
  assign n20594 = n2130 & ~n20593 ;
  assign n20595 = n2134 & ~n20594 ;
  assign n20596 = n2138 & ~n20595 ;
  assign n20597 = n2142 & ~n20596 ;
  assign n20598 = n2146 & ~n20597 ;
  assign n20599 = n2150 & ~n20598 ;
  assign n20600 = n2154 & ~n20599 ;
  assign n20601 = n2158 & ~n20600 ;
  assign n20602 = n2162 & ~n20601 ;
  assign n20603 = n2166 & ~n20602 ;
  assign n20604 = n2170 & ~n20603 ;
  assign n20605 = n2174 & ~n20604 ;
  assign n20606 = n2178 & ~n20605 ;
  assign n20607 = n2182 & ~n20606 ;
  assign n20608 = n2186 & ~n20607 ;
  assign n20609 = n2190 & ~n20608 ;
  assign n20610 = n2194 & ~n20609 ;
  assign n20611 = n2198 & ~n20610 ;
  assign n20612 = n2202 & ~n20611 ;
  assign n20613 = n2206 & ~n20612 ;
  assign n20614 = n2210 & ~n20613 ;
  assign n20615 = n2214 & ~n20614 ;
  assign n20616 = n2218 & ~n20615 ;
  assign n20617 = n2222 & ~n20616 ;
  assign n20618 = n2226 & ~n20617 ;
  assign n20619 = ~x234 & ~n2228 ;
  assign n20620 = ~n20618 & n20619 ;
  assign n20623 = ~n20620 & ~x362 ;
  assign n20624 = ~n20622 & ~n20623 ;
  assign n20625 = ~n542 & n1900 ;
  assign n20626 = n1905 & ~n20625 ;
  assign n20627 = n1909 & ~n20626 ;
  assign n20628 = n1913 & ~n20627 ;
  assign n20629 = n1917 & ~n20628 ;
  assign n20630 = n1921 & ~n20629 ;
  assign n20631 = n1925 & ~n20630 ;
  assign n20632 = n1929 & ~n20631 ;
  assign n20633 = n1933 & ~n20632 ;
  assign n20634 = n1937 & ~n20633 ;
  assign n20635 = n1941 & ~n20634 ;
  assign n20636 = n1945 & ~n20635 ;
  assign n20637 = n1949 & ~n20636 ;
  assign n20638 = n1953 & ~n20637 ;
  assign n20639 = n2749 & ~n20638 ;
  assign n20640 = n263 & ~n20639 ;
  assign n20641 = n267 & ~n20640 ;
  assign n20642 = n271 & ~n20641 ;
  assign n20643 = n275 & ~n20642 ;
  assign n20644 = n279 & ~n20643 ;
  assign n20645 = n283 & ~n20644 ;
  assign n20646 = n287 & ~n20645 ;
  assign n20647 = n291 & ~n20646 ;
  assign n20648 = n295 & ~n20647 ;
  assign n20649 = n299 & ~n20648 ;
  assign n20650 = n303 & ~n20649 ;
  assign n20651 = n307 & ~n20650 ;
  assign n20652 = n311 & ~n20651 ;
  assign n20653 = n315 & ~n20652 ;
  assign n20654 = n319 & ~n20653 ;
  assign n20655 = n323 & ~n20654 ;
  assign n20656 = n327 & ~n20655 ;
  assign n20657 = n331 & ~n20656 ;
  assign n20658 = n335 & ~n20657 ;
  assign n20659 = n339 & ~n20658 ;
  assign n20660 = n343 & ~n20659 ;
  assign n20661 = n347 & ~n20660 ;
  assign n20662 = n351 & ~n20661 ;
  assign n20663 = n355 & ~n20662 ;
  assign n20664 = n359 & ~n20663 ;
  assign n20665 = n363 & ~n20664 ;
  assign n20666 = n367 & ~n20665 ;
  assign n20667 = n371 & ~n20666 ;
  assign n20668 = n375 & ~n20667 ;
  assign n20669 = n379 & ~n20668 ;
  assign n20670 = n383 & ~n20669 ;
  assign n20671 = n387 & ~n20670 ;
  assign n20672 = n391 & ~n20671 ;
  assign n20673 = n395 & ~n20672 ;
  assign n20674 = n399 & ~n20673 ;
  assign n20675 = n403 & ~n20674 ;
  assign n20676 = n407 & ~n20675 ;
  assign n20677 = n411 & ~n20676 ;
  assign n20678 = n415 & ~n20677 ;
  assign n20679 = n419 & ~n20678 ;
  assign n20680 = n423 & ~n20679 ;
  assign n20681 = n427 & ~n20680 ;
  assign n20682 = n431 & ~n20681 ;
  assign n20683 = n435 & ~n20682 ;
  assign n20684 = n439 & ~n20683 ;
  assign n20685 = n443 & ~n20684 ;
  assign n20686 = n447 & ~n20685 ;
  assign n20687 = n451 & ~n20686 ;
  assign n20688 = n455 & ~n20687 ;
  assign n20689 = n459 & ~n20688 ;
  assign n20690 = n463 & ~n20689 ;
  assign n20691 = n467 & ~n20690 ;
  assign n20692 = n471 & ~n20691 ;
  assign n20693 = n475 & ~n20692 ;
  assign n20694 = n479 & ~n20693 ;
  assign n20695 = n483 & ~n20694 ;
  assign n20696 = n487 & ~n20695 ;
  assign n20697 = n491 & ~n20696 ;
  assign n20698 = n495 & ~n20697 ;
  assign n20699 = n499 & ~n20698 ;
  assign n20700 = n503 & ~n20699 ;
  assign n20701 = n507 & ~n20700 ;
  assign n20702 = n511 & ~n20701 ;
  assign n20703 = n515 & ~n20702 ;
  assign n20704 = n519 & ~n20703 ;
  assign n20705 = n523 & ~n20704 ;
  assign n20706 = n527 & ~n20705 ;
  assign n20707 = n531 & ~n20706 ;
  assign n20708 = n535 & ~n20707 ;
  assign n20709 = x235 & ~n537 ;
  assign n20710 = ~n20708 & n20709 ;
  assign n20798 = n20710 & x363 ;
  assign n20711 = ~n881 & n2237 ;
  assign n20712 = n2242 & ~n20711 ;
  assign n20713 = n2246 & ~n20712 ;
  assign n20714 = n2250 & ~n20713 ;
  assign n20715 = n2254 & ~n20714 ;
  assign n20716 = n2258 & ~n20715 ;
  assign n20717 = n2262 & ~n20716 ;
  assign n20718 = n2266 & ~n20717 ;
  assign n20719 = n2270 & ~n20718 ;
  assign n20720 = n2274 & ~n20719 ;
  assign n20721 = n2278 & ~n20720 ;
  assign n20722 = n2282 & ~n20721 ;
  assign n20723 = n2286 & ~n20722 ;
  assign n20724 = n2290 & ~n20723 ;
  assign n20725 = n2836 & ~n20724 ;
  assign n20726 = n602 & ~n20725 ;
  assign n20727 = n606 & ~n20726 ;
  assign n20728 = n610 & ~n20727 ;
  assign n20729 = n614 & ~n20728 ;
  assign n20730 = n618 & ~n20729 ;
  assign n20731 = n622 & ~n20730 ;
  assign n20732 = n626 & ~n20731 ;
  assign n20733 = n630 & ~n20732 ;
  assign n20734 = n634 & ~n20733 ;
  assign n20735 = n638 & ~n20734 ;
  assign n20736 = n642 & ~n20735 ;
  assign n20737 = n646 & ~n20736 ;
  assign n20738 = n650 & ~n20737 ;
  assign n20739 = n654 & ~n20738 ;
  assign n20740 = n658 & ~n20739 ;
  assign n20741 = n662 & ~n20740 ;
  assign n20742 = n666 & ~n20741 ;
  assign n20743 = n670 & ~n20742 ;
  assign n20744 = n674 & ~n20743 ;
  assign n20745 = n678 & ~n20744 ;
  assign n20746 = n682 & ~n20745 ;
  assign n20747 = n686 & ~n20746 ;
  assign n20748 = n690 & ~n20747 ;
  assign n20749 = n694 & ~n20748 ;
  assign n20750 = n698 & ~n20749 ;
  assign n20751 = n702 & ~n20750 ;
  assign n20752 = n706 & ~n20751 ;
  assign n20753 = n710 & ~n20752 ;
  assign n20754 = n714 & ~n20753 ;
  assign n20755 = n718 & ~n20754 ;
  assign n20756 = n722 & ~n20755 ;
  assign n20757 = n726 & ~n20756 ;
  assign n20758 = n730 & ~n20757 ;
  assign n20759 = n734 & ~n20758 ;
  assign n20760 = n738 & ~n20759 ;
  assign n20761 = n742 & ~n20760 ;
  assign n20762 = n746 & ~n20761 ;
  assign n20763 = n750 & ~n20762 ;
  assign n20764 = n754 & ~n20763 ;
  assign n20765 = n758 & ~n20764 ;
  assign n20766 = n762 & ~n20765 ;
  assign n20767 = n766 & ~n20766 ;
  assign n20768 = n770 & ~n20767 ;
  assign n20769 = n774 & ~n20768 ;
  assign n20770 = n778 & ~n20769 ;
  assign n20771 = n782 & ~n20770 ;
  assign n20772 = n786 & ~n20771 ;
  assign n20773 = n790 & ~n20772 ;
  assign n20774 = n794 & ~n20773 ;
  assign n20775 = n798 & ~n20774 ;
  assign n20776 = n802 & ~n20775 ;
  assign n20777 = n806 & ~n20776 ;
  assign n20778 = n810 & ~n20777 ;
  assign n20779 = n814 & ~n20778 ;
  assign n20780 = n818 & ~n20779 ;
  assign n20781 = n822 & ~n20780 ;
  assign n20782 = n826 & ~n20781 ;
  assign n20783 = n830 & ~n20782 ;
  assign n20784 = n834 & ~n20783 ;
  assign n20785 = n838 & ~n20784 ;
  assign n20786 = n842 & ~n20785 ;
  assign n20787 = n846 & ~n20786 ;
  assign n20788 = n850 & ~n20787 ;
  assign n20789 = n854 & ~n20788 ;
  assign n20790 = n858 & ~n20789 ;
  assign n20791 = n862 & ~n20790 ;
  assign n20792 = n866 & ~n20791 ;
  assign n20793 = n870 & ~n20792 ;
  assign n20794 = n874 & ~n20793 ;
  assign n20795 = ~x235 & ~n876 ;
  assign n20796 = ~n20794 & n20795 ;
  assign n20799 = ~n20796 & ~x363 ;
  assign n20800 = ~n20798 & ~n20799 ;
  assign n20801 = n546 & ~n1224 ;
  assign n20802 = n551 & ~n20801 ;
  assign n20803 = n555 & ~n20802 ;
  assign n20804 = n559 & ~n20803 ;
  assign n20805 = n563 & ~n20804 ;
  assign n20806 = n567 & ~n20805 ;
  assign n20807 = n571 & ~n20806 ;
  assign n20808 = n575 & ~n20807 ;
  assign n20809 = n579 & ~n20808 ;
  assign n20810 = n583 & ~n20809 ;
  assign n20811 = n587 & ~n20810 ;
  assign n20812 = n591 & ~n20811 ;
  assign n20813 = n2382 & ~n20812 ;
  assign n20814 = n2384 & ~n20813 ;
  assign n20815 = n2927 & ~n20814 ;
  assign n20816 = n945 & ~n20815 ;
  assign n20817 = n949 & ~n20816 ;
  assign n20818 = n953 & ~n20817 ;
  assign n20819 = n957 & ~n20818 ;
  assign n20820 = n961 & ~n20819 ;
  assign n20821 = n965 & ~n20820 ;
  assign n20822 = n969 & ~n20821 ;
  assign n20823 = n973 & ~n20822 ;
  assign n20824 = n977 & ~n20823 ;
  assign n20825 = n981 & ~n20824 ;
  assign n20826 = n985 & ~n20825 ;
  assign n20827 = n989 & ~n20826 ;
  assign n20828 = n993 & ~n20827 ;
  assign n20829 = n997 & ~n20828 ;
  assign n20830 = n1001 & ~n20829 ;
  assign n20831 = n1005 & ~n20830 ;
  assign n20832 = n1009 & ~n20831 ;
  assign n20833 = n1013 & ~n20832 ;
  assign n20834 = n1017 & ~n20833 ;
  assign n20835 = n1021 & ~n20834 ;
  assign n20836 = n1025 & ~n20835 ;
  assign n20837 = n1029 & ~n20836 ;
  assign n20838 = n1033 & ~n20837 ;
  assign n20839 = n1037 & ~n20838 ;
  assign n20840 = n1041 & ~n20839 ;
  assign n20841 = n1045 & ~n20840 ;
  assign n20842 = n1049 & ~n20841 ;
  assign n20843 = n1053 & ~n20842 ;
  assign n20844 = n1057 & ~n20843 ;
  assign n20845 = n1061 & ~n20844 ;
  assign n20846 = n1065 & ~n20845 ;
  assign n20847 = n1069 & ~n20846 ;
  assign n20848 = n1073 & ~n20847 ;
  assign n20849 = n1077 & ~n20848 ;
  assign n20850 = n1081 & ~n20849 ;
  assign n20851 = n1085 & ~n20850 ;
  assign n20852 = n1089 & ~n20851 ;
  assign n20853 = n1093 & ~n20852 ;
  assign n20854 = n1097 & ~n20853 ;
  assign n20855 = n1101 & ~n20854 ;
  assign n20856 = n1105 & ~n20855 ;
  assign n20857 = n1109 & ~n20856 ;
  assign n20858 = n1113 & ~n20857 ;
  assign n20859 = n1117 & ~n20858 ;
  assign n20860 = n1121 & ~n20859 ;
  assign n20861 = n1125 & ~n20860 ;
  assign n20862 = n1129 & ~n20861 ;
  assign n20863 = n1133 & ~n20862 ;
  assign n20864 = n1137 & ~n20863 ;
  assign n20865 = n1141 & ~n20864 ;
  assign n20866 = n1145 & ~n20865 ;
  assign n20867 = n1149 & ~n20866 ;
  assign n20868 = n1153 & ~n20867 ;
  assign n20869 = n1157 & ~n20868 ;
  assign n20870 = n1161 & ~n20869 ;
  assign n20871 = n1165 & ~n20870 ;
  assign n20872 = n1169 & ~n20871 ;
  assign n20873 = n1173 & ~n20872 ;
  assign n20874 = n1177 & ~n20873 ;
  assign n20875 = n1181 & ~n20874 ;
  assign n20876 = n1185 & ~n20875 ;
  assign n20877 = n1189 & ~n20876 ;
  assign n20878 = n1193 & ~n20877 ;
  assign n20879 = n1197 & ~n20878 ;
  assign n20880 = n1201 & ~n20879 ;
  assign n20881 = n1205 & ~n20880 ;
  assign n20882 = n1209 & ~n20881 ;
  assign n20883 = n1213 & ~n20882 ;
  assign n20884 = n1217 & ~n20883 ;
  assign n20885 = x236 & ~n1219 ;
  assign n20886 = ~n20884 & n20885 ;
  assign n20974 = n20886 & x364 ;
  assign n20887 = n885 & ~n1563 ;
  assign n20888 = n890 & ~n20887 ;
  assign n20889 = n894 & ~n20888 ;
  assign n20890 = n898 & ~n20889 ;
  assign n20891 = n902 & ~n20890 ;
  assign n20892 = n906 & ~n20891 ;
  assign n20893 = n910 & ~n20892 ;
  assign n20894 = n914 & ~n20893 ;
  assign n20895 = n918 & ~n20894 ;
  assign n20896 = n922 & ~n20895 ;
  assign n20897 = n926 & ~n20896 ;
  assign n20898 = n930 & ~n20897 ;
  assign n20899 = n2472 & ~n20898 ;
  assign n20900 = n2474 & ~n20899 ;
  assign n20901 = n3014 & ~n20900 ;
  assign n20902 = n1284 & ~n20901 ;
  assign n20903 = n1288 & ~n20902 ;
  assign n20904 = n1292 & ~n20903 ;
  assign n20905 = n1296 & ~n20904 ;
  assign n20906 = n1300 & ~n20905 ;
  assign n20907 = n1304 & ~n20906 ;
  assign n20908 = n1308 & ~n20907 ;
  assign n20909 = n1312 & ~n20908 ;
  assign n20910 = n1316 & ~n20909 ;
  assign n20911 = n1320 & ~n20910 ;
  assign n20912 = n1324 & ~n20911 ;
  assign n20913 = n1328 & ~n20912 ;
  assign n20914 = n1332 & ~n20913 ;
  assign n20915 = n1336 & ~n20914 ;
  assign n20916 = n1340 & ~n20915 ;
  assign n20917 = n1344 & ~n20916 ;
  assign n20918 = n1348 & ~n20917 ;
  assign n20919 = n1352 & ~n20918 ;
  assign n20920 = n1356 & ~n20919 ;
  assign n20921 = n1360 & ~n20920 ;
  assign n20922 = n1364 & ~n20921 ;
  assign n20923 = n1368 & ~n20922 ;
  assign n20924 = n1372 & ~n20923 ;
  assign n20925 = n1376 & ~n20924 ;
  assign n20926 = n1380 & ~n20925 ;
  assign n20927 = n1384 & ~n20926 ;
  assign n20928 = n1388 & ~n20927 ;
  assign n20929 = n1392 & ~n20928 ;
  assign n20930 = n1396 & ~n20929 ;
  assign n20931 = n1400 & ~n20930 ;
  assign n20932 = n1404 & ~n20931 ;
  assign n20933 = n1408 & ~n20932 ;
  assign n20934 = n1412 & ~n20933 ;
  assign n20935 = n1416 & ~n20934 ;
  assign n20936 = n1420 & ~n20935 ;
  assign n20937 = n1424 & ~n20936 ;
  assign n20938 = n1428 & ~n20937 ;
  assign n20939 = n1432 & ~n20938 ;
  assign n20940 = n1436 & ~n20939 ;
  assign n20941 = n1440 & ~n20940 ;
  assign n20942 = n1444 & ~n20941 ;
  assign n20943 = n1448 & ~n20942 ;
  assign n20944 = n1452 & ~n20943 ;
  assign n20945 = n1456 & ~n20944 ;
  assign n20946 = n1460 & ~n20945 ;
  assign n20947 = n1464 & ~n20946 ;
  assign n20948 = n1468 & ~n20947 ;
  assign n20949 = n1472 & ~n20948 ;
  assign n20950 = n1476 & ~n20949 ;
  assign n20951 = n1480 & ~n20950 ;
  assign n20952 = n1484 & ~n20951 ;
  assign n20953 = n1488 & ~n20952 ;
  assign n20954 = n1492 & ~n20953 ;
  assign n20955 = n1496 & ~n20954 ;
  assign n20956 = n1500 & ~n20955 ;
  assign n20957 = n1504 & ~n20956 ;
  assign n20958 = n1508 & ~n20957 ;
  assign n20959 = n1512 & ~n20958 ;
  assign n20960 = n1516 & ~n20959 ;
  assign n20961 = n1520 & ~n20960 ;
  assign n20962 = n1524 & ~n20961 ;
  assign n20963 = n1528 & ~n20962 ;
  assign n20964 = n1532 & ~n20963 ;
  assign n20965 = n1536 & ~n20964 ;
  assign n20966 = n1540 & ~n20965 ;
  assign n20967 = n1544 & ~n20966 ;
  assign n20968 = n1548 & ~n20967 ;
  assign n20969 = n1552 & ~n20968 ;
  assign n20970 = n1556 & ~n20969 ;
  assign n20971 = ~x236 & ~n1558 ;
  assign n20972 = ~n20970 & n20971 ;
  assign n20975 = ~n20972 & ~x364 ;
  assign n20976 = ~n20974 & ~n20975 ;
  assign n20977 = n1228 & ~n1904 ;
  assign n20978 = n1233 & ~n20977 ;
  assign n20979 = n1237 & ~n20978 ;
  assign n20980 = n1241 & ~n20979 ;
  assign n20981 = n1245 & ~n20980 ;
  assign n20982 = n1249 & ~n20981 ;
  assign n20983 = n1253 & ~n20982 ;
  assign n20984 = n1257 & ~n20983 ;
  assign n20985 = n1261 & ~n20984 ;
  assign n20986 = n1265 & ~n20985 ;
  assign n20987 = n1269 & ~n20986 ;
  assign n20988 = n1273 & ~n20987 ;
  assign n20989 = n2566 & ~n20988 ;
  assign n20990 = n2568 & ~n20989 ;
  assign n20991 = n3105 & ~n20990 ;
  assign n20992 = n1625 & ~n20991 ;
  assign n20993 = n1629 & ~n20992 ;
  assign n20994 = n1633 & ~n20993 ;
  assign n20995 = n1637 & ~n20994 ;
  assign n20996 = n1641 & ~n20995 ;
  assign n20997 = n1645 & ~n20996 ;
  assign n20998 = n1649 & ~n20997 ;
  assign n20999 = n1653 & ~n20998 ;
  assign n21000 = n1657 & ~n20999 ;
  assign n21001 = n1661 & ~n21000 ;
  assign n21002 = n1665 & ~n21001 ;
  assign n21003 = n1669 & ~n21002 ;
  assign n21004 = n1673 & ~n21003 ;
  assign n21005 = n1677 & ~n21004 ;
  assign n21006 = n1681 & ~n21005 ;
  assign n21007 = n1685 & ~n21006 ;
  assign n21008 = n1689 & ~n21007 ;
  assign n21009 = n1693 & ~n21008 ;
  assign n21010 = n1697 & ~n21009 ;
  assign n21011 = n1701 & ~n21010 ;
  assign n21012 = n1705 & ~n21011 ;
  assign n21013 = n1709 & ~n21012 ;
  assign n21014 = n1713 & ~n21013 ;
  assign n21015 = n1717 & ~n21014 ;
  assign n21016 = n1721 & ~n21015 ;
  assign n21017 = n1725 & ~n21016 ;
  assign n21018 = n1729 & ~n21017 ;
  assign n21019 = n1733 & ~n21018 ;
  assign n21020 = n1737 & ~n21019 ;
  assign n21021 = n1741 & ~n21020 ;
  assign n21022 = n1745 & ~n21021 ;
  assign n21023 = n1749 & ~n21022 ;
  assign n21024 = n1753 & ~n21023 ;
  assign n21025 = n1757 & ~n21024 ;
  assign n21026 = n1761 & ~n21025 ;
  assign n21027 = n1765 & ~n21026 ;
  assign n21028 = n1769 & ~n21027 ;
  assign n21029 = n1773 & ~n21028 ;
  assign n21030 = n1777 & ~n21029 ;
  assign n21031 = n1781 & ~n21030 ;
  assign n21032 = n1785 & ~n21031 ;
  assign n21033 = n1789 & ~n21032 ;
  assign n21034 = n1793 & ~n21033 ;
  assign n21035 = n1797 & ~n21034 ;
  assign n21036 = n1801 & ~n21035 ;
  assign n21037 = n1805 & ~n21036 ;
  assign n21038 = n1809 & ~n21037 ;
  assign n21039 = n1813 & ~n21038 ;
  assign n21040 = n1817 & ~n21039 ;
  assign n21041 = n1821 & ~n21040 ;
  assign n21042 = n1825 & ~n21041 ;
  assign n21043 = n1829 & ~n21042 ;
  assign n21044 = n1833 & ~n21043 ;
  assign n21045 = n1837 & ~n21044 ;
  assign n21046 = n1841 & ~n21045 ;
  assign n21047 = n1845 & ~n21046 ;
  assign n21048 = n1849 & ~n21047 ;
  assign n21049 = n1853 & ~n21048 ;
  assign n21050 = n1857 & ~n21049 ;
  assign n21051 = n1861 & ~n21050 ;
  assign n21052 = n1865 & ~n21051 ;
  assign n21053 = n1869 & ~n21052 ;
  assign n21054 = n1873 & ~n21053 ;
  assign n21055 = n1877 & ~n21054 ;
  assign n21056 = n1881 & ~n21055 ;
  assign n21057 = n1885 & ~n21056 ;
  assign n21058 = n1889 & ~n21057 ;
  assign n21059 = n1893 & ~n21058 ;
  assign n21060 = n1897 & ~n21059 ;
  assign n21061 = x237 & ~n1899 ;
  assign n21062 = ~n21060 & n21061 ;
  assign n21150 = n21062 & x365 ;
  assign n21063 = n1567 & ~n2241 ;
  assign n21064 = n1572 & ~n21063 ;
  assign n21065 = n1576 & ~n21064 ;
  assign n21066 = n1580 & ~n21065 ;
  assign n21067 = n1584 & ~n21066 ;
  assign n21068 = n1588 & ~n21067 ;
  assign n21069 = n1592 & ~n21068 ;
  assign n21070 = n1596 & ~n21069 ;
  assign n21071 = n1600 & ~n21070 ;
  assign n21072 = n1604 & ~n21071 ;
  assign n21073 = n1608 & ~n21072 ;
  assign n21074 = n1612 & ~n21073 ;
  assign n21075 = n2656 & ~n21074 ;
  assign n21076 = n2658 & ~n21075 ;
  assign n21077 = n3192 & ~n21076 ;
  assign n21078 = n1962 & ~n21077 ;
  assign n21079 = n1966 & ~n21078 ;
  assign n21080 = n1970 & ~n21079 ;
  assign n21081 = n1974 & ~n21080 ;
  assign n21082 = n1978 & ~n21081 ;
  assign n21083 = n1982 & ~n21082 ;
  assign n21084 = n1986 & ~n21083 ;
  assign n21085 = n1990 & ~n21084 ;
  assign n21086 = n1994 & ~n21085 ;
  assign n21087 = n1998 & ~n21086 ;
  assign n21088 = n2002 & ~n21087 ;
  assign n21089 = n2006 & ~n21088 ;
  assign n21090 = n2010 & ~n21089 ;
  assign n21091 = n2014 & ~n21090 ;
  assign n21092 = n2018 & ~n21091 ;
  assign n21093 = n2022 & ~n21092 ;
  assign n21094 = n2026 & ~n21093 ;
  assign n21095 = n2030 & ~n21094 ;
  assign n21096 = n2034 & ~n21095 ;
  assign n21097 = n2038 & ~n21096 ;
  assign n21098 = n2042 & ~n21097 ;
  assign n21099 = n2046 & ~n21098 ;
  assign n21100 = n2050 & ~n21099 ;
  assign n21101 = n2054 & ~n21100 ;
  assign n21102 = n2058 & ~n21101 ;
  assign n21103 = n2062 & ~n21102 ;
  assign n21104 = n2066 & ~n21103 ;
  assign n21105 = n2070 & ~n21104 ;
  assign n21106 = n2074 & ~n21105 ;
  assign n21107 = n2078 & ~n21106 ;
  assign n21108 = n2082 & ~n21107 ;
  assign n21109 = n2086 & ~n21108 ;
  assign n21110 = n2090 & ~n21109 ;
  assign n21111 = n2094 & ~n21110 ;
  assign n21112 = n2098 & ~n21111 ;
  assign n21113 = n2102 & ~n21112 ;
  assign n21114 = n2106 & ~n21113 ;
  assign n21115 = n2110 & ~n21114 ;
  assign n21116 = n2114 & ~n21115 ;
  assign n21117 = n2118 & ~n21116 ;
  assign n21118 = n2122 & ~n21117 ;
  assign n21119 = n2126 & ~n21118 ;
  assign n21120 = n2130 & ~n21119 ;
  assign n21121 = n2134 & ~n21120 ;
  assign n21122 = n2138 & ~n21121 ;
  assign n21123 = n2142 & ~n21122 ;
  assign n21124 = n2146 & ~n21123 ;
  assign n21125 = n2150 & ~n21124 ;
  assign n21126 = n2154 & ~n21125 ;
  assign n21127 = n2158 & ~n21126 ;
  assign n21128 = n2162 & ~n21127 ;
  assign n21129 = n2166 & ~n21128 ;
  assign n21130 = n2170 & ~n21129 ;
  assign n21131 = n2174 & ~n21130 ;
  assign n21132 = n2178 & ~n21131 ;
  assign n21133 = n2182 & ~n21132 ;
  assign n21134 = n2186 & ~n21133 ;
  assign n21135 = n2190 & ~n21134 ;
  assign n21136 = n2194 & ~n21135 ;
  assign n21137 = n2198 & ~n21136 ;
  assign n21138 = n2202 & ~n21137 ;
  assign n21139 = n2206 & ~n21138 ;
  assign n21140 = n2210 & ~n21139 ;
  assign n21141 = n2214 & ~n21140 ;
  assign n21142 = n2218 & ~n21141 ;
  assign n21143 = n2222 & ~n21142 ;
  assign n21144 = n2226 & ~n21143 ;
  assign n21145 = n2230 & ~n21144 ;
  assign n21146 = n2234 & ~n21145 ;
  assign n21147 = ~x237 & ~n2236 ;
  assign n21148 = ~n21146 & n21147 ;
  assign n21151 = ~n21148 & ~x365 ;
  assign n21152 = ~n21150 & ~n21151 ;
  assign n21153 = ~n550 & n1908 ;
  assign n21154 = n1913 & ~n21153 ;
  assign n21155 = n1917 & ~n21154 ;
  assign n21156 = n1921 & ~n21155 ;
  assign n21157 = n1925 & ~n21156 ;
  assign n21158 = n1929 & ~n21157 ;
  assign n21159 = n1933 & ~n21158 ;
  assign n21160 = n1937 & ~n21159 ;
  assign n21161 = n1941 & ~n21160 ;
  assign n21162 = n1945 & ~n21161 ;
  assign n21163 = n1949 & ~n21162 ;
  assign n21164 = n1953 & ~n21163 ;
  assign n21165 = n2749 & ~n21164 ;
  assign n21166 = n263 & ~n21165 ;
  assign n21167 = n267 & ~n21166 ;
  assign n21168 = n271 & ~n21167 ;
  assign n21169 = n275 & ~n21168 ;
  assign n21170 = n279 & ~n21169 ;
  assign n21171 = n283 & ~n21170 ;
  assign n21172 = n287 & ~n21171 ;
  assign n21173 = n291 & ~n21172 ;
  assign n21174 = n295 & ~n21173 ;
  assign n21175 = n299 & ~n21174 ;
  assign n21176 = n303 & ~n21175 ;
  assign n21177 = n307 & ~n21176 ;
  assign n21178 = n311 & ~n21177 ;
  assign n21179 = n315 & ~n21178 ;
  assign n21180 = n319 & ~n21179 ;
  assign n21181 = n323 & ~n21180 ;
  assign n21182 = n327 & ~n21181 ;
  assign n21183 = n331 & ~n21182 ;
  assign n21184 = n335 & ~n21183 ;
  assign n21185 = n339 & ~n21184 ;
  assign n21186 = n343 & ~n21185 ;
  assign n21187 = n347 & ~n21186 ;
  assign n21188 = n351 & ~n21187 ;
  assign n21189 = n355 & ~n21188 ;
  assign n21190 = n359 & ~n21189 ;
  assign n21191 = n363 & ~n21190 ;
  assign n21192 = n367 & ~n21191 ;
  assign n21193 = n371 & ~n21192 ;
  assign n21194 = n375 & ~n21193 ;
  assign n21195 = n379 & ~n21194 ;
  assign n21196 = n383 & ~n21195 ;
  assign n21197 = n387 & ~n21196 ;
  assign n21198 = n391 & ~n21197 ;
  assign n21199 = n395 & ~n21198 ;
  assign n21200 = n399 & ~n21199 ;
  assign n21201 = n403 & ~n21200 ;
  assign n21202 = n407 & ~n21201 ;
  assign n21203 = n411 & ~n21202 ;
  assign n21204 = n415 & ~n21203 ;
  assign n21205 = n419 & ~n21204 ;
  assign n21206 = n423 & ~n21205 ;
  assign n21207 = n427 & ~n21206 ;
  assign n21208 = n431 & ~n21207 ;
  assign n21209 = n435 & ~n21208 ;
  assign n21210 = n439 & ~n21209 ;
  assign n21211 = n443 & ~n21210 ;
  assign n21212 = n447 & ~n21211 ;
  assign n21213 = n451 & ~n21212 ;
  assign n21214 = n455 & ~n21213 ;
  assign n21215 = n459 & ~n21214 ;
  assign n21216 = n463 & ~n21215 ;
  assign n21217 = n467 & ~n21216 ;
  assign n21218 = n471 & ~n21217 ;
  assign n21219 = n475 & ~n21218 ;
  assign n21220 = n479 & ~n21219 ;
  assign n21221 = n483 & ~n21220 ;
  assign n21222 = n487 & ~n21221 ;
  assign n21223 = n491 & ~n21222 ;
  assign n21224 = n495 & ~n21223 ;
  assign n21225 = n499 & ~n21224 ;
  assign n21226 = n503 & ~n21225 ;
  assign n21227 = n507 & ~n21226 ;
  assign n21228 = n511 & ~n21227 ;
  assign n21229 = n515 & ~n21228 ;
  assign n21230 = n519 & ~n21229 ;
  assign n21231 = n523 & ~n21230 ;
  assign n21232 = n527 & ~n21231 ;
  assign n21233 = n531 & ~n21232 ;
  assign n21234 = n535 & ~n21233 ;
  assign n21235 = n539 & ~n21234 ;
  assign n21236 = n543 & ~n21235 ;
  assign n21237 = x238 & ~n545 ;
  assign n21238 = ~n21236 & n21237 ;
  assign n21326 = n21238 & x366 ;
  assign n21239 = ~n889 & n2245 ;
  assign n21240 = n2250 & ~n21239 ;
  assign n21241 = n2254 & ~n21240 ;
  assign n21242 = n2258 & ~n21241 ;
  assign n21243 = n2262 & ~n21242 ;
  assign n21244 = n2266 & ~n21243 ;
  assign n21245 = n2270 & ~n21244 ;
  assign n21246 = n2274 & ~n21245 ;
  assign n21247 = n2278 & ~n21246 ;
  assign n21248 = n2282 & ~n21247 ;
  assign n21249 = n2286 & ~n21248 ;
  assign n21250 = n2290 & ~n21249 ;
  assign n21251 = n2836 & ~n21250 ;
  assign n21252 = n602 & ~n21251 ;
  assign n21253 = n606 & ~n21252 ;
  assign n21254 = n610 & ~n21253 ;
  assign n21255 = n614 & ~n21254 ;
  assign n21256 = n618 & ~n21255 ;
  assign n21257 = n622 & ~n21256 ;
  assign n21258 = n626 & ~n21257 ;
  assign n21259 = n630 & ~n21258 ;
  assign n21260 = n634 & ~n21259 ;
  assign n21261 = n638 & ~n21260 ;
  assign n21262 = n642 & ~n21261 ;
  assign n21263 = n646 & ~n21262 ;
  assign n21264 = n650 & ~n21263 ;
  assign n21265 = n654 & ~n21264 ;
  assign n21266 = n658 & ~n21265 ;
  assign n21267 = n662 & ~n21266 ;
  assign n21268 = n666 & ~n21267 ;
  assign n21269 = n670 & ~n21268 ;
  assign n21270 = n674 & ~n21269 ;
  assign n21271 = n678 & ~n21270 ;
  assign n21272 = n682 & ~n21271 ;
  assign n21273 = n686 & ~n21272 ;
  assign n21274 = n690 & ~n21273 ;
  assign n21275 = n694 & ~n21274 ;
  assign n21276 = n698 & ~n21275 ;
  assign n21277 = n702 & ~n21276 ;
  assign n21278 = n706 & ~n21277 ;
  assign n21279 = n710 & ~n21278 ;
  assign n21280 = n714 & ~n21279 ;
  assign n21281 = n718 & ~n21280 ;
  assign n21282 = n722 & ~n21281 ;
  assign n21283 = n726 & ~n21282 ;
  assign n21284 = n730 & ~n21283 ;
  assign n21285 = n734 & ~n21284 ;
  assign n21286 = n738 & ~n21285 ;
  assign n21287 = n742 & ~n21286 ;
  assign n21288 = n746 & ~n21287 ;
  assign n21289 = n750 & ~n21288 ;
  assign n21290 = n754 & ~n21289 ;
  assign n21291 = n758 & ~n21290 ;
  assign n21292 = n762 & ~n21291 ;
  assign n21293 = n766 & ~n21292 ;
  assign n21294 = n770 & ~n21293 ;
  assign n21295 = n774 & ~n21294 ;
  assign n21296 = n778 & ~n21295 ;
  assign n21297 = n782 & ~n21296 ;
  assign n21298 = n786 & ~n21297 ;
  assign n21299 = n790 & ~n21298 ;
  assign n21300 = n794 & ~n21299 ;
  assign n21301 = n798 & ~n21300 ;
  assign n21302 = n802 & ~n21301 ;
  assign n21303 = n806 & ~n21302 ;
  assign n21304 = n810 & ~n21303 ;
  assign n21305 = n814 & ~n21304 ;
  assign n21306 = n818 & ~n21305 ;
  assign n21307 = n822 & ~n21306 ;
  assign n21308 = n826 & ~n21307 ;
  assign n21309 = n830 & ~n21308 ;
  assign n21310 = n834 & ~n21309 ;
  assign n21311 = n838 & ~n21310 ;
  assign n21312 = n842 & ~n21311 ;
  assign n21313 = n846 & ~n21312 ;
  assign n21314 = n850 & ~n21313 ;
  assign n21315 = n854 & ~n21314 ;
  assign n21316 = n858 & ~n21315 ;
  assign n21317 = n862 & ~n21316 ;
  assign n21318 = n866 & ~n21317 ;
  assign n21319 = n870 & ~n21318 ;
  assign n21320 = n874 & ~n21319 ;
  assign n21321 = n878 & ~n21320 ;
  assign n21322 = n882 & ~n21321 ;
  assign n21323 = ~x238 & ~n884 ;
  assign n21324 = ~n21322 & n21323 ;
  assign n21327 = ~n21324 & ~x366 ;
  assign n21328 = ~n21326 & ~n21327 ;
  assign n21329 = n554 & ~n1232 ;
  assign n21330 = n559 & ~n21329 ;
  assign n21331 = n563 & ~n21330 ;
  assign n21332 = n567 & ~n21331 ;
  assign n21333 = n571 & ~n21332 ;
  assign n21334 = n575 & ~n21333 ;
  assign n21335 = n579 & ~n21334 ;
  assign n21336 = n583 & ~n21335 ;
  assign n21337 = n587 & ~n21336 ;
  assign n21338 = n591 & ~n21337 ;
  assign n21339 = n2382 & ~n21338 ;
  assign n21340 = n2384 & ~n21339 ;
  assign n21341 = n2927 & ~n21340 ;
  assign n21342 = n945 & ~n21341 ;
  assign n21343 = n949 & ~n21342 ;
  assign n21344 = n953 & ~n21343 ;
  assign n21345 = n957 & ~n21344 ;
  assign n21346 = n961 & ~n21345 ;
  assign n21347 = n965 & ~n21346 ;
  assign n21348 = n969 & ~n21347 ;
  assign n21349 = n973 & ~n21348 ;
  assign n21350 = n977 & ~n21349 ;
  assign n21351 = n981 & ~n21350 ;
  assign n21352 = n985 & ~n21351 ;
  assign n21353 = n989 & ~n21352 ;
  assign n21354 = n993 & ~n21353 ;
  assign n21355 = n997 & ~n21354 ;
  assign n21356 = n1001 & ~n21355 ;
  assign n21357 = n1005 & ~n21356 ;
  assign n21358 = n1009 & ~n21357 ;
  assign n21359 = n1013 & ~n21358 ;
  assign n21360 = n1017 & ~n21359 ;
  assign n21361 = n1021 & ~n21360 ;
  assign n21362 = n1025 & ~n21361 ;
  assign n21363 = n1029 & ~n21362 ;
  assign n21364 = n1033 & ~n21363 ;
  assign n21365 = n1037 & ~n21364 ;
  assign n21366 = n1041 & ~n21365 ;
  assign n21367 = n1045 & ~n21366 ;
  assign n21368 = n1049 & ~n21367 ;
  assign n21369 = n1053 & ~n21368 ;
  assign n21370 = n1057 & ~n21369 ;
  assign n21371 = n1061 & ~n21370 ;
  assign n21372 = n1065 & ~n21371 ;
  assign n21373 = n1069 & ~n21372 ;
  assign n21374 = n1073 & ~n21373 ;
  assign n21375 = n1077 & ~n21374 ;
  assign n21376 = n1081 & ~n21375 ;
  assign n21377 = n1085 & ~n21376 ;
  assign n21378 = n1089 & ~n21377 ;
  assign n21379 = n1093 & ~n21378 ;
  assign n21380 = n1097 & ~n21379 ;
  assign n21381 = n1101 & ~n21380 ;
  assign n21382 = n1105 & ~n21381 ;
  assign n21383 = n1109 & ~n21382 ;
  assign n21384 = n1113 & ~n21383 ;
  assign n21385 = n1117 & ~n21384 ;
  assign n21386 = n1121 & ~n21385 ;
  assign n21387 = n1125 & ~n21386 ;
  assign n21388 = n1129 & ~n21387 ;
  assign n21389 = n1133 & ~n21388 ;
  assign n21390 = n1137 & ~n21389 ;
  assign n21391 = n1141 & ~n21390 ;
  assign n21392 = n1145 & ~n21391 ;
  assign n21393 = n1149 & ~n21392 ;
  assign n21394 = n1153 & ~n21393 ;
  assign n21395 = n1157 & ~n21394 ;
  assign n21396 = n1161 & ~n21395 ;
  assign n21397 = n1165 & ~n21396 ;
  assign n21398 = n1169 & ~n21397 ;
  assign n21399 = n1173 & ~n21398 ;
  assign n21400 = n1177 & ~n21399 ;
  assign n21401 = n1181 & ~n21400 ;
  assign n21402 = n1185 & ~n21401 ;
  assign n21403 = n1189 & ~n21402 ;
  assign n21404 = n1193 & ~n21403 ;
  assign n21405 = n1197 & ~n21404 ;
  assign n21406 = n1201 & ~n21405 ;
  assign n21407 = n1205 & ~n21406 ;
  assign n21408 = n1209 & ~n21407 ;
  assign n21409 = n1213 & ~n21408 ;
  assign n21410 = n1217 & ~n21409 ;
  assign n21411 = n1221 & ~n21410 ;
  assign n21412 = n1225 & ~n21411 ;
  assign n21413 = x239 & ~n1227 ;
  assign n21414 = ~n21412 & n21413 ;
  assign n21502 = n21414 & x367 ;
  assign n21415 = n893 & ~n1571 ;
  assign n21416 = n898 & ~n21415 ;
  assign n21417 = n902 & ~n21416 ;
  assign n21418 = n906 & ~n21417 ;
  assign n21419 = n910 & ~n21418 ;
  assign n21420 = n914 & ~n21419 ;
  assign n21421 = n918 & ~n21420 ;
  assign n21422 = n922 & ~n21421 ;
  assign n21423 = n926 & ~n21422 ;
  assign n21424 = n930 & ~n21423 ;
  assign n21425 = n2472 & ~n21424 ;
  assign n21426 = n2474 & ~n21425 ;
  assign n21427 = n3014 & ~n21426 ;
  assign n21428 = n1284 & ~n21427 ;
  assign n21429 = n1288 & ~n21428 ;
  assign n21430 = n1292 & ~n21429 ;
  assign n21431 = n1296 & ~n21430 ;
  assign n21432 = n1300 & ~n21431 ;
  assign n21433 = n1304 & ~n21432 ;
  assign n21434 = n1308 & ~n21433 ;
  assign n21435 = n1312 & ~n21434 ;
  assign n21436 = n1316 & ~n21435 ;
  assign n21437 = n1320 & ~n21436 ;
  assign n21438 = n1324 & ~n21437 ;
  assign n21439 = n1328 & ~n21438 ;
  assign n21440 = n1332 & ~n21439 ;
  assign n21441 = n1336 & ~n21440 ;
  assign n21442 = n1340 & ~n21441 ;
  assign n21443 = n1344 & ~n21442 ;
  assign n21444 = n1348 & ~n21443 ;
  assign n21445 = n1352 & ~n21444 ;
  assign n21446 = n1356 & ~n21445 ;
  assign n21447 = n1360 & ~n21446 ;
  assign n21448 = n1364 & ~n21447 ;
  assign n21449 = n1368 & ~n21448 ;
  assign n21450 = n1372 & ~n21449 ;
  assign n21451 = n1376 & ~n21450 ;
  assign n21452 = n1380 & ~n21451 ;
  assign n21453 = n1384 & ~n21452 ;
  assign n21454 = n1388 & ~n21453 ;
  assign n21455 = n1392 & ~n21454 ;
  assign n21456 = n1396 & ~n21455 ;
  assign n21457 = n1400 & ~n21456 ;
  assign n21458 = n1404 & ~n21457 ;
  assign n21459 = n1408 & ~n21458 ;
  assign n21460 = n1412 & ~n21459 ;
  assign n21461 = n1416 & ~n21460 ;
  assign n21462 = n1420 & ~n21461 ;
  assign n21463 = n1424 & ~n21462 ;
  assign n21464 = n1428 & ~n21463 ;
  assign n21465 = n1432 & ~n21464 ;
  assign n21466 = n1436 & ~n21465 ;
  assign n21467 = n1440 & ~n21466 ;
  assign n21468 = n1444 & ~n21467 ;
  assign n21469 = n1448 & ~n21468 ;
  assign n21470 = n1452 & ~n21469 ;
  assign n21471 = n1456 & ~n21470 ;
  assign n21472 = n1460 & ~n21471 ;
  assign n21473 = n1464 & ~n21472 ;
  assign n21474 = n1468 & ~n21473 ;
  assign n21475 = n1472 & ~n21474 ;
  assign n21476 = n1476 & ~n21475 ;
  assign n21477 = n1480 & ~n21476 ;
  assign n21478 = n1484 & ~n21477 ;
  assign n21479 = n1488 & ~n21478 ;
  assign n21480 = n1492 & ~n21479 ;
  assign n21481 = n1496 & ~n21480 ;
  assign n21482 = n1500 & ~n21481 ;
  assign n21483 = n1504 & ~n21482 ;
  assign n21484 = n1508 & ~n21483 ;
  assign n21485 = n1512 & ~n21484 ;
  assign n21486 = n1516 & ~n21485 ;
  assign n21487 = n1520 & ~n21486 ;
  assign n21488 = n1524 & ~n21487 ;
  assign n21489 = n1528 & ~n21488 ;
  assign n21490 = n1532 & ~n21489 ;
  assign n21491 = n1536 & ~n21490 ;
  assign n21492 = n1540 & ~n21491 ;
  assign n21493 = n1544 & ~n21492 ;
  assign n21494 = n1548 & ~n21493 ;
  assign n21495 = n1552 & ~n21494 ;
  assign n21496 = n1556 & ~n21495 ;
  assign n21497 = n1560 & ~n21496 ;
  assign n21498 = n1564 & ~n21497 ;
  assign n21499 = ~x239 & ~n1566 ;
  assign n21500 = ~n21498 & n21499 ;
  assign n21503 = ~n21500 & ~x367 ;
  assign n21504 = ~n21502 & ~n21503 ;
  assign n21505 = n1236 & ~n1912 ;
  assign n21506 = n1241 & ~n21505 ;
  assign n21507 = n1245 & ~n21506 ;
  assign n21508 = n1249 & ~n21507 ;
  assign n21509 = n1253 & ~n21508 ;
  assign n21510 = n1257 & ~n21509 ;
  assign n21511 = n1261 & ~n21510 ;
  assign n21512 = n1265 & ~n21511 ;
  assign n21513 = n1269 & ~n21512 ;
  assign n21514 = n1273 & ~n21513 ;
  assign n21515 = n2566 & ~n21514 ;
  assign n21516 = n2568 & ~n21515 ;
  assign n21517 = n3105 & ~n21516 ;
  assign n21518 = n1625 & ~n21517 ;
  assign n21519 = n1629 & ~n21518 ;
  assign n21520 = n1633 & ~n21519 ;
  assign n21521 = n1637 & ~n21520 ;
  assign n21522 = n1641 & ~n21521 ;
  assign n21523 = n1645 & ~n21522 ;
  assign n21524 = n1649 & ~n21523 ;
  assign n21525 = n1653 & ~n21524 ;
  assign n21526 = n1657 & ~n21525 ;
  assign n21527 = n1661 & ~n21526 ;
  assign n21528 = n1665 & ~n21527 ;
  assign n21529 = n1669 & ~n21528 ;
  assign n21530 = n1673 & ~n21529 ;
  assign n21531 = n1677 & ~n21530 ;
  assign n21532 = n1681 & ~n21531 ;
  assign n21533 = n1685 & ~n21532 ;
  assign n21534 = n1689 & ~n21533 ;
  assign n21535 = n1693 & ~n21534 ;
  assign n21536 = n1697 & ~n21535 ;
  assign n21537 = n1701 & ~n21536 ;
  assign n21538 = n1705 & ~n21537 ;
  assign n21539 = n1709 & ~n21538 ;
  assign n21540 = n1713 & ~n21539 ;
  assign n21541 = n1717 & ~n21540 ;
  assign n21542 = n1721 & ~n21541 ;
  assign n21543 = n1725 & ~n21542 ;
  assign n21544 = n1729 & ~n21543 ;
  assign n21545 = n1733 & ~n21544 ;
  assign n21546 = n1737 & ~n21545 ;
  assign n21547 = n1741 & ~n21546 ;
  assign n21548 = n1745 & ~n21547 ;
  assign n21549 = n1749 & ~n21548 ;
  assign n21550 = n1753 & ~n21549 ;
  assign n21551 = n1757 & ~n21550 ;
  assign n21552 = n1761 & ~n21551 ;
  assign n21553 = n1765 & ~n21552 ;
  assign n21554 = n1769 & ~n21553 ;
  assign n21555 = n1773 & ~n21554 ;
  assign n21556 = n1777 & ~n21555 ;
  assign n21557 = n1781 & ~n21556 ;
  assign n21558 = n1785 & ~n21557 ;
  assign n21559 = n1789 & ~n21558 ;
  assign n21560 = n1793 & ~n21559 ;
  assign n21561 = n1797 & ~n21560 ;
  assign n21562 = n1801 & ~n21561 ;
  assign n21563 = n1805 & ~n21562 ;
  assign n21564 = n1809 & ~n21563 ;
  assign n21565 = n1813 & ~n21564 ;
  assign n21566 = n1817 & ~n21565 ;
  assign n21567 = n1821 & ~n21566 ;
  assign n21568 = n1825 & ~n21567 ;
  assign n21569 = n1829 & ~n21568 ;
  assign n21570 = n1833 & ~n21569 ;
  assign n21571 = n1837 & ~n21570 ;
  assign n21572 = n1841 & ~n21571 ;
  assign n21573 = n1845 & ~n21572 ;
  assign n21574 = n1849 & ~n21573 ;
  assign n21575 = n1853 & ~n21574 ;
  assign n21576 = n1857 & ~n21575 ;
  assign n21577 = n1861 & ~n21576 ;
  assign n21578 = n1865 & ~n21577 ;
  assign n21579 = n1869 & ~n21578 ;
  assign n21580 = n1873 & ~n21579 ;
  assign n21581 = n1877 & ~n21580 ;
  assign n21582 = n1881 & ~n21581 ;
  assign n21583 = n1885 & ~n21582 ;
  assign n21584 = n1889 & ~n21583 ;
  assign n21585 = n1893 & ~n21584 ;
  assign n21586 = n1897 & ~n21585 ;
  assign n21587 = n1901 & ~n21586 ;
  assign n21588 = n1905 & ~n21587 ;
  assign n21589 = x240 & ~n1907 ;
  assign n21590 = ~n21588 & n21589 ;
  assign n21678 = n21590 & x368 ;
  assign n21591 = n1575 & ~n2249 ;
  assign n21592 = n1580 & ~n21591 ;
  assign n21593 = n1584 & ~n21592 ;
  assign n21594 = n1588 & ~n21593 ;
  assign n21595 = n1592 & ~n21594 ;
  assign n21596 = n1596 & ~n21595 ;
  assign n21597 = n1600 & ~n21596 ;
  assign n21598 = n1604 & ~n21597 ;
  assign n21599 = n1608 & ~n21598 ;
  assign n21600 = n1612 & ~n21599 ;
  assign n21601 = n2656 & ~n21600 ;
  assign n21602 = n2658 & ~n21601 ;
  assign n21603 = n3192 & ~n21602 ;
  assign n21604 = n1962 & ~n21603 ;
  assign n21605 = n1966 & ~n21604 ;
  assign n21606 = n1970 & ~n21605 ;
  assign n21607 = n1974 & ~n21606 ;
  assign n21608 = n1978 & ~n21607 ;
  assign n21609 = n1982 & ~n21608 ;
  assign n21610 = n1986 & ~n21609 ;
  assign n21611 = n1990 & ~n21610 ;
  assign n21612 = n1994 & ~n21611 ;
  assign n21613 = n1998 & ~n21612 ;
  assign n21614 = n2002 & ~n21613 ;
  assign n21615 = n2006 & ~n21614 ;
  assign n21616 = n2010 & ~n21615 ;
  assign n21617 = n2014 & ~n21616 ;
  assign n21618 = n2018 & ~n21617 ;
  assign n21619 = n2022 & ~n21618 ;
  assign n21620 = n2026 & ~n21619 ;
  assign n21621 = n2030 & ~n21620 ;
  assign n21622 = n2034 & ~n21621 ;
  assign n21623 = n2038 & ~n21622 ;
  assign n21624 = n2042 & ~n21623 ;
  assign n21625 = n2046 & ~n21624 ;
  assign n21626 = n2050 & ~n21625 ;
  assign n21627 = n2054 & ~n21626 ;
  assign n21628 = n2058 & ~n21627 ;
  assign n21629 = n2062 & ~n21628 ;
  assign n21630 = n2066 & ~n21629 ;
  assign n21631 = n2070 & ~n21630 ;
  assign n21632 = n2074 & ~n21631 ;
  assign n21633 = n2078 & ~n21632 ;
  assign n21634 = n2082 & ~n21633 ;
  assign n21635 = n2086 & ~n21634 ;
  assign n21636 = n2090 & ~n21635 ;
  assign n21637 = n2094 & ~n21636 ;
  assign n21638 = n2098 & ~n21637 ;
  assign n21639 = n2102 & ~n21638 ;
  assign n21640 = n2106 & ~n21639 ;
  assign n21641 = n2110 & ~n21640 ;
  assign n21642 = n2114 & ~n21641 ;
  assign n21643 = n2118 & ~n21642 ;
  assign n21644 = n2122 & ~n21643 ;
  assign n21645 = n2126 & ~n21644 ;
  assign n21646 = n2130 & ~n21645 ;
  assign n21647 = n2134 & ~n21646 ;
  assign n21648 = n2138 & ~n21647 ;
  assign n21649 = n2142 & ~n21648 ;
  assign n21650 = n2146 & ~n21649 ;
  assign n21651 = n2150 & ~n21650 ;
  assign n21652 = n2154 & ~n21651 ;
  assign n21653 = n2158 & ~n21652 ;
  assign n21654 = n2162 & ~n21653 ;
  assign n21655 = n2166 & ~n21654 ;
  assign n21656 = n2170 & ~n21655 ;
  assign n21657 = n2174 & ~n21656 ;
  assign n21658 = n2178 & ~n21657 ;
  assign n21659 = n2182 & ~n21658 ;
  assign n21660 = n2186 & ~n21659 ;
  assign n21661 = n2190 & ~n21660 ;
  assign n21662 = n2194 & ~n21661 ;
  assign n21663 = n2198 & ~n21662 ;
  assign n21664 = n2202 & ~n21663 ;
  assign n21665 = n2206 & ~n21664 ;
  assign n21666 = n2210 & ~n21665 ;
  assign n21667 = n2214 & ~n21666 ;
  assign n21668 = n2218 & ~n21667 ;
  assign n21669 = n2222 & ~n21668 ;
  assign n21670 = n2226 & ~n21669 ;
  assign n21671 = n2230 & ~n21670 ;
  assign n21672 = n2234 & ~n21671 ;
  assign n21673 = n2238 & ~n21672 ;
  assign n21674 = n2242 & ~n21673 ;
  assign n21675 = ~x240 & ~n2244 ;
  assign n21676 = ~n21674 & n21675 ;
  assign n21679 = ~n21676 & ~x368 ;
  assign n21680 = ~n21678 & ~n21679 ;
  assign n21681 = ~n558 & n1916 ;
  assign n21682 = n1921 & ~n21681 ;
  assign n21683 = n1925 & ~n21682 ;
  assign n21684 = n1929 & ~n21683 ;
  assign n21685 = n1933 & ~n21684 ;
  assign n21686 = n1937 & ~n21685 ;
  assign n21687 = n1941 & ~n21686 ;
  assign n21688 = n1945 & ~n21687 ;
  assign n21689 = n1949 & ~n21688 ;
  assign n21690 = n1953 & ~n21689 ;
  assign n21691 = n2749 & ~n21690 ;
  assign n21692 = n263 & ~n21691 ;
  assign n21693 = n267 & ~n21692 ;
  assign n21694 = n271 & ~n21693 ;
  assign n21695 = n275 & ~n21694 ;
  assign n21696 = n279 & ~n21695 ;
  assign n21697 = n283 & ~n21696 ;
  assign n21698 = n287 & ~n21697 ;
  assign n21699 = n291 & ~n21698 ;
  assign n21700 = n295 & ~n21699 ;
  assign n21701 = n299 & ~n21700 ;
  assign n21702 = n303 & ~n21701 ;
  assign n21703 = n307 & ~n21702 ;
  assign n21704 = n311 & ~n21703 ;
  assign n21705 = n315 & ~n21704 ;
  assign n21706 = n319 & ~n21705 ;
  assign n21707 = n323 & ~n21706 ;
  assign n21708 = n327 & ~n21707 ;
  assign n21709 = n331 & ~n21708 ;
  assign n21710 = n335 & ~n21709 ;
  assign n21711 = n339 & ~n21710 ;
  assign n21712 = n343 & ~n21711 ;
  assign n21713 = n347 & ~n21712 ;
  assign n21714 = n351 & ~n21713 ;
  assign n21715 = n355 & ~n21714 ;
  assign n21716 = n359 & ~n21715 ;
  assign n21717 = n363 & ~n21716 ;
  assign n21718 = n367 & ~n21717 ;
  assign n21719 = n371 & ~n21718 ;
  assign n21720 = n375 & ~n21719 ;
  assign n21721 = n379 & ~n21720 ;
  assign n21722 = n383 & ~n21721 ;
  assign n21723 = n387 & ~n21722 ;
  assign n21724 = n391 & ~n21723 ;
  assign n21725 = n395 & ~n21724 ;
  assign n21726 = n399 & ~n21725 ;
  assign n21727 = n403 & ~n21726 ;
  assign n21728 = n407 & ~n21727 ;
  assign n21729 = n411 & ~n21728 ;
  assign n21730 = n415 & ~n21729 ;
  assign n21731 = n419 & ~n21730 ;
  assign n21732 = n423 & ~n21731 ;
  assign n21733 = n427 & ~n21732 ;
  assign n21734 = n431 & ~n21733 ;
  assign n21735 = n435 & ~n21734 ;
  assign n21736 = n439 & ~n21735 ;
  assign n21737 = n443 & ~n21736 ;
  assign n21738 = n447 & ~n21737 ;
  assign n21739 = n451 & ~n21738 ;
  assign n21740 = n455 & ~n21739 ;
  assign n21741 = n459 & ~n21740 ;
  assign n21742 = n463 & ~n21741 ;
  assign n21743 = n467 & ~n21742 ;
  assign n21744 = n471 & ~n21743 ;
  assign n21745 = n475 & ~n21744 ;
  assign n21746 = n479 & ~n21745 ;
  assign n21747 = n483 & ~n21746 ;
  assign n21748 = n487 & ~n21747 ;
  assign n21749 = n491 & ~n21748 ;
  assign n21750 = n495 & ~n21749 ;
  assign n21751 = n499 & ~n21750 ;
  assign n21752 = n503 & ~n21751 ;
  assign n21753 = n507 & ~n21752 ;
  assign n21754 = n511 & ~n21753 ;
  assign n21755 = n515 & ~n21754 ;
  assign n21756 = n519 & ~n21755 ;
  assign n21757 = n523 & ~n21756 ;
  assign n21758 = n527 & ~n21757 ;
  assign n21759 = n531 & ~n21758 ;
  assign n21760 = n535 & ~n21759 ;
  assign n21761 = n539 & ~n21760 ;
  assign n21762 = n543 & ~n21761 ;
  assign n21763 = n547 & ~n21762 ;
  assign n21764 = n551 & ~n21763 ;
  assign n21765 = x241 & ~n553 ;
  assign n21766 = ~n21764 & n21765 ;
  assign n21854 = n21766 & x369 ;
  assign n21767 = ~n897 & n2253 ;
  assign n21768 = n2258 & ~n21767 ;
  assign n21769 = n2262 & ~n21768 ;
  assign n21770 = n2266 & ~n21769 ;
  assign n21771 = n2270 & ~n21770 ;
  assign n21772 = n2274 & ~n21771 ;
  assign n21773 = n2278 & ~n21772 ;
  assign n21774 = n2282 & ~n21773 ;
  assign n21775 = n2286 & ~n21774 ;
  assign n21776 = n2290 & ~n21775 ;
  assign n21777 = n2836 & ~n21776 ;
  assign n21778 = n602 & ~n21777 ;
  assign n21779 = n606 & ~n21778 ;
  assign n21780 = n610 & ~n21779 ;
  assign n21781 = n614 & ~n21780 ;
  assign n21782 = n618 & ~n21781 ;
  assign n21783 = n622 & ~n21782 ;
  assign n21784 = n626 & ~n21783 ;
  assign n21785 = n630 & ~n21784 ;
  assign n21786 = n634 & ~n21785 ;
  assign n21787 = n638 & ~n21786 ;
  assign n21788 = n642 & ~n21787 ;
  assign n21789 = n646 & ~n21788 ;
  assign n21790 = n650 & ~n21789 ;
  assign n21791 = n654 & ~n21790 ;
  assign n21792 = n658 & ~n21791 ;
  assign n21793 = n662 & ~n21792 ;
  assign n21794 = n666 & ~n21793 ;
  assign n21795 = n670 & ~n21794 ;
  assign n21796 = n674 & ~n21795 ;
  assign n21797 = n678 & ~n21796 ;
  assign n21798 = n682 & ~n21797 ;
  assign n21799 = n686 & ~n21798 ;
  assign n21800 = n690 & ~n21799 ;
  assign n21801 = n694 & ~n21800 ;
  assign n21802 = n698 & ~n21801 ;
  assign n21803 = n702 & ~n21802 ;
  assign n21804 = n706 & ~n21803 ;
  assign n21805 = n710 & ~n21804 ;
  assign n21806 = n714 & ~n21805 ;
  assign n21807 = n718 & ~n21806 ;
  assign n21808 = n722 & ~n21807 ;
  assign n21809 = n726 & ~n21808 ;
  assign n21810 = n730 & ~n21809 ;
  assign n21811 = n734 & ~n21810 ;
  assign n21812 = n738 & ~n21811 ;
  assign n21813 = n742 & ~n21812 ;
  assign n21814 = n746 & ~n21813 ;
  assign n21815 = n750 & ~n21814 ;
  assign n21816 = n754 & ~n21815 ;
  assign n21817 = n758 & ~n21816 ;
  assign n21818 = n762 & ~n21817 ;
  assign n21819 = n766 & ~n21818 ;
  assign n21820 = n770 & ~n21819 ;
  assign n21821 = n774 & ~n21820 ;
  assign n21822 = n778 & ~n21821 ;
  assign n21823 = n782 & ~n21822 ;
  assign n21824 = n786 & ~n21823 ;
  assign n21825 = n790 & ~n21824 ;
  assign n21826 = n794 & ~n21825 ;
  assign n21827 = n798 & ~n21826 ;
  assign n21828 = n802 & ~n21827 ;
  assign n21829 = n806 & ~n21828 ;
  assign n21830 = n810 & ~n21829 ;
  assign n21831 = n814 & ~n21830 ;
  assign n21832 = n818 & ~n21831 ;
  assign n21833 = n822 & ~n21832 ;
  assign n21834 = n826 & ~n21833 ;
  assign n21835 = n830 & ~n21834 ;
  assign n21836 = n834 & ~n21835 ;
  assign n21837 = n838 & ~n21836 ;
  assign n21838 = n842 & ~n21837 ;
  assign n21839 = n846 & ~n21838 ;
  assign n21840 = n850 & ~n21839 ;
  assign n21841 = n854 & ~n21840 ;
  assign n21842 = n858 & ~n21841 ;
  assign n21843 = n862 & ~n21842 ;
  assign n21844 = n866 & ~n21843 ;
  assign n21845 = n870 & ~n21844 ;
  assign n21846 = n874 & ~n21845 ;
  assign n21847 = n878 & ~n21846 ;
  assign n21848 = n882 & ~n21847 ;
  assign n21849 = n886 & ~n21848 ;
  assign n21850 = n890 & ~n21849 ;
  assign n21851 = ~x241 & ~n892 ;
  assign n21852 = ~n21850 & n21851 ;
  assign n21855 = ~n21852 & ~x369 ;
  assign n21856 = ~n21854 & ~n21855 ;
  assign n21857 = n562 & ~n1240 ;
  assign n21858 = n567 & ~n21857 ;
  assign n21859 = n571 & ~n21858 ;
  assign n21860 = n575 & ~n21859 ;
  assign n21861 = n579 & ~n21860 ;
  assign n21862 = n583 & ~n21861 ;
  assign n21863 = n587 & ~n21862 ;
  assign n21864 = n591 & ~n21863 ;
  assign n21865 = n2382 & ~n21864 ;
  assign n21866 = n2384 & ~n21865 ;
  assign n21867 = n2927 & ~n21866 ;
  assign n21868 = n945 & ~n21867 ;
  assign n21869 = n949 & ~n21868 ;
  assign n21870 = n953 & ~n21869 ;
  assign n21871 = n957 & ~n21870 ;
  assign n21872 = n961 & ~n21871 ;
  assign n21873 = n965 & ~n21872 ;
  assign n21874 = n969 & ~n21873 ;
  assign n21875 = n973 & ~n21874 ;
  assign n21876 = n977 & ~n21875 ;
  assign n21877 = n981 & ~n21876 ;
  assign n21878 = n985 & ~n21877 ;
  assign n21879 = n989 & ~n21878 ;
  assign n21880 = n993 & ~n21879 ;
  assign n21881 = n997 & ~n21880 ;
  assign n21882 = n1001 & ~n21881 ;
  assign n21883 = n1005 & ~n21882 ;
  assign n21884 = n1009 & ~n21883 ;
  assign n21885 = n1013 & ~n21884 ;
  assign n21886 = n1017 & ~n21885 ;
  assign n21887 = n1021 & ~n21886 ;
  assign n21888 = n1025 & ~n21887 ;
  assign n21889 = n1029 & ~n21888 ;
  assign n21890 = n1033 & ~n21889 ;
  assign n21891 = n1037 & ~n21890 ;
  assign n21892 = n1041 & ~n21891 ;
  assign n21893 = n1045 & ~n21892 ;
  assign n21894 = n1049 & ~n21893 ;
  assign n21895 = n1053 & ~n21894 ;
  assign n21896 = n1057 & ~n21895 ;
  assign n21897 = n1061 & ~n21896 ;
  assign n21898 = n1065 & ~n21897 ;
  assign n21899 = n1069 & ~n21898 ;
  assign n21900 = n1073 & ~n21899 ;
  assign n21901 = n1077 & ~n21900 ;
  assign n21902 = n1081 & ~n21901 ;
  assign n21903 = n1085 & ~n21902 ;
  assign n21904 = n1089 & ~n21903 ;
  assign n21905 = n1093 & ~n21904 ;
  assign n21906 = n1097 & ~n21905 ;
  assign n21907 = n1101 & ~n21906 ;
  assign n21908 = n1105 & ~n21907 ;
  assign n21909 = n1109 & ~n21908 ;
  assign n21910 = n1113 & ~n21909 ;
  assign n21911 = n1117 & ~n21910 ;
  assign n21912 = n1121 & ~n21911 ;
  assign n21913 = n1125 & ~n21912 ;
  assign n21914 = n1129 & ~n21913 ;
  assign n21915 = n1133 & ~n21914 ;
  assign n21916 = n1137 & ~n21915 ;
  assign n21917 = n1141 & ~n21916 ;
  assign n21918 = n1145 & ~n21917 ;
  assign n21919 = n1149 & ~n21918 ;
  assign n21920 = n1153 & ~n21919 ;
  assign n21921 = n1157 & ~n21920 ;
  assign n21922 = n1161 & ~n21921 ;
  assign n21923 = n1165 & ~n21922 ;
  assign n21924 = n1169 & ~n21923 ;
  assign n21925 = n1173 & ~n21924 ;
  assign n21926 = n1177 & ~n21925 ;
  assign n21927 = n1181 & ~n21926 ;
  assign n21928 = n1185 & ~n21927 ;
  assign n21929 = n1189 & ~n21928 ;
  assign n21930 = n1193 & ~n21929 ;
  assign n21931 = n1197 & ~n21930 ;
  assign n21932 = n1201 & ~n21931 ;
  assign n21933 = n1205 & ~n21932 ;
  assign n21934 = n1209 & ~n21933 ;
  assign n21935 = n1213 & ~n21934 ;
  assign n21936 = n1217 & ~n21935 ;
  assign n21937 = n1221 & ~n21936 ;
  assign n21938 = n1225 & ~n21937 ;
  assign n21939 = n1229 & ~n21938 ;
  assign n21940 = n1233 & ~n21939 ;
  assign n21941 = x242 & ~n1235 ;
  assign n21942 = ~n21940 & n21941 ;
  assign n22030 = n21942 & x370 ;
  assign n21943 = n901 & ~n1579 ;
  assign n21944 = n906 & ~n21943 ;
  assign n21945 = n910 & ~n21944 ;
  assign n21946 = n914 & ~n21945 ;
  assign n21947 = n918 & ~n21946 ;
  assign n21948 = n922 & ~n21947 ;
  assign n21949 = n926 & ~n21948 ;
  assign n21950 = n930 & ~n21949 ;
  assign n21951 = n2472 & ~n21950 ;
  assign n21952 = n2474 & ~n21951 ;
  assign n21953 = n3014 & ~n21952 ;
  assign n21954 = n1284 & ~n21953 ;
  assign n21955 = n1288 & ~n21954 ;
  assign n21956 = n1292 & ~n21955 ;
  assign n21957 = n1296 & ~n21956 ;
  assign n21958 = n1300 & ~n21957 ;
  assign n21959 = n1304 & ~n21958 ;
  assign n21960 = n1308 & ~n21959 ;
  assign n21961 = n1312 & ~n21960 ;
  assign n21962 = n1316 & ~n21961 ;
  assign n21963 = n1320 & ~n21962 ;
  assign n21964 = n1324 & ~n21963 ;
  assign n21965 = n1328 & ~n21964 ;
  assign n21966 = n1332 & ~n21965 ;
  assign n21967 = n1336 & ~n21966 ;
  assign n21968 = n1340 & ~n21967 ;
  assign n21969 = n1344 & ~n21968 ;
  assign n21970 = n1348 & ~n21969 ;
  assign n21971 = n1352 & ~n21970 ;
  assign n21972 = n1356 & ~n21971 ;
  assign n21973 = n1360 & ~n21972 ;
  assign n21974 = n1364 & ~n21973 ;
  assign n21975 = n1368 & ~n21974 ;
  assign n21976 = n1372 & ~n21975 ;
  assign n21977 = n1376 & ~n21976 ;
  assign n21978 = n1380 & ~n21977 ;
  assign n21979 = n1384 & ~n21978 ;
  assign n21980 = n1388 & ~n21979 ;
  assign n21981 = n1392 & ~n21980 ;
  assign n21982 = n1396 & ~n21981 ;
  assign n21983 = n1400 & ~n21982 ;
  assign n21984 = n1404 & ~n21983 ;
  assign n21985 = n1408 & ~n21984 ;
  assign n21986 = n1412 & ~n21985 ;
  assign n21987 = n1416 & ~n21986 ;
  assign n21988 = n1420 & ~n21987 ;
  assign n21989 = n1424 & ~n21988 ;
  assign n21990 = n1428 & ~n21989 ;
  assign n21991 = n1432 & ~n21990 ;
  assign n21992 = n1436 & ~n21991 ;
  assign n21993 = n1440 & ~n21992 ;
  assign n21994 = n1444 & ~n21993 ;
  assign n21995 = n1448 & ~n21994 ;
  assign n21996 = n1452 & ~n21995 ;
  assign n21997 = n1456 & ~n21996 ;
  assign n21998 = n1460 & ~n21997 ;
  assign n21999 = n1464 & ~n21998 ;
  assign n22000 = n1468 & ~n21999 ;
  assign n22001 = n1472 & ~n22000 ;
  assign n22002 = n1476 & ~n22001 ;
  assign n22003 = n1480 & ~n22002 ;
  assign n22004 = n1484 & ~n22003 ;
  assign n22005 = n1488 & ~n22004 ;
  assign n22006 = n1492 & ~n22005 ;
  assign n22007 = n1496 & ~n22006 ;
  assign n22008 = n1500 & ~n22007 ;
  assign n22009 = n1504 & ~n22008 ;
  assign n22010 = n1508 & ~n22009 ;
  assign n22011 = n1512 & ~n22010 ;
  assign n22012 = n1516 & ~n22011 ;
  assign n22013 = n1520 & ~n22012 ;
  assign n22014 = n1524 & ~n22013 ;
  assign n22015 = n1528 & ~n22014 ;
  assign n22016 = n1532 & ~n22015 ;
  assign n22017 = n1536 & ~n22016 ;
  assign n22018 = n1540 & ~n22017 ;
  assign n22019 = n1544 & ~n22018 ;
  assign n22020 = n1548 & ~n22019 ;
  assign n22021 = n1552 & ~n22020 ;
  assign n22022 = n1556 & ~n22021 ;
  assign n22023 = n1560 & ~n22022 ;
  assign n22024 = n1564 & ~n22023 ;
  assign n22025 = n1568 & ~n22024 ;
  assign n22026 = n1572 & ~n22025 ;
  assign n22027 = ~x242 & ~n1574 ;
  assign n22028 = ~n22026 & n22027 ;
  assign n22031 = ~n22028 & ~x370 ;
  assign n22032 = ~n22030 & ~n22031 ;
  assign n22033 = n1244 & ~n1920 ;
  assign n22034 = n1249 & ~n22033 ;
  assign n22035 = n1253 & ~n22034 ;
  assign n22036 = n1257 & ~n22035 ;
  assign n22037 = n1261 & ~n22036 ;
  assign n22038 = n1265 & ~n22037 ;
  assign n22039 = n1269 & ~n22038 ;
  assign n22040 = n1273 & ~n22039 ;
  assign n22041 = n2566 & ~n22040 ;
  assign n22042 = n2568 & ~n22041 ;
  assign n22043 = n3105 & ~n22042 ;
  assign n22044 = n1625 & ~n22043 ;
  assign n22045 = n1629 & ~n22044 ;
  assign n22046 = n1633 & ~n22045 ;
  assign n22047 = n1637 & ~n22046 ;
  assign n22048 = n1641 & ~n22047 ;
  assign n22049 = n1645 & ~n22048 ;
  assign n22050 = n1649 & ~n22049 ;
  assign n22051 = n1653 & ~n22050 ;
  assign n22052 = n1657 & ~n22051 ;
  assign n22053 = n1661 & ~n22052 ;
  assign n22054 = n1665 & ~n22053 ;
  assign n22055 = n1669 & ~n22054 ;
  assign n22056 = n1673 & ~n22055 ;
  assign n22057 = n1677 & ~n22056 ;
  assign n22058 = n1681 & ~n22057 ;
  assign n22059 = n1685 & ~n22058 ;
  assign n22060 = n1689 & ~n22059 ;
  assign n22061 = n1693 & ~n22060 ;
  assign n22062 = n1697 & ~n22061 ;
  assign n22063 = n1701 & ~n22062 ;
  assign n22064 = n1705 & ~n22063 ;
  assign n22065 = n1709 & ~n22064 ;
  assign n22066 = n1713 & ~n22065 ;
  assign n22067 = n1717 & ~n22066 ;
  assign n22068 = n1721 & ~n22067 ;
  assign n22069 = n1725 & ~n22068 ;
  assign n22070 = n1729 & ~n22069 ;
  assign n22071 = n1733 & ~n22070 ;
  assign n22072 = n1737 & ~n22071 ;
  assign n22073 = n1741 & ~n22072 ;
  assign n22074 = n1745 & ~n22073 ;
  assign n22075 = n1749 & ~n22074 ;
  assign n22076 = n1753 & ~n22075 ;
  assign n22077 = n1757 & ~n22076 ;
  assign n22078 = n1761 & ~n22077 ;
  assign n22079 = n1765 & ~n22078 ;
  assign n22080 = n1769 & ~n22079 ;
  assign n22081 = n1773 & ~n22080 ;
  assign n22082 = n1777 & ~n22081 ;
  assign n22083 = n1781 & ~n22082 ;
  assign n22084 = n1785 & ~n22083 ;
  assign n22085 = n1789 & ~n22084 ;
  assign n22086 = n1793 & ~n22085 ;
  assign n22087 = n1797 & ~n22086 ;
  assign n22088 = n1801 & ~n22087 ;
  assign n22089 = n1805 & ~n22088 ;
  assign n22090 = n1809 & ~n22089 ;
  assign n22091 = n1813 & ~n22090 ;
  assign n22092 = n1817 & ~n22091 ;
  assign n22093 = n1821 & ~n22092 ;
  assign n22094 = n1825 & ~n22093 ;
  assign n22095 = n1829 & ~n22094 ;
  assign n22096 = n1833 & ~n22095 ;
  assign n22097 = n1837 & ~n22096 ;
  assign n22098 = n1841 & ~n22097 ;
  assign n22099 = n1845 & ~n22098 ;
  assign n22100 = n1849 & ~n22099 ;
  assign n22101 = n1853 & ~n22100 ;
  assign n22102 = n1857 & ~n22101 ;
  assign n22103 = n1861 & ~n22102 ;
  assign n22104 = n1865 & ~n22103 ;
  assign n22105 = n1869 & ~n22104 ;
  assign n22106 = n1873 & ~n22105 ;
  assign n22107 = n1877 & ~n22106 ;
  assign n22108 = n1881 & ~n22107 ;
  assign n22109 = n1885 & ~n22108 ;
  assign n22110 = n1889 & ~n22109 ;
  assign n22111 = n1893 & ~n22110 ;
  assign n22112 = n1897 & ~n22111 ;
  assign n22113 = n1901 & ~n22112 ;
  assign n22114 = n1905 & ~n22113 ;
  assign n22115 = n1909 & ~n22114 ;
  assign n22116 = n1913 & ~n22115 ;
  assign n22117 = x243 & ~n1915 ;
  assign n22118 = ~n22116 & n22117 ;
  assign n22206 = n22118 & x371 ;
  assign n22119 = n1583 & ~n2257 ;
  assign n22120 = n1588 & ~n22119 ;
  assign n22121 = n1592 & ~n22120 ;
  assign n22122 = n1596 & ~n22121 ;
  assign n22123 = n1600 & ~n22122 ;
  assign n22124 = n1604 & ~n22123 ;
  assign n22125 = n1608 & ~n22124 ;
  assign n22126 = n1612 & ~n22125 ;
  assign n22127 = n2656 & ~n22126 ;
  assign n22128 = n2658 & ~n22127 ;
  assign n22129 = n3192 & ~n22128 ;
  assign n22130 = n1962 & ~n22129 ;
  assign n22131 = n1966 & ~n22130 ;
  assign n22132 = n1970 & ~n22131 ;
  assign n22133 = n1974 & ~n22132 ;
  assign n22134 = n1978 & ~n22133 ;
  assign n22135 = n1982 & ~n22134 ;
  assign n22136 = n1986 & ~n22135 ;
  assign n22137 = n1990 & ~n22136 ;
  assign n22138 = n1994 & ~n22137 ;
  assign n22139 = n1998 & ~n22138 ;
  assign n22140 = n2002 & ~n22139 ;
  assign n22141 = n2006 & ~n22140 ;
  assign n22142 = n2010 & ~n22141 ;
  assign n22143 = n2014 & ~n22142 ;
  assign n22144 = n2018 & ~n22143 ;
  assign n22145 = n2022 & ~n22144 ;
  assign n22146 = n2026 & ~n22145 ;
  assign n22147 = n2030 & ~n22146 ;
  assign n22148 = n2034 & ~n22147 ;
  assign n22149 = n2038 & ~n22148 ;
  assign n22150 = n2042 & ~n22149 ;
  assign n22151 = n2046 & ~n22150 ;
  assign n22152 = n2050 & ~n22151 ;
  assign n22153 = n2054 & ~n22152 ;
  assign n22154 = n2058 & ~n22153 ;
  assign n22155 = n2062 & ~n22154 ;
  assign n22156 = n2066 & ~n22155 ;
  assign n22157 = n2070 & ~n22156 ;
  assign n22158 = n2074 & ~n22157 ;
  assign n22159 = n2078 & ~n22158 ;
  assign n22160 = n2082 & ~n22159 ;
  assign n22161 = n2086 & ~n22160 ;
  assign n22162 = n2090 & ~n22161 ;
  assign n22163 = n2094 & ~n22162 ;
  assign n22164 = n2098 & ~n22163 ;
  assign n22165 = n2102 & ~n22164 ;
  assign n22166 = n2106 & ~n22165 ;
  assign n22167 = n2110 & ~n22166 ;
  assign n22168 = n2114 & ~n22167 ;
  assign n22169 = n2118 & ~n22168 ;
  assign n22170 = n2122 & ~n22169 ;
  assign n22171 = n2126 & ~n22170 ;
  assign n22172 = n2130 & ~n22171 ;
  assign n22173 = n2134 & ~n22172 ;
  assign n22174 = n2138 & ~n22173 ;
  assign n22175 = n2142 & ~n22174 ;
  assign n22176 = n2146 & ~n22175 ;
  assign n22177 = n2150 & ~n22176 ;
  assign n22178 = n2154 & ~n22177 ;
  assign n22179 = n2158 & ~n22178 ;
  assign n22180 = n2162 & ~n22179 ;
  assign n22181 = n2166 & ~n22180 ;
  assign n22182 = n2170 & ~n22181 ;
  assign n22183 = n2174 & ~n22182 ;
  assign n22184 = n2178 & ~n22183 ;
  assign n22185 = n2182 & ~n22184 ;
  assign n22186 = n2186 & ~n22185 ;
  assign n22187 = n2190 & ~n22186 ;
  assign n22188 = n2194 & ~n22187 ;
  assign n22189 = n2198 & ~n22188 ;
  assign n22190 = n2202 & ~n22189 ;
  assign n22191 = n2206 & ~n22190 ;
  assign n22192 = n2210 & ~n22191 ;
  assign n22193 = n2214 & ~n22192 ;
  assign n22194 = n2218 & ~n22193 ;
  assign n22195 = n2222 & ~n22194 ;
  assign n22196 = n2226 & ~n22195 ;
  assign n22197 = n2230 & ~n22196 ;
  assign n22198 = n2234 & ~n22197 ;
  assign n22199 = n2238 & ~n22198 ;
  assign n22200 = n2242 & ~n22199 ;
  assign n22201 = n2246 & ~n22200 ;
  assign n22202 = n2250 & ~n22201 ;
  assign n22203 = ~x243 & ~n2252 ;
  assign n22204 = ~n22202 & n22203 ;
  assign n22207 = ~n22204 & ~x371 ;
  assign n22208 = ~n22206 & ~n22207 ;
  assign n22209 = ~n566 & n1924 ;
  assign n22210 = n1929 & ~n22209 ;
  assign n22211 = n1933 & ~n22210 ;
  assign n22212 = n1937 & ~n22211 ;
  assign n22213 = n1941 & ~n22212 ;
  assign n22214 = n1945 & ~n22213 ;
  assign n22215 = n1949 & ~n22214 ;
  assign n22216 = n1953 & ~n22215 ;
  assign n22217 = n2749 & ~n22216 ;
  assign n22218 = n263 & ~n22217 ;
  assign n22219 = n267 & ~n22218 ;
  assign n22220 = n271 & ~n22219 ;
  assign n22221 = n275 & ~n22220 ;
  assign n22222 = n279 & ~n22221 ;
  assign n22223 = n283 & ~n22222 ;
  assign n22224 = n287 & ~n22223 ;
  assign n22225 = n291 & ~n22224 ;
  assign n22226 = n295 & ~n22225 ;
  assign n22227 = n299 & ~n22226 ;
  assign n22228 = n303 & ~n22227 ;
  assign n22229 = n307 & ~n22228 ;
  assign n22230 = n311 & ~n22229 ;
  assign n22231 = n315 & ~n22230 ;
  assign n22232 = n319 & ~n22231 ;
  assign n22233 = n323 & ~n22232 ;
  assign n22234 = n327 & ~n22233 ;
  assign n22235 = n331 & ~n22234 ;
  assign n22236 = n335 & ~n22235 ;
  assign n22237 = n339 & ~n22236 ;
  assign n22238 = n343 & ~n22237 ;
  assign n22239 = n347 & ~n22238 ;
  assign n22240 = n351 & ~n22239 ;
  assign n22241 = n355 & ~n22240 ;
  assign n22242 = n359 & ~n22241 ;
  assign n22243 = n363 & ~n22242 ;
  assign n22244 = n367 & ~n22243 ;
  assign n22245 = n371 & ~n22244 ;
  assign n22246 = n375 & ~n22245 ;
  assign n22247 = n379 & ~n22246 ;
  assign n22248 = n383 & ~n22247 ;
  assign n22249 = n387 & ~n22248 ;
  assign n22250 = n391 & ~n22249 ;
  assign n22251 = n395 & ~n22250 ;
  assign n22252 = n399 & ~n22251 ;
  assign n22253 = n403 & ~n22252 ;
  assign n22254 = n407 & ~n22253 ;
  assign n22255 = n411 & ~n22254 ;
  assign n22256 = n415 & ~n22255 ;
  assign n22257 = n419 & ~n22256 ;
  assign n22258 = n423 & ~n22257 ;
  assign n22259 = n427 & ~n22258 ;
  assign n22260 = n431 & ~n22259 ;
  assign n22261 = n435 & ~n22260 ;
  assign n22262 = n439 & ~n22261 ;
  assign n22263 = n443 & ~n22262 ;
  assign n22264 = n447 & ~n22263 ;
  assign n22265 = n451 & ~n22264 ;
  assign n22266 = n455 & ~n22265 ;
  assign n22267 = n459 & ~n22266 ;
  assign n22268 = n463 & ~n22267 ;
  assign n22269 = n467 & ~n22268 ;
  assign n22270 = n471 & ~n22269 ;
  assign n22271 = n475 & ~n22270 ;
  assign n22272 = n479 & ~n22271 ;
  assign n22273 = n483 & ~n22272 ;
  assign n22274 = n487 & ~n22273 ;
  assign n22275 = n491 & ~n22274 ;
  assign n22276 = n495 & ~n22275 ;
  assign n22277 = n499 & ~n22276 ;
  assign n22278 = n503 & ~n22277 ;
  assign n22279 = n507 & ~n22278 ;
  assign n22280 = n511 & ~n22279 ;
  assign n22281 = n515 & ~n22280 ;
  assign n22282 = n519 & ~n22281 ;
  assign n22283 = n523 & ~n22282 ;
  assign n22284 = n527 & ~n22283 ;
  assign n22285 = n531 & ~n22284 ;
  assign n22286 = n535 & ~n22285 ;
  assign n22287 = n539 & ~n22286 ;
  assign n22288 = n543 & ~n22287 ;
  assign n22289 = n547 & ~n22288 ;
  assign n22290 = n551 & ~n22289 ;
  assign n22291 = n555 & ~n22290 ;
  assign n22292 = n559 & ~n22291 ;
  assign n22293 = x244 & ~n561 ;
  assign n22294 = ~n22292 & n22293 ;
  assign n22382 = n22294 & x372 ;
  assign n22295 = ~n905 & n2261 ;
  assign n22296 = n2266 & ~n22295 ;
  assign n22297 = n2270 & ~n22296 ;
  assign n22298 = n2274 & ~n22297 ;
  assign n22299 = n2278 & ~n22298 ;
  assign n22300 = n2282 & ~n22299 ;
  assign n22301 = n2286 & ~n22300 ;
  assign n22302 = n2290 & ~n22301 ;
  assign n22303 = n2836 & ~n22302 ;
  assign n22304 = n602 & ~n22303 ;
  assign n22305 = n606 & ~n22304 ;
  assign n22306 = n610 & ~n22305 ;
  assign n22307 = n614 & ~n22306 ;
  assign n22308 = n618 & ~n22307 ;
  assign n22309 = n622 & ~n22308 ;
  assign n22310 = n626 & ~n22309 ;
  assign n22311 = n630 & ~n22310 ;
  assign n22312 = n634 & ~n22311 ;
  assign n22313 = n638 & ~n22312 ;
  assign n22314 = n642 & ~n22313 ;
  assign n22315 = n646 & ~n22314 ;
  assign n22316 = n650 & ~n22315 ;
  assign n22317 = n654 & ~n22316 ;
  assign n22318 = n658 & ~n22317 ;
  assign n22319 = n662 & ~n22318 ;
  assign n22320 = n666 & ~n22319 ;
  assign n22321 = n670 & ~n22320 ;
  assign n22322 = n674 & ~n22321 ;
  assign n22323 = n678 & ~n22322 ;
  assign n22324 = n682 & ~n22323 ;
  assign n22325 = n686 & ~n22324 ;
  assign n22326 = n690 & ~n22325 ;
  assign n22327 = n694 & ~n22326 ;
  assign n22328 = n698 & ~n22327 ;
  assign n22329 = n702 & ~n22328 ;
  assign n22330 = n706 & ~n22329 ;
  assign n22331 = n710 & ~n22330 ;
  assign n22332 = n714 & ~n22331 ;
  assign n22333 = n718 & ~n22332 ;
  assign n22334 = n722 & ~n22333 ;
  assign n22335 = n726 & ~n22334 ;
  assign n22336 = n730 & ~n22335 ;
  assign n22337 = n734 & ~n22336 ;
  assign n22338 = n738 & ~n22337 ;
  assign n22339 = n742 & ~n22338 ;
  assign n22340 = n746 & ~n22339 ;
  assign n22341 = n750 & ~n22340 ;
  assign n22342 = n754 & ~n22341 ;
  assign n22343 = n758 & ~n22342 ;
  assign n22344 = n762 & ~n22343 ;
  assign n22345 = n766 & ~n22344 ;
  assign n22346 = n770 & ~n22345 ;
  assign n22347 = n774 & ~n22346 ;
  assign n22348 = n778 & ~n22347 ;
  assign n22349 = n782 & ~n22348 ;
  assign n22350 = n786 & ~n22349 ;
  assign n22351 = n790 & ~n22350 ;
  assign n22352 = n794 & ~n22351 ;
  assign n22353 = n798 & ~n22352 ;
  assign n22354 = n802 & ~n22353 ;
  assign n22355 = n806 & ~n22354 ;
  assign n22356 = n810 & ~n22355 ;
  assign n22357 = n814 & ~n22356 ;
  assign n22358 = n818 & ~n22357 ;
  assign n22359 = n822 & ~n22358 ;
  assign n22360 = n826 & ~n22359 ;
  assign n22361 = n830 & ~n22360 ;
  assign n22362 = n834 & ~n22361 ;
  assign n22363 = n838 & ~n22362 ;
  assign n22364 = n842 & ~n22363 ;
  assign n22365 = n846 & ~n22364 ;
  assign n22366 = n850 & ~n22365 ;
  assign n22367 = n854 & ~n22366 ;
  assign n22368 = n858 & ~n22367 ;
  assign n22369 = n862 & ~n22368 ;
  assign n22370 = n866 & ~n22369 ;
  assign n22371 = n870 & ~n22370 ;
  assign n22372 = n874 & ~n22371 ;
  assign n22373 = n878 & ~n22372 ;
  assign n22374 = n882 & ~n22373 ;
  assign n22375 = n886 & ~n22374 ;
  assign n22376 = n890 & ~n22375 ;
  assign n22377 = n894 & ~n22376 ;
  assign n22378 = n898 & ~n22377 ;
  assign n22379 = ~x244 & ~n900 ;
  assign n22380 = ~n22378 & n22379 ;
  assign n22383 = ~n22380 & ~x372 ;
  assign n22384 = ~n22382 & ~n22383 ;
  assign n22385 = n570 & ~n1248 ;
  assign n22386 = n575 & ~n22385 ;
  assign n22387 = n579 & ~n22386 ;
  assign n22388 = n583 & ~n22387 ;
  assign n22389 = n587 & ~n22388 ;
  assign n22390 = n591 & ~n22389 ;
  assign n22391 = n2382 & ~n22390 ;
  assign n22392 = n2384 & ~n22391 ;
  assign n22393 = n2927 & ~n22392 ;
  assign n22394 = n945 & ~n22393 ;
  assign n22395 = n949 & ~n22394 ;
  assign n22396 = n953 & ~n22395 ;
  assign n22397 = n957 & ~n22396 ;
  assign n22398 = n961 & ~n22397 ;
  assign n22399 = n965 & ~n22398 ;
  assign n22400 = n969 & ~n22399 ;
  assign n22401 = n973 & ~n22400 ;
  assign n22402 = n977 & ~n22401 ;
  assign n22403 = n981 & ~n22402 ;
  assign n22404 = n985 & ~n22403 ;
  assign n22405 = n989 & ~n22404 ;
  assign n22406 = n993 & ~n22405 ;
  assign n22407 = n997 & ~n22406 ;
  assign n22408 = n1001 & ~n22407 ;
  assign n22409 = n1005 & ~n22408 ;
  assign n22410 = n1009 & ~n22409 ;
  assign n22411 = n1013 & ~n22410 ;
  assign n22412 = n1017 & ~n22411 ;
  assign n22413 = n1021 & ~n22412 ;
  assign n22414 = n1025 & ~n22413 ;
  assign n22415 = n1029 & ~n22414 ;
  assign n22416 = n1033 & ~n22415 ;
  assign n22417 = n1037 & ~n22416 ;
  assign n22418 = n1041 & ~n22417 ;
  assign n22419 = n1045 & ~n22418 ;
  assign n22420 = n1049 & ~n22419 ;
  assign n22421 = n1053 & ~n22420 ;
  assign n22422 = n1057 & ~n22421 ;
  assign n22423 = n1061 & ~n22422 ;
  assign n22424 = n1065 & ~n22423 ;
  assign n22425 = n1069 & ~n22424 ;
  assign n22426 = n1073 & ~n22425 ;
  assign n22427 = n1077 & ~n22426 ;
  assign n22428 = n1081 & ~n22427 ;
  assign n22429 = n1085 & ~n22428 ;
  assign n22430 = n1089 & ~n22429 ;
  assign n22431 = n1093 & ~n22430 ;
  assign n22432 = n1097 & ~n22431 ;
  assign n22433 = n1101 & ~n22432 ;
  assign n22434 = n1105 & ~n22433 ;
  assign n22435 = n1109 & ~n22434 ;
  assign n22436 = n1113 & ~n22435 ;
  assign n22437 = n1117 & ~n22436 ;
  assign n22438 = n1121 & ~n22437 ;
  assign n22439 = n1125 & ~n22438 ;
  assign n22440 = n1129 & ~n22439 ;
  assign n22441 = n1133 & ~n22440 ;
  assign n22442 = n1137 & ~n22441 ;
  assign n22443 = n1141 & ~n22442 ;
  assign n22444 = n1145 & ~n22443 ;
  assign n22445 = n1149 & ~n22444 ;
  assign n22446 = n1153 & ~n22445 ;
  assign n22447 = n1157 & ~n22446 ;
  assign n22448 = n1161 & ~n22447 ;
  assign n22449 = n1165 & ~n22448 ;
  assign n22450 = n1169 & ~n22449 ;
  assign n22451 = n1173 & ~n22450 ;
  assign n22452 = n1177 & ~n22451 ;
  assign n22453 = n1181 & ~n22452 ;
  assign n22454 = n1185 & ~n22453 ;
  assign n22455 = n1189 & ~n22454 ;
  assign n22456 = n1193 & ~n22455 ;
  assign n22457 = n1197 & ~n22456 ;
  assign n22458 = n1201 & ~n22457 ;
  assign n22459 = n1205 & ~n22458 ;
  assign n22460 = n1209 & ~n22459 ;
  assign n22461 = n1213 & ~n22460 ;
  assign n22462 = n1217 & ~n22461 ;
  assign n22463 = n1221 & ~n22462 ;
  assign n22464 = n1225 & ~n22463 ;
  assign n22465 = n1229 & ~n22464 ;
  assign n22466 = n1233 & ~n22465 ;
  assign n22467 = n1237 & ~n22466 ;
  assign n22468 = n1241 & ~n22467 ;
  assign n22469 = x245 & ~n1243 ;
  assign n22470 = ~n22468 & n22469 ;
  assign n22558 = n22470 & x373 ;
  assign n22471 = n909 & ~n1587 ;
  assign n22472 = n914 & ~n22471 ;
  assign n22473 = n918 & ~n22472 ;
  assign n22474 = n922 & ~n22473 ;
  assign n22475 = n926 & ~n22474 ;
  assign n22476 = n930 & ~n22475 ;
  assign n22477 = n2472 & ~n22476 ;
  assign n22478 = n2474 & ~n22477 ;
  assign n22479 = n3014 & ~n22478 ;
  assign n22480 = n1284 & ~n22479 ;
  assign n22481 = n1288 & ~n22480 ;
  assign n22482 = n1292 & ~n22481 ;
  assign n22483 = n1296 & ~n22482 ;
  assign n22484 = n1300 & ~n22483 ;
  assign n22485 = n1304 & ~n22484 ;
  assign n22486 = n1308 & ~n22485 ;
  assign n22487 = n1312 & ~n22486 ;
  assign n22488 = n1316 & ~n22487 ;
  assign n22489 = n1320 & ~n22488 ;
  assign n22490 = n1324 & ~n22489 ;
  assign n22491 = n1328 & ~n22490 ;
  assign n22492 = n1332 & ~n22491 ;
  assign n22493 = n1336 & ~n22492 ;
  assign n22494 = n1340 & ~n22493 ;
  assign n22495 = n1344 & ~n22494 ;
  assign n22496 = n1348 & ~n22495 ;
  assign n22497 = n1352 & ~n22496 ;
  assign n22498 = n1356 & ~n22497 ;
  assign n22499 = n1360 & ~n22498 ;
  assign n22500 = n1364 & ~n22499 ;
  assign n22501 = n1368 & ~n22500 ;
  assign n22502 = n1372 & ~n22501 ;
  assign n22503 = n1376 & ~n22502 ;
  assign n22504 = n1380 & ~n22503 ;
  assign n22505 = n1384 & ~n22504 ;
  assign n22506 = n1388 & ~n22505 ;
  assign n22507 = n1392 & ~n22506 ;
  assign n22508 = n1396 & ~n22507 ;
  assign n22509 = n1400 & ~n22508 ;
  assign n22510 = n1404 & ~n22509 ;
  assign n22511 = n1408 & ~n22510 ;
  assign n22512 = n1412 & ~n22511 ;
  assign n22513 = n1416 & ~n22512 ;
  assign n22514 = n1420 & ~n22513 ;
  assign n22515 = n1424 & ~n22514 ;
  assign n22516 = n1428 & ~n22515 ;
  assign n22517 = n1432 & ~n22516 ;
  assign n22518 = n1436 & ~n22517 ;
  assign n22519 = n1440 & ~n22518 ;
  assign n22520 = n1444 & ~n22519 ;
  assign n22521 = n1448 & ~n22520 ;
  assign n22522 = n1452 & ~n22521 ;
  assign n22523 = n1456 & ~n22522 ;
  assign n22524 = n1460 & ~n22523 ;
  assign n22525 = n1464 & ~n22524 ;
  assign n22526 = n1468 & ~n22525 ;
  assign n22527 = n1472 & ~n22526 ;
  assign n22528 = n1476 & ~n22527 ;
  assign n22529 = n1480 & ~n22528 ;
  assign n22530 = n1484 & ~n22529 ;
  assign n22531 = n1488 & ~n22530 ;
  assign n22532 = n1492 & ~n22531 ;
  assign n22533 = n1496 & ~n22532 ;
  assign n22534 = n1500 & ~n22533 ;
  assign n22535 = n1504 & ~n22534 ;
  assign n22536 = n1508 & ~n22535 ;
  assign n22537 = n1512 & ~n22536 ;
  assign n22538 = n1516 & ~n22537 ;
  assign n22539 = n1520 & ~n22538 ;
  assign n22540 = n1524 & ~n22539 ;
  assign n22541 = n1528 & ~n22540 ;
  assign n22542 = n1532 & ~n22541 ;
  assign n22543 = n1536 & ~n22542 ;
  assign n22544 = n1540 & ~n22543 ;
  assign n22545 = n1544 & ~n22544 ;
  assign n22546 = n1548 & ~n22545 ;
  assign n22547 = n1552 & ~n22546 ;
  assign n22548 = n1556 & ~n22547 ;
  assign n22549 = n1560 & ~n22548 ;
  assign n22550 = n1564 & ~n22549 ;
  assign n22551 = n1568 & ~n22550 ;
  assign n22552 = n1572 & ~n22551 ;
  assign n22553 = n1576 & ~n22552 ;
  assign n22554 = n1580 & ~n22553 ;
  assign n22555 = ~x245 & ~n1582 ;
  assign n22556 = ~n22554 & n22555 ;
  assign n22559 = ~n22556 & ~x373 ;
  assign n22560 = ~n22558 & ~n22559 ;
  assign n22561 = n1252 & ~n1928 ;
  assign n22562 = n1257 & ~n22561 ;
  assign n22563 = n1261 & ~n22562 ;
  assign n22564 = n1265 & ~n22563 ;
  assign n22565 = n1269 & ~n22564 ;
  assign n22566 = n1273 & ~n22565 ;
  assign n22567 = n2566 & ~n22566 ;
  assign n22568 = n2568 & ~n22567 ;
  assign n22569 = n3105 & ~n22568 ;
  assign n22570 = n1625 & ~n22569 ;
  assign n22571 = n1629 & ~n22570 ;
  assign n22572 = n1633 & ~n22571 ;
  assign n22573 = n1637 & ~n22572 ;
  assign n22574 = n1641 & ~n22573 ;
  assign n22575 = n1645 & ~n22574 ;
  assign n22576 = n1649 & ~n22575 ;
  assign n22577 = n1653 & ~n22576 ;
  assign n22578 = n1657 & ~n22577 ;
  assign n22579 = n1661 & ~n22578 ;
  assign n22580 = n1665 & ~n22579 ;
  assign n22581 = n1669 & ~n22580 ;
  assign n22582 = n1673 & ~n22581 ;
  assign n22583 = n1677 & ~n22582 ;
  assign n22584 = n1681 & ~n22583 ;
  assign n22585 = n1685 & ~n22584 ;
  assign n22586 = n1689 & ~n22585 ;
  assign n22587 = n1693 & ~n22586 ;
  assign n22588 = n1697 & ~n22587 ;
  assign n22589 = n1701 & ~n22588 ;
  assign n22590 = n1705 & ~n22589 ;
  assign n22591 = n1709 & ~n22590 ;
  assign n22592 = n1713 & ~n22591 ;
  assign n22593 = n1717 & ~n22592 ;
  assign n22594 = n1721 & ~n22593 ;
  assign n22595 = n1725 & ~n22594 ;
  assign n22596 = n1729 & ~n22595 ;
  assign n22597 = n1733 & ~n22596 ;
  assign n22598 = n1737 & ~n22597 ;
  assign n22599 = n1741 & ~n22598 ;
  assign n22600 = n1745 & ~n22599 ;
  assign n22601 = n1749 & ~n22600 ;
  assign n22602 = n1753 & ~n22601 ;
  assign n22603 = n1757 & ~n22602 ;
  assign n22604 = n1761 & ~n22603 ;
  assign n22605 = n1765 & ~n22604 ;
  assign n22606 = n1769 & ~n22605 ;
  assign n22607 = n1773 & ~n22606 ;
  assign n22608 = n1777 & ~n22607 ;
  assign n22609 = n1781 & ~n22608 ;
  assign n22610 = n1785 & ~n22609 ;
  assign n22611 = n1789 & ~n22610 ;
  assign n22612 = n1793 & ~n22611 ;
  assign n22613 = n1797 & ~n22612 ;
  assign n22614 = n1801 & ~n22613 ;
  assign n22615 = n1805 & ~n22614 ;
  assign n22616 = n1809 & ~n22615 ;
  assign n22617 = n1813 & ~n22616 ;
  assign n22618 = n1817 & ~n22617 ;
  assign n22619 = n1821 & ~n22618 ;
  assign n22620 = n1825 & ~n22619 ;
  assign n22621 = n1829 & ~n22620 ;
  assign n22622 = n1833 & ~n22621 ;
  assign n22623 = n1837 & ~n22622 ;
  assign n22624 = n1841 & ~n22623 ;
  assign n22625 = n1845 & ~n22624 ;
  assign n22626 = n1849 & ~n22625 ;
  assign n22627 = n1853 & ~n22626 ;
  assign n22628 = n1857 & ~n22627 ;
  assign n22629 = n1861 & ~n22628 ;
  assign n22630 = n1865 & ~n22629 ;
  assign n22631 = n1869 & ~n22630 ;
  assign n22632 = n1873 & ~n22631 ;
  assign n22633 = n1877 & ~n22632 ;
  assign n22634 = n1881 & ~n22633 ;
  assign n22635 = n1885 & ~n22634 ;
  assign n22636 = n1889 & ~n22635 ;
  assign n22637 = n1893 & ~n22636 ;
  assign n22638 = n1897 & ~n22637 ;
  assign n22639 = n1901 & ~n22638 ;
  assign n22640 = n1905 & ~n22639 ;
  assign n22641 = n1909 & ~n22640 ;
  assign n22642 = n1913 & ~n22641 ;
  assign n22643 = n1917 & ~n22642 ;
  assign n22644 = n1921 & ~n22643 ;
  assign n22645 = x246 & ~n1923 ;
  assign n22646 = ~n22644 & n22645 ;
  assign n22734 = n22646 & x374 ;
  assign n22647 = n1591 & ~n2265 ;
  assign n22648 = n1596 & ~n22647 ;
  assign n22649 = n1600 & ~n22648 ;
  assign n22650 = n1604 & ~n22649 ;
  assign n22651 = n1608 & ~n22650 ;
  assign n22652 = n1612 & ~n22651 ;
  assign n22653 = n2656 & ~n22652 ;
  assign n22654 = n2658 & ~n22653 ;
  assign n22655 = n3192 & ~n22654 ;
  assign n22656 = n1962 & ~n22655 ;
  assign n22657 = n1966 & ~n22656 ;
  assign n22658 = n1970 & ~n22657 ;
  assign n22659 = n1974 & ~n22658 ;
  assign n22660 = n1978 & ~n22659 ;
  assign n22661 = n1982 & ~n22660 ;
  assign n22662 = n1986 & ~n22661 ;
  assign n22663 = n1990 & ~n22662 ;
  assign n22664 = n1994 & ~n22663 ;
  assign n22665 = n1998 & ~n22664 ;
  assign n22666 = n2002 & ~n22665 ;
  assign n22667 = n2006 & ~n22666 ;
  assign n22668 = n2010 & ~n22667 ;
  assign n22669 = n2014 & ~n22668 ;
  assign n22670 = n2018 & ~n22669 ;
  assign n22671 = n2022 & ~n22670 ;
  assign n22672 = n2026 & ~n22671 ;
  assign n22673 = n2030 & ~n22672 ;
  assign n22674 = n2034 & ~n22673 ;
  assign n22675 = n2038 & ~n22674 ;
  assign n22676 = n2042 & ~n22675 ;
  assign n22677 = n2046 & ~n22676 ;
  assign n22678 = n2050 & ~n22677 ;
  assign n22679 = n2054 & ~n22678 ;
  assign n22680 = n2058 & ~n22679 ;
  assign n22681 = n2062 & ~n22680 ;
  assign n22682 = n2066 & ~n22681 ;
  assign n22683 = n2070 & ~n22682 ;
  assign n22684 = n2074 & ~n22683 ;
  assign n22685 = n2078 & ~n22684 ;
  assign n22686 = n2082 & ~n22685 ;
  assign n22687 = n2086 & ~n22686 ;
  assign n22688 = n2090 & ~n22687 ;
  assign n22689 = n2094 & ~n22688 ;
  assign n22690 = n2098 & ~n22689 ;
  assign n22691 = n2102 & ~n22690 ;
  assign n22692 = n2106 & ~n22691 ;
  assign n22693 = n2110 & ~n22692 ;
  assign n22694 = n2114 & ~n22693 ;
  assign n22695 = n2118 & ~n22694 ;
  assign n22696 = n2122 & ~n22695 ;
  assign n22697 = n2126 & ~n22696 ;
  assign n22698 = n2130 & ~n22697 ;
  assign n22699 = n2134 & ~n22698 ;
  assign n22700 = n2138 & ~n22699 ;
  assign n22701 = n2142 & ~n22700 ;
  assign n22702 = n2146 & ~n22701 ;
  assign n22703 = n2150 & ~n22702 ;
  assign n22704 = n2154 & ~n22703 ;
  assign n22705 = n2158 & ~n22704 ;
  assign n22706 = n2162 & ~n22705 ;
  assign n22707 = n2166 & ~n22706 ;
  assign n22708 = n2170 & ~n22707 ;
  assign n22709 = n2174 & ~n22708 ;
  assign n22710 = n2178 & ~n22709 ;
  assign n22711 = n2182 & ~n22710 ;
  assign n22712 = n2186 & ~n22711 ;
  assign n22713 = n2190 & ~n22712 ;
  assign n22714 = n2194 & ~n22713 ;
  assign n22715 = n2198 & ~n22714 ;
  assign n22716 = n2202 & ~n22715 ;
  assign n22717 = n2206 & ~n22716 ;
  assign n22718 = n2210 & ~n22717 ;
  assign n22719 = n2214 & ~n22718 ;
  assign n22720 = n2218 & ~n22719 ;
  assign n22721 = n2222 & ~n22720 ;
  assign n22722 = n2226 & ~n22721 ;
  assign n22723 = n2230 & ~n22722 ;
  assign n22724 = n2234 & ~n22723 ;
  assign n22725 = n2238 & ~n22724 ;
  assign n22726 = n2242 & ~n22725 ;
  assign n22727 = n2246 & ~n22726 ;
  assign n22728 = n2250 & ~n22727 ;
  assign n22729 = n2254 & ~n22728 ;
  assign n22730 = n2258 & ~n22729 ;
  assign n22731 = ~x246 & ~n2260 ;
  assign n22732 = ~n22730 & n22731 ;
  assign n22735 = ~n22732 & ~x374 ;
  assign n22736 = ~n22734 & ~n22735 ;
  assign n22737 = ~n574 & n1932 ;
  assign n22738 = n1937 & ~n22737 ;
  assign n22739 = n1941 & ~n22738 ;
  assign n22740 = n1945 & ~n22739 ;
  assign n22741 = n1949 & ~n22740 ;
  assign n22742 = n1953 & ~n22741 ;
  assign n22743 = n2749 & ~n22742 ;
  assign n22744 = n263 & ~n22743 ;
  assign n22745 = n267 & ~n22744 ;
  assign n22746 = n271 & ~n22745 ;
  assign n22747 = n275 & ~n22746 ;
  assign n22748 = n279 & ~n22747 ;
  assign n22749 = n283 & ~n22748 ;
  assign n22750 = n287 & ~n22749 ;
  assign n22751 = n291 & ~n22750 ;
  assign n22752 = n295 & ~n22751 ;
  assign n22753 = n299 & ~n22752 ;
  assign n22754 = n303 & ~n22753 ;
  assign n22755 = n307 & ~n22754 ;
  assign n22756 = n311 & ~n22755 ;
  assign n22757 = n315 & ~n22756 ;
  assign n22758 = n319 & ~n22757 ;
  assign n22759 = n323 & ~n22758 ;
  assign n22760 = n327 & ~n22759 ;
  assign n22761 = n331 & ~n22760 ;
  assign n22762 = n335 & ~n22761 ;
  assign n22763 = n339 & ~n22762 ;
  assign n22764 = n343 & ~n22763 ;
  assign n22765 = n347 & ~n22764 ;
  assign n22766 = n351 & ~n22765 ;
  assign n22767 = n355 & ~n22766 ;
  assign n22768 = n359 & ~n22767 ;
  assign n22769 = n363 & ~n22768 ;
  assign n22770 = n367 & ~n22769 ;
  assign n22771 = n371 & ~n22770 ;
  assign n22772 = n375 & ~n22771 ;
  assign n22773 = n379 & ~n22772 ;
  assign n22774 = n383 & ~n22773 ;
  assign n22775 = n387 & ~n22774 ;
  assign n22776 = n391 & ~n22775 ;
  assign n22777 = n395 & ~n22776 ;
  assign n22778 = n399 & ~n22777 ;
  assign n22779 = n403 & ~n22778 ;
  assign n22780 = n407 & ~n22779 ;
  assign n22781 = n411 & ~n22780 ;
  assign n22782 = n415 & ~n22781 ;
  assign n22783 = n419 & ~n22782 ;
  assign n22784 = n423 & ~n22783 ;
  assign n22785 = n427 & ~n22784 ;
  assign n22786 = n431 & ~n22785 ;
  assign n22787 = n435 & ~n22786 ;
  assign n22788 = n439 & ~n22787 ;
  assign n22789 = n443 & ~n22788 ;
  assign n22790 = n447 & ~n22789 ;
  assign n22791 = n451 & ~n22790 ;
  assign n22792 = n455 & ~n22791 ;
  assign n22793 = n459 & ~n22792 ;
  assign n22794 = n463 & ~n22793 ;
  assign n22795 = n467 & ~n22794 ;
  assign n22796 = n471 & ~n22795 ;
  assign n22797 = n475 & ~n22796 ;
  assign n22798 = n479 & ~n22797 ;
  assign n22799 = n483 & ~n22798 ;
  assign n22800 = n487 & ~n22799 ;
  assign n22801 = n491 & ~n22800 ;
  assign n22802 = n495 & ~n22801 ;
  assign n22803 = n499 & ~n22802 ;
  assign n22804 = n503 & ~n22803 ;
  assign n22805 = n507 & ~n22804 ;
  assign n22806 = n511 & ~n22805 ;
  assign n22807 = n515 & ~n22806 ;
  assign n22808 = n519 & ~n22807 ;
  assign n22809 = n523 & ~n22808 ;
  assign n22810 = n527 & ~n22809 ;
  assign n22811 = n531 & ~n22810 ;
  assign n22812 = n535 & ~n22811 ;
  assign n22813 = n539 & ~n22812 ;
  assign n22814 = n543 & ~n22813 ;
  assign n22815 = n547 & ~n22814 ;
  assign n22816 = n551 & ~n22815 ;
  assign n22817 = n555 & ~n22816 ;
  assign n22818 = n559 & ~n22817 ;
  assign n22819 = n563 & ~n22818 ;
  assign n22820 = n567 & ~n22819 ;
  assign n22821 = x247 & ~n569 ;
  assign n22822 = ~n22820 & n22821 ;
  assign n22910 = n22822 & x375 ;
  assign n22823 = ~n913 & n2269 ;
  assign n22824 = n2274 & ~n22823 ;
  assign n22825 = n2278 & ~n22824 ;
  assign n22826 = n2282 & ~n22825 ;
  assign n22827 = n2286 & ~n22826 ;
  assign n22828 = n2290 & ~n22827 ;
  assign n22829 = n2836 & ~n22828 ;
  assign n22830 = n602 & ~n22829 ;
  assign n22831 = n606 & ~n22830 ;
  assign n22832 = n610 & ~n22831 ;
  assign n22833 = n614 & ~n22832 ;
  assign n22834 = n618 & ~n22833 ;
  assign n22835 = n622 & ~n22834 ;
  assign n22836 = n626 & ~n22835 ;
  assign n22837 = n630 & ~n22836 ;
  assign n22838 = n634 & ~n22837 ;
  assign n22839 = n638 & ~n22838 ;
  assign n22840 = n642 & ~n22839 ;
  assign n22841 = n646 & ~n22840 ;
  assign n22842 = n650 & ~n22841 ;
  assign n22843 = n654 & ~n22842 ;
  assign n22844 = n658 & ~n22843 ;
  assign n22845 = n662 & ~n22844 ;
  assign n22846 = n666 & ~n22845 ;
  assign n22847 = n670 & ~n22846 ;
  assign n22848 = n674 & ~n22847 ;
  assign n22849 = n678 & ~n22848 ;
  assign n22850 = n682 & ~n22849 ;
  assign n22851 = n686 & ~n22850 ;
  assign n22852 = n690 & ~n22851 ;
  assign n22853 = n694 & ~n22852 ;
  assign n22854 = n698 & ~n22853 ;
  assign n22855 = n702 & ~n22854 ;
  assign n22856 = n706 & ~n22855 ;
  assign n22857 = n710 & ~n22856 ;
  assign n22858 = n714 & ~n22857 ;
  assign n22859 = n718 & ~n22858 ;
  assign n22860 = n722 & ~n22859 ;
  assign n22861 = n726 & ~n22860 ;
  assign n22862 = n730 & ~n22861 ;
  assign n22863 = n734 & ~n22862 ;
  assign n22864 = n738 & ~n22863 ;
  assign n22865 = n742 & ~n22864 ;
  assign n22866 = n746 & ~n22865 ;
  assign n22867 = n750 & ~n22866 ;
  assign n22868 = n754 & ~n22867 ;
  assign n22869 = n758 & ~n22868 ;
  assign n22870 = n762 & ~n22869 ;
  assign n22871 = n766 & ~n22870 ;
  assign n22872 = n770 & ~n22871 ;
  assign n22873 = n774 & ~n22872 ;
  assign n22874 = n778 & ~n22873 ;
  assign n22875 = n782 & ~n22874 ;
  assign n22876 = n786 & ~n22875 ;
  assign n22877 = n790 & ~n22876 ;
  assign n22878 = n794 & ~n22877 ;
  assign n22879 = n798 & ~n22878 ;
  assign n22880 = n802 & ~n22879 ;
  assign n22881 = n806 & ~n22880 ;
  assign n22882 = n810 & ~n22881 ;
  assign n22883 = n814 & ~n22882 ;
  assign n22884 = n818 & ~n22883 ;
  assign n22885 = n822 & ~n22884 ;
  assign n22886 = n826 & ~n22885 ;
  assign n22887 = n830 & ~n22886 ;
  assign n22888 = n834 & ~n22887 ;
  assign n22889 = n838 & ~n22888 ;
  assign n22890 = n842 & ~n22889 ;
  assign n22891 = n846 & ~n22890 ;
  assign n22892 = n850 & ~n22891 ;
  assign n22893 = n854 & ~n22892 ;
  assign n22894 = n858 & ~n22893 ;
  assign n22895 = n862 & ~n22894 ;
  assign n22896 = n866 & ~n22895 ;
  assign n22897 = n870 & ~n22896 ;
  assign n22898 = n874 & ~n22897 ;
  assign n22899 = n878 & ~n22898 ;
  assign n22900 = n882 & ~n22899 ;
  assign n22901 = n886 & ~n22900 ;
  assign n22902 = n890 & ~n22901 ;
  assign n22903 = n894 & ~n22902 ;
  assign n22904 = n898 & ~n22903 ;
  assign n22905 = n902 & ~n22904 ;
  assign n22906 = n906 & ~n22905 ;
  assign n22907 = ~x247 & ~n908 ;
  assign n22908 = ~n22906 & n22907 ;
  assign n22911 = ~n22908 & ~x375 ;
  assign n22912 = ~n22910 & ~n22911 ;
  assign n22913 = n578 & ~n1256 ;
  assign n22914 = n583 & ~n22913 ;
  assign n22915 = n587 & ~n22914 ;
  assign n22916 = n591 & ~n22915 ;
  assign n22917 = n2382 & ~n22916 ;
  assign n22918 = n2384 & ~n22917 ;
  assign n22919 = n2927 & ~n22918 ;
  assign n22920 = n945 & ~n22919 ;
  assign n22921 = n949 & ~n22920 ;
  assign n22922 = n953 & ~n22921 ;
  assign n22923 = n957 & ~n22922 ;
  assign n22924 = n961 & ~n22923 ;
  assign n22925 = n965 & ~n22924 ;
  assign n22926 = n969 & ~n22925 ;
  assign n22927 = n973 & ~n22926 ;
  assign n22928 = n977 & ~n22927 ;
  assign n22929 = n981 & ~n22928 ;
  assign n22930 = n985 & ~n22929 ;
  assign n22931 = n989 & ~n22930 ;
  assign n22932 = n993 & ~n22931 ;
  assign n22933 = n997 & ~n22932 ;
  assign n22934 = n1001 & ~n22933 ;
  assign n22935 = n1005 & ~n22934 ;
  assign n22936 = n1009 & ~n22935 ;
  assign n22937 = n1013 & ~n22936 ;
  assign n22938 = n1017 & ~n22937 ;
  assign n22939 = n1021 & ~n22938 ;
  assign n22940 = n1025 & ~n22939 ;
  assign n22941 = n1029 & ~n22940 ;
  assign n22942 = n1033 & ~n22941 ;
  assign n22943 = n1037 & ~n22942 ;
  assign n22944 = n1041 & ~n22943 ;
  assign n22945 = n1045 & ~n22944 ;
  assign n22946 = n1049 & ~n22945 ;
  assign n22947 = n1053 & ~n22946 ;
  assign n22948 = n1057 & ~n22947 ;
  assign n22949 = n1061 & ~n22948 ;
  assign n22950 = n1065 & ~n22949 ;
  assign n22951 = n1069 & ~n22950 ;
  assign n22952 = n1073 & ~n22951 ;
  assign n22953 = n1077 & ~n22952 ;
  assign n22954 = n1081 & ~n22953 ;
  assign n22955 = n1085 & ~n22954 ;
  assign n22956 = n1089 & ~n22955 ;
  assign n22957 = n1093 & ~n22956 ;
  assign n22958 = n1097 & ~n22957 ;
  assign n22959 = n1101 & ~n22958 ;
  assign n22960 = n1105 & ~n22959 ;
  assign n22961 = n1109 & ~n22960 ;
  assign n22962 = n1113 & ~n22961 ;
  assign n22963 = n1117 & ~n22962 ;
  assign n22964 = n1121 & ~n22963 ;
  assign n22965 = n1125 & ~n22964 ;
  assign n22966 = n1129 & ~n22965 ;
  assign n22967 = n1133 & ~n22966 ;
  assign n22968 = n1137 & ~n22967 ;
  assign n22969 = n1141 & ~n22968 ;
  assign n22970 = n1145 & ~n22969 ;
  assign n22971 = n1149 & ~n22970 ;
  assign n22972 = n1153 & ~n22971 ;
  assign n22973 = n1157 & ~n22972 ;
  assign n22974 = n1161 & ~n22973 ;
  assign n22975 = n1165 & ~n22974 ;
  assign n22976 = n1169 & ~n22975 ;
  assign n22977 = n1173 & ~n22976 ;
  assign n22978 = n1177 & ~n22977 ;
  assign n22979 = n1181 & ~n22978 ;
  assign n22980 = n1185 & ~n22979 ;
  assign n22981 = n1189 & ~n22980 ;
  assign n22982 = n1193 & ~n22981 ;
  assign n22983 = n1197 & ~n22982 ;
  assign n22984 = n1201 & ~n22983 ;
  assign n22985 = n1205 & ~n22984 ;
  assign n22986 = n1209 & ~n22985 ;
  assign n22987 = n1213 & ~n22986 ;
  assign n22988 = n1217 & ~n22987 ;
  assign n22989 = n1221 & ~n22988 ;
  assign n22990 = n1225 & ~n22989 ;
  assign n22991 = n1229 & ~n22990 ;
  assign n22992 = n1233 & ~n22991 ;
  assign n22993 = n1237 & ~n22992 ;
  assign n22994 = n1241 & ~n22993 ;
  assign n22995 = n1245 & ~n22994 ;
  assign n22996 = n1249 & ~n22995 ;
  assign n22997 = x248 & ~n1251 ;
  assign n22998 = ~n22996 & n22997 ;
  assign n23086 = n22998 & x376 ;
  assign n22999 = n917 & ~n1595 ;
  assign n23000 = n922 & ~n22999 ;
  assign n23001 = n926 & ~n23000 ;
  assign n23002 = n930 & ~n23001 ;
  assign n23003 = n2472 & ~n23002 ;
  assign n23004 = n2474 & ~n23003 ;
  assign n23005 = n3014 & ~n23004 ;
  assign n23006 = n1284 & ~n23005 ;
  assign n23007 = n1288 & ~n23006 ;
  assign n23008 = n1292 & ~n23007 ;
  assign n23009 = n1296 & ~n23008 ;
  assign n23010 = n1300 & ~n23009 ;
  assign n23011 = n1304 & ~n23010 ;
  assign n23012 = n1308 & ~n23011 ;
  assign n23013 = n1312 & ~n23012 ;
  assign n23014 = n1316 & ~n23013 ;
  assign n23015 = n1320 & ~n23014 ;
  assign n23016 = n1324 & ~n23015 ;
  assign n23017 = n1328 & ~n23016 ;
  assign n23018 = n1332 & ~n23017 ;
  assign n23019 = n1336 & ~n23018 ;
  assign n23020 = n1340 & ~n23019 ;
  assign n23021 = n1344 & ~n23020 ;
  assign n23022 = n1348 & ~n23021 ;
  assign n23023 = n1352 & ~n23022 ;
  assign n23024 = n1356 & ~n23023 ;
  assign n23025 = n1360 & ~n23024 ;
  assign n23026 = n1364 & ~n23025 ;
  assign n23027 = n1368 & ~n23026 ;
  assign n23028 = n1372 & ~n23027 ;
  assign n23029 = n1376 & ~n23028 ;
  assign n23030 = n1380 & ~n23029 ;
  assign n23031 = n1384 & ~n23030 ;
  assign n23032 = n1388 & ~n23031 ;
  assign n23033 = n1392 & ~n23032 ;
  assign n23034 = n1396 & ~n23033 ;
  assign n23035 = n1400 & ~n23034 ;
  assign n23036 = n1404 & ~n23035 ;
  assign n23037 = n1408 & ~n23036 ;
  assign n23038 = n1412 & ~n23037 ;
  assign n23039 = n1416 & ~n23038 ;
  assign n23040 = n1420 & ~n23039 ;
  assign n23041 = n1424 & ~n23040 ;
  assign n23042 = n1428 & ~n23041 ;
  assign n23043 = n1432 & ~n23042 ;
  assign n23044 = n1436 & ~n23043 ;
  assign n23045 = n1440 & ~n23044 ;
  assign n23046 = n1444 & ~n23045 ;
  assign n23047 = n1448 & ~n23046 ;
  assign n23048 = n1452 & ~n23047 ;
  assign n23049 = n1456 & ~n23048 ;
  assign n23050 = n1460 & ~n23049 ;
  assign n23051 = n1464 & ~n23050 ;
  assign n23052 = n1468 & ~n23051 ;
  assign n23053 = n1472 & ~n23052 ;
  assign n23054 = n1476 & ~n23053 ;
  assign n23055 = n1480 & ~n23054 ;
  assign n23056 = n1484 & ~n23055 ;
  assign n23057 = n1488 & ~n23056 ;
  assign n23058 = n1492 & ~n23057 ;
  assign n23059 = n1496 & ~n23058 ;
  assign n23060 = n1500 & ~n23059 ;
  assign n23061 = n1504 & ~n23060 ;
  assign n23062 = n1508 & ~n23061 ;
  assign n23063 = n1512 & ~n23062 ;
  assign n23064 = n1516 & ~n23063 ;
  assign n23065 = n1520 & ~n23064 ;
  assign n23066 = n1524 & ~n23065 ;
  assign n23067 = n1528 & ~n23066 ;
  assign n23068 = n1532 & ~n23067 ;
  assign n23069 = n1536 & ~n23068 ;
  assign n23070 = n1540 & ~n23069 ;
  assign n23071 = n1544 & ~n23070 ;
  assign n23072 = n1548 & ~n23071 ;
  assign n23073 = n1552 & ~n23072 ;
  assign n23074 = n1556 & ~n23073 ;
  assign n23075 = n1560 & ~n23074 ;
  assign n23076 = n1564 & ~n23075 ;
  assign n23077 = n1568 & ~n23076 ;
  assign n23078 = n1572 & ~n23077 ;
  assign n23079 = n1576 & ~n23078 ;
  assign n23080 = n1580 & ~n23079 ;
  assign n23081 = n1584 & ~n23080 ;
  assign n23082 = n1588 & ~n23081 ;
  assign n23083 = ~x248 & ~n1590 ;
  assign n23084 = ~n23082 & n23083 ;
  assign n23087 = ~n23084 & ~x376 ;
  assign n23088 = ~n23086 & ~n23087 ;
  assign n23089 = n1260 & ~n1936 ;
  assign n23090 = n1265 & ~n23089 ;
  assign n23091 = n1269 & ~n23090 ;
  assign n23092 = n1273 & ~n23091 ;
  assign n23093 = n2566 & ~n23092 ;
  assign n23094 = n2568 & ~n23093 ;
  assign n23095 = n3105 & ~n23094 ;
  assign n23096 = n1625 & ~n23095 ;
  assign n23097 = n1629 & ~n23096 ;
  assign n23098 = n1633 & ~n23097 ;
  assign n23099 = n1637 & ~n23098 ;
  assign n23100 = n1641 & ~n23099 ;
  assign n23101 = n1645 & ~n23100 ;
  assign n23102 = n1649 & ~n23101 ;
  assign n23103 = n1653 & ~n23102 ;
  assign n23104 = n1657 & ~n23103 ;
  assign n23105 = n1661 & ~n23104 ;
  assign n23106 = n1665 & ~n23105 ;
  assign n23107 = n1669 & ~n23106 ;
  assign n23108 = n1673 & ~n23107 ;
  assign n23109 = n1677 & ~n23108 ;
  assign n23110 = n1681 & ~n23109 ;
  assign n23111 = n1685 & ~n23110 ;
  assign n23112 = n1689 & ~n23111 ;
  assign n23113 = n1693 & ~n23112 ;
  assign n23114 = n1697 & ~n23113 ;
  assign n23115 = n1701 & ~n23114 ;
  assign n23116 = n1705 & ~n23115 ;
  assign n23117 = n1709 & ~n23116 ;
  assign n23118 = n1713 & ~n23117 ;
  assign n23119 = n1717 & ~n23118 ;
  assign n23120 = n1721 & ~n23119 ;
  assign n23121 = n1725 & ~n23120 ;
  assign n23122 = n1729 & ~n23121 ;
  assign n23123 = n1733 & ~n23122 ;
  assign n23124 = n1737 & ~n23123 ;
  assign n23125 = n1741 & ~n23124 ;
  assign n23126 = n1745 & ~n23125 ;
  assign n23127 = n1749 & ~n23126 ;
  assign n23128 = n1753 & ~n23127 ;
  assign n23129 = n1757 & ~n23128 ;
  assign n23130 = n1761 & ~n23129 ;
  assign n23131 = n1765 & ~n23130 ;
  assign n23132 = n1769 & ~n23131 ;
  assign n23133 = n1773 & ~n23132 ;
  assign n23134 = n1777 & ~n23133 ;
  assign n23135 = n1781 & ~n23134 ;
  assign n23136 = n1785 & ~n23135 ;
  assign n23137 = n1789 & ~n23136 ;
  assign n23138 = n1793 & ~n23137 ;
  assign n23139 = n1797 & ~n23138 ;
  assign n23140 = n1801 & ~n23139 ;
  assign n23141 = n1805 & ~n23140 ;
  assign n23142 = n1809 & ~n23141 ;
  assign n23143 = n1813 & ~n23142 ;
  assign n23144 = n1817 & ~n23143 ;
  assign n23145 = n1821 & ~n23144 ;
  assign n23146 = n1825 & ~n23145 ;
  assign n23147 = n1829 & ~n23146 ;
  assign n23148 = n1833 & ~n23147 ;
  assign n23149 = n1837 & ~n23148 ;
  assign n23150 = n1841 & ~n23149 ;
  assign n23151 = n1845 & ~n23150 ;
  assign n23152 = n1849 & ~n23151 ;
  assign n23153 = n1853 & ~n23152 ;
  assign n23154 = n1857 & ~n23153 ;
  assign n23155 = n1861 & ~n23154 ;
  assign n23156 = n1865 & ~n23155 ;
  assign n23157 = n1869 & ~n23156 ;
  assign n23158 = n1873 & ~n23157 ;
  assign n23159 = n1877 & ~n23158 ;
  assign n23160 = n1881 & ~n23159 ;
  assign n23161 = n1885 & ~n23160 ;
  assign n23162 = n1889 & ~n23161 ;
  assign n23163 = n1893 & ~n23162 ;
  assign n23164 = n1897 & ~n23163 ;
  assign n23165 = n1901 & ~n23164 ;
  assign n23166 = n1905 & ~n23165 ;
  assign n23167 = n1909 & ~n23166 ;
  assign n23168 = n1913 & ~n23167 ;
  assign n23169 = n1917 & ~n23168 ;
  assign n23170 = n1921 & ~n23169 ;
  assign n23171 = n1925 & ~n23170 ;
  assign n23172 = n1929 & ~n23171 ;
  assign n23173 = x249 & ~n1931 ;
  assign n23174 = ~n23172 & n23173 ;
  assign n23262 = n23174 & x377 ;
  assign n23175 = n1599 & ~n2273 ;
  assign n23176 = n1604 & ~n23175 ;
  assign n23177 = n1608 & ~n23176 ;
  assign n23178 = n1612 & ~n23177 ;
  assign n23179 = n2656 & ~n23178 ;
  assign n23180 = n2658 & ~n23179 ;
  assign n23181 = n3192 & ~n23180 ;
  assign n23182 = n1962 & ~n23181 ;
  assign n23183 = n1966 & ~n23182 ;
  assign n23184 = n1970 & ~n23183 ;
  assign n23185 = n1974 & ~n23184 ;
  assign n23186 = n1978 & ~n23185 ;
  assign n23187 = n1982 & ~n23186 ;
  assign n23188 = n1986 & ~n23187 ;
  assign n23189 = n1990 & ~n23188 ;
  assign n23190 = n1994 & ~n23189 ;
  assign n23191 = n1998 & ~n23190 ;
  assign n23192 = n2002 & ~n23191 ;
  assign n23193 = n2006 & ~n23192 ;
  assign n23194 = n2010 & ~n23193 ;
  assign n23195 = n2014 & ~n23194 ;
  assign n23196 = n2018 & ~n23195 ;
  assign n23197 = n2022 & ~n23196 ;
  assign n23198 = n2026 & ~n23197 ;
  assign n23199 = n2030 & ~n23198 ;
  assign n23200 = n2034 & ~n23199 ;
  assign n23201 = n2038 & ~n23200 ;
  assign n23202 = n2042 & ~n23201 ;
  assign n23203 = n2046 & ~n23202 ;
  assign n23204 = n2050 & ~n23203 ;
  assign n23205 = n2054 & ~n23204 ;
  assign n23206 = n2058 & ~n23205 ;
  assign n23207 = n2062 & ~n23206 ;
  assign n23208 = n2066 & ~n23207 ;
  assign n23209 = n2070 & ~n23208 ;
  assign n23210 = n2074 & ~n23209 ;
  assign n23211 = n2078 & ~n23210 ;
  assign n23212 = n2082 & ~n23211 ;
  assign n23213 = n2086 & ~n23212 ;
  assign n23214 = n2090 & ~n23213 ;
  assign n23215 = n2094 & ~n23214 ;
  assign n23216 = n2098 & ~n23215 ;
  assign n23217 = n2102 & ~n23216 ;
  assign n23218 = n2106 & ~n23217 ;
  assign n23219 = n2110 & ~n23218 ;
  assign n23220 = n2114 & ~n23219 ;
  assign n23221 = n2118 & ~n23220 ;
  assign n23222 = n2122 & ~n23221 ;
  assign n23223 = n2126 & ~n23222 ;
  assign n23224 = n2130 & ~n23223 ;
  assign n23225 = n2134 & ~n23224 ;
  assign n23226 = n2138 & ~n23225 ;
  assign n23227 = n2142 & ~n23226 ;
  assign n23228 = n2146 & ~n23227 ;
  assign n23229 = n2150 & ~n23228 ;
  assign n23230 = n2154 & ~n23229 ;
  assign n23231 = n2158 & ~n23230 ;
  assign n23232 = n2162 & ~n23231 ;
  assign n23233 = n2166 & ~n23232 ;
  assign n23234 = n2170 & ~n23233 ;
  assign n23235 = n2174 & ~n23234 ;
  assign n23236 = n2178 & ~n23235 ;
  assign n23237 = n2182 & ~n23236 ;
  assign n23238 = n2186 & ~n23237 ;
  assign n23239 = n2190 & ~n23238 ;
  assign n23240 = n2194 & ~n23239 ;
  assign n23241 = n2198 & ~n23240 ;
  assign n23242 = n2202 & ~n23241 ;
  assign n23243 = n2206 & ~n23242 ;
  assign n23244 = n2210 & ~n23243 ;
  assign n23245 = n2214 & ~n23244 ;
  assign n23246 = n2218 & ~n23245 ;
  assign n23247 = n2222 & ~n23246 ;
  assign n23248 = n2226 & ~n23247 ;
  assign n23249 = n2230 & ~n23248 ;
  assign n23250 = n2234 & ~n23249 ;
  assign n23251 = n2238 & ~n23250 ;
  assign n23252 = n2242 & ~n23251 ;
  assign n23253 = n2246 & ~n23252 ;
  assign n23254 = n2250 & ~n23253 ;
  assign n23255 = n2254 & ~n23254 ;
  assign n23256 = n2258 & ~n23255 ;
  assign n23257 = n2262 & ~n23256 ;
  assign n23258 = n2266 & ~n23257 ;
  assign n23259 = ~x249 & ~n2268 ;
  assign n23260 = ~n23258 & n23259 ;
  assign n23263 = ~n23260 & ~x377 ;
  assign n23264 = ~n23262 & ~n23263 ;
  assign n23265 = ~n582 & n1940 ;
  assign n23266 = n1945 & ~n23265 ;
  assign n23267 = n1949 & ~n23266 ;
  assign n23268 = n1953 & ~n23267 ;
  assign n23269 = n2749 & ~n23268 ;
  assign n23270 = n263 & ~n23269 ;
  assign n23271 = n267 & ~n23270 ;
  assign n23272 = n271 & ~n23271 ;
  assign n23273 = n275 & ~n23272 ;
  assign n23274 = n279 & ~n23273 ;
  assign n23275 = n283 & ~n23274 ;
  assign n23276 = n287 & ~n23275 ;
  assign n23277 = n291 & ~n23276 ;
  assign n23278 = n295 & ~n23277 ;
  assign n23279 = n299 & ~n23278 ;
  assign n23280 = n303 & ~n23279 ;
  assign n23281 = n307 & ~n23280 ;
  assign n23282 = n311 & ~n23281 ;
  assign n23283 = n315 & ~n23282 ;
  assign n23284 = n319 & ~n23283 ;
  assign n23285 = n323 & ~n23284 ;
  assign n23286 = n327 & ~n23285 ;
  assign n23287 = n331 & ~n23286 ;
  assign n23288 = n335 & ~n23287 ;
  assign n23289 = n339 & ~n23288 ;
  assign n23290 = n343 & ~n23289 ;
  assign n23291 = n347 & ~n23290 ;
  assign n23292 = n351 & ~n23291 ;
  assign n23293 = n355 & ~n23292 ;
  assign n23294 = n359 & ~n23293 ;
  assign n23295 = n363 & ~n23294 ;
  assign n23296 = n367 & ~n23295 ;
  assign n23297 = n371 & ~n23296 ;
  assign n23298 = n375 & ~n23297 ;
  assign n23299 = n379 & ~n23298 ;
  assign n23300 = n383 & ~n23299 ;
  assign n23301 = n387 & ~n23300 ;
  assign n23302 = n391 & ~n23301 ;
  assign n23303 = n395 & ~n23302 ;
  assign n23304 = n399 & ~n23303 ;
  assign n23305 = n403 & ~n23304 ;
  assign n23306 = n407 & ~n23305 ;
  assign n23307 = n411 & ~n23306 ;
  assign n23308 = n415 & ~n23307 ;
  assign n23309 = n419 & ~n23308 ;
  assign n23310 = n423 & ~n23309 ;
  assign n23311 = n427 & ~n23310 ;
  assign n23312 = n431 & ~n23311 ;
  assign n23313 = n435 & ~n23312 ;
  assign n23314 = n439 & ~n23313 ;
  assign n23315 = n443 & ~n23314 ;
  assign n23316 = n447 & ~n23315 ;
  assign n23317 = n451 & ~n23316 ;
  assign n23318 = n455 & ~n23317 ;
  assign n23319 = n459 & ~n23318 ;
  assign n23320 = n463 & ~n23319 ;
  assign n23321 = n467 & ~n23320 ;
  assign n23322 = n471 & ~n23321 ;
  assign n23323 = n475 & ~n23322 ;
  assign n23324 = n479 & ~n23323 ;
  assign n23325 = n483 & ~n23324 ;
  assign n23326 = n487 & ~n23325 ;
  assign n23327 = n491 & ~n23326 ;
  assign n23328 = n495 & ~n23327 ;
  assign n23329 = n499 & ~n23328 ;
  assign n23330 = n503 & ~n23329 ;
  assign n23331 = n507 & ~n23330 ;
  assign n23332 = n511 & ~n23331 ;
  assign n23333 = n515 & ~n23332 ;
  assign n23334 = n519 & ~n23333 ;
  assign n23335 = n523 & ~n23334 ;
  assign n23336 = n527 & ~n23335 ;
  assign n23337 = n531 & ~n23336 ;
  assign n23338 = n535 & ~n23337 ;
  assign n23339 = n539 & ~n23338 ;
  assign n23340 = n543 & ~n23339 ;
  assign n23341 = n547 & ~n23340 ;
  assign n23342 = n551 & ~n23341 ;
  assign n23343 = n555 & ~n23342 ;
  assign n23344 = n559 & ~n23343 ;
  assign n23345 = n563 & ~n23344 ;
  assign n23346 = n567 & ~n23345 ;
  assign n23347 = n571 & ~n23346 ;
  assign n23348 = n575 & ~n23347 ;
  assign n23349 = x250 & ~n577 ;
  assign n23350 = ~n23348 & n23349 ;
  assign n23438 = n23350 & x378 ;
  assign n23351 = ~n921 & n2277 ;
  assign n23352 = n2282 & ~n23351 ;
  assign n23353 = n2286 & ~n23352 ;
  assign n23354 = n2290 & ~n23353 ;
  assign n23355 = n2836 & ~n23354 ;
  assign n23356 = n602 & ~n23355 ;
  assign n23357 = n606 & ~n23356 ;
  assign n23358 = n610 & ~n23357 ;
  assign n23359 = n614 & ~n23358 ;
  assign n23360 = n618 & ~n23359 ;
  assign n23361 = n622 & ~n23360 ;
  assign n23362 = n626 & ~n23361 ;
  assign n23363 = n630 & ~n23362 ;
  assign n23364 = n634 & ~n23363 ;
  assign n23365 = n638 & ~n23364 ;
  assign n23366 = n642 & ~n23365 ;
  assign n23367 = n646 & ~n23366 ;
  assign n23368 = n650 & ~n23367 ;
  assign n23369 = n654 & ~n23368 ;
  assign n23370 = n658 & ~n23369 ;
  assign n23371 = n662 & ~n23370 ;
  assign n23372 = n666 & ~n23371 ;
  assign n23373 = n670 & ~n23372 ;
  assign n23374 = n674 & ~n23373 ;
  assign n23375 = n678 & ~n23374 ;
  assign n23376 = n682 & ~n23375 ;
  assign n23377 = n686 & ~n23376 ;
  assign n23378 = n690 & ~n23377 ;
  assign n23379 = n694 & ~n23378 ;
  assign n23380 = n698 & ~n23379 ;
  assign n23381 = n702 & ~n23380 ;
  assign n23382 = n706 & ~n23381 ;
  assign n23383 = n710 & ~n23382 ;
  assign n23384 = n714 & ~n23383 ;
  assign n23385 = n718 & ~n23384 ;
  assign n23386 = n722 & ~n23385 ;
  assign n23387 = n726 & ~n23386 ;
  assign n23388 = n730 & ~n23387 ;
  assign n23389 = n734 & ~n23388 ;
  assign n23390 = n738 & ~n23389 ;
  assign n23391 = n742 & ~n23390 ;
  assign n23392 = n746 & ~n23391 ;
  assign n23393 = n750 & ~n23392 ;
  assign n23394 = n754 & ~n23393 ;
  assign n23395 = n758 & ~n23394 ;
  assign n23396 = n762 & ~n23395 ;
  assign n23397 = n766 & ~n23396 ;
  assign n23398 = n770 & ~n23397 ;
  assign n23399 = n774 & ~n23398 ;
  assign n23400 = n778 & ~n23399 ;
  assign n23401 = n782 & ~n23400 ;
  assign n23402 = n786 & ~n23401 ;
  assign n23403 = n790 & ~n23402 ;
  assign n23404 = n794 & ~n23403 ;
  assign n23405 = n798 & ~n23404 ;
  assign n23406 = n802 & ~n23405 ;
  assign n23407 = n806 & ~n23406 ;
  assign n23408 = n810 & ~n23407 ;
  assign n23409 = n814 & ~n23408 ;
  assign n23410 = n818 & ~n23409 ;
  assign n23411 = n822 & ~n23410 ;
  assign n23412 = n826 & ~n23411 ;
  assign n23413 = n830 & ~n23412 ;
  assign n23414 = n834 & ~n23413 ;
  assign n23415 = n838 & ~n23414 ;
  assign n23416 = n842 & ~n23415 ;
  assign n23417 = n846 & ~n23416 ;
  assign n23418 = n850 & ~n23417 ;
  assign n23419 = n854 & ~n23418 ;
  assign n23420 = n858 & ~n23419 ;
  assign n23421 = n862 & ~n23420 ;
  assign n23422 = n866 & ~n23421 ;
  assign n23423 = n870 & ~n23422 ;
  assign n23424 = n874 & ~n23423 ;
  assign n23425 = n878 & ~n23424 ;
  assign n23426 = n882 & ~n23425 ;
  assign n23427 = n886 & ~n23426 ;
  assign n23428 = n890 & ~n23427 ;
  assign n23429 = n894 & ~n23428 ;
  assign n23430 = n898 & ~n23429 ;
  assign n23431 = n902 & ~n23430 ;
  assign n23432 = n906 & ~n23431 ;
  assign n23433 = n910 & ~n23432 ;
  assign n23434 = n914 & ~n23433 ;
  assign n23435 = ~x250 & ~n916 ;
  assign n23436 = ~n23434 & n23435 ;
  assign n23439 = ~n23436 & ~x378 ;
  assign n23440 = ~n23438 & ~n23439 ;
  assign n23441 = n586 & ~n1264 ;
  assign n23442 = n591 & ~n23441 ;
  assign n23443 = n2382 & ~n23442 ;
  assign n23444 = n2384 & ~n23443 ;
  assign n23445 = n2927 & ~n23444 ;
  assign n23446 = n945 & ~n23445 ;
  assign n23447 = n949 & ~n23446 ;
  assign n23448 = n953 & ~n23447 ;
  assign n23449 = n957 & ~n23448 ;
  assign n23450 = n961 & ~n23449 ;
  assign n23451 = n965 & ~n23450 ;
  assign n23452 = n969 & ~n23451 ;
  assign n23453 = n973 & ~n23452 ;
  assign n23454 = n977 & ~n23453 ;
  assign n23455 = n981 & ~n23454 ;
  assign n23456 = n985 & ~n23455 ;
  assign n23457 = n989 & ~n23456 ;
  assign n23458 = n993 & ~n23457 ;
  assign n23459 = n997 & ~n23458 ;
  assign n23460 = n1001 & ~n23459 ;
  assign n23461 = n1005 & ~n23460 ;
  assign n23462 = n1009 & ~n23461 ;
  assign n23463 = n1013 & ~n23462 ;
  assign n23464 = n1017 & ~n23463 ;
  assign n23465 = n1021 & ~n23464 ;
  assign n23466 = n1025 & ~n23465 ;
  assign n23467 = n1029 & ~n23466 ;
  assign n23468 = n1033 & ~n23467 ;
  assign n23469 = n1037 & ~n23468 ;
  assign n23470 = n1041 & ~n23469 ;
  assign n23471 = n1045 & ~n23470 ;
  assign n23472 = n1049 & ~n23471 ;
  assign n23473 = n1053 & ~n23472 ;
  assign n23474 = n1057 & ~n23473 ;
  assign n23475 = n1061 & ~n23474 ;
  assign n23476 = n1065 & ~n23475 ;
  assign n23477 = n1069 & ~n23476 ;
  assign n23478 = n1073 & ~n23477 ;
  assign n23479 = n1077 & ~n23478 ;
  assign n23480 = n1081 & ~n23479 ;
  assign n23481 = n1085 & ~n23480 ;
  assign n23482 = n1089 & ~n23481 ;
  assign n23483 = n1093 & ~n23482 ;
  assign n23484 = n1097 & ~n23483 ;
  assign n23485 = n1101 & ~n23484 ;
  assign n23486 = n1105 & ~n23485 ;
  assign n23487 = n1109 & ~n23486 ;
  assign n23488 = n1113 & ~n23487 ;
  assign n23489 = n1117 & ~n23488 ;
  assign n23490 = n1121 & ~n23489 ;
  assign n23491 = n1125 & ~n23490 ;
  assign n23492 = n1129 & ~n23491 ;
  assign n23493 = n1133 & ~n23492 ;
  assign n23494 = n1137 & ~n23493 ;
  assign n23495 = n1141 & ~n23494 ;
  assign n23496 = n1145 & ~n23495 ;
  assign n23497 = n1149 & ~n23496 ;
  assign n23498 = n1153 & ~n23497 ;
  assign n23499 = n1157 & ~n23498 ;
  assign n23500 = n1161 & ~n23499 ;
  assign n23501 = n1165 & ~n23500 ;
  assign n23502 = n1169 & ~n23501 ;
  assign n23503 = n1173 & ~n23502 ;
  assign n23504 = n1177 & ~n23503 ;
  assign n23505 = n1181 & ~n23504 ;
  assign n23506 = n1185 & ~n23505 ;
  assign n23507 = n1189 & ~n23506 ;
  assign n23508 = n1193 & ~n23507 ;
  assign n23509 = n1197 & ~n23508 ;
  assign n23510 = n1201 & ~n23509 ;
  assign n23511 = n1205 & ~n23510 ;
  assign n23512 = n1209 & ~n23511 ;
  assign n23513 = n1213 & ~n23512 ;
  assign n23514 = n1217 & ~n23513 ;
  assign n23515 = n1221 & ~n23514 ;
  assign n23516 = n1225 & ~n23515 ;
  assign n23517 = n1229 & ~n23516 ;
  assign n23518 = n1233 & ~n23517 ;
  assign n23519 = n1237 & ~n23518 ;
  assign n23520 = n1241 & ~n23519 ;
  assign n23521 = n1245 & ~n23520 ;
  assign n23522 = n1249 & ~n23521 ;
  assign n23523 = n1253 & ~n23522 ;
  assign n23524 = n1257 & ~n23523 ;
  assign n23525 = x251 & ~n1259 ;
  assign n23526 = ~n23524 & n23525 ;
  assign n23614 = n23526 & x379 ;
  assign n23527 = n925 & ~n1603 ;
  assign n23528 = n930 & ~n23527 ;
  assign n23529 = n2472 & ~n23528 ;
  assign n23530 = n2474 & ~n23529 ;
  assign n23531 = n3014 & ~n23530 ;
  assign n23532 = n1284 & ~n23531 ;
  assign n23533 = n1288 & ~n23532 ;
  assign n23534 = n1292 & ~n23533 ;
  assign n23535 = n1296 & ~n23534 ;
  assign n23536 = n1300 & ~n23535 ;
  assign n23537 = n1304 & ~n23536 ;
  assign n23538 = n1308 & ~n23537 ;
  assign n23539 = n1312 & ~n23538 ;
  assign n23540 = n1316 & ~n23539 ;
  assign n23541 = n1320 & ~n23540 ;
  assign n23542 = n1324 & ~n23541 ;
  assign n23543 = n1328 & ~n23542 ;
  assign n23544 = n1332 & ~n23543 ;
  assign n23545 = n1336 & ~n23544 ;
  assign n23546 = n1340 & ~n23545 ;
  assign n23547 = n1344 & ~n23546 ;
  assign n23548 = n1348 & ~n23547 ;
  assign n23549 = n1352 & ~n23548 ;
  assign n23550 = n1356 & ~n23549 ;
  assign n23551 = n1360 & ~n23550 ;
  assign n23552 = n1364 & ~n23551 ;
  assign n23553 = n1368 & ~n23552 ;
  assign n23554 = n1372 & ~n23553 ;
  assign n23555 = n1376 & ~n23554 ;
  assign n23556 = n1380 & ~n23555 ;
  assign n23557 = n1384 & ~n23556 ;
  assign n23558 = n1388 & ~n23557 ;
  assign n23559 = n1392 & ~n23558 ;
  assign n23560 = n1396 & ~n23559 ;
  assign n23561 = n1400 & ~n23560 ;
  assign n23562 = n1404 & ~n23561 ;
  assign n23563 = n1408 & ~n23562 ;
  assign n23564 = n1412 & ~n23563 ;
  assign n23565 = n1416 & ~n23564 ;
  assign n23566 = n1420 & ~n23565 ;
  assign n23567 = n1424 & ~n23566 ;
  assign n23568 = n1428 & ~n23567 ;
  assign n23569 = n1432 & ~n23568 ;
  assign n23570 = n1436 & ~n23569 ;
  assign n23571 = n1440 & ~n23570 ;
  assign n23572 = n1444 & ~n23571 ;
  assign n23573 = n1448 & ~n23572 ;
  assign n23574 = n1452 & ~n23573 ;
  assign n23575 = n1456 & ~n23574 ;
  assign n23576 = n1460 & ~n23575 ;
  assign n23577 = n1464 & ~n23576 ;
  assign n23578 = n1468 & ~n23577 ;
  assign n23579 = n1472 & ~n23578 ;
  assign n23580 = n1476 & ~n23579 ;
  assign n23581 = n1480 & ~n23580 ;
  assign n23582 = n1484 & ~n23581 ;
  assign n23583 = n1488 & ~n23582 ;
  assign n23584 = n1492 & ~n23583 ;
  assign n23585 = n1496 & ~n23584 ;
  assign n23586 = n1500 & ~n23585 ;
  assign n23587 = n1504 & ~n23586 ;
  assign n23588 = n1508 & ~n23587 ;
  assign n23589 = n1512 & ~n23588 ;
  assign n23590 = n1516 & ~n23589 ;
  assign n23591 = n1520 & ~n23590 ;
  assign n23592 = n1524 & ~n23591 ;
  assign n23593 = n1528 & ~n23592 ;
  assign n23594 = n1532 & ~n23593 ;
  assign n23595 = n1536 & ~n23594 ;
  assign n23596 = n1540 & ~n23595 ;
  assign n23597 = n1544 & ~n23596 ;
  assign n23598 = n1548 & ~n23597 ;
  assign n23599 = n1552 & ~n23598 ;
  assign n23600 = n1556 & ~n23599 ;
  assign n23601 = n1560 & ~n23600 ;
  assign n23602 = n1564 & ~n23601 ;
  assign n23603 = n1568 & ~n23602 ;
  assign n23604 = n1572 & ~n23603 ;
  assign n23605 = n1576 & ~n23604 ;
  assign n23606 = n1580 & ~n23605 ;
  assign n23607 = n1584 & ~n23606 ;
  assign n23608 = n1588 & ~n23607 ;
  assign n23609 = n1592 & ~n23608 ;
  assign n23610 = n1596 & ~n23609 ;
  assign n23611 = ~x251 & ~n1598 ;
  assign n23612 = ~n23610 & n23611 ;
  assign n23615 = ~n23612 & ~x379 ;
  assign n23616 = ~n23614 & ~n23615 ;
  assign n23617 = n1268 & ~n1944 ;
  assign n23618 = n1273 & ~n23617 ;
  assign n23619 = n2566 & ~n23618 ;
  assign n23620 = n2568 & ~n23619 ;
  assign n23621 = n3105 & ~n23620 ;
  assign n23622 = n1625 & ~n23621 ;
  assign n23623 = n1629 & ~n23622 ;
  assign n23624 = n1633 & ~n23623 ;
  assign n23625 = n1637 & ~n23624 ;
  assign n23626 = n1641 & ~n23625 ;
  assign n23627 = n1645 & ~n23626 ;
  assign n23628 = n1649 & ~n23627 ;
  assign n23629 = n1653 & ~n23628 ;
  assign n23630 = n1657 & ~n23629 ;
  assign n23631 = n1661 & ~n23630 ;
  assign n23632 = n1665 & ~n23631 ;
  assign n23633 = n1669 & ~n23632 ;
  assign n23634 = n1673 & ~n23633 ;
  assign n23635 = n1677 & ~n23634 ;
  assign n23636 = n1681 & ~n23635 ;
  assign n23637 = n1685 & ~n23636 ;
  assign n23638 = n1689 & ~n23637 ;
  assign n23639 = n1693 & ~n23638 ;
  assign n23640 = n1697 & ~n23639 ;
  assign n23641 = n1701 & ~n23640 ;
  assign n23642 = n1705 & ~n23641 ;
  assign n23643 = n1709 & ~n23642 ;
  assign n23644 = n1713 & ~n23643 ;
  assign n23645 = n1717 & ~n23644 ;
  assign n23646 = n1721 & ~n23645 ;
  assign n23647 = n1725 & ~n23646 ;
  assign n23648 = n1729 & ~n23647 ;
  assign n23649 = n1733 & ~n23648 ;
  assign n23650 = n1737 & ~n23649 ;
  assign n23651 = n1741 & ~n23650 ;
  assign n23652 = n1745 & ~n23651 ;
  assign n23653 = n1749 & ~n23652 ;
  assign n23654 = n1753 & ~n23653 ;
  assign n23655 = n1757 & ~n23654 ;
  assign n23656 = n1761 & ~n23655 ;
  assign n23657 = n1765 & ~n23656 ;
  assign n23658 = n1769 & ~n23657 ;
  assign n23659 = n1773 & ~n23658 ;
  assign n23660 = n1777 & ~n23659 ;
  assign n23661 = n1781 & ~n23660 ;
  assign n23662 = n1785 & ~n23661 ;
  assign n23663 = n1789 & ~n23662 ;
  assign n23664 = n1793 & ~n23663 ;
  assign n23665 = n1797 & ~n23664 ;
  assign n23666 = n1801 & ~n23665 ;
  assign n23667 = n1805 & ~n23666 ;
  assign n23668 = n1809 & ~n23667 ;
  assign n23669 = n1813 & ~n23668 ;
  assign n23670 = n1817 & ~n23669 ;
  assign n23671 = n1821 & ~n23670 ;
  assign n23672 = n1825 & ~n23671 ;
  assign n23673 = n1829 & ~n23672 ;
  assign n23674 = n1833 & ~n23673 ;
  assign n23675 = n1837 & ~n23674 ;
  assign n23676 = n1841 & ~n23675 ;
  assign n23677 = n1845 & ~n23676 ;
  assign n23678 = n1849 & ~n23677 ;
  assign n23679 = n1853 & ~n23678 ;
  assign n23680 = n1857 & ~n23679 ;
  assign n23681 = n1861 & ~n23680 ;
  assign n23682 = n1865 & ~n23681 ;
  assign n23683 = n1869 & ~n23682 ;
  assign n23684 = n1873 & ~n23683 ;
  assign n23685 = n1877 & ~n23684 ;
  assign n23686 = n1881 & ~n23685 ;
  assign n23687 = n1885 & ~n23686 ;
  assign n23688 = n1889 & ~n23687 ;
  assign n23689 = n1893 & ~n23688 ;
  assign n23690 = n1897 & ~n23689 ;
  assign n23691 = n1901 & ~n23690 ;
  assign n23692 = n1905 & ~n23691 ;
  assign n23693 = n1909 & ~n23692 ;
  assign n23694 = n1913 & ~n23693 ;
  assign n23695 = n1917 & ~n23694 ;
  assign n23696 = n1921 & ~n23695 ;
  assign n23697 = n1925 & ~n23696 ;
  assign n23698 = n1929 & ~n23697 ;
  assign n23699 = n1933 & ~n23698 ;
  assign n23700 = n1937 & ~n23699 ;
  assign n23701 = x252 & ~n1939 ;
  assign n23702 = ~n23700 & n23701 ;
  assign n23790 = n23702 & x380 ;
  assign n23703 = n1607 & ~n2281 ;
  assign n23704 = n1612 & ~n23703 ;
  assign n23705 = n2656 & ~n23704 ;
  assign n23706 = n2658 & ~n23705 ;
  assign n23707 = n3192 & ~n23706 ;
  assign n23708 = n1962 & ~n23707 ;
  assign n23709 = n1966 & ~n23708 ;
  assign n23710 = n1970 & ~n23709 ;
  assign n23711 = n1974 & ~n23710 ;
  assign n23712 = n1978 & ~n23711 ;
  assign n23713 = n1982 & ~n23712 ;
  assign n23714 = n1986 & ~n23713 ;
  assign n23715 = n1990 & ~n23714 ;
  assign n23716 = n1994 & ~n23715 ;
  assign n23717 = n1998 & ~n23716 ;
  assign n23718 = n2002 & ~n23717 ;
  assign n23719 = n2006 & ~n23718 ;
  assign n23720 = n2010 & ~n23719 ;
  assign n23721 = n2014 & ~n23720 ;
  assign n23722 = n2018 & ~n23721 ;
  assign n23723 = n2022 & ~n23722 ;
  assign n23724 = n2026 & ~n23723 ;
  assign n23725 = n2030 & ~n23724 ;
  assign n23726 = n2034 & ~n23725 ;
  assign n23727 = n2038 & ~n23726 ;
  assign n23728 = n2042 & ~n23727 ;
  assign n23729 = n2046 & ~n23728 ;
  assign n23730 = n2050 & ~n23729 ;
  assign n23731 = n2054 & ~n23730 ;
  assign n23732 = n2058 & ~n23731 ;
  assign n23733 = n2062 & ~n23732 ;
  assign n23734 = n2066 & ~n23733 ;
  assign n23735 = n2070 & ~n23734 ;
  assign n23736 = n2074 & ~n23735 ;
  assign n23737 = n2078 & ~n23736 ;
  assign n23738 = n2082 & ~n23737 ;
  assign n23739 = n2086 & ~n23738 ;
  assign n23740 = n2090 & ~n23739 ;
  assign n23741 = n2094 & ~n23740 ;
  assign n23742 = n2098 & ~n23741 ;
  assign n23743 = n2102 & ~n23742 ;
  assign n23744 = n2106 & ~n23743 ;
  assign n23745 = n2110 & ~n23744 ;
  assign n23746 = n2114 & ~n23745 ;
  assign n23747 = n2118 & ~n23746 ;
  assign n23748 = n2122 & ~n23747 ;
  assign n23749 = n2126 & ~n23748 ;
  assign n23750 = n2130 & ~n23749 ;
  assign n23751 = n2134 & ~n23750 ;
  assign n23752 = n2138 & ~n23751 ;
  assign n23753 = n2142 & ~n23752 ;
  assign n23754 = n2146 & ~n23753 ;
  assign n23755 = n2150 & ~n23754 ;
  assign n23756 = n2154 & ~n23755 ;
  assign n23757 = n2158 & ~n23756 ;
  assign n23758 = n2162 & ~n23757 ;
  assign n23759 = n2166 & ~n23758 ;
  assign n23760 = n2170 & ~n23759 ;
  assign n23761 = n2174 & ~n23760 ;
  assign n23762 = n2178 & ~n23761 ;
  assign n23763 = n2182 & ~n23762 ;
  assign n23764 = n2186 & ~n23763 ;
  assign n23765 = n2190 & ~n23764 ;
  assign n23766 = n2194 & ~n23765 ;
  assign n23767 = n2198 & ~n23766 ;
  assign n23768 = n2202 & ~n23767 ;
  assign n23769 = n2206 & ~n23768 ;
  assign n23770 = n2210 & ~n23769 ;
  assign n23771 = n2214 & ~n23770 ;
  assign n23772 = n2218 & ~n23771 ;
  assign n23773 = n2222 & ~n23772 ;
  assign n23774 = n2226 & ~n23773 ;
  assign n23775 = n2230 & ~n23774 ;
  assign n23776 = n2234 & ~n23775 ;
  assign n23777 = n2238 & ~n23776 ;
  assign n23778 = n2242 & ~n23777 ;
  assign n23779 = n2246 & ~n23778 ;
  assign n23780 = n2250 & ~n23779 ;
  assign n23781 = n2254 & ~n23780 ;
  assign n23782 = n2258 & ~n23781 ;
  assign n23783 = n2262 & ~n23782 ;
  assign n23784 = n2266 & ~n23783 ;
  assign n23785 = n2270 & ~n23784 ;
  assign n23786 = n2274 & ~n23785 ;
  assign n23787 = ~x252 & ~n2276 ;
  assign n23788 = ~n23786 & n23787 ;
  assign n23791 = ~n23788 & ~x380 ;
  assign n23792 = ~n23790 & ~n23791 ;
  assign n23793 = ~n590 & n1948 ;
  assign n23794 = n1953 & ~n23793 ;
  assign n23795 = n2749 & ~n23794 ;
  assign n23796 = n263 & ~n23795 ;
  assign n23797 = n267 & ~n23796 ;
  assign n23798 = n271 & ~n23797 ;
  assign n23799 = n275 & ~n23798 ;
  assign n23800 = n279 & ~n23799 ;
  assign n23801 = n283 & ~n23800 ;
  assign n23802 = n287 & ~n23801 ;
  assign n23803 = n291 & ~n23802 ;
  assign n23804 = n295 & ~n23803 ;
  assign n23805 = n299 & ~n23804 ;
  assign n23806 = n303 & ~n23805 ;
  assign n23807 = n307 & ~n23806 ;
  assign n23808 = n311 & ~n23807 ;
  assign n23809 = n315 & ~n23808 ;
  assign n23810 = n319 & ~n23809 ;
  assign n23811 = n323 & ~n23810 ;
  assign n23812 = n327 & ~n23811 ;
  assign n23813 = n331 & ~n23812 ;
  assign n23814 = n335 & ~n23813 ;
  assign n23815 = n339 & ~n23814 ;
  assign n23816 = n343 & ~n23815 ;
  assign n23817 = n347 & ~n23816 ;
  assign n23818 = n351 & ~n23817 ;
  assign n23819 = n355 & ~n23818 ;
  assign n23820 = n359 & ~n23819 ;
  assign n23821 = n363 & ~n23820 ;
  assign n23822 = n367 & ~n23821 ;
  assign n23823 = n371 & ~n23822 ;
  assign n23824 = n375 & ~n23823 ;
  assign n23825 = n379 & ~n23824 ;
  assign n23826 = n383 & ~n23825 ;
  assign n23827 = n387 & ~n23826 ;
  assign n23828 = n391 & ~n23827 ;
  assign n23829 = n395 & ~n23828 ;
  assign n23830 = n399 & ~n23829 ;
  assign n23831 = n403 & ~n23830 ;
  assign n23832 = n407 & ~n23831 ;
  assign n23833 = n411 & ~n23832 ;
  assign n23834 = n415 & ~n23833 ;
  assign n23835 = n419 & ~n23834 ;
  assign n23836 = n423 & ~n23835 ;
  assign n23837 = n427 & ~n23836 ;
  assign n23838 = n431 & ~n23837 ;
  assign n23839 = n435 & ~n23838 ;
  assign n23840 = n439 & ~n23839 ;
  assign n23841 = n443 & ~n23840 ;
  assign n23842 = n447 & ~n23841 ;
  assign n23843 = n451 & ~n23842 ;
  assign n23844 = n455 & ~n23843 ;
  assign n23845 = n459 & ~n23844 ;
  assign n23846 = n463 & ~n23845 ;
  assign n23847 = n467 & ~n23846 ;
  assign n23848 = n471 & ~n23847 ;
  assign n23849 = n475 & ~n23848 ;
  assign n23850 = n479 & ~n23849 ;
  assign n23851 = n483 & ~n23850 ;
  assign n23852 = n487 & ~n23851 ;
  assign n23853 = n491 & ~n23852 ;
  assign n23854 = n495 & ~n23853 ;
  assign n23855 = n499 & ~n23854 ;
  assign n23856 = n503 & ~n23855 ;
  assign n23857 = n507 & ~n23856 ;
  assign n23858 = n511 & ~n23857 ;
  assign n23859 = n515 & ~n23858 ;
  assign n23860 = n519 & ~n23859 ;
  assign n23861 = n523 & ~n23860 ;
  assign n23862 = n527 & ~n23861 ;
  assign n23863 = n531 & ~n23862 ;
  assign n23864 = n535 & ~n23863 ;
  assign n23865 = n539 & ~n23864 ;
  assign n23866 = n543 & ~n23865 ;
  assign n23867 = n547 & ~n23866 ;
  assign n23868 = n551 & ~n23867 ;
  assign n23869 = n555 & ~n23868 ;
  assign n23870 = n559 & ~n23869 ;
  assign n23871 = n563 & ~n23870 ;
  assign n23872 = n567 & ~n23871 ;
  assign n23873 = n571 & ~n23872 ;
  assign n23874 = n575 & ~n23873 ;
  assign n23875 = n579 & ~n23874 ;
  assign n23876 = n583 & ~n23875 ;
  assign n23877 = x253 & ~n585 ;
  assign n23878 = ~n23876 & n23877 ;
  assign n23966 = n23878 & x381 ;
  assign n23879 = ~n929 & n2285 ;
  assign n23880 = n2290 & ~n23879 ;
  assign n23881 = n2836 & ~n23880 ;
  assign n23882 = n602 & ~n23881 ;
  assign n23883 = n606 & ~n23882 ;
  assign n23884 = n610 & ~n23883 ;
  assign n23885 = n614 & ~n23884 ;
  assign n23886 = n618 & ~n23885 ;
  assign n23887 = n622 & ~n23886 ;
  assign n23888 = n626 & ~n23887 ;
  assign n23889 = n630 & ~n23888 ;
  assign n23890 = n634 & ~n23889 ;
  assign n23891 = n638 & ~n23890 ;
  assign n23892 = n642 & ~n23891 ;
  assign n23893 = n646 & ~n23892 ;
  assign n23894 = n650 & ~n23893 ;
  assign n23895 = n654 & ~n23894 ;
  assign n23896 = n658 & ~n23895 ;
  assign n23897 = n662 & ~n23896 ;
  assign n23898 = n666 & ~n23897 ;
  assign n23899 = n670 & ~n23898 ;
  assign n23900 = n674 & ~n23899 ;
  assign n23901 = n678 & ~n23900 ;
  assign n23902 = n682 & ~n23901 ;
  assign n23903 = n686 & ~n23902 ;
  assign n23904 = n690 & ~n23903 ;
  assign n23905 = n694 & ~n23904 ;
  assign n23906 = n698 & ~n23905 ;
  assign n23907 = n702 & ~n23906 ;
  assign n23908 = n706 & ~n23907 ;
  assign n23909 = n710 & ~n23908 ;
  assign n23910 = n714 & ~n23909 ;
  assign n23911 = n718 & ~n23910 ;
  assign n23912 = n722 & ~n23911 ;
  assign n23913 = n726 & ~n23912 ;
  assign n23914 = n730 & ~n23913 ;
  assign n23915 = n734 & ~n23914 ;
  assign n23916 = n738 & ~n23915 ;
  assign n23917 = n742 & ~n23916 ;
  assign n23918 = n746 & ~n23917 ;
  assign n23919 = n750 & ~n23918 ;
  assign n23920 = n754 & ~n23919 ;
  assign n23921 = n758 & ~n23920 ;
  assign n23922 = n762 & ~n23921 ;
  assign n23923 = n766 & ~n23922 ;
  assign n23924 = n770 & ~n23923 ;
  assign n23925 = n774 & ~n23924 ;
  assign n23926 = n778 & ~n23925 ;
  assign n23927 = n782 & ~n23926 ;
  assign n23928 = n786 & ~n23927 ;
  assign n23929 = n790 & ~n23928 ;
  assign n23930 = n794 & ~n23929 ;
  assign n23931 = n798 & ~n23930 ;
  assign n23932 = n802 & ~n23931 ;
  assign n23933 = n806 & ~n23932 ;
  assign n23934 = n810 & ~n23933 ;
  assign n23935 = n814 & ~n23934 ;
  assign n23936 = n818 & ~n23935 ;
  assign n23937 = n822 & ~n23936 ;
  assign n23938 = n826 & ~n23937 ;
  assign n23939 = n830 & ~n23938 ;
  assign n23940 = n834 & ~n23939 ;
  assign n23941 = n838 & ~n23940 ;
  assign n23942 = n842 & ~n23941 ;
  assign n23943 = n846 & ~n23942 ;
  assign n23944 = n850 & ~n23943 ;
  assign n23945 = n854 & ~n23944 ;
  assign n23946 = n858 & ~n23945 ;
  assign n23947 = n862 & ~n23946 ;
  assign n23948 = n866 & ~n23947 ;
  assign n23949 = n870 & ~n23948 ;
  assign n23950 = n874 & ~n23949 ;
  assign n23951 = n878 & ~n23950 ;
  assign n23952 = n882 & ~n23951 ;
  assign n23953 = n886 & ~n23952 ;
  assign n23954 = n890 & ~n23953 ;
  assign n23955 = n894 & ~n23954 ;
  assign n23956 = n898 & ~n23955 ;
  assign n23957 = n902 & ~n23956 ;
  assign n23958 = n906 & ~n23957 ;
  assign n23959 = n910 & ~n23958 ;
  assign n23960 = n914 & ~n23959 ;
  assign n23961 = n918 & ~n23960 ;
  assign n23962 = n922 & ~n23961 ;
  assign n23963 = ~x253 & ~n924 ;
  assign n23964 = ~n23962 & n23963 ;
  assign n23967 = ~n23964 & ~x381 ;
  assign n23968 = ~n23966 & ~n23967 ;
  assign n23969 = ~n1272 & n2381 ;
  assign n23970 = n2384 & ~n23969 ;
  assign n23971 = n2927 & ~n23970 ;
  assign n23972 = n945 & ~n23971 ;
  assign n23973 = n949 & ~n23972 ;
  assign n23974 = n953 & ~n23973 ;
  assign n23975 = n957 & ~n23974 ;
  assign n23976 = n961 & ~n23975 ;
  assign n23977 = n965 & ~n23976 ;
  assign n23978 = n969 & ~n23977 ;
  assign n23979 = n973 & ~n23978 ;
  assign n23980 = n977 & ~n23979 ;
  assign n23981 = n981 & ~n23980 ;
  assign n23982 = n985 & ~n23981 ;
  assign n23983 = n989 & ~n23982 ;
  assign n23984 = n993 & ~n23983 ;
  assign n23985 = n997 & ~n23984 ;
  assign n23986 = n1001 & ~n23985 ;
  assign n23987 = n1005 & ~n23986 ;
  assign n23988 = n1009 & ~n23987 ;
  assign n23989 = n1013 & ~n23988 ;
  assign n23990 = n1017 & ~n23989 ;
  assign n23991 = n1021 & ~n23990 ;
  assign n23992 = n1025 & ~n23991 ;
  assign n23993 = n1029 & ~n23992 ;
  assign n23994 = n1033 & ~n23993 ;
  assign n23995 = n1037 & ~n23994 ;
  assign n23996 = n1041 & ~n23995 ;
  assign n23997 = n1045 & ~n23996 ;
  assign n23998 = n1049 & ~n23997 ;
  assign n23999 = n1053 & ~n23998 ;
  assign n24000 = n1057 & ~n23999 ;
  assign n24001 = n1061 & ~n24000 ;
  assign n24002 = n1065 & ~n24001 ;
  assign n24003 = n1069 & ~n24002 ;
  assign n24004 = n1073 & ~n24003 ;
  assign n24005 = n1077 & ~n24004 ;
  assign n24006 = n1081 & ~n24005 ;
  assign n24007 = n1085 & ~n24006 ;
  assign n24008 = n1089 & ~n24007 ;
  assign n24009 = n1093 & ~n24008 ;
  assign n24010 = n1097 & ~n24009 ;
  assign n24011 = n1101 & ~n24010 ;
  assign n24012 = n1105 & ~n24011 ;
  assign n24013 = n1109 & ~n24012 ;
  assign n24014 = n1113 & ~n24013 ;
  assign n24015 = n1117 & ~n24014 ;
  assign n24016 = n1121 & ~n24015 ;
  assign n24017 = n1125 & ~n24016 ;
  assign n24018 = n1129 & ~n24017 ;
  assign n24019 = n1133 & ~n24018 ;
  assign n24020 = n1137 & ~n24019 ;
  assign n24021 = n1141 & ~n24020 ;
  assign n24022 = n1145 & ~n24021 ;
  assign n24023 = n1149 & ~n24022 ;
  assign n24024 = n1153 & ~n24023 ;
  assign n24025 = n1157 & ~n24024 ;
  assign n24026 = n1161 & ~n24025 ;
  assign n24027 = n1165 & ~n24026 ;
  assign n24028 = n1169 & ~n24027 ;
  assign n24029 = n1173 & ~n24028 ;
  assign n24030 = n1177 & ~n24029 ;
  assign n24031 = n1181 & ~n24030 ;
  assign n24032 = n1185 & ~n24031 ;
  assign n24033 = n1189 & ~n24032 ;
  assign n24034 = n1193 & ~n24033 ;
  assign n24035 = n1197 & ~n24034 ;
  assign n24036 = n1201 & ~n24035 ;
  assign n24037 = n1205 & ~n24036 ;
  assign n24038 = n1209 & ~n24037 ;
  assign n24039 = n1213 & ~n24038 ;
  assign n24040 = n1217 & ~n24039 ;
  assign n24041 = n1221 & ~n24040 ;
  assign n24042 = n1225 & ~n24041 ;
  assign n24043 = n1229 & ~n24042 ;
  assign n24044 = n1233 & ~n24043 ;
  assign n24045 = n1237 & ~n24044 ;
  assign n24046 = n1241 & ~n24045 ;
  assign n24047 = n1245 & ~n24046 ;
  assign n24048 = n1249 & ~n24047 ;
  assign n24049 = n1253 & ~n24048 ;
  assign n24050 = n1257 & ~n24049 ;
  assign n24051 = n1261 & ~n24050 ;
  assign n24052 = n1265 & ~n24051 ;
  assign n24053 = x254 & ~n1267 ;
  assign n24054 = ~n24052 & n24053 ;
  assign n24142 = n24054 & x382 ;
  assign n24055 = ~n1611 & n2471 ;
  assign n24056 = n2474 & ~n24055 ;
  assign n24057 = n3014 & ~n24056 ;
  assign n24058 = n1284 & ~n24057 ;
  assign n24059 = n1288 & ~n24058 ;
  assign n24060 = n1292 & ~n24059 ;
  assign n24061 = n1296 & ~n24060 ;
  assign n24062 = n1300 & ~n24061 ;
  assign n24063 = n1304 & ~n24062 ;
  assign n24064 = n1308 & ~n24063 ;
  assign n24065 = n1312 & ~n24064 ;
  assign n24066 = n1316 & ~n24065 ;
  assign n24067 = n1320 & ~n24066 ;
  assign n24068 = n1324 & ~n24067 ;
  assign n24069 = n1328 & ~n24068 ;
  assign n24070 = n1332 & ~n24069 ;
  assign n24071 = n1336 & ~n24070 ;
  assign n24072 = n1340 & ~n24071 ;
  assign n24073 = n1344 & ~n24072 ;
  assign n24074 = n1348 & ~n24073 ;
  assign n24075 = n1352 & ~n24074 ;
  assign n24076 = n1356 & ~n24075 ;
  assign n24077 = n1360 & ~n24076 ;
  assign n24078 = n1364 & ~n24077 ;
  assign n24079 = n1368 & ~n24078 ;
  assign n24080 = n1372 & ~n24079 ;
  assign n24081 = n1376 & ~n24080 ;
  assign n24082 = n1380 & ~n24081 ;
  assign n24083 = n1384 & ~n24082 ;
  assign n24084 = n1388 & ~n24083 ;
  assign n24085 = n1392 & ~n24084 ;
  assign n24086 = n1396 & ~n24085 ;
  assign n24087 = n1400 & ~n24086 ;
  assign n24088 = n1404 & ~n24087 ;
  assign n24089 = n1408 & ~n24088 ;
  assign n24090 = n1412 & ~n24089 ;
  assign n24091 = n1416 & ~n24090 ;
  assign n24092 = n1420 & ~n24091 ;
  assign n24093 = n1424 & ~n24092 ;
  assign n24094 = n1428 & ~n24093 ;
  assign n24095 = n1432 & ~n24094 ;
  assign n24096 = n1436 & ~n24095 ;
  assign n24097 = n1440 & ~n24096 ;
  assign n24098 = n1444 & ~n24097 ;
  assign n24099 = n1448 & ~n24098 ;
  assign n24100 = n1452 & ~n24099 ;
  assign n24101 = n1456 & ~n24100 ;
  assign n24102 = n1460 & ~n24101 ;
  assign n24103 = n1464 & ~n24102 ;
  assign n24104 = n1468 & ~n24103 ;
  assign n24105 = n1472 & ~n24104 ;
  assign n24106 = n1476 & ~n24105 ;
  assign n24107 = n1480 & ~n24106 ;
  assign n24108 = n1484 & ~n24107 ;
  assign n24109 = n1488 & ~n24108 ;
  assign n24110 = n1492 & ~n24109 ;
  assign n24111 = n1496 & ~n24110 ;
  assign n24112 = n1500 & ~n24111 ;
  assign n24113 = n1504 & ~n24112 ;
  assign n24114 = n1508 & ~n24113 ;
  assign n24115 = n1512 & ~n24114 ;
  assign n24116 = n1516 & ~n24115 ;
  assign n24117 = n1520 & ~n24116 ;
  assign n24118 = n1524 & ~n24117 ;
  assign n24119 = n1528 & ~n24118 ;
  assign n24120 = n1532 & ~n24119 ;
  assign n24121 = n1536 & ~n24120 ;
  assign n24122 = n1540 & ~n24121 ;
  assign n24123 = n1544 & ~n24122 ;
  assign n24124 = n1548 & ~n24123 ;
  assign n24125 = n1552 & ~n24124 ;
  assign n24126 = n1556 & ~n24125 ;
  assign n24127 = n1560 & ~n24126 ;
  assign n24128 = n1564 & ~n24127 ;
  assign n24129 = n1568 & ~n24128 ;
  assign n24130 = n1572 & ~n24129 ;
  assign n24131 = n1576 & ~n24130 ;
  assign n24132 = n1580 & ~n24131 ;
  assign n24133 = n1584 & ~n24132 ;
  assign n24134 = n1588 & ~n24133 ;
  assign n24135 = n1592 & ~n24134 ;
  assign n24136 = n1596 & ~n24135 ;
  assign n24137 = n1600 & ~n24136 ;
  assign n24138 = n1604 & ~n24137 ;
  assign n24139 = ~x254 & ~n1606 ;
  assign n24140 = ~n24138 & n24139 ;
  assign n24143 = ~n24140 & ~x382 ;
  assign n24144 = ~n24142 & ~n24143 ;
  assign n24145 = ~n1952 & n2565 ;
  assign n24146 = n2568 & ~n24145 ;
  assign n24147 = n3105 & ~n24146 ;
  assign n24148 = n1625 & ~n24147 ;
  assign n24149 = n1629 & ~n24148 ;
  assign n24150 = n1633 & ~n24149 ;
  assign n24151 = n1637 & ~n24150 ;
  assign n24152 = n1641 & ~n24151 ;
  assign n24153 = n1645 & ~n24152 ;
  assign n24154 = n1649 & ~n24153 ;
  assign n24155 = n1653 & ~n24154 ;
  assign n24156 = n1657 & ~n24155 ;
  assign n24157 = n1661 & ~n24156 ;
  assign n24158 = n1665 & ~n24157 ;
  assign n24159 = n1669 & ~n24158 ;
  assign n24160 = n1673 & ~n24159 ;
  assign n24161 = n1677 & ~n24160 ;
  assign n24162 = n1681 & ~n24161 ;
  assign n24163 = n1685 & ~n24162 ;
  assign n24164 = n1689 & ~n24163 ;
  assign n24165 = n1693 & ~n24164 ;
  assign n24166 = n1697 & ~n24165 ;
  assign n24167 = n1701 & ~n24166 ;
  assign n24168 = n1705 & ~n24167 ;
  assign n24169 = n1709 & ~n24168 ;
  assign n24170 = n1713 & ~n24169 ;
  assign n24171 = n1717 & ~n24170 ;
  assign n24172 = n1721 & ~n24171 ;
  assign n24173 = n1725 & ~n24172 ;
  assign n24174 = n1729 & ~n24173 ;
  assign n24175 = n1733 & ~n24174 ;
  assign n24176 = n1737 & ~n24175 ;
  assign n24177 = n1741 & ~n24176 ;
  assign n24178 = n1745 & ~n24177 ;
  assign n24179 = n1749 & ~n24178 ;
  assign n24180 = n1753 & ~n24179 ;
  assign n24181 = n1757 & ~n24180 ;
  assign n24182 = n1761 & ~n24181 ;
  assign n24183 = n1765 & ~n24182 ;
  assign n24184 = n1769 & ~n24183 ;
  assign n24185 = n1773 & ~n24184 ;
  assign n24186 = n1777 & ~n24185 ;
  assign n24187 = n1781 & ~n24186 ;
  assign n24188 = n1785 & ~n24187 ;
  assign n24189 = n1789 & ~n24188 ;
  assign n24190 = n1793 & ~n24189 ;
  assign n24191 = n1797 & ~n24190 ;
  assign n24192 = n1801 & ~n24191 ;
  assign n24193 = n1805 & ~n24192 ;
  assign n24194 = n1809 & ~n24193 ;
  assign n24195 = n1813 & ~n24194 ;
  assign n24196 = n1817 & ~n24195 ;
  assign n24197 = n1821 & ~n24196 ;
  assign n24198 = n1825 & ~n24197 ;
  assign n24199 = n1829 & ~n24198 ;
  assign n24200 = n1833 & ~n24199 ;
  assign n24201 = n1837 & ~n24200 ;
  assign n24202 = n1841 & ~n24201 ;
  assign n24203 = n1845 & ~n24202 ;
  assign n24204 = n1849 & ~n24203 ;
  assign n24205 = n1853 & ~n24204 ;
  assign n24206 = n1857 & ~n24205 ;
  assign n24207 = n1861 & ~n24206 ;
  assign n24208 = n1865 & ~n24207 ;
  assign n24209 = n1869 & ~n24208 ;
  assign n24210 = n1873 & ~n24209 ;
  assign n24211 = n1877 & ~n24210 ;
  assign n24212 = n1881 & ~n24211 ;
  assign n24213 = n1885 & ~n24212 ;
  assign n24214 = n1889 & ~n24213 ;
  assign n24215 = n1893 & ~n24214 ;
  assign n24216 = n1897 & ~n24215 ;
  assign n24217 = n1901 & ~n24216 ;
  assign n24218 = n1905 & ~n24217 ;
  assign n24219 = n1909 & ~n24218 ;
  assign n24220 = n1913 & ~n24219 ;
  assign n24221 = n1917 & ~n24220 ;
  assign n24222 = n1921 & ~n24221 ;
  assign n24223 = n1925 & ~n24222 ;
  assign n24224 = n1929 & ~n24223 ;
  assign n24225 = n1933 & ~n24224 ;
  assign n24226 = n1937 & ~n24225 ;
  assign n24227 = n1941 & ~n24226 ;
  assign n24228 = n1945 & ~n24227 ;
  assign n24229 = x255 & ~n1947 ;
  assign n24230 = ~n24228 & n24229 ;
  assign n24318 = n24230 & x383 ;
  assign n24231 = ~n2289 & n2655 ;
  assign n24232 = n2658 & ~n24231 ;
  assign n24233 = n3192 & ~n24232 ;
  assign n24234 = n1962 & ~n24233 ;
  assign n24235 = n1966 & ~n24234 ;
  assign n24236 = n1970 & ~n24235 ;
  assign n24237 = n1974 & ~n24236 ;
  assign n24238 = n1978 & ~n24237 ;
  assign n24239 = n1982 & ~n24238 ;
  assign n24240 = n1986 & ~n24239 ;
  assign n24241 = n1990 & ~n24240 ;
  assign n24242 = n1994 & ~n24241 ;
  assign n24243 = n1998 & ~n24242 ;
  assign n24244 = n2002 & ~n24243 ;
  assign n24245 = n2006 & ~n24244 ;
  assign n24246 = n2010 & ~n24245 ;
  assign n24247 = n2014 & ~n24246 ;
  assign n24248 = n2018 & ~n24247 ;
  assign n24249 = n2022 & ~n24248 ;
  assign n24250 = n2026 & ~n24249 ;
  assign n24251 = n2030 & ~n24250 ;
  assign n24252 = n2034 & ~n24251 ;
  assign n24253 = n2038 & ~n24252 ;
  assign n24254 = n2042 & ~n24253 ;
  assign n24255 = n2046 & ~n24254 ;
  assign n24256 = n2050 & ~n24255 ;
  assign n24257 = n2054 & ~n24256 ;
  assign n24258 = n2058 & ~n24257 ;
  assign n24259 = n2062 & ~n24258 ;
  assign n24260 = n2066 & ~n24259 ;
  assign n24261 = n2070 & ~n24260 ;
  assign n24262 = n2074 & ~n24261 ;
  assign n24263 = n2078 & ~n24262 ;
  assign n24264 = n2082 & ~n24263 ;
  assign n24265 = n2086 & ~n24264 ;
  assign n24266 = n2090 & ~n24265 ;
  assign n24267 = n2094 & ~n24266 ;
  assign n24268 = n2098 & ~n24267 ;
  assign n24269 = n2102 & ~n24268 ;
  assign n24270 = n2106 & ~n24269 ;
  assign n24271 = n2110 & ~n24270 ;
  assign n24272 = n2114 & ~n24271 ;
  assign n24273 = n2118 & ~n24272 ;
  assign n24274 = n2122 & ~n24273 ;
  assign n24275 = n2126 & ~n24274 ;
  assign n24276 = n2130 & ~n24275 ;
  assign n24277 = n2134 & ~n24276 ;
  assign n24278 = n2138 & ~n24277 ;
  assign n24279 = n2142 & ~n24278 ;
  assign n24280 = n2146 & ~n24279 ;
  assign n24281 = n2150 & ~n24280 ;
  assign n24282 = n2154 & ~n24281 ;
  assign n24283 = n2158 & ~n24282 ;
  assign n24284 = n2162 & ~n24283 ;
  assign n24285 = n2166 & ~n24284 ;
  assign n24286 = n2170 & ~n24285 ;
  assign n24287 = n2174 & ~n24286 ;
  assign n24288 = n2178 & ~n24287 ;
  assign n24289 = n2182 & ~n24288 ;
  assign n24290 = n2186 & ~n24289 ;
  assign n24291 = n2190 & ~n24290 ;
  assign n24292 = n2194 & ~n24291 ;
  assign n24293 = n2198 & ~n24292 ;
  assign n24294 = n2202 & ~n24293 ;
  assign n24295 = n2206 & ~n24294 ;
  assign n24296 = n2210 & ~n24295 ;
  assign n24297 = n2214 & ~n24296 ;
  assign n24298 = n2218 & ~n24297 ;
  assign n24299 = n2222 & ~n24298 ;
  assign n24300 = n2226 & ~n24299 ;
  assign n24301 = n2230 & ~n24300 ;
  assign n24302 = n2234 & ~n24301 ;
  assign n24303 = n2238 & ~n24302 ;
  assign n24304 = n2242 & ~n24303 ;
  assign n24305 = n2246 & ~n24304 ;
  assign n24306 = n2250 & ~n24305 ;
  assign n24307 = n2254 & ~n24306 ;
  assign n24308 = n2258 & ~n24307 ;
  assign n24309 = n2262 & ~n24308 ;
  assign n24310 = n2266 & ~n24309 ;
  assign n24311 = n2270 & ~n24310 ;
  assign n24312 = n2274 & ~n24311 ;
  assign n24313 = n2278 & ~n24312 ;
  assign n24314 = n2282 & ~n24313 ;
  assign n24315 = ~x255 & ~n2284 ;
  assign n24316 = ~n24314 & n24315 ;
  assign n24319 = ~n24316 & ~x383 ;
  assign n24320 = ~n24318 & ~n24319 ;
  assign n24321 = n578 & n948 ;
  assign n24322 = n964 & n980 ;
  assign n24323 = n24321 & n24322 ;
  assign n24324 = n514 & n530 ;
  assign n24325 = n546 & n562 ;
  assign n24326 = n24324 & n24325 ;
  assign n24327 = n24323 & n24326 ;
  assign n24328 = n1060 & n1076 ;
  assign n24329 = n1092 & n1108 ;
  assign n24330 = n24328 & n24329 ;
  assign n24331 = n996 & n1012 ;
  assign n24332 = n1028 & n1044 ;
  assign n24333 = n24331 & n24332 ;
  assign n24334 = n24330 & n24333 ;
  assign n24335 = n24327 & n24334 ;
  assign n24336 = n322 & n338 ;
  assign n24337 = n354 & n370 ;
  assign n24338 = n24336 & n24337 ;
  assign n24339 = n259 & n274 ;
  assign n24340 = n290 & n306 ;
  assign n24341 = n24339 & n24340 ;
  assign n24342 = n24338 & n24341 ;
  assign n24343 = n450 & n466 ;
  assign n24344 = n482 & n498 ;
  assign n24345 = n24343 & n24344 ;
  assign n24346 = n386 & n402 ;
  assign n24347 = n418 & n434 ;
  assign n24348 = n24346 & n24347 ;
  assign n24349 = n24345 & n24348 ;
  assign n24350 = n24342 & n24349 ;
  assign n24351 = n24335 & n24350 ;
  assign n24352 = n1780 & n1796 ;
  assign n24353 = n1812 & n1828 ;
  assign n24354 = n24352 & n24353 ;
  assign n24355 = n1716 & n1732 ;
  assign n24356 = n1748 & n1764 ;
  assign n24357 = n24355 & n24356 ;
  assign n24358 = n24354 & n24357 ;
  assign n24359 = n1908 & n1924 ;
  assign n24360 = n1940 & n2381 ;
  assign n24361 = n24359 & n24360 ;
  assign n24362 = n1844 & n1860 ;
  assign n24363 = n1876 & n1892 ;
  assign n24364 = n24362 & n24363 ;
  assign n24365 = n24361 & n24364 ;
  assign n24366 = n24358 & n24365 ;
  assign n24367 = n1188 & n1204 ;
  assign n24368 = n1220 & n1236 ;
  assign n24369 = n24367 & n24368 ;
  assign n24370 = n1124 & n1140 ;
  assign n24371 = n1156 & n1172 ;
  assign n24372 = n24370 & n24371 ;
  assign n24373 = n24369 & n24372 ;
  assign n24374 = n1652 & n1668 ;
  assign n24375 = n1684 & n1700 ;
  assign n24376 = n24374 & n24375 ;
  assign n24377 = n1252 & n1268 ;
  assign n24378 = n1621 & n1636 ;
  assign n24379 = n24377 & n24378 ;
  assign n24380 = n24376 & n24379 ;
  assign n24381 = n24373 & n24380 ;
  assign n24382 = n24366 & n24381 ;
  assign n24383 = n24351 & n24382 ;
  assign n24448 = ~n24383 & x384 ;
  assign n24384 = n917 & n1287 ;
  assign n24385 = n1303 & n1319 ;
  assign n24386 = n24384 & n24385 ;
  assign n24387 = n853 & n869 ;
  assign n24388 = n885 & n901 ;
  assign n24389 = n24387 & n24388 ;
  assign n24390 = n24386 & n24389 ;
  assign n24391 = n1399 & n1415 ;
  assign n24392 = n1431 & n1447 ;
  assign n24393 = n24391 & n24392 ;
  assign n24394 = n1335 & n1351 ;
  assign n24395 = n1367 & n1383 ;
  assign n24396 = n24394 & n24395 ;
  assign n24397 = n24393 & n24396 ;
  assign n24398 = n24390 & n24397 ;
  assign n24399 = n661 & n677 ;
  assign n24400 = n693 & n709 ;
  assign n24401 = n24399 & n24400 ;
  assign n24402 = n598 & n613 ;
  assign n24403 = n629 & n645 ;
  assign n24404 = n24402 & n24403 ;
  assign n24405 = n24401 & n24404 ;
  assign n24406 = n789 & n805 ;
  assign n24407 = n821 & n837 ;
  assign n24408 = n24406 & n24407 ;
  assign n24409 = n725 & n741 ;
  assign n24410 = n757 & n773 ;
  assign n24411 = n24409 & n24410 ;
  assign n24412 = n24408 & n24411 ;
  assign n24413 = n24405 & n24412 ;
  assign n24414 = n24398 & n24413 ;
  assign n24415 = n2117 & n2133 ;
  assign n24416 = n2149 & n2165 ;
  assign n24417 = n24415 & n24416 ;
  assign n24418 = n2053 & n2069 ;
  assign n24419 = n2085 & n2101 ;
  assign n24420 = n24418 & n24419 ;
  assign n24421 = n24417 & n24420 ;
  assign n24422 = n2245 & n2261 ;
  assign n24423 = n2277 & n2471 ;
  assign n24424 = n24422 & n24423 ;
  assign n24425 = n2181 & n2197 ;
  assign n24426 = n2213 & n2229 ;
  assign n24427 = n24425 & n24426 ;
  assign n24428 = n24424 & n24427 ;
  assign n24429 = n24421 & n24428 ;
  assign n24430 = n1527 & n1543 ;
  assign n24431 = n1559 & n1575 ;
  assign n24432 = n24430 & n24431 ;
  assign n24433 = n1463 & n1479 ;
  assign n24434 = n1495 & n1511 ;
  assign n24435 = n24433 & n24434 ;
  assign n24436 = n24432 & n24435 ;
  assign n24437 = n1989 & n2005 ;
  assign n24438 = n2021 & n2037 ;
  assign n24439 = n24437 & n24438 ;
  assign n24440 = n1591 & n1607 ;
  assign n24441 = n1958 & n1973 ;
  assign n24442 = n24440 & n24441 ;
  assign n24443 = n24439 & n24442 ;
  assign n24444 = n24436 & n24443 ;
  assign n24445 = n24429 & n24444 ;
  assign n24446 = n24414 & n24445 ;
  assign n24449 = n24446 & ~x384 ;
  assign n24450 = ~n24448 & ~n24449 ;
  assign y0 = ~n938 ;
  assign y1 = ~n1620 ;
  assign y2 = ~n2298 ;
  assign y3 = ~n2482 ;
  assign y4 = ~n2666 ;
  assign y5 = ~n2844 ;
  assign y6 = ~n3022 ;
  assign y7 = ~n3200 ;
  assign y8 = ~n3376 ;
  assign y9 = ~n3552 ;
  assign y10 = ~n3728 ;
  assign y11 = ~n3904 ;
  assign y12 = ~n4080 ;
  assign y13 = ~n4256 ;
  assign y14 = ~n4432 ;
  assign y15 = ~n4608 ;
  assign y16 = ~n4784 ;
  assign y17 = ~n4960 ;
  assign y18 = ~n5136 ;
  assign y19 = ~n5312 ;
  assign y20 = ~n5488 ;
  assign y21 = ~n5664 ;
  assign y22 = ~n5840 ;
  assign y23 = ~n6016 ;
  assign y24 = ~n6192 ;
  assign y25 = ~n6368 ;
  assign y26 = ~n6544 ;
  assign y27 = ~n6720 ;
  assign y28 = ~n6896 ;
  assign y29 = ~n7072 ;
  assign y30 = ~n7248 ;
  assign y31 = ~n7424 ;
  assign y32 = ~n7600 ;
  assign y33 = ~n7776 ;
  assign y34 = ~n7952 ;
  assign y35 = ~n8128 ;
  assign y36 = ~n8304 ;
  assign y37 = ~n8480 ;
  assign y38 = ~n8656 ;
  assign y39 = ~n8832 ;
  assign y40 = ~n9008 ;
  assign y41 = ~n9184 ;
  assign y42 = ~n9360 ;
  assign y43 = ~n9536 ;
  assign y44 = ~n9712 ;
  assign y45 = ~n9888 ;
  assign y46 = ~n10064 ;
  assign y47 = ~n10240 ;
  assign y48 = ~n10416 ;
  assign y49 = ~n10592 ;
  assign y50 = ~n10768 ;
  assign y51 = ~n10944 ;
  assign y52 = ~n11120 ;
  assign y53 = ~n11296 ;
  assign y54 = ~n11472 ;
  assign y55 = ~n11648 ;
  assign y56 = ~n11824 ;
  assign y57 = ~n12000 ;
  assign y58 = ~n12176 ;
  assign y59 = ~n12352 ;
  assign y60 = ~n12528 ;
  assign y61 = ~n12704 ;
  assign y62 = ~n12880 ;
  assign y63 = ~n13056 ;
  assign y64 = ~n13232 ;
  assign y65 = ~n13408 ;
  assign y66 = ~n13584 ;
  assign y67 = ~n13760 ;
  assign y68 = ~n13936 ;
  assign y69 = ~n14112 ;
  assign y70 = ~n14288 ;
  assign y71 = ~n14464 ;
  assign y72 = ~n14640 ;
  assign y73 = ~n14816 ;
  assign y74 = ~n14992 ;
  assign y75 = ~n15168 ;
  assign y76 = ~n15344 ;
  assign y77 = ~n15520 ;
  assign y78 = ~n15696 ;
  assign y79 = ~n15872 ;
  assign y80 = ~n16048 ;
  assign y81 = ~n16224 ;
  assign y82 = ~n16400 ;
  assign y83 = ~n16576 ;
  assign y84 = ~n16752 ;
  assign y85 = ~n16928 ;
  assign y86 = ~n17104 ;
  assign y87 = ~n17280 ;
  assign y88 = ~n17456 ;
  assign y89 = ~n17632 ;
  assign y90 = ~n17808 ;
  assign y91 = ~n17984 ;
  assign y92 = ~n18160 ;
  assign y93 = ~n18336 ;
  assign y94 = ~n18512 ;
  assign y95 = ~n18688 ;
  assign y96 = ~n18864 ;
  assign y97 = ~n19040 ;
  assign y98 = ~n19216 ;
  assign y99 = ~n19392 ;
  assign y100 = ~n19568 ;
  assign y101 = ~n19744 ;
  assign y102 = ~n19920 ;
  assign y103 = ~n20096 ;
  assign y104 = ~n20272 ;
  assign y105 = ~n20448 ;
  assign y106 = ~n20624 ;
  assign y107 = ~n20800 ;
  assign y108 = ~n20976 ;
  assign y109 = ~n21152 ;
  assign y110 = ~n21328 ;
  assign y111 = ~n21504 ;
  assign y112 = ~n21680 ;
  assign y113 = ~n21856 ;
  assign y114 = ~n22032 ;
  assign y115 = ~n22208 ;
  assign y116 = ~n22384 ;
  assign y117 = ~n22560 ;
  assign y118 = ~n22736 ;
  assign y119 = ~n22912 ;
  assign y120 = ~n23088 ;
  assign y121 = ~n23264 ;
  assign y122 = ~n23440 ;
  assign y123 = ~n23616 ;
  assign y124 = ~n23792 ;
  assign y125 = ~n23968 ;
  assign y126 = ~n24144 ;
  assign y127 = ~n24320 ;
  assign y128 = ~n24450 ;
endmodule
